`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
f+/ctYELc+/uhaDk9UPcPAJaXSQFIFZYBG60J8h0SeiQQmJRXrJaOeV3KVV/lgxJBX+Pi0uIoqsP
0dvvt0j0iw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ds8RnxyUdiC5UfagTnRdgf60gcPiiViW8hDU6PUQWVIFrIIkQkMyKnNB+w8Xr1qLiUBG5r4bOXXF
mErwm6JOoZIoBsQDC70o4vSL+APqLNFSv5xXApMJ8oplAbqfUWw9C8nrRU4CDut124eAXDPI5DeY
2JfMJZphm79HLBxzMU8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gRwcpx+s+b5LY0O8TRhmIjsPjqA3ufiQgXkVCZguAw8Z1suP9nPSCId7/spln53+f0/tJLCzfQ1D
fd2IUKNHJ4CCwxe5P3bfYOMwQGcGZYBnUI/rkBnbT4bLIULUKjdsdYIiFR4wj7A4r3rxdigXZASj
4bAQCWc/yTKuHPdOBkGm1xZsyE/cym0RYZGZH2+fxwCmec/mDDcJ/CpYhDoHMGEGbuBCGf8iBLWn
aeyZ9lCCeLqu6wdaCdWUNa54o6ZsntBpsV9wCPDRe9tE11ovPfBbXxn53PNK8XiwXSYMz8pn8OSy
qxbPTzZIACZ7R0Un42f8fBUIWh7tpxFHWyGs6w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nodK+3l/qqYipAuhJJUe0xOuCIN1x+TqZIbzLctg8etcdj4ns5ERwOiFTEWx4tFqSKSfiBrufhKt
yWt2sZ8CL8QG4oFnIznolrRNIehCN+4jyWbaGXKftDJd79ZqRspFhHLhD570bMSvSIgremGXk4v9
8wwP6uATc/QsO1FutHGO8KVpCzxvZd40lViRrR4PDuVgDCY+40pK6HkXuChY0nuCRXJET7H+tUta
9E+x1aTzVYUJ/1eoCVtOj+E7tu65BsmJ20dnWEHkyUeV1jA5W68X30ev0J7Hs51zJ9IR1Tc9k6oK
5cZGL67jAoPWt5mM6t5aS9518cZBqGf1oNIURA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
adHuDdS9NIcaGcdK+qIYLCeAIhoJ6/aK/3inFss/KwS901WcWdnwodtJYRl30WeSk1NA3ccYlgcP
qfRncDaW/cXj0qaABAOnK5VGPunMffN644DRlXhECkaoA/ySzb65JmiuN2S81Y++kCYraAnkSn1r
dHyKSUgx1u1NAyxKiVY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sq/klSwJOJjlA17FRdYxJ+Jut2VAUuMuo7xqgzJ1RKtGf6HYfMcvDsg7H1p6GKxKsxGzQnDq+TV2
yvialaGKR25jq3m+YqEvu4alVvAND91JWodFLGOnQyQ4wOlFINcRBk9iV4KuRcCu6thl6yqz+fza
9lJ0zvBITt2ks0M8BRMww70MNqtNWaJF1CC3Ni9vAu/yQQYVeSwkcK5UOnSxVuhiH8z04bmGbmYX
GiHOmU3jVuxhp2YjqPgDzrKbdsoqJhjCq4T6U3d0hobbkU3Vp5CdZdl/0SDjWcHHzcK62so6sjkD
SzhKe/etWPbsSxqUReKLZSO5LheXEkpPy9MNTg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YH2g8ybH0nesNjg6E7y8jBJXn8tIKyyE0livQIx7Re10TDRlzMmCmwkIUN5tlGSOGWmhLVQbK0g+
rKcGQQ14ncV/D+goyDwXomf/CSg8QBf4hEnCO7AC7l/rY6T9MCzXDi91k32Y9rgSa8psw1rL2tRP
V4n7LZWwLzpfKD6nULSwfOxlRujBnhDthCpfLG4IyGF6xIvXwGHiPKj7eN88s6/dLLx+cbAaF19O
87YX29ndjw5p6GNVK2qmLkTN6PXDG344nzObIwO0uqqA+FVVCZMMjZTL8g4waFPmSoYkceS61wYA
ixxKVaGor3lvI/QtRPUF1CQLzsC2AYuPvMnzBQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jvCTnMZdPEi0pS6fvoWdHBB+8zNm548wh15gSC5pcwD7WN9Y9MGIT22qU2zoAQUCxDDh/cCPO1Yv
ADLZ0UhpYD2GjpeuWT5ghd4+qHg/CkzJFC+ZVH8ykfyN62KFE3xh/MluLBCWRsCStmZJ0WYGWgUf
Z9tmSszFQIuvHIcpusuomjakCYe158ViTxw5O5I+Q+Pr5RKTSyOK+KeUwbQzEyKFWzqyleebXZA7
oqsF9JxaiyEYCepL4kzaHuS0svOYXFReS//cViwJO3phQKvtD4kTD6UUO/VVfK4cTr/eE4lDEGtp
k+LKlNS6OtEasR8I92J44GiANgTY6Us6Bt15Cg==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j5cGcfM8rqCCS6KkIv45MGGE7qR/xEFXp75tqUY+yuyLI98OR1gm3l5Igo0qt2LRcoEg4D1RNKOw
DnWeDNUo59EbHqHfiydR1fs4bfaSIqF6l3H1RQsLZBo4sI2WyMxSdByFFTGLb5Kt4TieIT75Psva
0GuLfhX8d2PRKhvO2rSVTOvN216IDzuy9UFfnJtMYeWnnhvRl/5WRu+Sz3OJbchfQVN3Cy4DX/Ni
ldwRLsO1e7pref4KcTGOk6rS1zTD9kPQmMdDuzqm7LeBRJWqvQm4c6gjU0r9BlEjqOi+Cgw4lVfF
uh1OgQ+uFd0WToDsc5z2+TxpMOrfyQgACWae6w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
UES+IZu64XTMkjqbaPltXET1OZoPBid+xBc0bRSFn7J8KxJ/pm1DLIcj2tEFoayryFgXrlB64R0s
OsKVk82WvpdsPRkuZkyn07rhrodyRmFGbBhN9NAQbYcXD2YZ0NPVxYe3CtP9WnW2W4zqDZm55raP
WQlKwcGTPFe7cBzaapbjcbaXtSaVbcJMQtFx4J5sV6VKJGwqapTRq50UDGaYufrRUF9635rw3/Yc
TYp80WrQYc/3Nbki0NTeReKlZpCkTdbb+IFJBdR2FJF3gEKIKkMvwKaqlVz6Ie0gTD0ivGqS7XCz
bKjwRvdXswDI3JEQQfRp7BnidRKcIx6q9pf5kJ/CkdQvOoJfqsy90ipPEzNpMdMC8fhSNz3yPJhs
T61l6R/S7n3euqfQBNeIGJSbpE0OUgXGs++OhsNWlmwXHcj0yoDRspmvAvaLvz1lbq+l8tsTCKov
JURzvR+NVAiXpeimkAuhPpaGtFp9J5tjEABD0Ia7ln7jYbPOgXVwdqTUhEocH8s1JdmoN3jPZJBn
II1dhuzXflhvHxfWFkeB2AHmsovc+MExuLcWwWqTuKUQ7VoAw/CfTTkR71SO9Wb1YIO1sRn1EDLy
qzMOOLMBmuITiVlh3MciLO8KQe9vi37UHUpBNz7o+a7DqkPNdFzk3XIqqJn5PYHULjeqap89WLI4
YMv+CfSNaAK5tqXMl1DSPLMgiw/LGQ3fwv8ZjBQ1sOi6RqxmPNV0LrIk+X1d+dh8zU0kmmB8u+e9
iOZ1MnvBea1+7Kkn6Q6hTy7E/ey0ZqpSEa7MMkpgvtOowC0fRYFkVJlfkHFm7ypNiV0iLNyIowqq
IhJR8NEhW6a55i8XD+ZfnxKx+nXIYj3DeyJ6eFzY6RFbhLxO4lNLmZVv29RfBrCYSESHEeFYJNWQ
BbUOaSP7xxgrKKOUJSPQVWPEdq1nKxAiD6s234uS6jm7+aw9dYbvkhOULlsyFDrQhL+DQP3EbkKx
cCyR9wdRwOHqsxvKEcXQ/jLNRo4i9IVZIeEzX9qmvtLWKVC4LQ54Dg05g+BLoMxTQa22x0qmeA+I
oprvwhBLp60QaOxvA/9UdMoiFouT/mxyVWlksYD61cv7I308S2omD8KpNtsItGuoFsdat2rC8kUm
yThdbMOBJVCs2cdJz/+m/ozgkEfaiYni0LwAJdxK2OKCFgOWYuZUjSyZTppYrH1BjxWBRNndsJCL
rDs1l930FhqsDyiAGc7KuQfT1pRK0RikHWIQw86sKtTpOfdNcn/E4IiSWXiCo7n6k5+hLX78Cz+V
niJn+EDyliwvkqnv8i7IN1pUNC0Ge5MD1oc1GYfvB39vg1241iVJxvosmRfCbnarY+mUGtQj/Zmg
PQJwnLWiNpmm29tKpPvUPKQc9+VvGEckGg/XsNr1StJxuEsJgwFen258YJQhtS8+RoPLjmSBSIG6
YdZsKcjeiunjZC6vE2S4aMZi8vmpWBmwJTCmwkp2h5oa/34C2gu4vLb8w76FkI1qq2omDP6ilfO/
wrkVyxt8PLS529agM/SPjNaEPUvwsZmYLyhV24w1w7D3pf1f4CSW/VZGlWabXzZbCV1Ra8EZWv+G
HXe1msgYyE7XpWuGGyIZK3clFmMi1xqIsVpmDZkcScG9lPFAr4hPE8aNyXXiuxM+BifHASjPrasV
S6tHBiztC57ljxkEQB3sUGSH7mWQuKzENlYze0hwoqMtj8kxJa/Q3MWM/KW3hWq4IC+cZgu2lu7M
BTB/AdhfNUHle2UQslqUwZpbjUVkYCNVRgmHVvtHWu9Ejf2rePZKhCXz7EbBRxd/HBUytqpeQpTX
5cGwUOP5OLw2fEMjEl3kLAhkU/oRivxtE/iDlJksxEwWiL9twYw6yagy+H1A0eFUjtgqchHM+Md8
u9DvEmwwMjXkzFiOL4PH1PYZc1XnFE9AUpyPXDwouUZp5kMjZmd7LHjEfWYaHg+OzQgj0MVWVn6b
6VAyhvEuONsPAeaSp+3Du3eKUDtwDB/Qc5PjgVDYkxiroJ7hrtgjfaSQ9+2HX9w5cqlOMVb3hFiV
LBnDweKQNb4py01Cy6b6rpiSSNLWBzpwB5dMWJkMnJA5UA/hy9mhkXVkngcT2B3YEu5TJS6X9izx
fsBf/KRLsW14LzT3gHqElcBR8tLRYiWPk/t9FQVYs+QQI/frYam2CpWRTcyp3SmdPNoLcAscrBYq
0jEfu1Yantel+J5cF/9XAmFg83A3mGw/3Rgaj6+TC7QiC+56MhD0awqQ24DE9S/fAKeu3A14jPQs
vVaiM7H3/jN4pB8FryrnlX43I6rMsEtsld5irrXk8w9tbfEFSziAuT2cID3keppvc/T2hDqBm2Iv
4oy9x9gWbOzQsuLcBJ321DxlI7vRMtYUzVu8+O3XjC2o6TZBHdESdh10o/nsaPooEuD1uITe6dC8
KJk9phLM5vvdDpxzLLZzGowdPLSa/3GOMAXodtwmDOHbu3t7JCTPcfk9CGKZwvw4WP45IOpoc2Fe
atcY3NK+u8+B80zEjwtLYxFcvHzqQiAyMTkOvMIYW3/1e7DYmf8sXQSt++O8LKr5XAfYHYzV/gFe
YtoqUHT2mVhS1weFpZeMUZhz+AOjO1IUZn/iWa/S1z0uZ1qBWRFfcVxwwwoGn7wPEMkN4fxn+pp0
58pICdOH6G7bDIFOVUWkzhW2PHG6ik0PenLvtbcvzBzEFSWyfhnn5ktDh/bsat+m7XbfMZUQ4uQl
Mx5YO+YNWKWPjWAGuO0AYEZucZ994hR3ZlGfOaOVzEy5dkB2Yi+AherCGpigQQRFR1flmQdRT9nF
t1AMKGmALPRSnQTtVhYckqkLipE8U5A4JgUrAOO+wqLJNhfIi0hkrnMlbjJDCEpUL6/9vBJqy83r
iTPBpMwIgPmB9qYRiLhqpFe7BDlMDPCYVP14bXVt64Y11SegzRqC3+OQfPY/JcKPf7O1osYH2VDK
bN/6sRAvRyu51uexIfHKR0mA+GfDDdT/xrNEZirF/rhj0vWULzDVLuDyWxkR045M8vsgirB9NRvx
LLvwl+y8LPLur8WIGCLSUMYTaecjSRzk09O6x8ubwDlxn/EfzYcuUE19ZpI0ibtJpL5WsHqqABnM
UGCFyM5CqBQE1Uj8RLyRV/MTO6c5hTq9c9sriu98CCS8WGzvoBzmC4ytdo65UHyog9bo4Cgllsmw
eoMlTV7O8o519OQY3ZVZlSpP6b76w9JfzvHNuQWFGaJaqC1PiJBW/rdVCW42FXOKShXxurXakhNg
fArH3hdLHs1mdu63beHfe98vQuBnYP5Ft0n9XmJQECXeQrCl2//BsjL6DJcWzhnXKfdXbe3r/hdC
8KSW/LZ9921eQvr49K0Qxjh4mPVdSrJ2oXF5O/Omp+YKMOEX8NfuBs6ZajzhsmmN9lfHl9pfTzAK
TrxPLsr6rhidA4dkG83grK4aJWeGa75cPC2o+aCkwLZOGj+JxUFoEXcNSg1/xqUNGPthJI+H4ghp
Ln0OBYYhnSMNAm0pDUWYP3ZUkJOf+pdmwK+crw1gn+un63xXytrIAWTXRkJtB2OThEW5GGp201ji
rfSl383SGUx7AMZuiU7E87prnsVSJIgmm0jBEtbKUiKADSVcDVV9KgaluFytFdTL3XmuwVaCvSZJ
zrAx/YQ2nl9gsb2pjUPKBvb4480L1WWtVy0ZQAo5ckcXAA//w+ac4SJ9sFO9MIYfGKdqWhr1GcSc
yai/CknrtORt1wCb+6anfpdU/kmO+na8trn49V4KN1Updu1PkmoTcduNVtkD8GtYOockhJHPRJy0
dTQmmslT1fzN37YViA73jMu/H70+ByTQJRq1rhjTzyBqrAGQ8B172J1sBUj5M32VWmTeR72MrX2O
wtl3Rso9eZCpXysyIcqWSigtJmxRTyEKHY/H3mmCAvhtALqLkXZinnc0m9vNUkRzmjwxf3wtFU6A
GxU+q9fjiZiHZZobXIL3ZM2xpbhTG/O1Zg/M5oqSyLzVV7L5CZl5qpR2nw4CreYKcehPb2AIs8f+
8ahiTnC7wMpHlMr9fa8Fd/nRwMsXR+6Th5a7ayV9H+ZD/LrAC2qMP2Tt7bGxbdkoy4j2DKKwdS73
Oc+YGt3JMCrekM+JBKagWccSrDpfrCeYYr7SKoZ0c0o3aQhD4AyTnhuT/PglSDwYjHAiL0lir/3o
jDAUIA+frkiV+aynvheRTB01pgOO8ZBPEJragdDtM5vVYIBwZbTkhNY6DRfF53m6s3+RIIU/HwbP
xIf14LJCWFMJuPDKu+PagtRt4UafHSgDwE23WuY4a8VHMdEckROBd+tk5KU5/ydRN/T67YuXYE+M
i2NJ0feEUepQ2djNYTyAz5LOKTmgCZUL5eI9oz39T3UxpBrGn6m9zU4Pmw7SMM/Q+X30D3U2/JeJ
4vTgy48mOTG7IjJbd/9kjrrGBqH4VREr90hspcGsx4Lsz6rcWrtofC07V05kWhrMOATRTGLx6rno
pMDLD9P03FwGW/+/3B13ldpCk5abe/d9zKGNIMRKqwgrY9pa1w5cmx5tYBK9v7DLtNiZNkeaClzw
GIDow1woI4uBHBpoXlrQ1PXrxEGpWjm7GuB8SiZRn6wgvY5N475itU0mS2xg5WRlz/0kR4APkf6o
DwyElj7393uyTK7MBVMfSdiwAs2B3QiJ4Nxm5GC1G9UsewaZyCGgs07zBCwb9UJ8z7XZmAH6zrPZ
HAsl6P+fyreUQycBOazv1n0YzXbLpSP+daiF3buSIUnp6n7ZKGtejotYQJo/ssCq6Ktx5UL0J2DL
ANFB4t3/SSnD8z4iFTVAcQp19cQO3rpp8Lyq+QNJpJD51u5kHy/W4DkbOgt+uRtB9Z/MGsOpy/OA
JChF2iJZvhQNXVAcv/Ug187Vk/YCYoxnK5uLWjRxCDeTMFRo2iAcHziwnvgs9KOqquDnd+6ZY/hg
1oqZjAqzl62RJNwOEzi1aYaKTibsmFnpWRyTk0MUs5aupvY3F0kbZgBdxlsHlz/7R7/ykbZNy5Rv
6BG4VmdlQOKYJBxU3QozHSCXMpQywYpzkiU9pJinrg1fUyfBjbfZxS/BvlKSdN6yxcNqLBhfubGX
xDm//zOwaak9fffFYS/tNa4Iq5b02TyPPXmu4KyHHwXV7hgFbcq0Q7nWwQEVd2M76j1ejl2xODj2
yhf9zpuOJs+Lj2Kr8JkvcoVCGuH+LIKkpDXdml1QvmnO8QqOkEqBGV+6kdZmfDLXwNzFi9f0mSb3
nkJ/0E1x2M/pJpsj8wIYET/Ce7JRTKISccFCScyyV2WwDK0e4CYMqrcXYIvQ/MOf9lomYtYEgmFy
LjfeYVGrpqhpMNljzn7VO7mIFkkzkQW/Tccm5c3PPeU07pOD4INtl9dxiwFPpmAewVxaBitTKylr
SlN4lLRBw4aTtbQs6a13BX/6D6muEEA/dZWHhxQzViSnZFPmPb5BW2vgMdtlhgJX3F33pD/4Qf8O
VgV5ubY1l8cIAn//E0j+rDrhGyb8BFqpC6rcZQE0OgOKONzfZx7gNB8bwgSAmxdxRf69V2TZby/H
cN6IbullrJ5WrsFsMe0seMNYESYdI3UdtbMKJkhIB0X7EuD41belyFaCXzlhX7isVwDqNG+NU3NF
HT1QyCfZFP/13Ob3Gzc9Wc8qSPzjblOC7RJxb3LI+IUR1HjEJWjsFDB+oLLBf8izVpK1dLCAqvP+
XeHjIAj2EEZfl4imVvOAL2Cgbo9yuyp1S0ZPoWXyl6N2/n+suQbCX4qo2+OYwqiTGzfD+QpD+mn0
+cDpPHZVYnSeNY9e5OE6FGsxogg0QuVNFnMmUTI3fu5J+N87j23xkLhWcSzQn90wNwI1m5FHmn8t
8p4HFJiDv8p1s1JOfg7vlmJEXNnFq/i4OUGkzdHrKTrYpSf+IAB5DrLvQ0oqe9qEEMztJWaZMFps
t66c8daSkpXz0qTQsBB4Vv5QElLFkQFNf8rGRXGws2fYMTFUUlAbOxEUN5iwdL4vzHnRrmVzBjfj
o/YqH2p8BRnKj2X7P1deYv33zD1cxCt7xNJY0BVz+KtSqgmCWJXYl5vw28M99kf4nloDluzD4Xu7
Q1me6i6qPv0x1/gj7j83GqRjysszw7sgUQVUPkBz6sHc6a3KkotgqPIkk417ewhCwE1YAe90ZjnJ
lFUivKvEscNjAVb10vhr9UkTTxmR6ehaxItP/lPNeOfi2zih8sqPKGAHZ7xJAMF6p2+TsIEfxEnD
QLzuPB560KMsGOkcFUEx43qQ/pMI+7+QZJKr+dcxtPB77JeaEoaIbk/3FNskyg7TJlxs6/tAHRDT
OUi5OoIEpiNCvcq5uJYWk0M0f0cBiE3DpAYMFC+JksAYPza9vSXC0fBEJeQyT2uF1pvE1egIm3yq
hDCxADH8oKyXLwAluDvlWQYt7fXcmG0BSaSI0e+9zhChPmHCVm679bVM/hx69wDWyRG7xT7lnppg
FbLYKhoG71XaK7cl12AutDpwWNdYn1KwTqH0/v7G618zTcPbFMPJul3PfmoTN0EDMCeUVLQ7vBUG
7V8nbthgTLo9TGVQM25m7q75aHaAbKfdUpaWfdru8F7kdPZXE9VjC1MLAQqYmvUhnyJDWKhrXkGa
5ik0JEDE6MwSMkBjC2wthwIthe1MRyOk2EhBj7v01B9YVuJ4kRAAGMHF35o9qW9yXCLnHXa05Ism
rGH0Hf28Pk0AaOFylrinqwdMlzH0+A/urMD6S2g+Cx87cbzORR41QhG86DgNHCFd+a6PPAy7baai
IV+3TYesLhcTigup4cMWKEkeY3HFRN6yvRpMvra9gJ8QAzol/aaGEA1hd4/rt9gPGOM9tyj7YVtu
Ahk0IWTxsSyuXJItOKO3WdiN1aA9pLzxh0QG/JPqRpHNk4fpMXIEvT/a3NNAhxsHem49GCqXx0I4
UmQLMALIm2hlY81wEocCroc8Z/hFPd5ypHUWnC0fi+vXKCCXGwg9eTqG9gvxYVvu6XpXefQ5Uf8O
PqRDn7YcUvDbZziYSaBewYfsi5Ynh9IPM9PKFTrDnaPJ5wZwpNCpgO1YkHCbw+yENKAiePEHIDKl
+5cBBlfd4EM/5NzahQLK8/nARf7bGz9V0NAUcRDL0yQ9e5Ypb3UnbzSrZIBusZjzD6ypGmiEBzIb
ezX8awC0CPeZYE0Dh/JWm7MFr8yS8aQyT5a2JIrMAkAqPPPKgthzD81R66HLqb756c51jp4cX9N4
jkTWayRoxaDqIKhoQ1KLKnGV2JgaVpC2zb16MNNXiNd0iFyDC+P1umlBZ20p9U2Pz7Mrhis9YjPE
4phalzTEJq5YZtK0Zyk7rHy5A6hAGShAcXyCV+/yd+vdHX9zlLbjsKQ9foFJ596FGGkvUdoIXlIX
KOSkhQ0uB2ci04PLJCh3pRguz4chTvwxyL1tse6Qox0SvQU0bVHoVtPgwuK7CQ9bbitolnyoEhjN
XAJsoADTCpnzP8LGWoSdNKxCBndu9mLAyAdq9wu1QJwcss1JvWLnR+IxdcKmMZnreW5V6sta6A9c
E4PIj58TlJ0hpVfDLkqGtgZejBPX6l+QucMrDOTVzl9q9Ue41VGGblZFeAkpdlMnJOVNt7bhn65k
ODj8DMnMc2eZfCkI+bR0FcsSjsyXDz1bZrVB7GUSzPaohZxKl6JuT3yOJZIp4S/5Mv9DBXMJHuBT
kp8X1JawQZccFF73/J6lOY8+t1OwP6WgqujPILJVfrv3bfhDZ9wTG0gvtWFpq7+PuA9bu7zDSBAI
smHP4iubjlk0eEYIUw2qJ0QPN44fGtsSgDqiu8BWyg0Flmy5/9yiycTRUEjWMfqg2w0dgSm81HUO
5GZAfZzpljXGZDysXwZVkuUp/JxUhZ6C1wehE6WIntwEomBCHXCNFhrM04in5iNT2FFeB+ETadEa
Z6B02WC6dzaKOR5JFu9Qt58Fd6XB2wXLWF0+wnPz88lCHbiRMDDdo/8mcyG0ldgeM+8zbE1bqsvK
q/PU7avI/fj8CmC/eau6Xn5VWJ+baTtgtmUWL3k45y40z84JEXOVYBagd//rGBY+tda5doZhtuiz
xEsfz0C0oGPRt1svfqrQBelPHuK+rDEh3aE/6pvf0N2+/h2xatkXsLWRrYXTyA3qu7AGNbkrvXNC
lBjKcSUUe8XCYvCygcadlUapKaID2z6XKuP9osahDAT07ireCBNQ8XBnUL8ob2emPKxfVSDPN0cg
SInkx8mawLXQcFkZG8CsO/p8AJj4xXh7viGt5zWHiaY5YIrqzPZkO3kX0xc6JBJnlf9N4zl+x1oX
wOkl6bA/KnG79cGc2/dqgAwB2vaUUXPsj66JBSoBAPqbf3ZBP1CV+KxIOYEWvsKmPejp83AerNux
UnPH8Zav7O3PJDW4/0CsLlqL3xTR8XtOgpTev+EWJzSB8yUoQpMl5hLNJdvKSEnYWPFLS5Acj9bl
t0+A/exbqe+1wd/6VbUOCZM8JeVCq/zSwH+umsZHySdWW/0eWcn4DiIs7r4NKCXc2aFAlkQz6ngn
9ewmrcHrnb+xTdaoHON0GUDCQ4T6omANUjwpjJHQB5J5r8sq0TKaKbzp6zOPWq8WXrmPzvGJh1B/
F28VF7DvHpxkG22VaOI8vyzIy9ptnJH0aPmDIwyQwT5I7U7q/4ZUdU9Kk4f4q4X4/6nnh0f93sq6
5tN4HiGuGBrl8vmLdQ0R6QFFgYRc6x3cQ0+fBVYatERuVRoayBv0Jo+rmOvBaCZ1o0SqambKtGsy
L9JNQYSTKJmEY+YTmZA3EowSUSMOHltlWhnOsZi2bg8SYVxpBB/B5fideW6t3kWbz1FKIah6Jwvr
VALL4x7WvkzAlTkWzaooM0cqky/J0W03yinqxBCyk6HXsas/Wq9uLM2qRX4rI0OLoRZjkedwdL3S
sNgiup7lnqvtPIXhZTqr+8/AfAhRSTrcwPMZmIFvVj/py+3B0a2IUpOqdDFlLYimtPzL/gbCDrZK
aj7cqI239ejRc/OuE2s5Ny2JFCQJEcqkNhAWSlmNlzynUKyRhPK/tSnKwuDwmOi/hd/nbuUtVbpl
dJrmNj+Wz0UGM1aYdrhDmacEvaCJRNso8A1XJmx/DjJqFJpq35TlpMPhAkseapgUdD6dnbBflVRS
uXdHv+3S/TuWVOwslNCUOHtAeSr9RV8rj7Mz6XEadB+uzq2T31rMt2QEtFEzgPfP+c3mLuh7BKo8
sONuV8UjsuSZsnZFMtrfY1y37kR1Y4ly02LF329OH2s+pG4RL4ZVKTWyEChdLrS1XnBVnZ03sgme
e3Z55qDyYruPAbtyeCX7kMKdyf6f43P8ruNT/0bInNACjanOsBOe/+CNbVwGJgIBsY9il3OiZ7Ae
amV5xZH4CzzJcTo9KTKGgGhwFMxMVgSdCwfZfQL5LQx8hpZm7w+L77YhPzVxlI9aoRQST61bHm7Y
aNxy2aaOVNSfu0QC0h/2PFxQTHWXWlHAFQ/i65hkNJOIUPUz/alWWtrnlLOp0E5X8nDFWPxt5Ivr
EQepnxxFQqA21a9vpCvvR2xA3YwyHcsJmcfpZDqAN/0Vu0oZyKHsG1UmsZ+o//YaU6DMACuzrgot
FfZpyuL4eTqJ+DqSwzP924PjoQizyYYdNcCVsbVmVS5pgrWPaQUs/ZLUe1EXqDuPq7NT6ZXE4WGB
LcIUAip5I73H6za+dqKnRHGkRrj2ytA1BsXWLC9u8jT+FzcQZYw3u89YntVKQp6nJ0DccajsiYOy
MlyBwjXkXOSVRwhC80GWBo567u+PdZZJLbI+HQB+7nX3Ju0GDZw5d/BxsiOuClwfuUp9dmY7UDjo
EzFax98Q/Md92lvy3NOdKwanLmmxPcC+DsEugS5Q5xM3MnB0yB/rnEFYM8S1p/zPfpItKQwwJAtk
tMU4SsZI1G0QZ9YsfV0F4AmRVACHAhvT21Z2GAbNqbr1qZzysjQbce+GLdVI5R679HNoUtLkOQj9
YQoaLrhTp8SIHIQuaEAEYAKskvNjV1XhtcPIqVR2jVkcl/st3QrbJBPx5xtcE7JIKH2muM0sIRLL
32iSzZ1kOKKC5nMuR0nBSBoaO1laTnpgf4lGIpCd+U717aMUTEgDTqAn0pQUjL1vHMWtJqkMxyAZ
uaA1fpx+TZTHZvwJY+GoyXOVJYx4KBWS4/l8+9rzOc+o18ywW5qotsABZty/jf8kzhlB8LbB6W86
p8pLTY2QAN68xKfnQIrE/+F5t8gq4OsRoQf/7MttFqVeotUOjdvL6fhl9JklaADl4n2AduDmS5iQ
ohHDdSykHicH4LuCglhktshidkOq5S4zYbUahOtDn69M/Ss0jtN91ZRyx++XLASxKbJ9sWcNKnwX
Y7aY9bXkHsdT2/s1n5onHa8FfoEMR+M4y0A5OFuY6T7Ml5CL7nGWdztaFu8YSeAQejvlXCAmPGIt
L05HT5IdAqAvCh86iTR7JNgtMf10wW0AidY9GX7Rx1HJbL2gQNwgG6n+5A7LTrTAxre+smgncLsU
WL/dpD12deBq7br2Imb55BTgYMDuy4h8maUSpp74bdq6hfpFRLpdoPuX/oc0pSPNRcP1ZZMCTsFB
Gnnr0hZVaRMjIwkrGk43cu3SsIYZcIWnePvKAgr99mq5TpI+r1MGUotZz1wlxVt1XKbRSEpOsVB4
69jazfNcB4zvgEOpZYETFx/sgf6nqZ6MQUiiWlOTFCwdW+Xdq+ID9a57cMT/6CyvdiW3q88/NH60
8J3zNxzWfsl0XyWgHLf01CsNneCnuQca3OOg9Fut4L0Nkuzv7An+nLqxyya5adEA8eYN2UNn++mB
cd27mVAj22T8lGIU6hBlZufdUvZBvgUlja49mdvJ20QsgSo4RBUH0Nd75D+JXA0oPmS3npyIClAQ
ghgK/DXzoCN21iH8jxUjx+7o3h+Kvjr0isYSMfgHutH3JMFic8YcwXEDughB0N929Q09R9UGWUjl
OZdeZpZxOzA9+VxKoGaoRWw4LDFb0CFt4/aiLblMqFhsKlmdfHloOO3ukFEidaoX4ak3L7Fge757
rnQU9Zlx58CQlL6ooUTOA7Dn5hWMZC0zfQAuKiWl0RtkeZ02BGW95pz4qr0C1sHFkqr1S9mU5+RY
fQMmyK1Wdnc7jqvkAOTlWRNwUiuM1NHPvR2ey9Q7rxyvpIisfA8xdNrHohUA9dQ4qv2gqgYW56IK
wbbuqeOtb1Thqdqz91uyPFXRG0WfqgUFHVv/Zqwen4mYXpZkdnNeo+y1yn9ezFi2pxCXUP3pU0WQ
y3b0yawkJwNyZznc7iXqDSvPFo/3fzwx58J+8BpliEes9gjVyGx673j92DbMQFBhQW+dC2knn+JU
NwaiEO+FmWvC3CaY5TYyuSfXzJzM1YgU69jgHGKlUwDG2e6LPiggQ+OgJcFPjnQ/lVfpIg8Nl2fv
xvb8WuMwuEJhq4XZS8wgok6tyP9p4wkxMJzDXN8O43S7LVzFFVyT5WTBGlukXTnf2Iu5Yl1PCaz1
qot89g9EOhMN3jMrJTkTjgeZkfrKaLZ/yoqpC+EeDMaGMATj0x+vXgAa9QpsKWTkENyfLNIKkAn4
yg/gBnwBhx/vE6Q70uSFx743S/wKFh4RHb0WZTRu/tkRORq/bL35LPE4gnFE2jD35T8ez2PRGk5L
tg9ixB8mF8VIM32oQLzSLzwifEYm4FYBKhfSPLYEgcaCVbDWwUCuRdu2H525tZj2CCRl0nVgx2A5
hl5810VY2B7PVBDJiyy9m2Apw79T+BRepJkZuklyxO5bvIngNKXGEAtQSIWyiziqquLXP1tdhUGQ
Q2xd5Tf508DDbYA7yUiPJlm2Bj9GaARWhWby1yxchnjfvzx76CDRnwVMRMiVLmUMJ8hHAvS00oiu
Ra1BR9WlfWqDm5B7YnNWMsoznrTO+W/UOSghw2LIp3FJuFBl5TLmGonv05fGvycyFhmWgjF2OLyn
Dzl9uxJRe8zDoTOPyBMl+6ldBf0n6op6TzNRkNwJXlvyNdrz8mHdcbHB8HG9SOpSYDyqO0VjY8Wn
Ks1/g6HbfxCGvyiTO078WHQpdmJbY9kB0In1zCr8kq7JoVOu97MsWSKIYMNwgotiUrv+n+VcdPQC
BaTb7kRI8lJKMfQWswXOKO6VCIYapaFnNBma1Fdyd8by7ok0XCHFtGsBIIqY09NWf4t+83un21I0
Qhe/eKYpT0TB3x7uRnZ8W355aCtg30D+70r7MBWigF7LOS4IX3Ohu1pQl41qDSTlFxGb1bTS2EIr
ANa90MnkPBPPXw2j+CDmvtyRG/7WCDkWwmVhZXu1EpjHfdRAYEQe1gNORvrUsffVk9mzGSjnanBv
ncxD9UtIh/yw7pCKY+Iap0C5yvcrDl8fzkWdc9cNTZQLQD/uKoUCO1aB1yXFRxsp0n2PSwWMKllu
LHSpfPtWYywiIyiEJFEz6wF6ZK6T87gWv1uBk4CFV1VrHXJlqyj/8jNsyL0nWXI/HYgODQ7egsGW
PyedVlZx1ScBbD3F6HEDOYnLkLII9YPiWtag+FZPWfnGG8/pYSXqDhFQcXdoE9TPa09ah2CndG5Y
d68mndUvqNVqTotRxoSJFTYQwPGGaok8QPlKLLx5jtGp1lbKvwBmW4U4PaCqFe+jiRp0nIpSLCHL
jBJLzkkAs3WgxC/1/L1o3fSaYNfOq7vVRzT9IW+zpn6pibuVYRtIHXt8x2443SS0E+WtIC9ej9t7
akfS/jO1oOkUengYiUZ8LMftHSXtfYu14wlVfCuFF9cUac2jXwvZoQ5tmdRmwz0h1vqWT9toE1rf
EOn9CBQRasrtJ0EdFA5gP14uQWjxjoQFtTaXrsKMOjJ+YCp966RyQfrFzXsFvBHz4Q21FEoWmurE
rUvCY51/qbnpniHY6rbCA0tJP8fbysuqm8n5rzZp4ijGj+6Ov7JHsEh5G2kL85z/LEsAkfmPh28M
56ursY1Yh/IpLKRqre5oSliz3vYLioeLltwdjVIHkqu/DZBGh1J1A+GdYJUALcv3yl+Xt+A4ZGeJ
T/+RhCuzwl2aXXKRNpJQ1Ojt3ZKo4uSApkdFrWS9z20Rll3nHW6530P5w81PUgMxrw7jabtdYKmo
1Y83SLPQLNGpgZgBpeB85t4A/awZ5MXSNA1YCVKD2hbTccAiVMDucg1eZ9IebRr9nv6ImgCmc3Yy
2jFoYXnctNmYfnWNTY2SF+QS7VMcUDWBtwhSLSSVKBOGg9hfoRK5pwVjBXsqoAo6R53+86DDAhE1
cDYAanNLQYFA2JAXSSwpWvh2J0FAGT+RKwtUiqVH91kbXFCFbjo1GnnOHkbekUuyOYVncDAKeSdF
uKz0TuY08hyJYWcGP9Pj79bSverFmoWSsMrWMxdYmpbNkkkfwz/pLpfaEKOwCv35ZcgGyHm+iXpZ
BhiJwhlnOONV1zHn2eegSqFnj0qzFCwdNzNxuEplxNYDhXIDgo14L7oyxK/SENQyIfgs1kUHScob
iP+UyMsSlZIorUtflcV/5jkkNDWfW8Rs/rbgm848JCOJVGEs4er0/q5RQCEECE0RIpv6zSasURQi
47D56jmMhDBBTYBSsKLD7k4SJtgv2lUCxv5VWxGohXIEuqTPb3Dy/OF35ncZLG67bOajUd75TLhq
cJk1hoi4gdq7F/tBxxQU6t49cVsXLMO2PzUGRoeZVjOSFUEUgUerIuORIMMHleXmbcg2zZlC4vsS
JL4LElGATJC0DfgRfPJIctdWxXc036A3oGgu0/dpzGgKKPoqABje/dUN2EvavFETFkcl1CCeuLrr
GArS05dw57Ef/JA9TAr9k33wGM8N3XNEIlJuMjxWMDvxSjNrQjiZ4EfDRthZYxsirpIoSZvZZHra
ow7uZgPfahzrS+6E/8aPsHKXsUOW7G4wB2zx4DsmsMfyr+1cvEYYwQ8/V4rgif7/E06hMEASDM4b
8h+lDjt/YqHA2VFDUI/p2VbysHAKGdUfDb2qTI7Ya20S4rxAf9gyatdsA016J5T976YJg2gRvqBO
gbHHF52gUgIFtHm4tzFLj5fEsbMv0nHAq5LTy1QHDIXz4x2lasQN43Dn9XfOsN8RJ8lE/LbnKzmB
/UdIjicCq1g3Im9d4DxcB0VqcP/xgfJ29w9Jrf4dz8mycf4my3+RCK2z4euOCVhAiubjhojFvzmY
06/RQ9v2FfSFNcA2VwLQ8ZBDim0Q1pvjkY5I/1PpcW9ZLqtDTicpKynf/Yq+QQNd0YsVRtCo+bDd
FYefb5biInlc3MIcr3yC7i4zUblqbvbHOUYBHkZOGkBOlQ4MHpKl7HxJvLoAAl4uc3k15eyxpZln
NAFlualv41ziphaYLV3tL9IfrlVyXsheuKron0Mn0RDA0sHgrW7ce7vy5qge3AVCLFxneuGHq7Sl
FAVDuoWESiIhl3btXKYFB0abzz75TcTSL3ZYiHG4Ox46dnV1I2yh7TlZ+41LALoF+zJVLWSeodZy
6sB1OPWCp/DR9rm3qNurmlNK7G2G3hS9C9YlVpLqy70EUlGWDu/0BbN/fRmcfs1IQFL96p4p8A/X
ZMKTqfK0rjtOe///x/dDRz4x6il2jEEyzr9OXANCOeAOBzs/+bbh4NHXQU0aWKb/DrrEi79iCGeV
b7eS9IF2IQbCqFpH+W0kK5WQ/vnoJE9iKGv3xRsRFTpem+ZRM8HEgwINlWrOBlW0p4GEBQ29ZdTp
iLoUXy0XklWSgKnVY3lW24gxEmjjpliKI9OwPG6VSA0nAljrHXZvRqfLoor6Z4KDV59jYJ+/najC
2aYow48o1aYl6kTvvfkQJjXb9HTo0l1y8eN+MYKCjqFduXeXgk2ttWJax2I3wIBR5GrC1rSgJZsI
jslHtlkw432EqHyeDOhebc5O+nQQe4TtXzJX1DCVml0ux/NnMOq0xEFWRSn+CBv69opeSlB3OvHG
/TjIhsAk2SO4FFh6mb1nszooQ84qkdJPKgOaTM+oPryNHcKCNgq0GJjeh0RPrnIC5C9Uxs39UdlR
ujpr7/nHS4TVq5nJT1qkrgusE6s228RSSbb6nMjaGnYUb122EOqcM/QNkFp7sNNXThXl615qcyzG
2jLNonCngw2EQaXCCVVvpAtrtkahB57UQKc+AIt7ReH+3OI29Dx0lm2mh+BAMLzInNHLKDGNFIKX
kIR5YAHLlsgvtFYL1YK6SnMGLcwMgCKmBINhxhy7gF3vlDKhD1ATSFVUo0UFT0U72OXuoQ9Wwh/p
DvnCDf6FZFyDr0nqi+8BDQd23SSuWqYKEQ8fJ9SeCZ+CpeIjLsymy0E9lahBVovhyXhB+f87wqws
gN1uj5DeH6bS/+I9nCxZjVDowm4emaC02ssA1b+8LtHAgQB6zRYnKjrXHdvRBu+Vdjdx+j/W3vGC
/Gkgenl3adQDnisMVL8uq6YM8ktgiXQ3JRVXBmEWxb5wHxuyV5tGuRHJXb/fNc8m2hAzO1ZTZxYT
G1jkWsx3nNVfJjfuZri4mXmxO9Evy1aBMFYbRyrfW27tuRdY2MyPiwemiGdNHqt8K60zjdxmA9pn
DI4R4ueMazhXhJEVmjgpoH8Vtr6NkQHLSJcwLVr1WjEd1Ty97kLhl11NcdiepHBuPljYHpRGc+sh
foWsleXeJhsiWThLs95NCd5vSrrE32IaTZaLgKCdywGcieTwX+qH2MEVNvSd1W9l7t0OzGk4+HvZ
yAP7flSmlzhicmo5N/fIOfS7kTMKp4WGv4Fyy81hNtEKRd2YShgjuh8o2cT6VRcXZ/NF4QtlUAks
ilbu09E+fjl3tySrSjmAwLUWsJS90RL/pgVq4IHsMMBkasjQPBTLX+DSDGxFlIYatkLFaISPLnao
N1FezcmWh3QHwhhfUESrwUdPoUffmEvUYt6bbT4s61LVYU4SOpoS8n8EtNOryPwhKSY8ZAGvwjOu
x9gZIeGsNG1tPpWo/zdE1yonMpMAmUGFb6njNpq0evORLmFv78qC8Xbo/6jeUdIwqO0xS1omkPhH
RggZJdttQTXlGYuECW8i6ylgDQzyZWCLKFryLgNjim1nh/QEtN8zNoCElKjDQyrEzmgg8y3xRYbZ
EdB1l04m9y2XPslkrm+H7W8wuIfr9PkT9in3QXtI/A6sKqtsuPQDxTn8yhDPBwpqOSH9AX5HpheF
foJa4XLBvQ37xGuMs0I8jyf9hP2T4QnUrOvYmo0Y+RQWMk7chKNLvilDjSz7ikud4wiiz83a1TOa
8lcs6m0udAqIsTw1HZ+RI852qpqhb9zsW2hy4Yd4qmHJkl4VQvSFEf1f7q4uw5D+Ssuckg6bjoG/
ReMOcmRXpMdL98Q8bOX9O/x+JzswbxmwO2ua8N28v9IBc+fHimn8OrrYjepcbWYj7Te1NeFSFPwn
Bsq2w9ZE+OW8kPlre8EoiVXFA+KKt8oGipWr4qIlzm6MLdKfvZypysPa+/h8p7rozLx+tLIn7rGk
8hVTkd9FbEC/FWGmJiYHE7xeTXrfvWJ6PzUY8dfG5rnmRXVOiKJ0cHOVgbCAx8088EMpxHh5DcbV
+lhG9QDSlgYWntQtMxB/QAdPdH9AK5gUYkbxwLdk67H4oL9PaKOxx6wz7WSEQHPDJM8isQd3h062
llcwFlDqksyBmF69ogjNqVX+KJFgAV66EqKy9XYDNCPpD7ERz7El33adf0/6Y26el5mDeRdCB7hW
EL6znhkB3/WNT6Ptsn+HW0YXmHRo1LCqeTfg+GDCk5pJwT2Em3Jzuznc/c0UiOrs4Qoyxf4vCAC7
kzy+qMNBU/JCmC1XCVYMI9bxClEMqyEKmltW9B62RII2y1PwpSXCdIpXMXdTOvDo6trUljT4x0KM
PHwxAEXAw9mE85GhsqAlUZyKXg1R2HIgBOay78jsifvzb31dGmuhouq7cPCc6N0RoYiWkDWSM3eW
68mcWj/3NkYpkE0kT2ySamgMl/iClEAwU37s5aaoRkNz88mHZtLDpLvS6KZ8qLW2mNR+Vr0IBPCN
X1FXeIif0qRxYELgQsZnNy9heGRqdquv8iQf9EQcCD/xgi6nPWrKpodNosLl1aj91p9UbqnBCzpG
I/yvnRBK6N8st4qAUZYxz3fP/8cTKKqrHpteDi4hG/3AfeNkiKpHy4b6mwTr5Eu4xbc7dE3jhH8U
fLnPbuhGI5QX0raBEj5faFJvAkHpTPb2nflz4LzyCeFmrwAdRsmVH6IdgNbJG4jHJU6PZmZlnqZH
XKe+9J013yQTSCqhdNodmQ3HR2Zj46DASoenMtBjP41nO2oAOnrc+z9kDIyw+AiH0dsjfj4VJ2Ts
+hhXutFuWqxQ2faybNzSgzj/eOGDGb3d/ES8xfCougbvpzY4chCbImiSwTKXa0RgOi17FKAsFIPy
YigMADkrceCyqRcP07Sff9K8uUdk+2+L8d+cTEU47PgSK1Fn8D62fe6yGYm/6Ff/vEFP09TF4CpI
5yybxfnb5aDdJa0Xce+ikb4JLD28rTugTgFuhMIZQ7eynPdZMrahKzWb+bbLdWDSGPc+5cwKHfKL
8aMoUB6hZ4N5LNXGwO/MdgeTPt+pvBL3eYj8NA9h/E0ojZu1v6mIV84eF0NhoBNn4YRSVb2wTU7n
Ta0Yd1BbihswvZ2faMDlYBIgQRmJEjv7lYaar3fMdsiuMRLhtJJIEZL8M/USJz4GV4r8mfY0lYMJ
44BAmM2h2FVnSWiOHypNG23tp7jaNsvEdrstPN19fYmE5p8rTf9ipRzvUoO/i9GLIIcV2m7qK1Pl
FhWaqlzWFZHGCJDEoBxa6jy9QCUFeRoDonUo50T/AFZkLOnYqs0oHec8PlXipCtl4jSEzMXIhCuV
yfc5w22cG0TaL1YA/BWjH6GR9pzORVthUSd8Hne4jgMQBpqbTXbOXvdUlJcrqLIZqAL54S0fMP4Z
f4bPLqyJKCZbOzn0mpdlGXnMIA4F8zDmTRg80+3wIYeg407S1u8wPy9zTItFyUaMxaYbZPYFqnfF
mvoCqdH3lDu1dXiJaWrwJPg27zLuUdtezYSbD3isLZH2X/w4n/Xra9IWPOmD8EhYW+3JtyosBZ1s
p17hg2uvdGmcKqZkkXG5g0RAAhIqBwOBPDLmUHMZvNI6+kga+s8jk3kaE2nmpdt7naC9GNQSBBnl
rlr5BCUzSkVDK3IfvE/S4yezBWzZT2HKQDjv1b6EhUeg88Cx9La0jnfsEm4CR83Ch6ItRhds1LOP
zmJNDtctZnVz+lWwGNdw5KFTmormDxLJD5X601317dbW+Ri84+ZYaV9bNw1PL4w5B3Gxa1C7jIqM
DftGwwlMYMCtCCqdIoK+sFpwCoDwzy/Ru5qBKSgcFkLSaKtPDKA6uaYAgr9XmM4TycJc/kKAdoUW
5zbl/amuiG9pwIyJEddRUJcKvx7neBqr0IJ6o5hY63B2+XkgQeLwzSyXR1wz5eFXUrI4N0xb3lP7
FuDUGXzD2oxF5mBdQwK9eb41Z8ZSfYHoqctSgKb0vfmouTdybwrO5nQY5VreS1mH8G7YyVOtdoBW
nOlpzGEpRTMSKDdGahua/TtR/kMA315IqsHLy/0S3jB1RSUG5zxPfqqFjdjfyqw7fqCgss6ypOJP
yvApLfJVRSiDLqq8salDC5tfejltojRQFmzW91SpVrALFLh97YFsNa7/t/Xv3qNPqMpicioeMkzM
aCJocHSEqScMGJDJ+J9Q8ep8VKB1IAwC/2FpI6eFc7iam+YAMyuhaoUfSZPRDK4UmqEPHg3dj6Io
3j5k1NmhtKgq8+Aumj43+vJR/UiPKq9COQY3xwhOG5gPwuNAtQxH1ojvX7hkWc2bBwOJW3Z64fBv
x2vm5cy35HqkfWC0Yl9zeRYy8MOfPfXf5bOhxAtUzASGt+3eIm1zjgIHsJjxXWbJMs/ovoM6oKyK
Su8/tHxngqxmE/5qgZDZmR8bTWSvKX8AdnWETPLXDqAQG14Yur4T399K26s2GVmbr07Di0Wfs4yt
AXO54O19QGVC5eVwW/yqncu3+NawXGdBI5DQIGNJWc/3I/CaH2r/D70liJctOPcdTK3JofnRB9v2
CBoRNZK1LtUJ3fY4V/z4kKJfhOmG8jYFRubwl2DmaG9jkw9ZQscOc6E5dUZ3cPsmPAtpjU4AIZNz
hGdcGL5+f7IhkI+LvmUuJbMPkC5O0IIQXRsBqeAl63jhu19JLTWD10J/tsjIkX2h2LRY0PFhtt+B
nulhGh/Fs14RqgW3fdgmi8woZU0Fl5J+VrkCM8DbkbX1gTbET/cXh+QQ3mkkNxZyBQHZQRu1xkMI
y69fNspunBLnyW3u4Vu5fZR9NAmIEUl+u6fIbXlygdIuHrEMWUL46ipZ0uKEL8MzCYcmkSAS7Mzo
nRjSZvbhcQk/KtK3CihthbOOuv/tpGUwabIj6zQSdBiHhy7P9FJk7Hdd6CNk4v02QMyd357rWxYV
M6ZCW0Y2gjaANhqp4YFzgOPWMwkVXi1Tli44chDEYF1bIVvMNw3fIgoNAStU8s97IpfETqrS7BGX
X9s4i9wP5Giwagi4MDVrdLsPqMTDFsfHKN8FPCWe676C5AKDzdthHQHcsne3//u5CLBmwSSAYbyw
AY4ej9BQRgtmtnSByiwSQDw7sJAKVuNR5p5/Vh/G/lOUv6z30xZJHC8rge0UBX+pQZbYjyjnTqbx
b+ITDX3uwOsSj/UAgnZyXGdFdFO9AIiq7Hw37An+ni0MQ+pyu1cIgGr/8xxjPnx30kdJu7Q9aKp6
TR//ZpJrTXwVapc4EVsdb2Tf+O8Kgx6nM6k7TpW+Qpr165M0cNVLRHzvuLe1DCuVGLuR+p/ny2+A
SNWPyT466Jv6ZNH2vGySl9sW+qbmSjWFgAZo2YEvoZ5EveSmvaVWnve3NdHJ1c2+lsOKQlOfDqqt
nkcEj7qL9D0FDleQqTH29b6no73yizc9CnxL0ZqI0DUDBsLULX2fx4bhW2ocJe2uahtsdAlDr8Ae
4b35G6mnRT6sc19fnSynRC2CYYHV0qm4Mjl3ZN2iLURdvhGfyC1iDGt66xUt28PmL356e9KRjaUR
dq03cn0cyQEEb5EbGvxAcezBJ6nqcigd6G8kdrbFp2Fs6pL4LAki8yHT3Q7grpd39+zSxwdux9EJ
BeNghtuvuYxm1kSRXEuBZmgRrJk/cLN1LQHoOd5zbJwGCC7Eaj6WpLwXDJCZjRS+WmtEnZHVsBQX
87jAnqyVcbeQtE8dXMz18oWpD8yQNvZ+VKBY7hsSE4L5KUJxywxCtmIsoxpWrcbzPsIH2iFWkdVp
clHVFdyOpHvpg6ERoncXNSrE9nWEeMEdaxbIIMM5ekhCSwDSKkhZHQTjSa4OnUlYk8jP4bxHdFPb
uu1AY+nCbd9upgiX35rOYJvzEN9rahewuOY3VwSU4BQx+50mMSKARzvME3KpSoVXVEx3RyopJ/MT
fO/kVhXXzPIY6bFa81ve9SKSHQNMfyrgEtYDUx/j7CotEavy7Qum6MOHeBBuNNf4bYBC4enB+/Bt
p9z5lI3LQzkiBRFY40MROe+DR2GEPq6LDEAKOEXyM5xNDHnGv4KiqKorqrIHtCkQIs3YD9+PSDrE
Jy2JjXo2ksfUHyt7QdJXy1YVYMB3cjfT2U0WcsIQu7dalqTUTsTKAPhypjLB7IIjaYKCejp/XIa1
hdhGwQuy7N+n5QOFlxlvybxRm6hIVPtN/v23FvuuR/T+L5OK8NYh88NyxCuMyu5sloRbZUAE406O
5cParq2uKSt7ySdZYxHxT4hhUaY4fcP+QVbRJXOsIEF08VcY//km0AjAJi8ESe4V2/O7pxwXZ2hV
5AK2J1DUZZATyGbmV1Hgj6cfJeAMf0LJyfyCksbf5MstKzf/1tTNQacSvhU3AherbF5bh5UziyJV
nwHWHsjRXEENo0yCpHcQ5+E+P2ZKBjFAT3mFOj9SQd2geHD0pR7BUzrH0QmMRt0AjY7BGjrSqdQa
ZyUnyNy/Nl8nVl55/65Aufm9TCqLpRH1ioIfGBd7cSyWmvkeVDDf9RxcrhDnRcRUTOOmPYBsLpuU
0cKN+FP6/q3uaCc6wOYTo/C9D1JykYWNo4Lyscwyk1bvZ+s+cXSavVWZmEKEBzb+sSzCOdyoVxyc
L+jPrbc6WmH+ZMjb/wE73RMJEBjDP74D5SWpN3q3S887npIHki2VfCBhRXQlDVWJo6MJ5Mg/Lm7P
BYhrW47nqwJax5zmFPELuiOP+IzIPdT43aWvWV0aCOxkLViXjF074WrcTKMg0QZHx+P93Oro3Qjk
VAFY4J8DxVWDQIsgJYV3dDxfZUZ+HdPV0GHAVAHkJXfO/VF1baAjHpHclL6YaidVy0nnVdSer8b/
Oo5TUt4/7vAlq3PPkv79OgmUEB3Bl1ILgA4rlvFQgaoQE8R4uKr1MdJvKn+RJCM68IhbKSjFPupO
Fr/1AMCg/+yS7c+OnJK5KCXLF360pXTIJ/lASs19+ffdyuJ2ObMmXPLLl2sWTnLkSfa6Ifq11sGO
A1HqvpsNkVsDDgXMC4s5A4Ly5p/NZYQDPOctxewm8naitcMfbK7D/FOo4751AbEv9VEivlJKKsVk
8GSGp8JmkSgJ7+DTt+a4UI2fwgDYpFc5MjTX8ZPSNK+l2wGWVcEX32JY5GYogA139ZCZBYC1Y8TI
npNyPcU0Pc+woRW5rHOmPHWNeSTsG2WiA2HEq2touCScox2bzlr/m8pw7R4NzEoyN0SbF64MkOur
BxQJYnsSIx1k4E+m9QuE0095DmaneW7n+33gtKrprTi2/biQowvEqMv+m1c4TKmRH1bRwwWs5Wxg
w5M4k2CJ7GWoUyKIY7F0u8ijaZDGWONYzbrdDPRjnVdKkG9ip3tlsicJsfHZ+B6vNOjSLcp5csf8
CcIl2wy55be32X+HyrVyYsQLtKrYSHX0jjhP1ZVBf2KnzC4q/3nuSqaFUCAKL6YX5BOik+ChUXEs
QKnhhmwm2GX5ZDcsqsPC1ReUcVRrXiTzbhinUYKWg9RFIa5qb1L4GYTYhpFbPrimCFC4d9Hi2IzQ
RyHJ+8T6TCjJHA5uZ3+ULQk1eQ9T8DGFgaDvWe4kg5CUnGbpcERu+c4r0noTKylU5bQe8sKbW8da
BgERT26sIgwmW0DricivxsTojmhSyASqSacOFOH2U4Jhlfkt/bjtP241+u13dS3tfzz7uKxWEnfM
gWmdC0fUSJdi6Sx2MVUk7UuOyi/EOVXfoFk2qNDj+pHCR2FyNy3qjjH9MipOHP1GpgtY83QID+c7
CUveYXIprW8uPTxNMUFsJFuPor1gNpfA5b9jO4fkw1zpZSxaFCYDHMtuD4MXc/tUnfGf+19aLO3B
6rI+EBbXB+NWg4uLxz89B8A8jl0UB10I1OBSMc9e+HNmw05546jzyHb0IjvAguA6PFtqy6BHiMAB
0Nqj6Pg4KHXKyBqWoQ6o7qGj0ZtG9xGphj3qsT2NQ0RiEPtyz8TUKp0GfxUuKwxQr0Ti4BQD1fvm
kIk3jHupMrGPG+IxZBJ2gSuEHO4cjUXh6IdMt0QKySO+LoNN1BodmdHZDxObcUnJFKpuwsRqKpOV
Jum2clq8wse0VGf5bIx2XU3JqNcii2Mwuht9Wcxc8pjzfpLCZJbTmyzFw63O3xhPfwXp4DjeX3b1
IXiW7fzbBZOA6t9aYW5gYihUXNdoIADnQGb3sp8bSqwdY5eLb5ifvNi+oZwG/xQ+Z0IAHSlxPWti
Y5z6tkWY0GbAO/yOWhRpJUwYatyCQnyfn9DFgsaqNnPs/PNfIKWzAW5aXXtd5xf7eCKzTnQKbsn3
Ts8yz4/FEGTah4udjaZOUwzaNxR68oRdrKA/ZK0b0g8ooABd8rjuqwiVkXaQqlN4nIp+WUxhmR14
koz7STPFNpRguoNYoX5vexfL24dO4Vumy9NVvgWpJ5pH3HvZzzU7JkpmDCMOHsSOoL6aGpAgnBek
xjnNEw3C9Coj73sam0/0NK9lSsYLxJHbnvoXi/X2/e1V3KMCmLv7ahBdPIMEdQ+DnYSEn6GpfSmz
uDweUJbTyNvCPS5OOmcTRCxkFtC2f/tYey1G+E9R585GBFPyRx0zKVH/u3uKYq16wKPEp0Q2zL/t
9HILnmC3mGCIFoNK8tXaOfrNvUcGUKTHYsZuYpFkV5Uxly7s0O0rZt5SgU89vFhC1XfubjXZt3+B
p65x+O4lGXoOnD9ySpN36LmQ5tMEAe0TuwvGXWFgRy44o6gIxdPO2GAYn1tSiGjG0puK0amNpNug
DsD4bA7HCJtuUeaefAMPic7dmaJyFzJn7ZQLoknOpLZquJZWuQrsN+6tOKEqXK/08xSusnOuZXjw
hj/fWJHAfSBIgkzm76sqTMr9FjJYwkF+WdbQcuO8Ww6uD15wqZwfvtvLVudLnEmzSDD9Hxpc95JO
cG3Nsb4cc0TfAvJ2N1kyRUNW7Dov/o69yYBXU9pFasjN0bUwQuq977AMrlqudIqPJY2rYDlZjwPx
IV1h2lQ/yBQbeFjRq1/5vx2Tdb20Tyb/c4AOQjepR0+Ys8dMntgmna/7x/qP3kGUK/dHQQjBVxmI
7s0ee6Fq+0lGTqhjkqLqRYSL4vXyyXr616f5VTPMK1cJBS7QmZXJcG1dg4McwQNhJiyXk8bImj2X
UyBGafuF6G06PE+JpLeUYpHkyCVZHV5H6IT8tEtSBT4NKg1J093LAetJFpL4Xu9WG5S4EbWM0r4v
jC7ijEPecfXcCDllquX2czhMAdavpGKG1hALQkzL9E72w+pGnQ84eSxJQqbvURd2WYKXdJ40KA51
oUUcx2iy9w+0zDN+JQ6hceLC9cAR2cQH5Wt7WZeAcLVRtNl83iNE+nLjhXweUDBaPDUqXMXVI21R
D1+wtk8K1TAbOdQLBsVCPK+mBHAJdKkVIEf2YzfWj158mg5TJnjhPbAODP0eSZxn3ghE2rD39LpG
WwsR0fjiUb30BQQx4ssLjsYryxCvs82mnTrXtoeRyxZZfhv16dZOvmffuWcnKm5QSuf3NXUT6J4O
n/em3Bsx81Sff066O2Zl1ruuZTk4CQKa4Crm80as06pvCxk/dhpO3w28eE/WRDr/ZaaoOmiIUD+g
tEH2sUpzEJsPwfWPx+21svL0yRXTrgGj3LPNIZzzYwJAoYOiSwUJ9pBFW95kbzb//a1o6OPXZEUe
oNg1rpJ4IQox7oihnPrYATSP42f1UohlF4B/qb67Vuz59V0trHGdcRfGg5DJrQ3Kx6/kznt7+YCO
Hdn5Wjd76dsArXVQvyYe81ZyIsyiCTkoIkSpLaPaWotpt1qkiGmT98C9PbcWeLnRpzLOiOhH0BVY
LJcVvVe5aV6dUKJVgZPJ9ZE1GxWyYugZSnLfzDIDMdCRg+UYXCbflK1JWMoJ21lflW/7i5YzhUBa
Ind4NmssuFLh/VmdeNNxAKukrRsyk6vlnOx1Gssf6HobvHEmMWBXSYW4HPa/ciR37astaxBUnT9M
ImrObwr2YuzjF52yYEL5u9D8io8moV1PtjTb7onR6sBhBYOFw3QGpLvs41pE5NV4SKmtXTd+O5pr
cnIYxtyIXhj00JQmEqhUfXpUGt8iZjNi4MRpgtWO5gG5HR7ZK+sei0szgvJgpUUtNZOStM/WkqxL
r5YYeT+amaB/UHuObSHxSKtCkbuoSwq22CxiwBtA7/1KQ3sShZhTCCXbDlbXVY8fWh6oh6mEZ2hq
lk+P48LuQDvzhgYPVt54ZL4v1MUA5PDMDL76dz/O9JpmCfKisHXZChhLmWCM9jLVKEBF2jbXhyWp
VRl/+Ryc0LIxCMTxB1zzQb8VN7C4X+imVYfbkwPSsFf4dtYNpIplAdJmaDsEgdongx9T+2YAWOCr
tEkjJCOMT4fssvEJ191wNsDwrH57ukDupt+2sjqkcUGRdSzbCk8YUgKSLC+DqtXGXZo3Z5F3J5pS
mPX2PNwJRyP9ZUJKjKscmrvXF1cF4pJHBRVjROmaIYMRW0WjO9fDnTKnqdrJyBq8M0YCHfyBQCO6
gKiPVwZVLq7JwUn437/e3mcQvbsRKZ2JUviZkTmCz+40PEdlg0u3b2ID47qe7vYe273TGQy9l8gV
jQlxrFluQrmOaC7zz9lceAQGtGfFtLB3fCa3kK0GOE9ZpCW5A72iQqGYT3j4I4I+415PJbzNydLx
EVR2/gcqetUIO+QQQrSZ/hbQNuathZJqcOXVPyH0oLJlaeoXCvjaQYFDaTx/yb8dsUKel5wK+qRL
2aXdDAj9JzOeB/AI6m2sVTUoLO63nQsUewH8LFRhbK6LcyVh/lM/HRVINiH2U3jSEotRaRPFJGlu
iiNH7z3TJYyoVxO4N4OQP0KToRAyd/2G5UEFgs2QGfzgsaN9CmFlRdbWGDGHZHicJfVVCMPjvK5Z
NkmO+/ZVfG1a0PDFEWm1OJn7sZW0H+U9i88ercQIWF1Fi4xZXh5a3sQFdWy8JL6l0IJfica2cYgJ
JtF8yGmf8nsW1nrFxD5pqDEgpMmJY487uEng2wN7hHpDHV1eRcO+O4f71lKwsvF6J/6M/UVQU/4n
3Qi6sMU4IVRpAFfedFlLJfYGMkAoYiKIXImUfwGyj45uutBvCZTK17SGoCzEPHr1pWURaS7rPrVo
EjW+vVNPnDBrr4LAm92+lOrGuCtvOXSFcaE0YVwqby/MaKooB5fNPElW/a0PsY75gqQbK9fQpJSF
4OFceBjZVSpx46GlpZhk5ouigIumTKw+CN4JrLYfRIMwmmUY0RG1PPW6Y38aIs0lG8lPvUBo8D4d
1u84Oj38GWERypr20OsuUz+9FP3fMpUB2QCHjr2+bxhT5byo29pbDOrAwjxoU3Ved2GQV52R46zp
zUrAyZXcCEG64sMh5sl1ayftdtyi+uFoj5z+/yBIHsbVQNzALBTWTQawse6MvQ1uecEK+ux+7DNJ
9clMEmI41N9pxi3wu+limYBBFBGlnVJRZkAuxNIH1DWh2K0K5EnLp+bYFDxHUQYUOgx4LLyJvnB6
cl1OgurAlcUC1wpKrqoeAR4u+wcqnD51GyuWoN+SK0QykXqHRo4Hxr+0AY+4q5VJeyFd3n0heqf1
cQFFjooB16DcsCi3O9PqpZdAUaE8524dDtfNZpp2wYU80UobHtx+WO3DEvXVlFnHJEjkt6ofUVDA
7hG7GH77PA2NV3C8pBEcBdeWWZA6WYTFo0Tp/W3IL/cT8FjBDYkpHlwVQytJzg3NEhnla0Hb9WbE
pIOdIwPJlmj6U9+o+jpVe6fIvuM8Um+lGyeq8osivl74GNCdO2iGSkNiR3IXQ+aHwmQnH4ATWtm3
kz6lEtZ1pxg3zJYoIWTAm1mDjqhQJEq8UkR5/HUt9Bezaa+IzGdt1jXNFKJLtbYvmyd2cHJFRMph
jJGNFp4lM0fctpXDLvIlBqCrarjctJOuJLQTfnw6DsJhYOk2e3UXmQDc8L8n4EyD5zy5JCldGnfF
kXFSV8wCm8RxafiNZi/60cgyqNIhSSpCFEmChD+YPdeGsM3dcCWF6g95oGe701c762RR4FCfd0V0
R5O/2YU00Mj/GgzqwgbcvpOasgq22mgifiPW+zFijLx3JWh+d7xHxkuyMel+N1mgU0d1QOlBxOl8
VhrF3wbjnbc45ItdSqsOtJNfAeW8L2JC4KcN9o+UOBkoqbDTXFZldM1yMa0mMhIys8S5PlLyQVd0
E+odL08/xtl74zEw3Fe7wmLgYh4XfZWcvvKU4QfcsTA1/KvjX8S0+gmUKA4Lu1fsn/6X+Fv8pt1B
Q8zX5r4Vq1+A3mFPYzIj3nqcy+magNmvMvmE0pVR3sCZwNJCbi7CfrqIwYMIDz16VTGdhJrV1LU6
YPp5fBV+tAWyVPJu179cDOPA2EGJ24jRQY7eKsYobrT58GJbLXGvPJiJTXk4PWwt2itRDxbyzz0I
2gmcfdSVrm1DFV2us91+dCBTI41WQT+2NkBwykgWnM1eJTWownrvetLT3QiFE+YggRZCzUT3KTgg
24yEfte+OK7RlBbDnp3R5oWx74DQol+iOnJuToNRuStgWu7f0AXVEbtolikD87HNXgsjKmCDNJEB
D4v7fqhMeVPpdIJhy1eYmj4xCOOn5O/rirE+DLKTyWnrZXHxHP676wlU0/JaCCq4VClMObriWEeb
cQuhhIB1nI9u7RQrjZ/lgSRIt/T7rUth2F6CV7o1GMVtpOH/P4Qyx1YUgvTYBII94ftyHypI9N3p
wfne5ZEGAwufqkxoMwHEaJPDLvx1b3Bz5z/Bk7J9Gbpg9K3YtoBcV30Nge4VRqZxKtbUc1M8g+Bg
cunmN86HFNSOYqpBLnirUCR75p4xesDlsx4dsD5iGadRt2JLMUtkjCRKYmIZFGU+ha1hdkEpFe+6
aOP6H2rm2QldBfL77k8rOdOZe/IK7cNqh7KGLJZQwNe0Qwlg0JLn/QO3yJMLPPo4SpTaQ4OUbql0
cNDcsi5lNYP8AShhRkM5ksYUs8kjQIYu4/bsj0v2xeJPKVO04XXtSLpRNKhfdtzgK1m45yOSlNlS
lkP1BmZxHZZZeoFpgjBdzyTB6OTbaEajb4Gdkg+x+QckrbH8w9etog6OpPtX+nA+a67/a83A1FFk
ExJbBjm1f/6AO3YIdfNScGQZp1UWd39W72FkmCusgvD15B/8fXKkafvqw/IUSAim1tQDYT+3s+i8
2qVzaTYZpKpEUh9E9VlAwR16n/9nZRlAvtYui7YHnaSpmzlhfIPxFwuG5IV1H1opU6AY6lZM+UfI
xH/0TEF5WRSH04fWmo182Wbi0twF/GiRFUWITmY0z/bgNLBw04wlGynfziT4wkfDu5UXbckU+c7u
DaqCbkW6mHRvHZyCgi4j6jWECaXdgFl/KAnmgFM+WJ2KgesizZEoffpnR6LMYeWvAG28DoDHboR5
Msdz6mnmHHA+gOBHDy9z7kmZrqTvcCJdlo0Auh13Vil4kNlK7d+TW7mp/cJB7MzRQXLQTNlgDsZ9
0Mva6SLxJGvrBIA86oTa2f/htM+6iVtIoiAvXBZ+ZU3GUQymKvYlMkEvTyPMBtPaSgPRjUQyOE72
OTBJRICpDHh0LbCWhY07bbMIfMw8pOsGnILkKhc+OSdQYD8UCLHtAC0nKcqGBQVkubWYBaTxaRQq
idjw4k5ivf8Xp4HRG9id1mK7yo/L35r6bhGX24ffmOkeXUHslbayf7lJPAItunK55kD8i9R1F82V
BYeesfcBSe1ZT5ZBilF1KXBbRHtFbdIWvtSE6cWusqirLAeVzflKyVmA+NnxfgkZFc2BOEHazOb3
lk36HuUALYgAXTJ1Hs/qfSRbKMjWF0fdkg3WNAKu7Ht0mWa98vZyLF3DA3qCjkahCnhjY/eeOZQV
iVz7ZwESh5vYz2/1IYa/MsNE7R8uMbFQJ7UJ8Fb0vh1KZ/nlD7RBr/5qYmCUGjcSA591UrGqA6R+
si6Bb4euGzrFpkTZgoE3pktcEHMlLU/6uFUiMNf3z8WFmYHo8QnCVgPVf239bwnTo6T+iBVmHhGQ
+sadY8R+jrH727wjZ9/dcd16RJnL8re+wMGUhdhcGRMQPd1a8siH7DxOSApOzrZeUnYhIAftzR2p
Sj9qzoIC/eMPJNZ6Cpr8/YOhNzUkVsrNFOaIWYKdXlb43FPvgv5NLOIBqJoHPCJbj5plf7IrBfDq
lASUTtLWMO57pH9rC6fcF+JAHidOmJV3IYyDqNxwRBsJukkhooUwvgY6URYOcJ1sIwBAU2oYCft/
cXYdVnPxRyfweq8rnv+MPuonNGzQOR1b7eYls8MRUchcB40T7Hqk0SZ/ax5rJoMYFM48HUZ3pnIR
XLlumQNosuhjBeT41Q6q9ZuiTvaCHHh1qH9777AM5aHltowqiIWCpro3e/rfWD3q1l25JdMA2Trs
XY4cNy1leitGpYKpM4uodoTO8EWsyM64eJgJbnxojJM+tsmezpQu9m1SuA8G9HiENkqi2aooEkS/
PxirTDbtN1Qas1zUlji0Tqu7iYXiDUsfmXLqWYcOHRPoZ5MJ/gU1z/eFH7mJaOo1GneCwwMoUrLc
KA5138fCKeoP5Y/fGQspYw6ODgohF2oxoMIfjNoW8Uxc0P5dkw8ZuAyQvKg2ytl9RYMi0ahOm44N
VWF4AFfDL3Eplag3YjwQLSSmw2NsbgzA9khow3GjCDQKrV3Vl66MiD2rwUl/i+tq9FHW0C8UA7+w
cV5yUf/6Zbovwh//g8WhWWl7mY2L6SBcKr7gxBb9PwzY1Lg6whLZlA3Lx9Jx0bm4PlW+iz3l81gk
c5RzmanZjHWP6YLPqTrhKsHcLVtrC1Gb0gQYvzRLVZ25Nv0JS+AUoBo4l2OY8s+xXvcU+JqhsDHl
h0RrE9UE2Cl6A3l4em3RgjZ/zJmCczHvZcv0vHT3gT7Ky2gmHis+yhyuTJNZaCMWHqKx8v4bmGGh
wRAvKM65Y8S/aTcI8vx3fVVzIekGFumlKr1xN02zOvpO6PXMFSQvh8DMRG/vFy8uhZgXPTJ7GK6/
hkR6ke0Sj8+9zgaDd7Hy682saj5w9OudijHMESZ5OoDCbXQy9qUvOAIyTKrCAApHSlOjBjoJMFrC
59E6ipv+uJtwb0M5k24SxdyVh4eZnz1H3SWvSEGq0ohWTof7pwn2xoAuiDDty2NygAyDu3TXtAab
LnvuWxPpEzb6/kea5XL+k4+n9sIz7xcX6Gr3mZT8Y0qgHo+S3azKFofq8UvGlg3JV2oinwhgiucw
lD4Jl7VUfOgsaFokKA5TPK4tp9wYn6NZtMsgK1JzPrsd19NSBTdNyKH6iquhYbxXcwtUmnrMkCn/
pjMCr5cVJmAAQ2lp/yhKgl/CUjxDWt76/fLQ6glE76uQ6VYnFuhSNuyPGidxGPp7EKiV4XqCaWFX
oLSln3GgkkB2u2CbGGJIZkr550NuRMqaG2O7NYGJPbtK+sK26oM9zjLw4YFVx9UldlCVAU95UfN3
9aRWuJ5mnXzZMMQfvG6rEZK+ayskdRf8W18r2WT31Zw2ABMXFv0VQRH20RwzRWHZKxmHfbxnFPCX
7mfQewgVc11OiemopYB+EdQOQc3Mn2xtOR4H1/78ja4gfkM7cGpc+FgOV56rZe6ktxA+T42lzHR/
rSNpXjJwcgrAAWAJgtGaIe9mWQBYXZ7hslxJzViAhRWboGxxAXG22TxBKBNL10ztcZ3zkB+ZNev2
UyZz342HZaJz6ipRyNgbRwvX1olhkIXN0w+RZaRlkfYfwldt2TuEuSY911X2fXIiIpDrLd1Y99he
TxFEPZZDzoxJi1xxNeWWb9TmHwC0Piiy/+l2GKT0VctOOyGsiTkPM9/DhIJTwTeVY7VxO1ORc1kq
Lm5C1vZzDvnH/cGy5tA5d2Mxp9EFNx/Gv8hkLTBNGc5vAbTBxHjFNGlkeB4EWaDjYdu6h6Ob6Mwc
uWYkS1Tf03RiMMGWi9BwCziTtuUqcqDsI8PrzBba0K2DUa8CBOtsj4C+0Rh7dEDuJYN0S+pxpejo
6pVFuQG1X0B5GM667/noMvLL3vkZTBPuLLFAit6eNN5yjJNWhsebKqLr/Tu+8rXk1HlGqIW9dIk9
QJLRMivzhrqNUyfzPENwTe+b1FVqpbQdIlpnDrGiSXQIioAeSi0lfsNU3qTGuE+IG1i40ZINMeHi
7iXYrvDnc/UmV2AqvN7O6ItYqId79B8Q+Dykyo9h42tDzm3i4m0sO5DEJF//WlU7FctHdMzhMV5l
dlCCabQX3YfnXCsWd6tWfIIK60YNJ7Gj7wHr+IhWrFDJekmui31fFtl6ZJJ7Cc0dOL0cUPNK0+Ua
RFsbsyLB45cT3+qqlWiADh5hFvha/eNdhSb4zJWn5mQiCltd3m/zoF0dcnx6B2omMugXhL1PFur7
AFo6Vjs1fVvbDJD6sGcpovnGfwWVdgZXiTvNQJWKlz7AV5K492+t76jkxw4TvabdD3zMnlUz0V6o
jXmCxz1JX86fu3S2DicOjk9iDPKVlzrqv+36+/nkFU9OpQfZJT+wwMj3RaYlOLWwvH2rAq4Pr8uS
f0rqJ9Gnvawbgw4OE8z9IxTIYZV+A36jwxxOLvFpdxUkJjQucRhi1npuLmwQPHw73gh3i8/cZWNN
PIiFNoGbdeK9VKye2EqZdqfmKply5qgZpBtdJvpw0Gc5KpFIbk3jnMmzG36y7PEo92lc74z2dfNd
2ZNwEFIdvNnf70YnVoq7qMntfoTBnfgQV39KNW1nr0KbKFtrMHwoo5i4hZOrgJBCwW7x2G3IoRzU
CiaNA6OmMfFbsD4JFl42idyHk7VG/cxmRohNkgeFs6LwfR7zWBgNG77co5RyGVo5KUql4iEtunQl
fwqeHtNfo+mDxihDSnSM74YTfcxSVEn+3bSffivXL9nKWG6j/wFeVpQUkK9w6KF/wmqgCd9vtort
n6nswn26dHw89Nh1gvewWqa0gpFuy4Hi+UMqGp/Ex+lVHL/hso6BkjwU2/q0sjXRBIuPZbIbUI9W
x6AiliXpeZmzBkgDtpjz6KXIJZ4Ms2NvZFGXU/rwfNDlrU1tYVffKuDCj0oIQPZmXlZ2gWkx6Jkt
XfiMe4BHuTQvQPmcyG8NviM46eS1yElkyhVnV6qLR2vuWyE3B8kad6imXACm4Zt4T7Vb9f6HAfvO
z6zyv/2tMaOpSj8sv2vWotuQAdXsaGVIZsXvq4wYdp3uaBNAnoymrvqzUhMGUFpZl/yoHni2sBFN
HtU5tSkzshrmE9abNdX8LGWEf0nBvvcjE2IYkS/m7SU7dQKAk8Rq99AwowxfJwhuNec+uzdH2eW0
JT61LPjDuDXmS1iGM+B8I6utiZb9IBXHg8aGnGLUNR5Sdjja+S38/ybD5K3egaOhzd94kID6PrXH
3IIGrKQan/G031aMzy9TtnICcwVtLgibtpJYQWRk38273oW46c2gGarjDudEbWQVGL5aHUwS6PVZ
K4QlIT56blfD8tBwJCyZCV6niTlzn6VfDrAQ9+kV4XiZ4zpIDBtF8/RPHjOnJCEmQonjDoC+zJ7K
zKDL0Fx4Z01Ns5rCEgACjO+qaFI3Dbs9Jci1gxzi8DUeQ1o2bA+/zN2fORULRz4bC4efeny+TJnr
OLuqzZFOaJlAlSffGpLJe6qR86wQgXDGollqyqcqoe7bLySO8Ylu7EK+bpAtSbynGAu41tLarSrY
SSkHI2mKXXAodHJP2TxuYs3ZKlIBoaXWgghxYpiDne7vUehOAE/AjdUEQMYCNAApVx+bYM6zDWP/
HgXp2IMJAdFCxdBoqAWaA7zMUABZ8bFQV3Glq35iKnFZv6TbfNs2BdMknS8alJwFzQrPqUj1kWo5
zg5+p1j6RVTVzCmXVbO/AbcpefOtv6nq2/oxSqmregP3QifUvAWcSyVw2esc6aZZcTmxeFAE0oLF
bYsjd+8LKab6xHDlSU7uAan8EQCg1xLViTJUpMrn598iIzEriAfkvqpkNa2h2wPFOPgQf98RVfRZ
ktqNz/8K1UnsKJEXyXS3isFAVm0IXvF2F0gRuWULkIO0q0/OYqTcVIJ7UFQLatQKZFmY0LxO5W6U
6/Ti9IsBHtuBIZumRSCTtGQSnS5NGovWFIjJoUrrUQ2dPEQ2RJ+woCRjYP+zqdDg+TrcMZpKpGOY
G4dFVZZ5GfRl4feJ9mhzTeYe1LOw9C43xCqQGdIS+48WfnypkNlq2UX7H8TF9hp/Z/YzuVpWOSBr
zUir1KxVynUA7NCcVcBbXxqHhTCTXDbmWTQCDOGNtqIndW/1wD02R/LImPUTwh9iaAIc2adFEl6k
WKhLoJJfIPEKCDjvAi9iHZqkE87RY3p8QeGUBLjsJSdDEExz5GXQaE/Q/GWwM7Fir5aDAbOQgdqd
KMhzVhNTjkeLAZIU7NmDPHuW3nNahKewJFqMkyzAS1pk6z7Yh3TPRXVJp13KuJ37zz7nmLUkABUN
A51MQqZQTJz1E6exFVrHR5EmOcYtuQ7d3fQj3ELeZyhXA5Wxh/aPMlhWBg/Egyg76XmknMb50QW4
H3n8M1Q/EdhNsBPKNbijXV5sG1TvIPjdSqOUcc4F8UgG9bTemu3XNTV7Bx+OYd+FfcX0D7WSsdsj
IXPejthw+blOgz2RotNGNnktBjCcSXqdwobs1A/7nT4L4GeJaRlGdf0xyeVK+x6wwgkCagtKfEW5
JXtJ/CjsI/+7BU8Jums7KT1STVa07bp4MGb3NuTP9nwfOGd4+OEa1zwYQ69kJB23tsrtHBp4NoqV
JnXRFE1lhVb0NQ4jcK9aOFCmRdxW1v65eyUaAFI56m1XMzgsuLpamFE8cJVlekXayaXiQKyhHP0t
XTi8sXlnujNsTQbioY9YCFjQ6tdIMbEl3zHvVEuJD0miwVqWBnH2FIX7gOpS5UC6XefT46j468kl
9LqDd4ryO9eCUXkCUsduMjHiYmbX6qDS8WMw/Ss7s8X0EQuI+ID1U2X+o+lcJtrW6iNVAPL1RNra
in+YseZ/ppsbeCfnXbF0+EU4nM4j4k9sfhOHzsiO3+5ha90dVABFtx3cmh0fuuyueshfHX81Tktz
+gCZtvYk2MmLxBCfnATnH1pkauk8G/+J8ACzX+r5XPIFbZuOZYyJRayVPOba1DdpqUJq4LxhdeTI
NxchhC0YZqDHsnkSmSX+lxDWa8qKAeU49gbHmqhWQF+784a3et5pE50T2Mn5tw/r07gfx4kvFVjt
ajs+MB3nIC90d/jaXzFbaF8fwpZLScSLh+nGzyUOoFLy9gGG3teYr0P1QSTHPKn4Tx5Ou/wFyOvB
+8i8FTJJEgIueMNKRmjBWTDkGdzHnmO6XfPlKeVet2SgwMSobMK9ZYkff8A0+Zj/zJecm/pVrZRp
+mB3GC3QOVQFAvRqBWLwXr3AhrDbqSIKUmJdHwGS5VyvagNMU60HyXs+nSA3WINtRuwdGVQdGwBr
RD6zpaCHRiC+xq8/j1xSGZ/TFHveehuN2CD1tPgZtjOg9/RTVgwpHblfZKsx78oQ4BMxoDC/iBbh
z/Rpxt7CcnLBEyc4eeiGRYQKx1c8mXPUkK4Lqrq/LZhzOTidXR+w20+Al3V+a9cyrTpUXHo36CRW
eWKdz67pfQecyNzrfJIuOMUVguokJW3wUvJOhmXKtVzF97tieJIhr6RVTimXFEA3MekEEs18q7dN
dsrediJnV/5ms83AIahB3Jvr5/c9SOkuTEedJMHhHfLCkeBPoSQ3ufp/Ngb7bRk0rVFUwXsTDy5i
83R0CY86rMqK9olCxb9ojfj1PBXXX7azoIJaYCRHz1Lp8XhUgkX9+bIQEmGFEhMnKj4DmkYR4NVZ
crj8ujJKBAy7cX1rZDWqDto0XT+kn1KDkFzzaY56vbohm/cvnK0SdSfUSl8kc+74LHMmvYFO0gml
0/n91kcDc0HiSipH8KcB3neP1YOSwCyMdAjV8EFyf72KxCklqJZ4B9ar7HZuza2uL5OVnmRF+fhv
MRidIF7b02HVFkIRNHvjK3u5KBKp0oDc/zqWs/dLW7RXDrdoQpl27dBzb/0zxir7E2LBowI1xuHI
JqwwQyBDGbWwLRKQ1z0NwlH9KC6EHbvglTGN93ujxKSN0JkGk9Qi62BkGQTxUbZ9LRqq92UZab2M
ItEaJQ9R2XHPTKgzvzFI5VTKBVFCT97Ogfa4upfN4rqMPdfx/0aijwgjJ1ppCK7Hwdn8MOwji5Ka
Qfy/fTKUszdQrSsvy/RLJ4aQAQ0KSB8Xolb9sRWa9wWRLLMU102bWKtSklI5qRq3aloTd1fyqxuo
YMghBk+ORrVUgaWsUIMADUgJB2ol5o1hjfiMfcRqVRyFOVG+JP8N8L+bkUeBfbQ3VVPTKnk7TEhE
HeinJXYujeg8NuPnpbPoRFIfN1ZI/HZXFDQIfGnp7p6WcxPPVJKCuo/R8FsfMyqHWJJGmVwiX/XY
TiTkv8pfMvlNT5UGVDWsMFsgg/dsZLGqeTzunEzaiNe5YUJcI1PP6z1SJNahIf7t35rPG70ncleq
uwpjUx+5yo3VPh2VtsM2t0LwLyL7wknk23Ksx9ol4DCHuK0gYXOamjhFtlxk50yRSuG5l7+Rqymu
S1FDgHLV1CKI953YYDS78oQVbH8eQyVkTjOLSD60JJqjwCNy2SEny0yviipPFXNtliCNzvVnDsRi
yjrnGp+bgCcn4HnBxCxRPxX3KX1RGwZYXVyaxwDA1QAwL8ab8etDLg7gECJ8q9QN9d2Y2yKBnHvt
s7hiROC56perv8Z7y7CtcrgKU10/mieqj0lVIGr84ehNVANcryvdag2bTJNIBImK04Lf3Gw/SiDx
q4ZKT+9wn+yIMQuhcHCtRD+ebp9OwppPMx+vRFy0wtsVi+jSg6P/AKDn9H0v6y7F6JR1uj5vel50
0p5CQ3WPU3lYjEfly5AHYCoJW5Xvb2QDDPIUPcRudNOTGjGlAOkMYg57ZMC3J27JvnoPFFKyBAxc
d6gF7A9phXRtgQ/+sqMzqfhucdQ+KmtmRrTZR0hGFkR03CGNaTEPUSTZc80MU5IZUBWz5l8vZYh1
nyt71PJ3PycQgZ0V0ZAFHkpaYwkZc033xuIfQ2VH5ezHb4MdZje23LhsTY7ilJjGyHGUOqkMCA6G
0+SERjBnjub8/K69NWyg/1IIK3wUO/7uRBhUWbhq6+0KIvjggszUmQ/uxkAbCVDnSJoIKL+4oscr
yElTr3ppzsXyyiC00xxZ4ryRyu4z5QWE8Niai/sTixojpWe483qwngPOlK+dfpTzTLRL71euQKON
QGagQQH2H/2GJmMLLeJMwFo0Cq7i7IzQh9D9bjM1eyoEdvzJoFYhPA3dQk3qqcbs7+ixZ+g7LZ2D
9TcVJkw+C+ZD4ZVxZit3DqAxFHJaK1LmBjdYM7At3ni712Cf7yfOPzWVMhjqozj4es6Kc8dcfpNh
Zd4039GPW86ePv9wXwh/MVw+stnJBq8LV/7910fBpLzXM97wxllQK4/JBEQiTYZmsUJIQX+uU8jX
5pLl6F2Sr4zlikxg2IlmcCrGS6SUADfKmotDAWp79Nvg/repR06WmS1swYeAENM15FelX2lqwikb
YESevpD2CYhnMqa2l4xSVujUTFRu9vZ9i7XMIj9cjPNOo7+vAsqaN0Ep466j2GcF7/P6j2ipVLYR
MP2rH0x7jD1uazr82ax2tNReu8CisAqyE93wdiAEZcm3Kk/fB22tlSkEihoeNh92DwLJu7sn4Ogd
Dgdd5Dw2WVhGmTAmECZMX1jb7lJHgV/w1DRrzg/e41rQLorzoGdO9tAYwZ9npCbzQCCy5MfyxPg8
C32z2YEu3iF76fU3BnhXvZxbxvPzbGS8f+4FHggRfmN3XAglSGll1cwzufYnQb992THE2CtamS7N
T71SP4NalQAPP/z8f8QWc6j0LFvc3q5aElKq9JuxLNO67sOLnYGtzFDjIn6X3G0PzW4Vm2fD4/81
qZOhaXyNfvq8t0DwHjQOedV/TXoi6ajzlHZH004okscDnoZotqAjI9c6oKtQuzK58qiJZ1hVXRUL
pFsbQ1lUGu52fsKQfDC80YSvxBD4Qvm7IbvfQ6OSI4ajAkrqCIu0HEsK0z+kXKaFWrWvqPPnwQoC
+6RrxtP0q+w81xtF83eAxGu69PwxB2Fsfx53r6UD7FY9Ht7PI2B928Uem8KMA333cd7auJDZh+Gk
q/45LDyXsQgbOk7TaSbKYHmernP/lSDRaABxwy8L/qAkGDddiWzJzqIEAdbxTEP6TdPhXnichHmX
iiarxzrZ9u2VF6WG9wuO7RfCvFyoSpvqLzyLqbm47TwMZnw71jeKw3Tjc3peeMRmBUXpD3zRJIu5
5yYS7pcQnE14eACYQIjaAGpOBVqJEWpz2jDD4fcg7C+eaWYvVNFF8PliA9WumALKQK3qoajPZP6c
+UuzNNkWg1BMDLs7xtrl6xDWCcbS8j7B4c7MvchF6pzOq2XcvGYVwFWJk6Av0UE1JqGp9JUkpnsI
ZSLIhEBVKh1lHRXIFM1NCziDLZaxz77y/ONiRsiA7RjwN0WYQVXjnW3foV8TuG/4SrUyG/i/xCQP
EU1ZqocKIsUA2RyFKME5VasmylbJNi5uJ62FFNmgyvGlIIwP47vW40DCIbJx/wGWyZ5xoZ3wa8bl
d/QxNbQKDllbvmFEnH4oc6vfq/XDJnheT2Pi+7CtSJDtdAyjWkiFLM7GJZA8CGk3FSjcYukiYK6q
5b6jHU/ft8ZtoIF64JaQ9cDKxk6d/L+72i85VtmdP+dYJTndI6hV+sU5PvAsh/3+ExpOwLLy9pY7
b/KTZyGEzNwiEuxsadsaem6naJ1IpZ2lm4snDZFmuTlgG6OQelHv2ypxvNczXSVNySVpdchb/Hjo
5xEKvAG7M0TdZQzNyvORos4wpVnBIMVNnuEtYPr7pLgoEoyGftF/G1lqO5YkS+7Z2QGpNnriV99y
8Gyq3eei9ek3og7lH5KzuF7EgjVLZXj546xwW1Qy2aIKm5iOs2Uq+gypOK9EwCjyquX7nw5yKco1
I0ofohTRxGltD9Bobm9SJ4M69E3HO0p/Edueu1inCfJcWA75FUrxCSYt6tH7VMjdikeS4Z/FRowH
11722BerxaNR0wZdepLbFEyY6JHBceQ4oIlQSKmnaHlEWUMGigTfucYIFRMIcuACaMMR3PiHbGnM
e+VP/dBId203hJzT35gX1EReqZCEQQrSgAo8lUlZlF/h4yhhyS2OlIma9uUYiElINrRQCPi2zzhP
XlC4a/2Jx0I3bCE/i/w6eleZe4awiiX6OeTSUzSw1PW3+DtBimJbKr6LD9QFZZACnmnn/wyQPmkR
9OdkP2oe6cRwAxDHtUIoUC/uso9KM5ex2yPi3FbFwdt0lspIWnJM0DrYEww+8apDHWJIZu04Nnmr
ZdWPItwCb2KhY5qFZgCN+5hJodyBYS9cVR7VwBoi9lRV+Yq7poIZ3dkBkPgI7rzrKCNDr3c4R49p
QjhdtIKzWGxw3nsBZTWW+y68Wdmdv0z5PxrmrSAA+AbZLbETuBBTzjHAFPR4Bl0FyHG/ObEF7z3O
RcGPjhMyokrTCp95YQL8ZEBk829JCtZlPozZqKQ3UAHTcy85FtHCr9XIkwF3tQ6ExChjId5PclO+
XXZsJkGQC8ZZwdRAmEdbeMet1Py78Wr2dPp6opE5AxYxiI/1cPDfyRZQtj3iONkwMOl8smGqQbGq
xkum7hHNi1azAgiwgqYhuSGe3ZxH0ZBA3GPicQ1+es2ZwqerCpoZWPI2qW/3zCgKLFzFICXxPBTA
eLrHQe5dzAYA9ftxY35XBb8h8ofWJDvQbdRuRhBMaXTlZ2TH88iPpctkwG+Jb6HYcYB369ta2vzw
PZyKa5WPUXTo5fyZF/YcwgSYhpkNQ++vMJUE3KYuxwOfIJF75siilcdsh7uJj3IFRa+TCtQgJxQL
GEUSEI//r6ql3644TeGThkcJ2S5NTEOOmbSvqq99Ub6sq03fNSxqohXzJIpa6i9lkt5tE+j3D1lX
wiy+A401Xxb4Ltg/0Ecakh9Ze69NIUZfu7iVi6GtPPiO6VSwQlUV/B8pUz1e+oKhQvQWu50FzhGG
PcTamU+RdYglft+9NukpRXFOu15xFVug3wRxbLcX8r0Gne2Z2NDUcxnCEdhjPjgm0lfS7l1nPLvH
pr+5hfd3/y4cvottS/M0bTLVAoiVpLbIrIGUj/U890oIIRroq8ZMArg8FLL1Mbz+wCIjNqwsyNVk
i4Ah96ok4pnzCkG+OcJwucrR2LRlBmkPUKeBOCry8lJj6L4dAwPk6ZR/buO/kdSOf1Bk9VgUgMnd
ZJybjgdPwiw/q/l4nStqxH1L05ZA5R2QfzXMT9D0hOOF4jP/BTEUqFQXorkQgdFsY5AOQw84iJHo
E0CbaAaaxcBzkjppHMhyW17NwldPaN+HL8IG/E1xesdvmRo8FPSHJxgOTmwHzs7oBne50pXQVLOL
dJM3rI8FnNu44VQAdLGA1+1b9dY7CYG8d0xFCfkGJEIn9poc1sa6gNB6IT3lpz299uCA7dIuYifD
UVrYaB5pt2aocDNoShmSwnI58Zy++kJ970bs/0YbnI17MefePv8n4PtOKuizUp2ZS3YX8XPPRgoK
tYvxlKltSLuQXngqjy03eQ6YPJSfctOEvC+47/moXfQ/81AK9DrM2wm4Ja1Bqb817wC4tM0U7pih
5U8KsORUIfhrVoIt3AMAZ8KJr8SyUgqvNbwJbICQhrXPf34b07uYf24PT1k9WiXFnHjVLGpiXHQ4
DJvfZGTaObS4/BEi8dmhbxyoa1iiJO3EtwTM7qsABI9RqpmWLn/1c1UFhoyOAW4ylHF7G+v0Cs6U
7wbWVkw0eTmZGp+u03vjYt2IAAc5MQSP9leoxyNYSiy5Z9dpI72GejfKzhGXpPZbHKE9NCP9Lpdv
vQGF6M0Ef8unWtsmyLnJall0RePX7QSlzg/ntpwom92iJSBRgIF1V1IXwIDYXrh895o8Cambwx/T
4+MFZfd/p2RXgNcEIAjPniyd/1SBA+ebtyGYEtDw6EuXQ4usbrn+hR+p4+xzJnu4Xi8As2LLuK9S
9c04UumWcyhLW9CrNloY19hAIln3471GFXZ+Xwk3ObzV0TOPqgs04WRXVr4sHSuouGcr79xKpInQ
zzjQ7PPZL+Sv8V2CW9uFE2USCsIK+bsuNgvd7Zn7fbcDdGfBob2gDaZDLv9mFCl8zkyiNftJoOT/
XXTJcGqrQWMUtgkpyzqq0/X4ji5yhNTOnisexh94nQ1jYD4Ufk8RD0IUxm8/+oAuxU0aUk6OvtEz
55f/lM3+aT5o3+zxplO6OmTQlTphcIMpvwwqkqwZEXB3fmDE0R9uoVv/E7g8mpbQAKCSYuLxoAxF
Y/yda+Tz5UFNN9v2Vt2RU4dkuAXRqo8MuDad2IjXBaquoSSqPsX60YL2+pxMQEisRFhWttdaCcdt
UIz2Qroat3vY3NBWpXhvydc/k/edudnhaMZIFUAsJQO87RCkMCw07F1EWD2GRxhNnXQaejhsBBOD
L0qA+ON8eL7Ddz7lAsfDW8o+y8eyOLpRw/n5F6IJkwCDgCC4ZbTNsyp1n1XJU3Vs7DUDTLlaZk3R
ph8feb0DkieKvg5DEbB17Pm7LjXDyJ5AFNzrWdPrh6efUYW010WbziXNgE7kHlzA/w/3594euEPe
wsWkCCQD+GIpZw1Q2XA4DEhfb+5zG8kq7Zr/jVHZ/7+dH5tmact8LuoDhQP28s0Ra7XUVAIUtTva
rRLWhM9Xh94x3JT96D/nL/Yx6CXRNVPzXF1y4xtzl8Hx+RbjrIXp/MKek+qY1A7DACZPshyDmucn
Z1EEuBsf6I1S9XSWdOMurgYPb/BHn0SB1nfX3as+qaYc56LDBp0kke14oXfMbLfHsgMOABj8R1g4
aZ1Xsj2hMMu3D6uq3seHdA6PT7U0uP9LrEm+hiV5oOk/iHHmD2xo/MkTFb+pI6tmTMUn5q/BepzE
Ekn4ggI3Y+d33vpthnsIqbQrK6zC5ceyccj3bjdr1MUGXuN5RGEaRzY5lfNAf2tjLcd9UprBa0bh
OTiWnt4/rYoPgoTp5hd9cn46fvfs0bD+VwrTRWDEPuEjx9xwJ1UwyzNF9iA15C/7pLeW2d92JdsA
ELI56OosKRbwAx6BJ25U/qnCcGmbzUA0Op6pzoLkf8xsI0gdBddYW92qFT/pfuh4dHm3Zf/E3bPo
HQ8WKJEZqRO0kQ/Wf6dTCfr2Pay57W7nyXUUelfYfuz4R3qjS4Ahq6MBkDGraTxZlMSWXURq3M4F
ZaBxYCieh30eq9EeYPcmYOMiVlmu5n1CWtWP9x08/mxsQ0aW6c0uJEiT4DFw5wqmGUVuZ3comzK+
xFNTPYSSKu4q5yftXBKbflY/IlAHdYd7DUXwlygR+vA1fbweO6pizU7XCde4kOW2fCoFMYvvPAhC
Mx2UFtIA0TFeTBZyBU2iRXENRDZ2oBncWYMLv1a7+u2G/Ixync0UBC/oDIqcT4LRjy4hr4lte5K3
h+sNrXj7zUHroqgHlzbDsdZGL42CKgrI74Eod3xg4KQMe8OzdnoRkLmOstrPRldnoudOmjE9vDU8
Udjv/J0LX8f7tHur8acx9l7Snhx5bJMZSDmBN/7E+rJ7UsVOms9NTgdPvTqORHzmoCuF3h7SxOEy
O+poN6Yw6sRwNFCZ3LkuQ/XHBtQTySYcd6ew17JtfAKR6eFKZ8/798MALxuLxIDgdYFCd1tn44K/
9bP89AJbG//KJPt4E+uoEuHg6o6fe+INeslQ2Gud4QIA5BB+7DBdAAGJVoY+grEW2b6k0YDy1RM8
7KgEUf08PdQW/PTShrpiwLnscwufjibMZzTGc5ckMXHt10HmUP5/KNiQpgehJ+YMrcAumvWhLQSf
C2qf9PgkA+5WwILZxop34MnFoREdUcalilgVC2qaAXcE9FJ5JV6MaRkL9Fz7q96FHD3QT/AAr1hZ
8WakIB8w9cv4v7ryXltUAbfp2aIgQLveCDRNeMzpWtFAunL/HwOjSuBAo3m+ClAfDjEF2Vycxyky
81ZbOXEcXdNHm0PvUne2wY4U9huluOzoyNwo0XbJGd0IRgbnh5YeqhE22zAcEE7bXfW3klrR4PlB
qYfsGtHFdqO5ACDcIGoeYJgVcmrq95nIjW/O8crSFxnR6zqLVtyYtetoyyFbmNSGVhevmjA1qZ0+
pMf60xn6yHXZIlxEIF1LheVSCLD5upbza2qGz9zfmrtCTzqkQI3zAAFea760HHAASJfn21uXKVsh
oB3/jwoqxjlU+8bsmwZGO//cC6RdVq16TIzXel0hwb9qiozyrMh+yJX3uyeag1ybg8ezp+GHbRFE
o2myb16M9Ji/9fWuY+Y0G5eQQQ5ZFwFxPAgoPGH7gDalizPlhqEKn1G0/LbnpMNuuPbc2G3wY8r/
5JoOPwf8fvFtv8QdzYx6lqG1JuMQe2KOm86Yz0B0w5JHUbnkGD4ye50AAK2l3iac3SPfAow+02WH
mHtoGhgXUE+37iRlcYzt/ejFnpxmeh4PjSQB6PTAqI8wKwJEjqX6UxFPEL6Cn9BciDrdo2jS5yhT
wnVY/ss9C2LJFkKB3ld8GAtE24Ea5aWbZY8FJFcQgT1/fMAUjMeUUzo4x5MIBJL7qvfk/jvVARGi
Ev43lUrvbuCZWH/mxkNr5Haz4NvqYR9Oh/MV64qH/scSJSrLreIpbZ9pXNVtFCT293hjgT6eSwqA
ONIMIh8HvjOb/vE6nXltN1f9gwAQWF6rZkkDPOzsoNIgVFQSSb3DJ60IguOnclvlANplzB+P8IVe
HNunEBhdHR35acejc35Wbn2NnEuBGB8Vg+p54O6MlxnCfTtJwTeqLP+Un6WVOum1qY9maVCohY7D
NFFSKZjkossOhwl7YhpVmxiw35lahrSzHGqjOjDSU1YDNCYSwCccJ1ztF6fJzi0raoDjSlL2r/9A
VZuccwG2WkOvm7GpkpGhbQmW66bdNCF5vkLapM61A0zjhsA75fdq3criGycnFnBfsny7Y5A5VnBB
OAGMGkfox9R8DHResWXjRfC09rvsOQIFtGAuocJzbobLPvFW3lnAkFXLSlcHkivq+j31w/HhUwoP
RzxFx+FC49LQPU9uXHlB53tAAoc6Y9UzLeK2sPm11d5ScCxDi0SLc5hD3fmoLpXwBzKIXfJ2J+y6
iutIvDLJABOU/+1G1th+rTJflIR9+ufiXwQkZWrNulxiQSDZyqRJC79uhB47gYImdFGE4aq1rJDf
tEH20pfr29B+5aHBsOK9y4CvJhk7kQkIHtgZBTUhk5s2gX5W5Fh2zABj3R39ZXaiwWh8sayUhOsQ
7z6fP8fr1rZw8n6UdNmpFSdM7trAgLpoghgdDP8cy6bcVxKkZL2RR9l8KnthLbKOrCVMX1fPtLe8
N6ujxvQ1GLhhiQEwCqKUpuWG4o0lSzRr4g7NJIw/jo1H7ijj+IBp647eYiaBC4O5s1orXTwEHyS/
Kb0Ab/iTpuTeLx+z8/5VRZbVCBxGwTydHyVV+erSFBJ13a64Jhfc8Gp8wzoKfyCrCM5OGk+TWcmB
pM1K7VH8gnaqsYme/dud3fBKwzOWyCYHqtCnBP2Uxn59F0exyTLWhxXAWAOtIYMk/9D1XoTPdY5B
SgSCjg5uvC6P50PxWVq/bPw8/y1UunzyuP1eDZVYmPHlZWN1Ru8FzWJUyvRZ+rx3XfdiozCk0Ej3
U87kPBZoSBz4UCs7bvnPN3LqFbR4W5xjH2vLNk5zLt1Ge5Rtvd7KzCi/We5cM5WxAO0zcLC83hQ5
WpDUAW6qkRSXf/BTuBUyvW7V/anT+FGPrLUHxyzbdqzw2v0yTwpKvZ+tUJi63FRnfdOY1869/RCE
EsjLJrB9f4LjLWCRnxPcVUiQkPsdJcNN1GZ+reJlVm6iDySKeusvJ3O/YMBhhZK/vVolPQOMl+n6
9h0HGLL9MJzVgfmyuYKY7zObvz5rTc66Uka1iC6hTnRGoyPp+1knC6TttRcvnUiKSkclnGKWsdYX
sAONIs2wR7n9N6+/1LauWLEOBj49OZDzLhqlxbXU6BNdyzlhNu4R48CiMToIx7ZHWjr0zO7474P8
0N9fw3gP/MmIfTEPbE18J22dEpwrTJA4+mjop3aC3qRTRGnAEO0XJeA3Wc4TiC9OqJpuRh+teBBv
R3uDMMkH7CAUu4skLAU7uni4xIBZeVMyJcP5glk1B5VrYPBK+uvjU7Z2KFFIHkoe+D7yPxh27Jps
5QQE5Vk/dOJx6+a+CBnCQs68qEDyatFnGI4iG9ODoaRB4QnvM/OmKSVlklOqtQOol9PK4pppaEfg
bYh/pGDPYyhdZR5VSvKeaIUB2hRsOPs9QMQ46SKvo9OKqc5dln1LMiGee5s6+tKDHatpzKeDYEsL
7jZILUxX0xn/2V2lBX9yKsKrGgfUJR6cVLBrtfRZgf60qCvBOEc2SPYBc72JmkHyayZFiiCAq2wH
V80fXBLAq7E1ooRl6KvjwG6YD3VWM0sDbqM/XXFz6PFtXfwaOgAR5r6yn/WpLzZPLylZX/0VWlFW
mRECBMxKfdGzvrabcFPttEnBYNN4wSi4oHSucFXv12O/XaOiNmanvYbzbQTc1dAVnzGJjsIVngBp
DJWnUJIcdKgEXKg7Xb4yL2r2ifs2p83K2VMpgdmn2INBJNPhUh6sRMlhI5kMo4YWLScugkrjSPMx
MCdWDeiexz13Dq1okEuXITRx5dpO15kM93AlYQ3R40+lCQ14YFea+mJa1xKCtyu+GBI75P7N7x0C
LbM/ttshZ3eb/7IoZQvxPIUgRI1UQx/IpOKE+3FNpHg33hyuEQWSR+TG3oumIEWqYbFPpXgoPzGd
HA2f/RC6LdizlY8rv0sAXsYTcVJI8nuPjOjcdDi3OfJlfcvPOnBggUklP1kVV3etr+tFRYnlQkI5
7EOtgo73J0jdMorDZfzXVhG8h4/T3VsYwGGCnWlLnuNPpUCwPPMSuAdhU2ycly6RJt0MBio3lsE6
ywzKWkBd65vEuj3mz3Gv1IKNYva24i61RsoaFoXY7PJ+5kizJOZnuvEKf1RiARxcDh1GPyXZv1DH
x2k5Ozg9oYXbMfg4dex5iXj0ku+3s6F5Z75iP3aifidwCYuf+mlqnBXayNKah3Gs4KZ8lN0tjSYG
UxU5ZCP5eZ3XPld3fCvVlu+EXFafrArQxhu7Z1L2zufP0C43DbjponxG/r1R5JfXabANmtjPz7Eq
HqIDXap3HdOitOL6TR3sTBQolSOj4WuU4pesE2Sup7FfHJnXlkIJWpi4jIxfFtWjJDXORG1DngDg
3gffiKcRXfd40WXUXPjQsrfuGLnKW+APqxt90lfDBvsD5yZSEfNfS0lx8uHRoYbhest/JRBtfF4X
wyKqALMM9CBa7yNiImOeFNtkKlm5GMf5zPWy5gGvC0AD4G7dkIIcPqd1db9NYd5lnud6kAVAWPXb
5jOg949N0O4dibXcJoTxa7KASVuPRWBp+90SjzF54z5ywOwfDBbut731xcf/PuVP8aA3NXqsictq
ot6jCPbEOdfim4kO3NGB9X2n8SNIneFca+tW1dH0/4KiAA85tvgha4/nI1ybdOmSY1qemlYucMKy
DRPGjAmX+384VoQlbVMeaI3IpWF39yXZ7qeC0N/3GD06OrHKwNQKcLZRzNaxrPPDQxsWpmCJ9Ank
G498feMgIxH2kTKvi0CoiKh36XTc6L1GQTKEcKit5n0ej0xrjzdqmSie3/n5zgP3ZCzhcQY9eBKW
3aexnuoZ7W2HcRUKZwEcFBVLwyZ91wLB+G6DAQmcq3QYJcogDrokmZKElV2KDqQDJcMuATe9QEjv
DqUsKHYzhXhCswCiBYkjwhGPUq8X0eoK7RRUYy50gm7mS1dq67J0Pg6WXXkXwTw6KIz+/aHKXDL4
HfHz8NcOkkLp/FK/7JGXGvpRYs8WP0Go5WTKenn9WQPozthfp4+Ew+vYgTdQ54FyaUfpwUkGFhiE
85Aubqw/Aq1sv9Lw142r+qPEUhvt2sDwCEH/LH9dJ9eYgKZGbhmf8R4ZcXoYvZjKXfI5hX5Pdg5P
kvzMWPCSb4Ttyzadpygc89jr8zutUeUN+Ww4m0NJXGmXXwJIrCFGBFvgqD0Ir/VGz1vKkxgNz+ZA
q6vUAFVOgCbM1sylH9Dk6uwkzBYo9PLpmQ6+8zbo1+rKF8C08+uY2MOB/TwavPQq51FOba5wzos3
BKpDmjKJ5vtLPecP/eGGaz6S5ubMusaDmFsNsXjRzAXMwhLyvx8NOdjQp7+Hzsd7w15k6N78sNf4
HIuBxANkER6gl+tZfTWrIcnwBnYqlT9WQGRS/jHxxef1A5910pmh8wW28grXicMNW5fzYOf6eqlC
kDLhjpXV0MP0Vc8/hOi7WIQT3NIDghvGMI6Q6Mr6t+GOiBLoJFk0m/AgfM57O2UIQXkHOR2SG8sl
HO8d8N3ZCtne11rCg1/qiLTndhtRK+g4aGeBbkpS9L6h3J6aUwHou3I8Jm5qMpjtdpUdcQwNCAqi
QfWN4UWI+36P58+VxFaHFgyC/zTs2CuiJVNNxb+g5+lTW+yEpNcG141K7MWcqQvyTkQ9Ze5ArWUq
oq/yDvbVGCt5Ni8TbYBrgJOeddbopQV5L5CifXMtKE0rdkE5BMZPxGHHOKdbagjemA0JKVfDJq1i
h+8j4JK9R1F3Y1nm0SWIBqibZWuhFLVDbwO1zPYs0/i+M7ECrNb0dGFw8ag+8vTgIcvxRZ8nLvyP
cXh+i+SXt6dkv+MrSmH1En0l5Ir+eRy7pZHO4uhmF8MqYHtBVRGyKH3ufu3kzK6BWXE8QXIjY/HI
UxMcXJM6Q+Q+Y/B8OeVft6BgwijqCHKgp2s3ulITu7Afj+hVbFb6DcC60hpHhetxuJfursn3HlgD
sf/DAqOyJwySVPN3MWROcZ1jE/fo7Ibw9Qzvjzqrq2hFQgS5ycG3cowKxS59QMoKOy+b5Yii+0Mm
J9xttkO3n96t4DRpwjhHTRODOvRephkO0ZOW/xQjOTO6ExTORy69Lltmsrq1o8CeTS9PY8mmescu
YfBqbVB0+qH/IIETWlYofR7HaRrP8OJLpf67LkqtW/xE0bWQ8de2utZWQhbkrSzzwLYYCVhB4n/R
jpWnWnBL086AgZFZyvVrvsztLB2azX2r0loFBx2us7L2U2MGwMhHeOsOli0RoTZYMJzO+Hquz3jy
rgc0F+tlx034nZpJo16WbsQjODkN6Y9RXyt+f0oXNMgJE+zJLsxkvC2sKJ2zzQCghVFbQvs+8WgF
w82dsfyQOsooglFjwZ1M5BMav03S3aJ/dJzWtcAEBR2MCxl00sipwxUGcGIaB/FQJ3CQ7/jSAho2
9SsIn/ryNdRNnP5SHDIWFZRb8Y5UmXQOJUof24kXpBDlBDZGXDLC0zIEq/8BoWYZ1q62yzwPEe/r
VZVZbnI6mg3hDpmRWDhzo3Xy3lUzeOaGc3SQwE77HvvpMNfmw6qBvHt87GWJBycQH9eCc53QOS9c
LMey6XkpB6orYEiOjGf0uyosO/bovglTFakV/dDoCylTJwASjnu4ZBC2bWAzLR6YLDpcGHU8inOJ
jkayJLSrslr+oysX8I3YkIj3h7B5mbgWqPPf99oUUKWgYiWB372UMWWqOX+sxjc5rxop9cf+io0D
qEo3qPtjKIShvkzUCNgVS8oiijQEyxEpsJi4QLT88WTc6qFwaO/s2FEQy/6YtDYEDF42LFaqn6Lz
+GLMHyjKx8LWQ9B8n0noaY4Nqmj8mhp6AhI0xL3IZWJfSP4dOox9cCDq1w+UPVuko894uoOCo92I
skJXB3s81aYth196F+sHghf2KWjn5ZsHeCz4UuiS0P36EXArZEfAiCFtRWDDqzqP+W/MZrQwz8zS
Nw1e4ustwLRV8I+u3F7mqfc6NuSzg+nyKApldLx/DtbeiXYVw1cHAQXWChZAhL/4BnHtda8+U6Hw
v4qQJVclGM/uJHYq2O5pai9VkneMFSMUo+FV8jf+BAVU+caFoU68+Drc2ywQeUsE5aepp3lBqrLs
jYm1lHJUiSGTBh3p0A549IgjIoz0c/PBL4ZClo+oyliT6MlozFKzZnWdtKXOTsrkKmj6Wn2RZq4Z
SbyTJaLfZzVCdUTJV1YIUFyRN/hH4OpGLRcpIsF8sPINQpODiEtKqSOaOyVxVYncOgfI9k59nlMM
6FzSLILwIrmO5Dkv8j3NWh+rFBfUAJ4bHlMw4DgJ5XdRGBrdpqas8jFsvmGA+shHW+/0z8fgzM/5
OMHXoQ5qKQx7+YIHdf21Ogy031Jy67YSSy3HslXiNLUyFlPl+XF2sNTOOFxP7kX+Dq8xEvUVx/SH
UUvA42vokQnS1KjLr3liDsxENDOI3fVUtcd1zrWLEf+KUQAatmmHuEmOkqLBCTukd57B784Qgg88
zHO9BudPfldPe9YfvbkM9IofUA4kkzEkj5YEKhkrvh5tLyVzjd3rKiiBpbB5dgeHEuKACv/hXFlL
RimVFsDynfTsA9KtpoJ825miUofaAzlS4StGegBySGW/U9pymniYBXq1rZatRY7lztAfrofdznsR
oFhHRrVGgSS+t2yEI084BRTgiFeQ79OguAxK5HFFS7U1/WHcEaolSR+S37T3h19lpAqSZy66KGIH
sqYM0V06Yrc6Ku8/LkpAjh79xLL5120fTPnKYQVZhVk1ZG6YjS6zaTp+0Yx9c39Xj5iJnIQ3foU0
2rfSVWQCFZnP8KjJA7dnPnLQJWVjgqMRY9wDiJ5auEH/FkBp445eHdmgC1JJ+qjPSKNyBofYA5aO
lKob+PdvyAusMZxS2GoEJo0YmEY9HIcKesTZ0kW8q9Ma9BwXvPXiZInCuYwCYDxR98523gCpgCFb
cFUnm9qV9LIuSG19SL5gumXBW/t6CVfTpRDImzL5ZFcZ/+RjtxsVFKCOB8WY3MwS/PtLsyGIFfyU
zmYm6+4sEgPc5MvxZDNSGm6JQC/T0zuZ+QOU47QNTlTZl9fJOJt6vs5d/yau09NN4Oi4GThG82ya
+fysan0exi56KgK+9TGEuddTVz2yUaW0bDb39yz5xH111kRbcLhtcOzSITCrzgFpBrg6nb+vdj+Y
Ku84oXyEkC/xyAKQBX3bT/x9ewErdUUyKOj7PcQ4AJCzRkdHgtv4u6P7PdmYkrXRsj0lXLRE5jnV
NEXe1CoHFgl4I37bc4tj6ePN7WRaTR2mJJuXpehXyNFlye7TpHStoVH3NVki81qW1kMZGZxYO+0M
ObneRteRfGtDj+WqWEaDOYGaXzvlTQqLkp+PfLh4EmXtifIQrN/4Nnvw3FniRnipXzNqwenC4DVh
6TviWuFBaHZLyD9KgFHYga29YVtv40dS3FSiCy18uFJD8sDIWwDz4GPKow6++nYCdMlu60T0Tz6E
Oug3r0cEJ949jMAfO4++Z0xIDdL1VxCOt/F80w42Ne4Enfc/RenZjurG5PZfJpscv3yBM0I3sar1
gi6R2eNBvEkkj5J6bF5ofoYcGRTI+1MbcTYNjXH/BYteWU6LXqUrhHCD1zF/jtPYohSd8Brmcp5Z
QnZfT8n3aFMLLQm8v6j3dpw00uPCZECqqVAJ+dn0Kmw3QSd4grWqvfXZayr2jfnfBxxaEcRiwI/3
7LG/syDx6yXE9LEk8B3zyml2fbtYzwVBQ2Uak87ikpHuEzY0RFYg+UPY8LkngMfJi7AnTdXpAWt+
5IpUcErClvDzoZ4K3Z3ERO0fsc3yHOpx23C8YdaD3KqJDacLVVwuXjG1OogUh0jxLVXdviApsfMn
4V1FNjNw4g7pPqWGt2UhO0LKC2uf7UO+XnfCarkT/wxS69SjNJybmfRZCa1tXtMKTNqlUAGOjJT7
5DSYtnEhFaRAef9IG+smy9F+jnCPYMnh/kTc7g8UA4e9GxV4Iq8rTO8ZWU59d+svdrJKY/ZMCSwy
HuJOha0Mdf8S6rMpCCJutioDU/X40zK8wMhAn/imYiK6T18wxbaOQo0+4grmUzGb3y5LUNQZeLJd
flBXzwdYg/ith4uHmTXDUw6V3Vd1miJmgg3CA1WTekk9hAYsDE968ZrImfcyrkQ2BpxVW+KsDU/r
LV1jYyQmnm5ocGjjd76xvpf8q3SflaMWAXj3qYweYzCzY5DIXnVsKMqiqPXEp5KTbYCbVB7YoVyg
x/wmMOgASewZefj6J/t1mQQCVBd+2Efhvdg7dsGSbVtV5lIwRrniOAARSyPfBRU0Qu/wANdwKekA
42HV//LQDSmYk8fX8siLLCCK/UHXryc4LSomh5lFqGNqOJt0Qruv0kuktyHoD6g8ogc75x1/zS8e
ZMDHmOBEQ/vNPWk3z4+dn4QxTvf4te4JzKhs9mjjBPIl8W5YSNm1A47qp4F/+P7/VcVeO9c9HKAY
GtffU1sSE9KW9eRY7hJiJz7wtWbRDkHdMtD/L2LHhCyaEz2DJxXqItBLdAW8MaAO/QYdqcbSuHTY
XybZ0xsxIwXM1QsW8v+zH9zkz0ugoBEmJDZ59exlcQXitJa0fnEAojKm8TIiqMFd0yIRdfJ1l8mZ
DChBPrX9RCvPropFpKTpXjvSx1+8bOhji9a4y3r6fLXOr9ztUMkCPWhaECkypTr6NhgtQsPbZ9iA
zNi8FS378w7BURUyXTYdfVOr/eyNrpt/YCNJ6GkpHns2prfgsDupJvRLI2SUx/N/m7LHuU3AIIAf
CLN03xyO2BmN/doB49FChZo1KQLM8FZUVM6b0AIjTmx/D9mVG0Cjxl1ln1yErv0pK+yCQfm8Dy7k
WhuGkfgB62WFU6K08/nS0KPLMuXadUDaLWNszHiJRZdN8tVxiItUTSyTSozFaYHI3N0xD/H7L/Sd
xJD04EzjqQgN1fFvlSDQr7e66YdQIGYwt7UkobXF/zFp6rVe5PZhDn84AYvm2d2jjvds5oOboEXo
YrrZAK5PuYN/M7CySaFlzcjnuc19Ejb4I+9QzRg8/gaMUy9O31e00ALhVJ2HjSFOjhii13l6iiX+
TRZI6CH48xDOAWOXB9A8RM4HcVQNt2VQ5N1uAle3zBU+OjQungIkLa6mZb639ulooelZT0MFxGTK
Mn55P9O9qc8zXlPziUgDr/fvtAuxUcoLxRKEDxgfUxSYoThxS8SFBLCsuMxcMHyjinnsc5Ddu4+f
ztslKJkd0ZVUQY4YNrLWYyRb/FZLihdX5hA5HrlQsaifIOBZFfEhbbFbECj8tfgYNPjIB99HpaJd
kQMiPOf2kvU3pXYnt0Jb0Haj4xDdPg9deMPFOnMk8Gu8E/eDtbsVTIv++uuojHHVzNifKmJWQk4h
/oY/KZRYHKzd5MzPXOVsiVgkpgp4+puP1EfPaPHW1cPxE9ilflBQbDmSqdAgdVONKVajhmY/Md5Y
SazgsKth0PVgcGuhLSBQr1WF1EEj4l0ULSyEwjwsfx+94vBjcWsMmiTyEYE9eVDWnCTzFpzqPTb+
Gp0+miGhd5Gnoz2qz36FIT1A6oUUrHNoR4D2BIaP93+SE0suDY6neAqzZGxXYxtrOr9f5+G88vam
48m07ig6iczd3p2M3Gu2zq+8XUQ2ecQhLDRK29+dhu/1e4tVqy34D39mjZfpwA3+ZG3qauUOQGQP
7CufoeYjGh6ybDaHkJRXE5YoblkZgsLAXYsk0doBaFnYcX6bdn9RJN4C7SP/VhlroZh8XwT00lg4
KIU8Z9mJRNAhq77SrpgMhsNDGKaXX+N1WhBzf3zZirwJJB0So1Ap2fUJzbAjRMFsXcdf3SMFRD3Z
7tttKLfTm7Mfoku2x+m4SPi4XAtkZOkXHlyGSloNgrGK5l1G9QZx1P/gmnu5aUVhYkfFYePR9U2+
LejncpvLccU66sgJaHVzvA1w1ZcMOudLFdGhILGbEJF8JejtnhRD9B3r/RR5S7xLUdM9iVcXAVCi
0XO8nOFh5kBffpXk6luuRtxi6Nl9yjyVjaXnN/iN+oEavZqTR56FWPraSbu5crGOuQA4yxs2q2QH
CVCqzbg01eRjRqFF+EqJuIW8SaFAKmLCGovn7POTEVLwXCwt08CfO01yih8IweNlIg8gjCk/4hGb
0MQP10muTDOEr+xMccJ5fO7Bi/HERNGtjFG8tb3D/uJnxIj49bcMoPVuxnU92TD2+CjHfLiM3ROb
Hoz/J81E1XWPMApEsDf8fkn/KZP+dNPQcsf1zs/bt0GgJ7ArRMI6L7x94GOrwv5gx1zLHrqXAxJ0
K0/cpfc+Ag+qVVZjgj04uMPoGsfkfA3P7TYlX1cFRrONJokDWYmVOIDQhaz9eIUEe1jbP57VxS1R
je4nghLocVS8AoRtMdY/Odmd1FrP3sThSOJDGFSxJlMbhbSYqW+EaZ+jTdh4L36glWmrmLIB3CST
7oNBDfIxo++447cliJ0QxkupKHTpwjMiIkpxSPiDMy32FJ3ft8j2pDrboJ9wouvWmdYC6o6KQIV2
Wn8hMpxxvSm169zn9H9pVsa691cwIVQ2WQkkIRG60IftUclsyAlqu18a7Na2qMsWc1ClTsY6ah2x
1LVKWpiakAbFNh1KSx7RwXeZdEqS7cENJsZm5wG0D9rEYVFoPqWLiDssPGE/5/FnY1bKPgjAP+vF
1ir58henGzBYENWgzOXIHAr/5gPkKKxlXbtcm4X8yVb6FxfBpme8OmDIrbq3NuNaz0G+Ye2k0dAS
3uX6YPN2r/sCEJJLufK4xGtmn6AM3FRX/C0m+bJWC6vLD0zJd/0xzsHiwl+Gc7fAh6toM7FJc5Zs
UIltwNG/ZsvMoMZORNRLfHbmSADEmhh8Ggqy6pGj1RJHMH13zqhuXcldzZmmpdkC/K+GeW/HE4pr
uF3F9DkOz4FMgkWD5HQO0kYhki14MTCKDtjC2/mogWRDcOBJVz/xpLeuEj7PFIbuG8Ik6xhsxpkt
kPxVuKhHnXBYrEBOZ4Ho/NZn4GNRkmupVY9StULBqXRSN5WLsxBb5GMXv/KnmDbsso9bv43HYKrO
C1pMk7vE6ltWKdcHehV5FQ1XwgL3VN9rUdehWhrlXBVvP3JwJMG87NQKWNphsTA2qiK+O/kZhkYJ
EDqf7R0Qdo/TJ07+vtXNszV1jCcp+h7t3LbRXWAyxSTazgnotk49xtvxMsiR2dvzGsnbvJBl0ye3
zUClLykL/c46FOWFr3Ad/tIprJMgPmCK37h9oWvgyja6c+gROFqLfu+lsQug5yF0MpbuAEA/TZoM
Iz/LbHk/BPbFcukVmVmf3dXYKjNP3CBDHIb749WYlPJN46H9jEYT+rUTTYJB0UgF8FmBc1/mpHFl
Ls72NFXxu3jGwOiqDbjjXusxpwBHJ1kTWxkplRHCYATspt359RWTm5najoD0hySrTojmYB1o3LVU
4XKy/8/Gp5cjwlRb73vPpQiRF5UQFA/vb9BRQ38aY2fn16aZWY5y6x2QMN5TQF2Ls4JNmCvo3GY7
bri+nI+wEVdSgyAl9+bIJR5/2EypgXPxMWXKE2M3cUFRYLEa/fNrOYHMf8tCIlypPovB3PHc3PSo
njth2CBgpdGSO7rMHa/e9j3Sr3EwNHytB3/LjMpviW+kVDmtmnxgNMT9DRwIjvRi3pjrC8Lc+86n
THJB1ulG1MnBWFC0+DB5tWlHEttCKUf5GJsb7BPzACs+6NFcBpiq1pm8Dsqb9LlD2AZpxe78oDey
hGevaI5k0kDjNzXj8yKpWF341VZacFeZOuOltkFbQOvY3j8rSEMXlKwzrL1EJSAEVI8alpQlUvo4
dSJgPl0LAKPaoQjQwbESlUIEwk9YFminOLN0hNU7QYp4EL2ocEKEEGfn6sSvCojgpRuq9VQdNxLa
JyZS19KjJZbHRFbAtsILYNz3zyf3Xxf8H4Nt8T4/hRAp40//zezGiT0a93oTJk/zcuNiZU8v8hem
rsnFJ1ya1Fpm1ZT7c5KqJA3j3zdzazOi1ZEJT16UldVTGPWFS8N6yBJnc0DqtRvcr0ljisTY6o3m
LRXSOAzepKNqjGwlhBTH+PHh4SF3b+WANLFaVzpEhAEmjUap4qi8BfLZ6e/9MfrrU+TlbSl1Cb+o
P5+n66Dq/FDbsWK2zrUtzjsOuKG1w0Zu2o7eS8gbqrl6SRBbOFVW247Zqp0LLB7Wf/kMnpI3uR8q
o61BzDcP06aCNeE4WMlpFwIyBoPo+0TgjZW59DIQ4yo/7bWg7zZY8DlRwmOAkp1c/uefU9Bl8Ann
buPT4m2JGGY8OhvVxweJjdbzpgHNrXsQh7ic5zmZpxFL0FjxQpaaPwHTsNHIGfUJjOHcnjrkJ3C9
MViB//29QmlS0C/itRKVaRsH9T5e36g9V+1bbmoTAsr92deh7qyjoAmstP7h5RF20fUsgZx8/ByZ
uZ6xa1f4onuNnbMWYq8iARQQc7CdF6a7AxhLXU03Kg500RZOJzPF9PxpXVO5E+3IYnuk041paJ7V
QD504mhiQJO1JzBc/N563RQA+dYAKt8mRLYLTvxvf/DLIrwm3E+oaHPADpZZcv8zy20vlGPrW6CV
UFPNWue6UdQSsogRQBSr8BbfgcwViPz1u51e0vbj6WQEXj1KhVjq7jD1l2whlm04OyYXMXSqCPxb
+CNQNbeQ5CkaWHSlTIrBVJuQIBfEVck3Eh67ldT0orIjqvD3u2EL4lj2+GW2vZBwgKhb1yJv/uef
zjOGJ+Xgtjx7kLGOQbO1QD5HWM1PK2CpOiszr48j2G6BSyeC1lIcEXSjS/sLFyJcxes7d++kw9Qn
eInpSyBMxfBJ6X5PNVUfAfoRnQDSQbGWsEIG0KpdP17W/pB+wJ86ithQdPsYIwJyVQszftvuvjBl
cLgSHjmW5THDn+dakRqZwCf/8gtqyNUmNrU6ZUq8klskiMoFai2rZLs6rdQd7CkvgvOq3NgVSKdQ
EZFZ06Rz6GwEfH6EQbbW/533TsSgO+mkqGzPKwgVVTBnfHNn7CE7KaWR47HzwWM7V7Mi875qqgic
mQAZc1mjoY+VITa08G/4ZZ/cE/J4zRWJXNOlRvkMLpCjjCZ2AhTTAoBV3uzhUZNyvp7U9WeqByKZ
g5807S0jsctZhDsW8x3a1HmyDz6U/CO7D1I8CGIsz8meNuh2/f9rR6xgF/3Dj1tJEWQBATnovNWy
h88yOJqfR+brFQcXT5TjwS+sXQPkiS9Qh/WkeEcKD7oAXCkd92cNt8AETQvsXXaerCruL+zPJ/RV
CWnGsuNbsfrpO4nZJcXdffsC4Cte6zXg8qoienidOYzaV4/UyB8PeLV8noPQvedDItuVINDLFz9M
vlmGLxgOfDLQObGoKMApy9GdIxaW/JUGY54FYX6xqoVlWw0eMRDrwWjidYYweXpCQW9YR3HsS31W
MZXiJO5ls5exuWW81E7tzvYbopzpO4aNLOWKBN6FO/1+kyz6T0tjhXVbBHYIIQtrR0hF0mRk+pL2
5Z0C2ompVH3YJQVshl0mtl4/wnJ/kK8IIOEeb1K6RQ/nKgvoUygJhIXzuAS3Viv8oq+RuU9Np4NI
c4GQRRwyYfF10brDplZJSY3o6p+ZpFEWMhm3K5KohogstuNYHd9MAYX4e7V0ZZZ3qWTqG1QX3ckV
8a8c/keUzCYKT2jOrbV9OoapDjQJ6+dwzIXe++F6gSGjCgKbuOQlmRnlBR7ZGT2t8HJ1S6aLQHnX
LlZ365YypWg9Q0Z+EptK94vybK9IVsoreyinUWPmkm718+JNPZ4bxRWTBJoa/mPUcJ6PWDE1+EEq
v+yKzYkcPtD1vMN1adlhT8SxVGBwjg6BU9ZmRQ/C0wfd1JBKoSMNOH2+Ug65gaS7k6jyysRPy/SH
ENJEQrAIa5h3lnCjBNVoIUGRAW1atMdVripRx/marRrwL4a7TReEhgoofM26f+Wo7r+Xxn5onsQD
2k4gsOSphdc7e2bSiTCaQvmKUMoTGFZlmTsDRZ7ykAVob86n5m/pQSreuwxdGT0a2Yp1zi+egukP
pfzmf2tHjOzbhtAwQb1hwyetUY8zEunHoJxlIX89obJ9QSeQqoQKIQOYcL705TxafavyahxPcTJY
IT+XWAx6Gac3r+YhBePvpeFneZmrVn7gm2kk2ytntVaX21MjaftyG74q3KwTwd37L54T1cd9kmB8
slmOACBh/M4GeSHCa+G7XB2dNULa3uIGyIBGsOXPJ37CmOnlv8axOo00DNFbreYpQzLyrjhklCGg
FAyaZdZLUHP+CMNgxH0gyfZm0QCSOoX1bDGBlQKVNTkvA/s0yFXlCAJFoAeD/rQpjXuIfegJes9J
L3KfNOosK3WTepZeZtp3W+ZHAsD7FVyZ0JnJUUgCeE93Tx4ArP/68pQf/7r8rH/MV2j75C6HAfMz
UC7vcziJixpeEto+gCwceURJCGGDeWX70wWIMfl/CSD4o0CVHg8yvyCi3E0isnx3oXgVjEJE+eFK
IbHQ6IW46d7o1gRRCSi3JSnFa3l/A8R9uRJY49JniWgp2wJa3erxIzkvnv7GxotItaC87JoaD4Mz
/lndgl5GypCtfSVGb6Y4jn8URMhBCCHQnYRLoKhcsbEpJRf534K5iCowdoKj9Pd3Xl0pnsjcTYDs
8pKWsFZXcggjNA34FODrjmLd2K/o+iuOdR4DyFcfb/K/oceRg0vlRodhEieetIb9J2wq1CtE+iwf
gmNhcutRc8p1XDFFeexX+evW8yvxgcCkwoDtF3U0IRNBVdaMLM6hTCvBqBfQOS6wGJ678UxU1n7f
0XkDg0hEy/IwDmBUs9G3P5mcK5XRMU/9Gq7KPSl0oDGeEayC+QxxLZg0rnwZyT6nQ7mYKtXhqluu
TPTBMpPlpo3XThDFGEB6BcukzBNB/Ll9rOxrgN6xjBtPaLA6OWIUYbgDbVE6wo9eqh20F5r8HsSv
O955oAUa24ptYE6MHh9K/NamgjMGEUL1eKJe6fgKsvgEuKxNNohpc8PhXZrz7EJb1S4qUD+hKGiZ
e/5M8DThD+mEBf1Uf1hk8frUpBdgFjlljD00pEc3VvkZ/5HenRiyAuX1RtIrp7fnHYwQEXsqlAmD
zZR+nf+w6J0eOOrRtJ0EJ1KwZk11xH0IGI9rWCI1MjYtDYFrrv8zns+tkyfZpfl79MzLNKSMZvhS
J9A8mE9FFp4/BChhc6PDkdbdWvsoQnHDSu5FJOmRmVDiEY58yntoEsVEiqsPKv9av9aU7gZJwgfa
W0N4DuqOo265C61lmLMu+GbvwKMNyO7rE0hoHajc6qEkv1iVhunyctbiH77ez5d0v71p9EiUfiJ8
glZbAACQh1EPYY9LEqdMXr9MFBqOjHhzVxGA5nlddS4fFqutv9CqOHrAeMlzliJmcX2TCN6cr8Z1
5J+jsG3Z55eCXFSl7vmP5bvxmkDWKUntuN0HzcXYhj/oHsi/AL9ukhFP13nCcbu/tedIBjdEAimk
KmHz7mEUr6GU1RbWU56/8rOB6NxJnH1x7LkBGc19KpLArR+Vb7qmIhzLGQL+LLVxvzAo7dZtJPvy
NNAWobjYYAYtQoH280LcDQAoslrHQ6Y9bj/2Ck0Lg/7XhKqL0cNcXB1aYnvkXRJABw91A7Blw1KG
Ag0od1426G8Ex4Yg4qj8+tJ4TgZ8whrX+w80/8qZP/QQNmW48K2lZMiqYq7NrXwatZTmdpSATD/Q
yFedL/B7jglmTOBhicn3i+sIf6yauLanryZ2DAqivI422ZIo2Mi+fkzoaO4YjVSyAbFOxve1ewpn
C/t1A1r3dzL6hfIrTzr+R0PkMJLnCx4XU8QVtUQ/kI+tdZh7S1pCXrsRAQyGRGhCEBy8H1lhzc2I
GUrLQMMZ8/Ny5RHBqZX4f3KWxBSwep5xHSEizJt35Uh/pPLkCXO3QrvKvv0VC90PROriJpNexrYx
e3nG0s/ARvqBELHssgZZuq1l+P0EmQ73dRu3SoGAw5+Ag0VVfWoZa+R7vRmohJArOTtTzgQ+YQFQ
aUrZtel507qlV10AQcD7sPAxh7dgo3HI1NV9JrIaaU8hOW7FY5a83cDUXS6sLfvxYvH1ocO3eW2I
98JvUAUKdES44pRP+QImAE0EyayZi1kroPPqut56Uc7TOREtq42z+gzGfKXVYBMvNb8cwbeQpKYQ
ia9kkimUW6qKdKN9vp1hvxfjwg7/gA9tYzcHqLKnjNEee4jXMvnhpmqd6nlLiZK+9jFzVy1ivDBe
aTA5GKSiM0sTZW/7LuWCfLTOJyPkhGtYih+6uVni4zSnJ2nh81BKZ8rBv3CPjrOd0+UjiOLldFCF
/pXg9on0lM+CYHt9iIWmw5wyJvYMTZAdrNvtMxBXiRYXlTUaZhc8BxOg+3ZXikqQADKmGl2RoxJG
FeKg1it0WcF+ohSs0rmIzJZMPp7KL+rII5JkzC23ENackOlQ0oim0hyaZcpZAeSHZHScOzj3f3ky
QVr7higKdf5yGFuNeJI4F5pTkfgH9dFUP9RvI9Zdq58wfFapls3RIldOATX5EOBij5wzgw99Vhco
xvFI9fGZtrrP7skZ0w6ch/IpJGgSltqJ7wRHzJTtUNix9DXAL3SFFrZeSdgrblcR8FmJernpUqHO
HeKf38XcAspBJzoNodjHKvaZ1DFiHwldwCKKMeznrTU5kcHdHBJbDuIOtEIa6y7oMRZYohgEiIJT
N7dylz4dJ864xG9tL/JAi4uGhrBKSQ2XXrt9AmdFk3Z09aa6cSQguIvUxExRzeeVeSePxMFzw+iU
pyvTlwvGEfCt0/Nd60bp66e0XwTonV/Ibw1XmyjWr/f5W3XDhVg3oekY4Hdhk3iydb07sG1DuOQf
PZ4HFnLMn6Fajia9LzagfN03ugLNl54zLZPJ8cT+jCdtXvgbE9V7yGRGOOapeY5ujYT67U2dk5sB
sWpUsyqabXijO/v3Tlh7iwqugzCRQWgnb165EyLlx3VCAkxGCGm1XbSw2mtTSrULHjJFTwCtry4a
p/BeuK4OpABGdhvcC1wCZ8bqVDHnTpcTM9T6JI2csgt+ftZ48moVUSxbkUJTYGCM1OiUewYDkdse
x9Ez2FYcTY8bG57FT5GKMBdNo+VFP4ixQEdqxU3cpsZXbGkIKvBltLXSYTqIYREGpuBIiKp+gDq2
fwyGwoYcHMr+Ko2ebW0RylO1W0h2if8eQbWDEYNfDi/KKYARTMhVrqrOYR48UqFTrQsThAuODvRa
c3sM/WGTZ/b8WaHuRTJ03p/CZw70V6vQlKUA3KVI0vF+jnUptQO7fu3MyA8T2a0Y1OfdddWjr11a
JA7OsQU0vxEdY+6OtP50qzznIRUQ5XYwfQfUjCz86Ysb5nY4HCybGKyn5PJhUulAsRrE8MkqD+1v
gvCwD9atx7v9rQiR2PtbamtAPQtXt1R9CIFwc/x0YJhkIlQJi9uO6ud0AP4b4vzjTd8S+8AqxlLL
Ux66y0fJ/7AftXMYEwc+Zmrs5bMBhbMFbmLnLioRVqmjGWCNbuG0Y75K5c9NS90Bu3FShaCRUWx6
GZta316nIda9GMi2Kub3d5SaCHZ0Rx9V5zITKaJJkq1G9Rp7s8AAsdrhoeqJUZFLGinszR1UadP7
ifO81Wv6QgUCHPIiFscOuDoSv5/rIsxjFo4bqZAW1z58WgzfuqbnX3dXRF9XWTB8USHSg5ipR+If
Gr1VutQUtGnV+URLL3IhuAGmBaLASK8cAtLnPrR2ehxuRt8hoJzOsKDjTM+WgcOan89FRKPrIyyk
c3YDCLF/um8sijrTCEPaovY/C/mwjGB51j6ejKkiqpTQIGRsKlKc4dNkwLN0Q6wKzlGeC86NZ3Fe
HypAIfRfZH4E1PPuT+RZiNDJeTghq2JsDmaqMHbti0HkMQHNXLf7IkTn2NuM+Himci62G7erlhqc
0TEU5Rh4jK9fVLdGfwdOccvBIeqVs0FHLbL2EPXgEmhzXZLA71/lTmjyrIZ2MehlHnHtvJrImpi0
g+PihwJR6lJ1LNPRVK69fywDhF5f80yaw0tBK9n3R+N96o7YuN2yiAL6nqfH3CwBdn/xS164nRD0
r/6MIZzKpGn19j3l2UJVow/DIvFjMyTYa7+KICLWZEzsCmuDbHsMhZqkA2lI+CnLu+eS2saGRpjL
JDzcANbboi9md4q9je3nxVf6mveZxJGQXAZA2DUprwslRfOcESEn/30kfOY9MZjPD0CtJUEzvBhJ
gO0b0m75XBEhSYT7Jc1riYslVqjr1aIyFjE8cV1U8sOBIVqmSrqtpbZN0bi3DiN/kNOaARpqe32Y
AsLaAgMti0FD+vb/qgKKU20jtENUR/J81Nn/I+gBm/ITDVDUmGOWSK8lac5EexaLGtirTo/5ao/q
xD1nnBec7evvJPb6UqRseNoFT7RrVbVPaAtSbSDwmX0Zt06Fr3rh04w4ldHJxI4F5y4txmQ1T2aO
cVYnmtYl5D01AMdnaR2PDsVx0LoXzabrSmqBVh+ajnOZI2MVEWB1v4Fp+c7d1yQIbcMH+IdcCi3Y
0WcVN9XyiWOY2GkfNzPHNhWH/K5ujK+pIQzHXtat3yzER/W1rAS9GayI2p37qgTt848X6LMJqqcb
7nniQ9NqWYxMUr6nez431YXYjhBFMDXZbnBT4ljEch7BUHpcrsaVgn/wxjItBfgM+qH05IeKEHrC
EskR1wLlalUrWjdiU2N+784NZGbERfi3q4QRHHReDGGcpv3fWq1VZLugOV+1kDXqcdklLY8Gex07
dAlUvgnQeTgrRRnnwtDUl2DlD4WjAjtG3Shg3UqVAxCwU1WyOm4+sh+sPYAg/9YxEvEMZzqL3AKe
JLtzaOcITWixPGsJyNRlXAIPNpn91S6zUMNAiVw+COc6wxjwwotq9r0+GMYVR0xO5Zfh8oSzzdYX
QdSjctbpXoGWHpj6mzB6kaVfLfO/NBea4WNCEGHluTKU3KrB+q5TGuuHv+UvTVV3cMm4jSiLXQDj
5CmcxdfW+1ZyM+hpm3eQ3vFmyJWSJTV0GAhr17gTodhqGpGCImBcfB1ES2xwZN0l6aJ40fxS/OMi
TRPfRhO6/oJwmFY8x12o9Qe7Ph4/mDuSr3JSxpNcmEprn212piOnCy8iAQDx7fwwCNbn52OUSAx5
5sVvQmBD3isedZv1LdQCXZUwZ+WlTB7ux0bfyWfJ6Dh95tr/x1edDN4cwX4dYjheIlYBYTE4WGRV
FZdwMHOSgXMf8TB5dBTzCopN0y3eY1Zt0JvD0597T6MTO0CiF+43neFisCRQ/eOEPqu/xfzuQdUx
BMlyfhUiF7WiFeHxl/z5m4Ar75rJkF4nL+aCaNLV9TBspHRfFpMKMGanmqd7H0+TpD2jbfG+pkmQ
lyHqwiLlaAM3eowgYk9h2hreKdlm84j7UBzwKdVjkIDO/5tTcuakEG86KUrq2+inHRV+cptyA+06
BUkwcmhDDfIDVqcC+rNNC/BO7sVjFtDH/qu8jMKZjH2vkV00ibs4PHbyYljU7Lws6SfugE+bgURd
hjmx9hB7qieuV0TmAz5SmhUi/kEDGQEzshupMYWlVvU97jAjU1yHB2h9k6I+UY7duILlUIN7A9H2
gveen/0BsSo+iZvGP/MhN/gDZ1i3tIlJKDljfMnrmXzgYOvOJon53mvhJVCEtRXyKKUirtliQsW8
hwU8mEqVZy9TKAuSeVEc31pFDThVG8Tfw/+gVBD5IhXotJaiBpNbZodoYAXGE5z4AySrj+0x/zj7
AJbVK1x26xKLAh47bO8xfg1PlbyJ22iUPq43DKdnOTBYKlka5RTaiwEzF/mHJYRWEoB+BfnDe2Bk
PCUH+LAfqugdXF3w3EZ587cb3Yo5094F3fvSK7gDVk/ZtYuVjyUjRoYxi20NA/OMHHEADxSB83VC
pY7aJQ8UJ/mFVYCakqF7W7RKBoN4ZRb1vEei8FVLAKCUdQgnV6ChiauITYLu7DRdPxSZ7qx4rdze
M8BIXrZ04jWDfmJS33iC8qKqfLcvnpqxrHC2o9rN/gm4E+BG1TypJqeXIKZl1qDjyRdZFVaJ2LL8
vg1ZrhYO1SgEqGdcHtsR4p1kt0ESjdkms6U7xsKguwXMosgLd/XPg+jDxulO6kU9O9hmJPJ3gmT0
O8DR6n9RZofTg6DEeWiM5JmZW3Kk7MNs6yvYgtTJ9v4wFCuc5tLuzfze7PqterZWLnP3o8K4lwvH
vj2f7qVNRd6aS4iKKNziI+kUFhcpHDUoWhUX0T71LbEwLDJZuzBRpSZN91tTT1oSfgRWXkZUBGYU
bbyn2onM1BdaXC3lwmkoQr1gFTRUq97/pjKT9SLur447uYjgrxg3QSg23sJLXK3Y3PFNmjpZTbmR
pP65LFhsJDthExeLqg3WwDKFo/9OSqMkKfWuh/2Jd66QBzkPlrApzYw5jNVLE1J/2zeGW58Mn2nq
yCKcVeGKU8Q1rRtZMBQZ3yKdmr9y8C5E91Q041qXlHoVQEq1dmP6hrgJTGmEAFqyW3MuAQeQkhhI
QIl6OKtt3sz3gAjv5fhKoL4gamJGARrcikSHYeAdVjn9SlxreNpjluc7wE32zFFiMPuWsX7OHpvl
UdDbw+hHGEQPQo+rKh2SMw7d9JEGqZKkA4SK6EUbNp7yo96CN3liWw2KQKa3TUPsvvYGXYRA7smX
uuAj8+/mnfX+GTeKbsPD0AXb7psw7mvgU/fuKTT8ndLb5wmG/fWddiX/NXNOBNQHmA40vZyFZ5JL
4omwIsEC6DpcSSmT6RpX5xRQIEwfCd3eMfpLfaz41Fu0ftaFV5C+1iWl3kST3dtQ5WRopZo1I10r
hC2QHoGc+g+mmxnSt9escZNQRfBVcYAhDEOI/BLSpAvwKeAWFxXw8Y097iuDnfcn1+NDiiT2EWFl
29rF2ALX6heKzTwlUGZqwV20pAqe0yLZXL8q1onpl43BPGLDe/jiWRFIJSylA4Iu0yTMlW5z8QI4
fZ200IQb84/WlFAfpVXW2jmrb+AJTRqiunTLS9hmN0kgWnLV2BXVlCN9jqBKSSMfc/cJHKqbxOhj
ROliN6e3ykoVskTcQjgeYZkTb2jAHs3MWOl0a0N/sak+EAHhdJ1LpmSzz37q4VkQJCkSG/vQ1aDm
HSNgvXyUgot3JUWoBsfblPfEjgbtempYEizHodL5p6s44d1Z3rQz2qWSV3cz23inFHafQKWgZ1hW
sAoULBYnY3NW08R1aC5ibaT5R5eEyB53gr59AMd7uV59ovKQZIsNm98LBjfh6KpzjrLOZYhX56jo
GqPpLRXE/pSdiJ8d4C86UrX+c5g6h8rnIjjV1C5hJ2x66bRV1aXWLydATQAaHkqvsn5iMCB3Jqna
igUUfL6LpEt+E295PjrOEvw54dkBgxQ0oD3zWdtlE+AxWDiuxclimw8Li2Y4L7gVmfqGKZslxYcy
OQRCAyKexwueIzWrifCLVuoLk2AUghdx/13Jb2i6Bem3pEHfyRdP13SOgQESWUsxoj8s3UKU7L+e
xKmlmTpSzBBQMs88mUptV0XNxNmcaI8ekBW0s0j7T2rXezehcmyX/NCP2WF9XHFzpfTLvPCtmFxb
R9idNdDH2YSjowYRc1atBt5xE1wJWvJg71GcOjU8PbsbWIik+uMxrsmfPuiqfG3HjK4HGjag3YAF
1afIdnHuYpWkrSC4hNOQC+SQW0Tpo9MCCl8/FHEYLsO5GofO/pXtA32iAFhjrq9JaWFB6squQ+eB
qtgjfNf2bfVy+jtYks87MOBSyFUReAbd/Qg9avyfd1/bq60LUC8dYbzxU75hOZH6GxA/2rd4R0u0
I12utKsWdoCkaIq6/tu+GrXv0g2V1BidGe7dQaNam5wi97pRTZv8rOsgFvPkaGPQnreCdJAtIRx5
MDNX3ViKS/YPo3FRBjaMs/MlB6Qxl0zZaGCprhDIKrZiKw8T4vIKEVVqt8peskiuJD46sBtbWUTv
4QwKzWI84m/jA7b05/Bk2siU79sO7F3TbvM+6nn0iGsO8oeHu81M+f+lErahDtO2iyqycZ0c0R7+
gUYwjB4/bWwFCxX47Jw3Vf5ZEiSQRhyZdLR2Fv00z0WxpuqFAMZVQgs19G4oyZ474lcwXllBeOZ/
qiPt7gsTrdkdDfaR6Zr8BNYEV9jrpeVU0dwrCUlLspjPz3zhd33VFDbL5dNkSt1RQXwnBa+0hpjL
7BtapJDewZrxlD9XxnnCwVndGEnON4ZqDeoJqRIxnETD0/sfxhqQcMkx+I05J1h7w8R2SKdgWTHU
hulsTN7lIHN2Ep7LlvxJJWyYBPmxPpuatUrPA7x33L0hc4uekHEUtl9gla9ZIz5Di7xqw3GxvzR7
TIa6uAF7hMy+yz+JWg9fzZzVYeV8eD16ng0FLkRipC0y+1xXP7QZcKplZxwmVXS3ZfGzQ82YQIq6
n6GLn0why78kIUhs8AJiasuxRnnFOkBOT0yrlaspbg9j/ycuTFQ/rtdp0poXCtdb6kpFthcEPfYx
9i7CYRqPfU8Mc7YMIpjSvZCEAIvMp0Fj0vfsaqPkBarx0u9rDKiXPCiu6qNfQRD8c4x/Gm+ZEGtm
2B7107BwS5CICVHeQ5n/FsMjvyFbEHR3SSEUP0e2f9YoSUmRGxf6Q7Q27x2NvMRvlGg9icv5Sh5n
v7+bBcnX54lfgkAlgr+asuA7khaaLQbmTiRQIlzzNn5mZ7uw5g+Ig5Q1HGpmrS6xhLlv7QDjTGw7
Zsv97/7IXGBbFxIDsAHWeDreYDCpqXXhF9Ogtsb28BKRQZk+LuK4QjAZ3+5QsX4aCYLZQuwISRU3
wyXqcUK14SN6bmZWm2fGzCUFCUhm6K7VORuuEoBqlwNZiElYd/dVDloSS+1k9xnfcijOJFor4hME
7CTLNk5+5O9f6tGl+dxFpPjIh94h7T/UoIuh53oaLmGWCdpad+GXHzHZ66/nDQVJFUmPxTPwfHIj
xKyk4ytKkIoaOZG5CNEqqyAKhmqCZ68B7Jp6ihzt6j7gF7z63lnn0SJ1hmwUGFB20d3oATwMp76c
g5D1AqSxDc9hvwiCvY8D9831OATvNE79k1RAT1CzjH16PZ5sKqKplPPh39r7y4vC8JOr2TViyz5b
jJ6PRGaSUgC/UhwLBISTldykzu86Q/JPEmDVqhaKQdhqoGhPHaXAauFeP9tKPcOXscszp18JJLBy
Pp6ykKPgLbOAdKevR7DFaUV45fReW1iZQhorPkZQCmSFnX08YtVpKPDt4PDncVlR1KHUcLmG5ii3
cCoPNY26rK2MSQ9ewPHWqzzw+GTNAYXmCMk7OvkYFZPPpuAeLEPOr9VKa6AklcjwipOJI9P0PUta
74bkk+7Jh2rgX9osXMk9iyVG0wXdVQahhtVEHLjYWsuq6ueTJNVBibv4+dUdpIMo/ESno9b5f9iM
YstubwUT5kvJnQUIR69KbmVgYw6GcBez4Hu6TIktEyQj8uN92rgKNWPa+wVdqR+9YKXoJyA6ePOK
DaOotgYlfnBf5F5ggdf9AU6Ev1LUYcRSK6P9+oc/pYQE7JefKz+5NPDi+4icI1z5LPtNq1vy5FBe
sB5XpNrLycweoVKI7ybR6jQwTnNAggi26KHd13yW31W6Dtj3Rg4eU1fS4EpI5m01yV4hoRaMnLuZ
N6fzUxl/HiSoluehHqUyYfY/7CPyae0ByMcvWueAL934Z8sxp2csRlaLamaukzkqtjvMkvxp33qa
0ou1o+8zLzSMepYiihwv9Wzr3jDOxgWhE9SrXY5d4FxoIzI9yGG8894jVF/tqLe1ak4BZPHRh7Z6
nFeOzOx9Hjt/zQC2Twu3vG27Jl6ceAJgIKjJAFGZyI2LUbHIiE3yRJtoIKD3TKE6roPDLUJLLEs3
GJkFW0rk8feqPEGolbxr2mSGEf7xmFrH7lVQlOsyxOyOshEhak61IQ3utPL8B2reSfnbpF0WWNp2
hXb0omwaV4AfF+/wkGqD+vbpD7zYx5k7ZnLSwmvzmMDMZg2lvnJ48/F3g6uJKp7fJxmg2aNIMir5
cid5anpBzoSoIv1vgHClaGIa9a5wBkGn53O9VCmWkxeWHWTg3ANIXze4Yk/CZ8CbNymWJS9COjYT
pWJQng2nH/hdJ6aD2n9aXkFh04RMUUD4i1W5D9V45Ac+XMW3YUmrQGuKEmvIm0ylCrTwCTQ+Gqmi
68DgofPbEII8ulJicJT21Vot1L7b3t+biLu6LiaZWPrlr7bmyyLeLbldUYnp6YI7SA3ILj1+vhMD
tNH6B70FiWQZ2Q0+L7/mWF5uvapcSjK4nGDHIP520pz/QOrI9tl39RQxCO0e9qFXoejJkgcgw+gp
yiigNC6Rs2/DLKKdLpcV0WZD39KGDJb997HPVzpiz5Uv+etJAlYcq90Ty/bHAq9RoalK8NpxNur8
k3xtj5UoHSu6uwmjISWwrJ0JKcS0EANtgb2Ngxw/sTslW7pvJBLZDRBJG2SV+JvOrOK72mmss0SU
4lJIh7kgCJ/gJpjQvrlxMqlYR6QJHyBwHtU8Aoqh/NXeINiSCukzeY1nunDFCH1CWZsF3yd6vm1K
CoDpYJhNo3p0T7gJqmirUWUH5/EH8SyALrOZT59K2WM2T5QtrTsUhPo/JvvReS9IpW/jgZgRmmPo
IPli98q5PGWfmUSRIdRNnUyt+eCasKlbBLCgHejmFCnLip0vItsXWsEGi0YIsRikWffdnj/TvE6V
CE6E+3mRSnxrPEEw9tR7h6vc6t8ygFZQlDyZ0s26HYirjhCD5JEu5kig69Q+PQbnmFQz229kH+u8
Hmyy23DFavkcT7VFr22Slfecabw+6mAyd9aGqVS/OlXqNNB5PRw+thQ7lVMNBf0pgR7/t8Bn+A/1
xFTboUpVktXVxK6DWSCPMRnNGm2Yk5gncNvi5rxjaZxy0PtgHHbLW/1aaplaVVMmDIHRohjP2G5u
PYWCy5EHAYZQZqkDsbwDK/PQNYFq/wBPBxmXhYLKQJxFto4mapV/+ueRqrVBuXZgwpXR8673SblO
iVb/mXMcBMJ90ePyl+XZPXBkPnnWDaOAVJbBpJFYtg1DV+JiuXW/Pg+CYb+eVplXVzC/kxyoR7bp
EDcta59msqr8oPKZb5sIO+0ZxMGfCtFYSCDILJNKxe6iVaVJ+hkNO+ETx9RYW09aanCgY/r8INkf
KPaCvAMFWp+M+3ueA5lVT9xkqyEHnsHWBt0o6X5ZkCGcS+ycE/jLaWLyjUHwQFw9riwQ43CIW+8y
SfbwfhKQqBVAXY1jEwWbN+pifh69jrxRjIak5HB7MnqhgOf4Em0KKq1vH1YwS5z8tR4hFAvPf0i+
43cMiQRoRRtrr+P0C2BEbN4w+ixjxhruisJbgYj1v+Ga45EsZ85f7VUQWXBp/dXmRiu7+B2f7dPM
W2OLb57SpizNwiJuXUAKEmrsmZ3JMSfKu1Mj+hurV4mtayNWPYsGo+ZOqh6Q6E2vB/nHJqm/JQ4I
3iIgY/ePwqijMz/bJi/ddNDAX2D9VXTvSB9FsCp42dObnkwrmmG0064UCeB/zTmfDRubiJL+Rfoa
1f95IRGkZhKuLdp3D2HLWGmh80FccPIrNV4+6MLUdWU4FqTWvFdfY5CWN/gp/YgTPLDl7QMYjwPd
HiUCesUqgt7zrpVXLFsjO/6xw8BCgwD91nHAgYt8o++nUw78cabjFiS3ZheUytdsDWcSCbZJrX9s
2h5pBDQ/QKWYOJ68oEQOeE6dqpBcOzXmrgTjo30gqO74VGXiGf95CR8yE2oS4j9lguLVIMs5DaHF
TaYNpEAiDMTEXUqGXVCFgQhO3/70gAUujiexQRwtxLI/jVZftVZaqFtieIHZ+ST8hGlMJPW7VYJ4
u2PTIOCfmMe7m+MbChLn2yoREYcjk/55cCps7T+Bn431oahc/lDUqGDizbhJOfb/FNyCPA8LckVZ
3DjKslVSKIax6yNplTWeYFbiItSrWyKL/F+XDm6bBPzSidEdi/aKw4ej6VtNRBHsCg0DKMqsewDT
5y3WAfoLPNNZSRv0WKLSYGr6iLUKiQKlFTNS+9ZHtLcdjjcm8pjKxsRiXriu5+IVwZ1+ATlG8AJz
/cfI//HOk/hrjs1kP9o0TzXe53lnRapNAfYvLfXCZwxan8dE7l86WN/sUGhDjOYsa5mbsUbTHFzg
ubH2VtypDyCG9zY2TxzhHsF8cAX/hrX0c2qH5eqRPxAp94uiHw4X6gfIZbOowBmRbMd3GcSjIGlP
BNzmuK+ROHZrSF7p2TvvC7TAtKJ84zpfDnMW/EUwmwlp35GLnZHpJGgSlE0r8gDgfkMfWRrnwsQo
9DFlywS7mEEWzdFZxYX5ReGM1Gp20N/nHRqZwkG6abL2VwW27+FVcAIz+LarWgKJBpIcMEX0HkTI
lX21LwxOexhm4vevKcrcoeZulwy1NaYkFEKm55V/Z9mxSFK2DVClsnA5ST7x68UMmtUYHjXTw9mn
u5nupn0ce6WhMWamIvO4wj7q8LCmTNkbh4Tb+Ka2s4ekx+h4Se5aFMSrt37e23GcYt5xkzPF8zAX
kXc1l1fnkeJnx42pqdx0t9UezayZh4KOKgt+uceZ1lZWeSX1de7Yukm8XNGy56G9nTT2UOqh5dba
zRpSYo+LNO6IrG3ifkhIBuVbC13izQ9fQx+hj3+kiT3XfW3q610DURrw7Upkwo4+5tEO0MItUJAC
U0FIKkVfDpJ6J8HQ+cxSdGRQ+shJjRvsazbwmXaLHXvOieLVKV2KgzHeB6C4pSTWXXzf7qxGDmxt
TkG/eah4Ac70xFxLK8zJNT1tGSIHvpJAcrFI3kA9ijPMp4UIAGtohWMaV6CDpf2d/R5xCM3sbBub
ZnlqwTnlDDXgODVFGqOu0WNlRmXPkWS+xzXBb7xfZvBYAyyUK1gtMaNWj9hr1ycyCUSjjCRZ88UQ
iHHUW6CgOT9Nk02LqGldNqoj00nYXuA5pmzZDd1RfdQy7CxkieMUIxgV8jw7RRSllFf+uVx0F5F8
vRowKgAZpC1yArXx/Lp6nw+YuGkyig33XloRKSwmMrO1JY70n6uu+qthtNXoAPcEqBfWGmD8XAvk
PruNMifvsTo1Yw0891E84Y+bQS7kHyYorxxZBn3MCktjRowfiCyAnl3Iu0ckbTQKsQzzo6B182aN
uWXQYHPqaKmWBxsZYHL2ZkkqUq24DAj6io9F06CXdzq3JwjeV6VhOjAOSgEdsTmQQ9rUR0r+jsTm
hs/7KTtiBEt2DLbZFSbBFAgvn/5d8urgsYAv2tfP88vQe+2b1KGALMsg134ef3sAHyXpJPNztxXW
igLgP4zabSxFN4CCjQ6oT8pDqJk866gR1ZWYVg0cd1COzpY1+U47FIgsyAI8OlsCmqh76yeY0pD1
airR49h7CZL8CrTd7HOQOVpf+bHinEzAxIJen80ZmDkdJ+vjJP5EZRJPqcGWJnF3YQK944Jp+c7x
ZEBvuejHWXvraX3a8YAZH1IpCVPXSbg+oVcL2vj6uGviJiiv1/6TJoAwFl+gv5biQtc9HzrLK5YX
1sRn48TplmfguxitR+se3bGt0/EVfL6MgGrvrp18eF2lPm/NDiww+5ITNYUMTInec0GjEa7q8Jws
4/HObNmFtX9INeUXldSkIhzzPSul3tjHkWB4GpzJU3ezeqtybDbOAu2lRbGXYV4lPZLOrcwWog2/
7gnLaaWxybzdyBBcR7AFHhTKxmysMjFnsZR2h1zNhxpn+DgMlCjiwV/SCyVWqIHwUoML8xcDDPIv
rRiafBshc52d6/H1zgO7VJabrEUKyzumpjVLtIlep0+fUOVPVlOHEaRPHwng1oME1i1lLKWUmADd
Mwp8XF8RJKtI6JcXsmNGIsZdv6cYyf43YdipWs44kywkH+uokHyJvpAxvxaT8yqN4RT5CVj7PYz4
y8+KXfpdN+PQJLIYzKhz516dRwf1NEnrvy8AFqEtE6Z+0RKzRea/tC0Msh2m2bPi8XiXATwn6XKA
EyPp4iNnkzpIdDQHg8DGyjbiKB8jV2/Efbz3+eabqzkfurCsMrSG6aNQqdBk3pDxzZ8NtYeIEp9D
kr9iS3v/hkrHlwcljECU3XPqErHo9ZLyFFM2j5wO4k4+UBGb2Vx16i0gRVifysjF0RftGj2pVazM
tEuFcJBAOYFkmoxHHL0PlgwxkflbbklfjM5GSx0sch/4La+CV7aU8JDQ2tNYlosKkJLNo/UbdAZA
Bb1yDZx4XMaqinZz2agUi6BVjrG2AcN8SIYGj3I85r89azpub4rJ/DTRhqgebM5j1gGJXbhDOMzo
TAFJ4pB1LhPnpufc3anZf9+dUTi/3clicwNc8foVSmY8ZDRSlC8PfheFKgScFnKwFvbw8GSzAufH
T+yOaoM7vAbqcd2Z2dx6azKbK0XdCcJ80cPEAVQYkRQjZPo4Sqrg73y0lEUofudJNILIjR4KKRm7
kH+E/HFGPtd4YNV5Uk3GbwC3fToK5x9u62oBFnAUO/J+iS64/QYEN5plVy4rS92zVG77WUUBh61D
5NImiZRD+GKxX4whaWSDSkKwHKUAooBVMqXeC7Qy59LCJYzNtYiHcxHh8BQFmXK3+tQbuFcTgge/
9NLaZee2mxwRMfY4BNz8osrUtpoKBvHSFswnKXT5gNMCb9arW1s7PVk6AiaJmN5RVU7xkCxUpurZ
9LI5gO2Ct+2VWcB+A1gR1RXhVh6it4xvM2f+OfJgIl3vYmrHYOUhUEtlsQoUX/Z8cZjAy1d1xNyZ
DKP5NC77/Of7pN2ZS59lliBLVCPA4LdI9q2GiL/TD+OTb5OfTJi9+stAHAavC7Ll2hpXcFRemgTx
La4Lo0T5InpvL1BY3aQrambAQHfoERWic/Ba/ebQhfpO9rF1lE58ZfCwlbVlcXiIPRxLaCs4fm4P
YP4SDeFYiOsZ2izdkxDCX/LdMBbhtRlPmK1V14FYt5RLZ9mmdA6TSnu9DaQibD/s4aQVIoFa2XTU
vfqlC7S8rtZ93EIbZVLRtEwdS9BHsVB27lfOdbOOLv1KlNgb8y7XnLsc6eWdx8aGPENVTafN7jcM
kj3sM1TsCgaP65RoIKWIDHhjBhNB8cejmrzyfEOUguuTugWXH2YmSvNu5hd9ccvQDbE1uM9ZEYke
VUuInA1727aToeiSCtbiNKDh6cUe+JDdDx/+8ZKdVSK7pFEWCjWB+n9eqFUQemZ4XXhMyldwdIFQ
daVx+vDntxp1pb794j1NDF1u+G1YyCI+rjOdOIqFr64KO4112623LphmOtrTkXabndQOGoEjr2JN
ISxaMLd3Nd5IZmC3uE/rcU4Ayxjutwao9yZmUNCKvqgECexgFop5jjr6d3aO3v//WjH0kQNry71h
7s50Ni5teVa8Rkxz2vvSVXG1GhKogfVdFqiaWd+DZ0sMJG22E9K1iDoFZi+MRUq0FHisVewX4jfI
7WDoKEWTRGj0NZH3KH288dBd9FWiRqNPAFaRFm1HkR89RmiOxl0fADsPax8m+j2/ABC8DaN8M+d4
5AC0Dqh37DKKFGfjQ1chaJwP1vugf17dJbUXUceqM/Ppo7Fj+r08yHEmUB/iG9qSdOy7Zkbh8DmW
3jBJwI1mA7DA6DeZbTYRCc2X5DtGhke9pxxeQH7IvyG7ace8ygKT3k0LIaQ9Ev2nQeoi0SwQ/d8o
vUTJjj2J+puemvC+9ucM7WrEzhrwBh5iqrvTxiJMHVvHztdsHp77eTI7jFGyTlLCjX9+3qJQOWvV
DLFdfzjVkzVHMiUuFjsXWMe4k67GymUwdOjwe8Q5f/RTwlghm/fVOkqvWNHmKeD+zsWHWOw7RyTG
oYi3+HtNesdFNRyDOtOG1CKIpPQRPZ/3ed+dM8j/M1k208p7mn5tz0gxvJbctKBj1cItbDr8U3e7
n+Xg4RlFd7Mrr1hfGGa1iS7+x0r9vTS2rkTG8sLCDu+rN00ZCjLvtSFjfEkUl8b22gtK/vJW7mTL
pR26i1oFvKm8Z6Wpu9FEAasBiOTdQ/drK0nqCw9djumQpDL2wBu2/OFFIS4Fav3NRqhFWgxQlYr+
sOHrFYeNJCHSsgqdoneWEfcCOFyROlaoquZvVrZzYJjMAbTsX0+qLjJYmohEchBu4R6lRyCRXXPH
/Q7zeLoERsRluTCuV8zdhzmrcZTTt9On+Num25nHdnFidi+5DX7aDkA+sm1mhW8Yd0710SIXVMnr
sdyGdmRKKBksdfWFckF8S6o724eUZ68lIHZ3qNfBIRmUZgdFSIztq/CTCjd8OkBYO5mwPxx+V41r
+aZy05HVdjEEOmZFy0txF6J5KizXsStR7yLAclayexS78kq+xzGyoFDZzOFcIRMA76hQ3IY1BMFb
LkTd/hnWiKe6uGNHyYAUgRSTVkyfEQExIEtOVRR+Cf7JtCYenIf5dxHJhKFU5YWpuitx1SR3azjJ
wHB9UdkWL/2Yg7etMX6GmsdG+ZbjYST00ZPlf/WJddiZ0zAvApkrXK5T5+O82jOS/RvGDLL00rCe
q6O1Bu2ZKlOnqMI2FKKU38zPIz3D7kP3vMeKD82TcqhoYEaL6d7jREMIEpahfvu1Le8nKa52xl88
tJo2OKLm27Srz+4in7XXOTWcRYyM+7Fqb8RU1Yl1aL9MxyWqH3KE/KBNJsQ/ujWNjWYbKmFlbaKp
GmurqVrtwy/dJWooelbGSlqplQtCPzrEs+6OnX2ixC9MsAOa1kmBvWflqng/gOfXDbWu3I96I4DQ
dDwu0mqDSWAQUg7I4fyCb/OjhiV9/3/1OATxLt8JqXKp/MgbN2bHlfcR8CqD4NQ/2t0ogRU6m+/B
e7X8bsIqIqWGZvInFgPaQV4Il3AN1UXtW/+1efwgZUX1Ku1buKyyw8He5a64UhH2n9pQLDtrtdAJ
heJo75z0A2M7I6jtN/IItdgKWhV69A5r03Z40AttvZE1497y0DlY71KHTIO9j5uSrwjj1UL4ytZ6
1Zq5/fQOdXVdthsZVzba3qS6oh8VcY7tNQRMSJl1azScevDoPM97elKNiw7/pC7KBCfW35q++kxs
Kr/Hnqq3SUmVpSmZVMwp4mE9veBNgFEmnQD1isO1UlPNh14Gw/+GDNUxLO6+0paILj2HM8aKxihG
agvfaKUfikcWAAf0v156nt2102h4Eu7M8K/DV2J4TJ76KtEG4O16ET0s694me53rPO0I53+dTFvQ
4b45/yKg8dTDk0wJspfl/KdGHKvmbf9+di9MKkRj/1OXi4dcETMWmeJ+p7RO3Vn+MZFYUrZHMtnT
Dm+wWNQcBPyPHy6Cx5mkQBLHSokDbhaVaVkA6wKsJ7mC8iiZ71iELRpi0urB/TOtk+/iJXZaYkbL
IHTJA+IMPgBnK0Wh92jpqqa3ipg2f+BOBswQ08U5lk2oOI/BldEm8iMdDhLtRKdv05XIkZzfO0sz
tuZZchSBNgkjXF8MMCsI0ardj3l6UnjKGx5wOiEdaXfXXAHjITlPpHhj1UzYNjpk3ZBroYjvv0e4
PBaEWwiCQTZyLhlbmE4qZfUKKIGu6IhSOfKQ95bye11ISJJbF4NKhGkS2RG7fyAkQiL7usz3MP93
V/YlPPrmbGWE0uaZxgkoG9qG9H2NC+yL8HORrl7lcONCuCVn8nnjplpnInLbOQx7SfeO4GnSQhZO
AOmV9gnYoo8A1Rug4CZK+hrC5RYSmwrYTkleEK4jnFyE6zuHntu0sKi1yM15QLyaxoMgc6N+6fxw
eDBvYaESyd37r4qy6HTME8ARioIxa11jcGeX3G4MGoDAHjG1iGYUQRKAENv1YN+Da17Y6PmCRsa9
9oiGk7z/vabooEyOrwqn5hInTtcr6lGFXaY4gXKBJcYztXvGXRWlPF8JWzxDrtNTGgFTMkbkkwbX
cCQXT6Xn18pAHsffavc/kSQvkYOFLNwPy4LkSX/HCc3MFEB8Dm5eWvlxsf/beJ3+AFZycF2Jdfdv
YO8xU4oTRCXLTqP/d5f8aQWnbK55WPtT9UAwozMFyU9PxOQuZYsY0tGYb8eiQg8oA3iO1YfpImdg
aHcHKmSZEb8BBi4ySIohrPyLjL75cg5r/DbZJjT2YCmOSn76pztZXeH6nIw9urHd/vj0IkRGgCkG
AnbA6KWMHHMcD8kvcEBounH218RINph+H/1tCKq2HnfZa9AerWm/Fo5afk9KD2/M7HPf98Wf4m17
UWEBZu/mygeB2iHuDkPvVqv78q+KFPWiCX6NyqFLxAZlqMtTmIitOhMJZ6Q+RwFfIqD+dsRhFYkk
lSEheafQZz7oQsOOrhOHuEnF4qFrvxhMvq+2HcSzt8Ll1NnOAu2as8G+ep6hdshDDcUyyLGHgOgE
m+GnxzslhD5s8SRzTOeCtfqF4xY51zRDQZwkX05dyrgex4hI80YnmQ87g4+me+j2hRsQFQH+mbhl
p+11J/gpkBlXxUhlqC0bB7hZJRcijBd16R5u5SBJfjfSNE9BU1iMZYvmulxbCe0J+vBKa7+tDlEU
+QCD0WUcCHgWg1yK1APLABOyfB5LST+Cv/gqci1mEcNkdq9wWt9RDYeIgadSgXnu5QvbO2exHOMM
u+LuUcAjD8CQtZEh0dBzYGoSosDaxH38uY0GPTOjiC89wgW0Slr95BSr33Qgqva/t1GYuk8ycH31
5H2El0oo0NEblqcrJJP5fPP1GIG0Z5EYvjYI7DIuT2uWghnGCm0NZ18u3sjElNOYL2rOl1x6j065
esIr2FWeb+mo2/A8zxvDNEw34BvzEq+6B5Uml8/INvFhckFsZopWgZB6JcrZqmEOt0wQ4y43JFjc
jv6dirdAaSW+3Y5PkpAVLjYTtixlV7koh2mc7SzplxZdy2+vQvObB51qswopsiSeaYpORykg0PEH
lkiX1W7QARlE7I1bvyT28aBBix97YeP+xy8Aw0QggXgvESSvmll5KbenbUVenRULoWs+NOaKbQtm
e5lSGwBUlG68hjnINsExdl6hOpau3L9owrAFW83R/CzNRMrFdQ44K9cROdSpAhsZ1qyOLbHLNCkI
vtukhvRaszNvVLhAMzR2/J2WiukIbdCJHU3m40xnrUiPUP48mfl+khpndes/bmfc7QxBXrdKoRcU
SpO4XJKSdbFu+KVTXdx0YTaf/0yAixQ7DwW3Fs7lMzcuiHUymVB+srNsFnCM/fsjul1cPYhOvtQE
mAkur2wfxqjjHmpW8ipGdv37zUmXpMd9XFvDBqVOygWj77P9eo0zFbZDbAKRnVTlqv4C64d9crPM
1dlY0ntDpliD5f5bfl4emmxGwiKsdOGnccks+O/HoD20Dlywyn9ednOZARd6qfytxAkTc2zAuFO8
snaaJM66jURhzWaBQxg1Md+w3SEyZ+xhvvB8/BOrcbTFxIumIbsQsasHH90V91+H3Z4nJGXcSGIQ
X6SegNhi60dtP2tRlgsUO02C+5mrFUuic5tjl8+H6V+9nx5dngj2dvQ597Ii4w3L/qCkgwrYcHjH
8UJb46S/UCLKu7MPI/Pv2bmrNCYsGUTUKXBrH6LbUSictvPw4Fg1F8LtApgnPc7Ey/dRRbDVXHEt
QthfQ03YnhJOY9xGP1/4dLJLVmsAIt5GZ2OgNMQTHznPFOMgSENGOpHI3oIPnMvVpycbVOUA7FYq
j+jzgp3Kh7befkV7qr2lvXdE9DW2AAIMBcfIbtLp7R8FJpg4nJhGgp1dHBH0WLmo34eFbf4NbHNK
T3ESaJphsjcX03xUg5o5VDPpwVfQ4O+PaMOtbnXU81NHZxfLZL6C1lK1xKb24mh34SI7JmiG67/j
Tq6kdT91c2gHgxkiMSKZtK2qjeX9ngZD6oChP4eCAWJUrH161KuOdYGYn2FJWBBgMpN6Y9o8Rl6N
QexLV6bjAMNuqqOk/jw6wkGMn7e84xt2DoZm/R9ulfufXQTcAeUP2hTvkUQHybqAC2og3AkH2bBX
GqSrN2Fqt51c5sqcJ0/T2yHOyzWaJsVr7lPxB6zotk4xOTSG8MdqJXtE/f+iXWUAnhEpxo34NFFb
Aa3fP3XMj4Lgzk3Octrq3bGkqwNIWbRa65+56NY0DvM5lhCQmr0vQhStywlrF+vJGiY6YKlxOjtT
abW+H2wt2nHior5tagPcDqI+HOYbg57aJYU0PJv47+rBxZa/cNcKXS1Aqci7pKiRQgjsVvM8KbjP
KPMV/8X9swz7izL0BlILeeWDZLGL4KXhfNyOW8C8/a1tX6gUTHGxtzr2Rncs3f3Io5P+CzllMrMJ
ucwtN5wyJNObJLCjJieIjpO1RHa9NQGUiBxGJN0pIREkDFb6vhifbt91YAUBlecT1R6FRkL0ozhC
0xiXsSitdx5xu+QhaJQ6gjW++lgnJnUUycpltShdAmn+L7RIfn6bZ+so7HnyG24jchXs5M4rZ7Bm
kJss1wrclCrj99gzv1XvF7TQfNeKpEgjbQfibTaTkFk0+C4GJEeXcMmKEUwyQXMZHIDXo5svF6In
Jez47iEbe7pWc3/73Px5yL8P0VBXgDRfP219ZKy54flipdiwSU35DWVFGXIw2bQycYPgDI5ZBMdC
TCBad9fje3zVRvTPpXvK1p3EgV5AaZIgg+mkjrd2gkLUPIBFtGjmVjked8bIcgHYX0GpGBgJHX67
af9K/fsIMXknTBDokbZ4g4XuzttA7ZobBWXAKT32uArmsUQQnGXjQolhTCxXRJ5zWW4pDWhGNHX5
yGFEBQBO3Tnw4Qx7jhHdn2Taq7453+knyobmDcMO4Br3GtUK65IRnPwwkjsQoeLm46KoxLnzhSSW
Mt80ua8jgmrY0PtJPrlbcEhJMoujfnlg/gn1W7frTP34PbZLspwFL0gFkMMooG9CCIIWw2PEqUYJ
boVCGCnDjO1tNZa2CPLJDdwmsjB8M7GxKre7HDwk+SlGHyar69rX5Nx7h8XYbewjAc6VW5eHGQlR
GcJ676XO5wqkth3b3ZsTzdNqPXBgjnDryaKSdXbubcFhoqtWHUSyxZY8sbpbbxAE0Bnp8nUypqwy
rYas+qBZuHg7eiFaK+YTDfOxSn2zER+HXoLMdYYzoqsShwBBI7zCgBwGGZXR4MS8fTSoAFtvyUiy
1dPD+UNYW9kTCkRO2uJRtYBTnykjy3d4Jxdr8n6ycXLLoq0Mg0sQNyBNw1ldBy8YLdyypNc4s/ld
Efg81/8TdUzmoIpJxbq0wUwOXXXuTWIXLz0kqceI9resmwi44zdhOuT4fBZJC4Ve8tGDRkb2JbKW
AruHazb7B3D5UKnGvW6wVRKKLtf6Ro+aooVH8PXz7ahLpWoY2edfd0dQA8rVlZkQ3/O4XQWFmbwQ
Yt94Em6Q4GZ26oThJqmluv9/Hhc5ZRbErO4Hs4Ef5ox/L2UF5Ufrlr9fglm9tMIpvYeNJzuswIFe
wM/OVyHIOk1AQLRVqd1n2z7EyTR7e0qrJBoj9wiGxUKYr7T43scAfH7z8zOddbvdRPX6YloJL2nq
hxz/QxX1YSyvy8vkoN8kZrTmvankuMTuSqsFihyXkvxAbdn3JIqg4oqVO4Fzgxi0jpq0ZeUmZS1t
aS6Uqo8GtYrkpPwk3PriFbvc9uL5VfQNVN6ihaw1wIsgV0S6DsJCYXyEJ4RoLXuk6pGb7OxkmVBN
JZVKCYjtqvZriobeMvQz2c/YEqwPO18G4AtdkhLhQU6ZeINvwMZ19E/8FX2eBGAyabPTsfh1t+I/
1J43yf0iuX551rc5jjb1Q43W08wCTuAYc+wiE/+qMmYUZMpYMZHW/DHPM3bNnPnn9jYlL04Zb83T
P6jWWluESfSC9WXCfFhMzSuNs1023rWvbE3xeoCuswftB2hetZH2Zp5v6SQm6tckVGY7eN7jGo05
268Is64M7trNNo/UCRLM9zOGXFaSrwC1VL1rzx69aAzrWQ00qyK8NtcjPhxkmmnL+u7HLUx9oKtD
17wVaf/f7bg3OPxyzocxCSk3aXRCBXchG6hA0jJpmn1DcX5yy+v3/0s6GoD8moL3ddsYEgZtXVx1
a30DCCTTcOndiRCrwaJtpqnUXDZoRrB2nvzY++/UyTNokA4Pyf6zEKw0NdjwsL6u6eazxfP1yzm0
9M5cFouA/IkDptwqPmkKoeNXT7yXJYD+fEkxtHd0ziUve7TDkwTmoT9QMQzRihnTLDgkx3itL576
pDiKKpCBCxlRut0M+suow3gm8TBvWLnMH3lHGlZuaWzwKBQgc1cpG0rWqTs3J8e/HNBXJsRba7FE
6aNCjVlcmzALJWw1TX9Eb21+wmFTJj21P0CFtb2nHlgae/GL00o8/M1YX0tBzcd3Xrc/klJ13j+h
OXsP6u1LtSYbDJsO8Vp2TfVEt8PCbEmlWb1dxv2b763nlBr3OkwGqljK+YdHUMWEFRDjvIWXsA1C
J7Mw2GPiW/B38Xb5Tv1ZbBYnV6dF5a7fheEk8Y687MprB2gcc6PJThZaeQ0idy2iUvMAacdsMrV2
lZphimeuFKZLR7cJBHuzg1MKywNmScaczc9y5o9ohcFpuGzPSxuh6JOq6Jyk8AB3BNk06DmU+gFa
cmT6e5buzsy5Qtcq6VtAUz+DZZ3o2wja728MvD8s6ndhbGYu/CojyQ3NO5H6yft7TmZFOyuxNyVC
gUpvuoGlKhTslJEtsSkEs/r1qqCJHpiuKQsb0ZRWcYnt+V/vw8NbTgVTZwD6a1qEAjli1FxaflzS
55NY18L9Co9Z0KpgJUR8U80w3Gcw+8AetSigw7pWt2SkmzjPU/n+oX2wXuQOP7XaoGFFfMGZwgkx
/WL/PtXfIdlF35jBwwNnOdsp5THBAR5UxEjheKAXq9pCSQWQnM618Px+PzZZY6+UMB8suTwzv8WO
1YsuXkZtb+Gevf3FlYXFPdbLRD6hXH8QJWgULDhiV14110LTLML1904783OxYy8JKW5MNWuKtw3H
BClA4IG8gVFiaEqZgzcXF/Xka6sOqiCKUVhFElfKjX9Vn1xk3JvNFRFnFcMVrHU3uuv5MvNOObAk
orrrswcIPrBj2O8wXm0RovFOwrxGoZ3XTc96hHHCr8QZtehmXgic8NCr9kI637YCiVXLtMF3vYXr
DcnURZw9KLgNlNbpOMx0zCbG0POUcmhi/ffi/wZ/JgSJ6GNwRYMQ7fnUeqltEiMU/aIQc+90aALC
AdSjkhav4oKge8zgqvdBx+ddd6SIrm1PtdVumjiw5Uzv69+hjboV0x3Tow0nv7OWX1PsLaLfFjgL
sctyR73rriHMTlY+BbiEJRVHEpBFHQvQe4N9HBfhsTljmPxsuZeE95VNrAs0HUkOOkzclqC6KmAw
bXms4HvoEaq4lL6jIIijJZN2dIp8dJDTneJqflz4UEidN+mqn25jYWjediEFdYQq5GuYJznfInL+
8TfpU52UCyQPWdqgcdOdzulJLW74w4lYOaQw0tO86iq8luWi1F5nKTC/7pRoJZEuhOivehBtqshX
T9LRHi5Poqk8MRtYo0yD/Flnxuxi77gqq5qVYU1rU6U1ezwgoHqT7QSPxZJy+W4n0wLVv9zhFFa1
gDlKDnl5+RoCw+nvRX6Muj+Vzuu+U6St+KCEfdCMT/N6UmxX7S0C0inLwszGuzgX/fgt2xy+ndH9
NogBSoMmSHUaW2c3MWQWmc7pK1ngntQ2XfRbj8NUQN8QXa6qIfgZhjMbFYjmUUwX7ag5zjGMz9Wx
IOvIldqNDcq2FGSMFVApy4p8IoeHi82FIYDKN3NP8AARLQ1R6OsfsbzDhaCY4FSmqTIorBMUk54n
Y0L/j3JCFWcfVixk0pcBjWgT/7AyU/KeOP6pXj8X7KBp1fiRla4LNBRwFuJCO/U/9hVsw9Hst1CR
9e4oz1W3JCwdsLoNV01BcI9R55ijIi5FguxmEOasRKQGAmOXZytTNO99yzMrNN4cA0HNFn2IvsBY
oYzIraZdcHt7FD/DmLxFFDHN3Eq7VrRtJp8aM849GXS8UW4tff9T1OHePTNjhC92znqHg+ZZJJhi
HbAY6oEbbFTOFZcKtk+JzigE+dD33NHDwWnQB0QTFpTca94uvcV4lxJ3A29gejpWybWD0wZ5cYyn
p+7u/aTTwmVjjBaBZnpwiStyBBF/CzC/dUu+p6yBNfcWAwL+jsNLvaCvwUKssbdv3PqyRV08eB5P
fQhotxyR4TkyBq3WBIcyvBzrOxZGjPXQsMkyLlFlk0fP7e/2zFB7ozZtVZTZCLT7ByyIBkoVe2qT
8y6eSD7hokPyn+QwcxghJlXkCEhkpFPIv/lbpuRqGPbcReVz9EXXy9Hhc/gh6itH0MeO/K1U0gET
hNVWNKVBOkp1EEoec0tE3wtWJ+ppOj0P9sS7PQNVHXlldyjxYgZH6tKh18U99RxaWuJM6tokRwvg
twHvKl1la9K+FofVonANoilcXaVnQfwh4VvM1m7mRDermk8X3FMvXU+cP27ZvbY/VBUf7klWVVGu
ocXi5gPsRDyEAKOVUlEPThkLfamImun7k8he093UzkhLwUxDkxpe8nVtmsw/u/7/FfdzqVfume42
WBNa2wsKWizU47D4tR3/inRvmzukjNbSQe451hPsRCaAc5EXkC8FQlXVsZASRGw6j9QkNe0KbB65
8tOaeiPK6IU0bRewiLZanniQV2YVQhy5IQI4FtYaQ0f110HQ0YCTXpJr8NJN7asavMhHyVHQV3nP
clVlnN/MZyOGwD49j10fj9MimZ5xyBwdb3pbt6R1ahWPgRo6xdAVYhHc4/rsJqRguMego7Umjs7Y
WdEPf0Cr3RNkJnweexVvXhcZrPeW1cGUh8VWkAypy1JJaQt7zo4AKYn4/00f/3hiDZIYEOWc1Qqz
Fq9unuxCocXeo4+bD5rygeJGQ7nQyF4vJK06sd5sm+kxkhTlgnGmt2xWtNW2z1+ykGfSSsgsIFa+
wb6oxjXdDxd52cYrBxVAMf8ueRfUcozrRtma0vNPdZwSq+mRIEAeU0DBMgJbIjVtuHl7kbPN14td
n0mZSTJW2jIYzipbebi3lSs177QHCtVwz3ltimp8C0NrLQHbxxRjS+4x3kUq/r1BwdSjeQmM1OnY
ES+BMp3Oon3sTQYCOfHVKtk4X6LZOmoX7/YC2+f2/23z6Y30NYVzN+/jsqDs2xRWjKwpqLAPX/41
AkA9Xrr9z6oPw6h5l5cZ66a8KHU2LLqBqdAF2U0qxe/ywzHfisXPsMzmbZRawsXgpbiNWlHsBXBp
t9+qic+BRfww4wNWfzE2+Kx8gmOY0JGby4aN+r5vehjxN7BRtHPwX8A2gWky5JSavXQXopE1X8Av
/4lyuDqBOhtAoCu2gG49LkvFKkJbSR2JFvQZSLb4xS1ZNG47LgY09skoGS82JvPEGmwq4C41UXrx
xN8gET1sFaDTSt9Kd2Hb0TBkzJ5gySXtRTCYZxXWwXk1ILsV8uOTIotSB6ZzHeXg4x3pPA2tQysS
Lc9QBqD0ZufaUXoJ77Zct4/HTSfb12Ew83xJtTq2L/I4DsiTJtGVWK2mqACC7looitqc50L3qkDN
xVjp92OP2XhSrgc7JeANguedDPEsynpz0E0IDUi8Id4DKUYv7c9zfM9jPsyFJkRj7ghaKjTfi511
gxYwkDaEU2BdH7/LWcdfs5d5PSgjmq7weB00TTB4L8ziF6ADNyaKtzJbS7RbB8WCaWFBB4cpwP0v
rg4mS3mYo+Vl7xurfx7yuOUsb5+2DUj5ijNB0llAsZzITxexHu02i11la46TAOQqcj0EjEphX9AS
zsd+/ldejr/0SmBOvaH8i75vyly5/Xtg2Kmn6pj1Uia2DT/tRD89T4AFKCScPAcx81x44SIr4xG7
lLl0ETSOclppgQH5/OftGCckVyJlSnDDXvBo3HB2LqGN/OcJt6T5DDSG/WSvZQFsDjyivElhbAVq
WQqasevYuxctTFXerFkZwAqQSFZ9esomUF8yOjqYAUX8lvrZ+EskI/Z0Q7CNBxPVK2VYgLd4d+mV
c8DICO7haR/ECeY7TVCGtDRcwLTy5QAX7UBoRon60QQUbTjX8Y8E6vLked4w6gXfiuAEQ0MQUbmR
CLLngbsbMKXPBz88oM0Sx3vIlKcY5BbzTIPOBxCFMh9GVq1ws5E2pg9+dEMC4ltoa0MqLTG2hdBt
8BGDwllGU0YrMo65tPFEoWA++yuYh6BAsBs9nimva6XFbsCnjPSce5CLFMYm/DsQTNy8xyHL6Iv7
Qn1Z/EYMrhAOA+kPGD9WYkP1r/p/LdMhN2qaafhbp9GDVHE48zYTsPqtTZOD+3fnD14bj8fqeNFd
ye7D8gK+AXiLtK6CVY1+XNKdm3tbG6mv1t+oLzlXmyELzYe74OEmmSU16ab6ztEJzR2ywecsaimG
UtQTv1mmwqZc8+IiU25hHbXLTozyW0Du8lKUQ+Vome2sn7VkcAjz4TDChbVrRf/qB6T54of636ck
ypvYDjhTRkovylFxndmzY4UhzAwuMK0WGQdZox8vdFHgy+cFhBkWYl1WyrC4jUX2AnNBcL9vKYUU
jNpYM0PenjvZs0Ya+3a9qHRyYB22yh1yAmTT6eUos8/wgWrHZlj1VT50yCVrDCDPIA3CDuRcW1OB
O1oJmAJGmsni2xAgJvQy7cBcjBe/P94OpNDZosQKGD6/hjm23HzYPIiddUONrXDI41yDk6Rb3qqe
xr9Gie3ftpQVZW1MDGBmneTgk3144KAM5AnadqCK/4mhtY7sAyE+VjdMspg8kMVTX3hjkCgRq9h8
LQfolAfS9oqPhJBzh6MpCXzRMK/m5KL09rhqWPp2VrEwprLj7dVAPxV01qSub4c2ht7slB8xVYC+
SdUeZJjlCNm2vS67l9td1KtFnbuycha/zzR1QXUfQ0zwwChXvehD9tBSlAwAmkPCuZE6my3afMlo
4V4oTG3CI6DD6b1QAnsGU/N96vwEe1aeuDsvW7q21YZbjfB0+ZHvS0eJmOwRydZyKv86PH7+5EBl
QmcqGzWM0w7gUj6lIQNBDlZcIQRZplfZK/PXdox48PoHeEWOcCGz6cucfiSEOa5QJcc/vAr5YQZ6
wZL+dphHjpKSzC8tBj8B2+Sr+0DMzS9ImR6qadCk2kcW6fFApRUBQroDpnDnxfDRA7jIJDh+FJk5
c3CxYwTd2CMMwIVxBBvkvW5Y0X8Hs2h68eHRV8QaH75Xmd0XHnX+CTgadFbsnaMDN6tcMXZnTA63
aXCBDClIIegvF7AOXjOU3N+Fja99FQdwGjbTSr5sTsSyETp+u4FIQgZx9UARLixyKaM3Eeq4ERiO
5BtfY+v+ucMTCQLUXv/gCtX4yQhhBq9/9AbfJb4SdmKz7JYF+f8R5bOJrnuEK5GvuNL6GbeTdd75
ZWzru683Qf+YCwd/JbbQpUjvepq7PJZdaGMEFZ8/9KCXEKSWWb3yX1589ak/l+hBfJ3SvhaLBJ5Q
xPyMqzCOPP8s6Dp1fk1+bntX/roYGcsD0dYSFheN+M5Gx/+OznaudKC9M6kSOcXbuSgJSeYyVEsh
e5kr4s75GUq42g5tn1vNz1CeZn3VAWBY3dTM8c4WVT946O6NNRQTBkwHdKfN/+VwnFBNN43ZYOFE
OEOyCFBMpTkotDv19jMU1HODHnmQV198ZMO/k3CYr+nW+nplLrJ8WW4xj1j6P5aH1TQoJTkTzy06
SIZOQ18VP4rQXVTAsSOIc3VZpfoIXk5WIrb1BzC7ePPqGLVEM46NPgJfglaQxxxy0sIn7dMgXxzv
jbjk6xkH7P6mEs105ByiQ2sC8z/Kq1J29F7YPg4TvwptAJRhxg3M1oWHyL5XABfjUCLhv8w0siEo
RXIK+jh/yrEtTj33LCh7j1Nzu9zOQ9T3x3QN3BUKKy1M1d7GqzMJP4Nv1z4JRlG83jpDA0lt9mUY
2eBlXYnNyjdYAF7/ieuPTuag83UBPy3tYOlAsyJrn7kF6qk7sJAyPyG5dPz2i2RENg1lpIgqlCpp
A9vfTYthxMfY/tzyZIRQFjbDofYguhYn8r2cjABDoDyjGj8Q3jEpT1tBy/yk+5GPiybIjs0nL/lI
PuE50pXmuYTJAKskDUWRW5Y9zeWr3SfbLA1lim0chpIuiepbqLhXRjDMhlZs8LwAkRTypORYSmYE
0AeUCi1GDdUlfA7xwud6+QGNVj3Xcaophid+J/bSWEPYu4gldLnKF6bxNu+2hyQFJZiacQWsnikX
wu7TU/KQdMFgGcc9T/NhLXckEon06xmW2jTNZrqBID9lKhcwC6evflNQyoaK96XCGDplFT2Mqn75
7gdsfWmp0eJfqIA+RDHFXquqBULRIu6Z8PGM3ZVI8pwtrsi5v9KwdpSLgk+jkVsruejNWaQhVnKN
nIvs8YPXfPcCdFoQs6rdn0I5+/cExVFXREGG7+DBNfXSyQJvkJjK0tFNOq59zbbwhDvS/YuylaEK
XwXnIknxyUxIcqicOLZElX2LJbMa1n5YpihppkySRIzs2KC7kJG8LdSUSXWkEWPx2DxUBbDU2veH
tLbNYB7k1SLPyPu7XdkkK58DC7A2AfbB4xZLpvarA3VvzmrzbKnSWyPeBDZv9BeNXbDnxNa89w3F
jLB9MU7zCYyjn3zUGqwgUkvXTBS1xBdNtEiLjLOr7JmL73Wu1xHckQTEstepdsnvySbVopr2jgvI
Xg3W+/V05m3FnMCsRqDuOGwtr7CrjGK5oB0dS6lo4SSCe4RFN3yldOrhsGlPxEEmUmNdevAJDsUM
aqniXz7Tbk07WXry31XLbnyyfYnW5xD4nVHPyg+hB0ibdC/065r8vW40uisOrktBVGnd7FYR/NR8
SGMf5xSS+KIniwnkssN6b6md0yYQSYILX4E08kSn+uOuVeuRu8xDc4BrgsaSLThHlVPhtd+WX36P
WbUfT1zva2Vj9zpqYXvYuM1StYbnymiQQowCc6eFJPWwskdc5aDak1wE23CAn9k+fBUsCdERokXt
eIXKtGLUo7/XSQNm1ecNJ2tjVV456hbFzMboWQXrPLA3ZRZHDr6LoQIneI8HtkHdR1zJo97d04De
98M6BPvzpcGdeQc3ZrUipyBnpp7SWNNjzZppPeQERW0xlGGKAeZsykr/SdxR5eOPWkL6AQMVx58A
rRQqWL0n8ggCl6ZMbWWmmEYjiwajZfeQX0X6S6kIqDE+icjoiicUt+oinnU13uxHVFOurmuVOBiY
qBL9S2JlrQwOjYGR8DyPZr7qRtTWflM8c+q7CSqcUwE2fR1cyj9pixGfHS7xba7XUoly5HKV2Ne3
EKcGKZlfbyZen3pUcqiaFHbRtoHPlFpseZiJMTheOBRb7q2nEpOWkAp4ltrvtaNMX7NdIc52ztfv
Iufhlme+vfEiFXkuDLc292evfmrXeHxJ++BFl452CDR1OCteACLrS7t513H62RrMKoKi19ysQ7oo
UYrnAo4kIoEMaHod9ah63943Or0ai8a9AzRlyeB0KRO5Fw5avrnsSJZrclCxUEd3E12siDjegyVR
w6s9cUvkpZ7ko1abYngSazZZqjHLg8GjDfpNYF2pRak9QR8/M9eiefGuOgozvymLei0AWmtcAu4t
y+moQfbKT21YNmUELyYs/9L8Euah89QR6/wz6NXswXNoUqvnujqmzvVP73T2Eh7cvrVlFcrxqHvA
XpY+5mdph8tmzeyf3gOs4ya+QU4apGtLFswn7FbLO/+Onb3YBFVkPSCA9sg2txSsodaWi19l1hCE
oW3PpCNPLJ9f9IhCtY2VJYkIhTxS/6fPqiBBbbvHdpYbTwVxvGv6ItsTCHoB1S//PkVzP7AAG0nP
Z+Hz3LcJ4q7WhA6lePJHDXvGtskVp+HaH8SO4Vl1SCQiOKS8dKuiOn7sLxu21eebcSqZe0VGNXOH
q4DWBCG9QnZpkPwaicHcHnCjLiDRCNuNZFkbd1W7dFRcoUI0q7dIk9wNHMkWMOYgtj0DbeaqWeha
rRem++NfJDLgCqUWB03nZsmZI6kUHfMHMIqCZHmY41Lr4AnUJWOaNOYeRAJtQ2IoqR+oEdwb6dW2
+TzMvI4UMwuCpwIRlJ801PfvEUziafEVw+DImWEBMbPjISrkxM1wKro5fxbHX7uQWt3eUrdv7xXF
0Nv9yAtkyTf5pBuhLTZkFom+4e7w0kycD01plrjVIMyTSASf+hW+BRbB3YJennqizFwnobmIdnak
Uzs+PG0kFF1gYwgDPWijE+ZSRxunrTQUckJ2IuZuZvz9XJ/MxNG9q6Bxh2jNKIK7LXvTl/EHK5vk
P8b4sPwDDO/b6xvFzuwM0VOxbZ9Wda6OmdDu4PnpR78R8AdkbMeWd5EMuFolRdyYxu7Scskge/JI
YmBXR7Xbvyf9QktX89M6TVq3LgP+r/mMrenQ6i6Zff3u0U/i1X+BCyA0zod/3xbbNPTHq/zBM6rZ
XvZysKAqwhO6fwDd6HbpQEIr4G0ZRJ8IbBW7W3nhcIxcQ0b/ELOl6wtbzNDZciEG56CJDG9RdkBx
HRCaKOP54eWoCeY9PnmOwIb0WcL4IMGsEMqixZJw76pQg25V6cSh1Ja6DEU7UIc3yBQ2MSCBNzsA
Psd06V0ggmsKrToDuEeni9pV4WQP+jMjH5mnjV22ypofPkCFdbqNHU3gzo3zfE/In4e6+XMQ2ydx
DknPu+bKvHfdCEY2Q5JJ5++ZK+HEQXWdwroAxXrt28UPhcUvG4dXmVP1AepcOzni410HPhenWdna
EmoAK9NfL0GcHYmCrS9ZfRRsCBt7I2WGyRCpiqQovPmsRmynunS1ryyUqOXYtq0YEI/slKXFwqm5
RwPNFf7f/EOLaAldqyA3fDPIq0pBoPMuYfID+TejB1ztTCqUI6cyCgO82FlsR85X6nifQy+tiImI
wVqHf3LhPAOmS6yhMgPMsA7ic6uKOZFrgnULiyNv6q4YHgLg4WjJ/Wyc7U/Qx/he06AFtUNxiOFl
F3o8hktWgIM+Gw9oN14Ro9aIWXrI02lPEgJ2fhwCK3Sg7WOaDuLdU7C2d40YFCpfWic2uC4D917k
zd6y5RZCcCF59xpfW27G79OoMatelbr8UBGxgvTmYB6LGi5eMjru6QPNVDrehOJHCatjozksglax
utZ+p9Jon6jW869MibZzAllXjlUr4H9UmMpJp7AH3vcysD5f5lGnldVphHbc+yvwfyWjGMyE2gOF
ArivWbuvyWsqHcGdvpi4ggomi1OYpknc2wySSmX0uhX3tKg0KfUgacyCXKESJdkBW0KMInBavtEN
f8axis3z6MBSuKC+2uKJIdxyvdCbNmu9h9TqhYNyMeUVY4bMiHQOeDjrKjCu0biC3tIbpkxcmkXq
shl7JUpOpguEfkS+lVT6n6D+E/oKRIPr/YhWrYbH+ejA95uDhE+QbR6ovHC6iI5uSnSWGA9gWAHV
oKF3DY5edSXq8l7MaevOt5VKrvAAz+a/v8FtQk4YV857krVE5HMJbZMz9/r4nfP+u4heg67fp6OG
boMJJbDZzNPrLsBVNmJKw4JFRDFE/t1pQ4a7odY4CSFHkAmGKrQoRzQmhYyrariT3E3uT4JB/Tmw
wiaDpWq8pOhXoueRMvpKGYY3ldGMB7tXRPIZGK2oljZ29diJ2BoQolrWpBJsI2y5+v6O8GoLKyQS
hUmqhgeNGq6JUy4RMOmnnWpVQnD1YGwKdjN/Kclo2s8sGDHX7NIohdGgBOu3MX3jsrr0vdUGEbny
akm7BkBnl0hwLg0nvXy3LXsxNRrwR1qRtk0HjaZRPrMRLmVCyol2PrxR/du2/9fkWBNfGQ0oHnAu
YC11ACX8kCzSfFj9h+f60iSK68UC9kuEeOL8UNn4xkiNy++VuzYz/Rbbetq7bVKC20fCjuc+JkJg
E4fD+GJNcN9qftT3KDvB8an+o9D/+3vpn3fFUgPCUx7hWmOV7gpQ9MQ7BUgJA4+Tk0bmicIgNDi2
+mrsHiOPoTCWdBFr1ctSP5jtrqnhF3SvRa/oRsMlb441xvLWomxvDoxpb1fC2Bc/xk+QpMpy3Dp3
R3AzlNGEcAKJrQp/7zrdS4zfeGBhQhnwZubncTX38f4z6sOBGOHPY7u7SygLWy002DR5bxRnbYgR
OZDS8pHs+g/OkItZegBV3jcn5ThWig0xzWw/V4xsW2hRxUhFfXh0y9p49f9PKmFb7iMsZeoVP2Xk
r73Nj0kn8jwBt1/HuHZjWIHensSptvpjT2h90aBoX61jANAHZ9xpaINowoz/ZFXk7jMEycUSuizU
PqghnvDdW+8ixexNql6l00hMDuxmfzQ12o3A83NghvcslnpkYfQ/RMc6TSt65vwtMNpHWL8UlWFI
sFgKDthtx7uqktMB/bgFq2P9F70+VpSffaQzxlqb8+CY+Skb4yFz1VR912ChuW/OqxNI4Y9c7vox
uP3SPcZ9040iR0EY6Kc9kNufA4Q90gPUUudJ6hyiX/XLpYzMqjirm2lTuAw6e2vvI+Xsm1r6Q8fG
ThFtC/vWCNLxFym0NwX5i+tEwDP7PLJpyNeQhFNGG3G3/wvowMCot5vncTb8IWV+EJUfXrdaj9C5
Zj1DXjaJCR6wnYyq14fBCE38K5JgoQsiSbM4yP64V4K3i2Dod8k9XP417mBNmNAG5ZknAjocUARr
F1qhTG1QcTnTHIvgGv3QRmh0KYjYDmWIZjTzQmcG+sxvkB1nTc0CgF5zYEf4tYFh9ATPdr+T/PKz
Z+t5TY05BHwOYdcWd8w4VfUzn6rSYOiX+Ggib9zcIcLGFF+whKoBdLNd2R2lPViI8+2sPdreG6v2
q4B6Wd7HkNvPLAJyqgj5z5SQfXykThy8DhF0vrg/zCr8ONT/tlGKUUJs8uqwwV0dfHqsOjdGTL55
xPaEoU7IQ/msLh5qMV4HmQIWs1j2JZu5WN3KLE2i/AGEVdO1KpQJj4aYqviMFj3jw5X39WeIfwsU
UK1+ZSprJVwIWeseHfsnS1W6rHArKzcpi0VTJA728Geldq2+U7FU/zfxnuplKaQZ2P9/HkXVXpEj
VO2xiGdA4aqrmk8ZWbWPuA73k60szxlYFbJGCRn0DF/PUN9VHqP2KzF+mT0QuWzKFxg125bkYGPD
AV7X+Qo8eyQT9YOG9D9CLxuxb+qpuSE9TgWAY3kfRTPZGKVoWSGaZHXK4CEAj9Kj+F6ID3B6TxQd
O0uh37bI2u+S+n1+7K8ppJWkjuhWw3b9ebwUDuXyRhWFv3icI1mQMid6wPZ6T+Tr3tiSeR4DO5Kr
6BAunHWIXlru5N2MipYi9ayPps2RaizZ5mNU0Wu6FuG3ktVJoSoGs1c7hQ9QTDKvmXnOhqzRtDkC
zARmljpmwojxQ1y3vQEibur8TAVw1hYJAo7hof9QmwMNqN1WiLtFO0kpSSoHVTyqu3wrL6jDRZpg
KR8XQ3hbQ45CnEQgIhFv+m0ZSQBC0g/lAMOUuKZwppGGbMc8ZgG4fOWdlHIKLJ1kCvzi4bTw65Pz
lFbm8cJjzTQazg4im0HpTPGj3xBNEz6rPp+yJsn7rvPyvvoh9N9bTjmEMBhlzFa6BLUmNU5RcYnI
qoTxwoGwgoTshXhliA9nq9U01dF440sxM99xMAc+7kntJGgY2ctFdIagDORHoE/ida7wEKoqMPK8
qlkWkQxXmSa05T7M/asOCKoJNZQcNbyh4PAXt/yjmY8NEF1kJPWt2PWgYHzDRs7LiQQNJT4+hytS
bLRihBIukTjrCcXxmdacmQ5y1hVXXyzOstu4LQN3nNYh+tg1JngeLd/MwwMPzZBF8/Kkq/KcIK7V
RAp2cfe1QstQ15NImR9gafnb/zC5qkkX1Z6GAtLLe9rW7YwLBbiF+WW01foheFhVdM8ujV2BZ2/v
jSrBDdZ/d7aUXHqFnOj4sh1Qi7TJ7hKlcLDpJfFLDscjR/D+5FNTQxsEpz1/bLPOyyYAcNDyuJJJ
G9OJwAJ7VbMz+ydCYqnCH8lHcM/dMmywPSKlfkdoBDkgG9MTRuVkR4D0NgJ5kmhPXxxCKiP/WNXe
hIy0Yi4c3r2Fp7KsnNkx1H7FTLcfdHRCM4Jo11etPwEAeexAiuzwco8pRTWtiggVE5PMTBXa6cRj
HMON4cjWNGsK7l7XQnUWjpB1yU0aLWTcpeORDHe5NpHfq3oAoAwhUjYyumkbtWFyLcWhYFVjXt9k
iWn+7GBRonSnwNZtDrXbkcndz6xtKajLutMv+TBs52qa3HgDxD6VnaUZWNhY0Uhuje1AMmEJAaSK
+2t0XlaBgkyxYXsbHmDT9a4cCEMfvKVoyjJnJR/oK0qH2+rzh9gDEexMTjkVRjYRSqaT17PfnHJS
5ZpnwlZeQlB4KZwXLBUBHKrWeuVK41D7D4PCDeF991+ecZRpdRNCgTPguoAOyqSqgSaE9jGL/mfd
efmJL6tAj8io+Q66+rIQbXXQ8zcz8I7GtGnFLhBB3MADDC4ovx2YxFWX6rvOjdDTHB6AqF7Z+Vns
ZC5+vBo8euZX7EuMRcpOaipWeWqRsIESrX/9kcfF8goXIS32FI4NNXHFpHi/4SLzzs2g9fAGQqpz
xvWxeYSbvl+p0DTz6uDk5cNhfrdN0GwX+5rgE4TY/wjnq53Mic/RjXANhfKuxIpPmDVTFSJX1rNG
ArQ0dedWi36QeFcroBlAsafi+uqWYdzCUnfcNCdTx8LTJk5RD9/U0GuuQTXfmG6B+1mtH/Aq74Wf
5WhY9y7EnPkORrWQz1kMDtcgr5T8PmYyWlrK88FYgBC3q8aY1SYWdwmjv1YGFMShqEKNy1JQDHQF
z7eCqoixauYNGvz+xBe5joHao9u/HhJkYtkNgjaijfAxua/PI9D4Ct5vIcK741l7xowCcb2jY0KQ
wxwW5ljP/S+y1F4EW/gCduTtIof0/ZIBcXtyLuim3VxnwwLfI4lBYmyve6byG2XQ35/HL5+eoCmx
o1Xa4mjI6Jg3PEBAU1ZPhqtnrdQ7gV8fdf3IYQG7mKMhX3BXA27HG8BXaRKPgu1wFqtWrEFGimha
/bNbQZAex6rX94nstFv6MVWUBupaHRHrWLCSJ3cm0ZeH4hGDBv6LeZkbP/RpvjcSyrqxpbCF0j8b
nU+eliXfxIJBGxRKXODTWrFi8ywQol4aaetiXbpUOy9prn6PlHbrJxu7FFSaKJBfz+YDeJM9qvzf
aFDWzxA6Z3IW6B+NrdOlerhHnXKarfEATGhmEwBgK5kiqOITjbkfoCYug5ItSaCIMfp3TbGfzQbO
4sMjxzNBHKICrQ2vJl6LiC68tJmzJnVhD20hMB/hunHmPM767bzXI0EgtfgA1opVbq7vwWQ/C6tA
eBLR2uEND/R1MUa7pl66WrnwGA9iJanxpmTipLTIvplnccOgFjjQShzHiJkM9Uh3DbUE5kaEOhal
5Yi59ft1ArPSdkhf74TOAxD2h3fdSWfPc0uxkR+rHcXKzEdI4ljW5DgUuW4ktfS2OlGfpezmQXDq
fp68s+tsa+uyTSc8RuzoaFmeiaG8ZtBTJaKqIFOebSuh4G5ovZkpDQtj0gG23dw5GRD0B98uUP2I
MjEOybXComF4+q+h3dpzj2xd56VDhH0oJxE7l9KCCEFm3P3M2v9RA0emEruQmlFQ/mkbvvYKBd1z
ml2fVQwByCkUwSPBd0irpF9SSOED6wuiAoIeN4fs9J6HxnxpsuDSlCSmUc8NGHrSFf+OD0/jnXhY
yr7qgGNGgyKA4usQnHm8T3Hj8nr1LeW3UI84NgB66WBdYyfwJTU6T/qQgVAyV2zyqMUF4grfzry8
8Z+QraVbrBHF/p56XXlXx6nT3ATiuCWv2ox9UL7kZN1TIgNqtKhRIFJk7/3Uz3XqMVQYyTWxgCo6
pNj1frfgoGrO2nQDmAcMJUJ0FIenhbsXgEk20ZsjBR95tMeOo7RUedGsDpJq6OBLXoHvWG8GDaxS
IbpywZeOnbnyWtu/eL9UZN3VkWRr3zRKFKRKTsYiUCtaXVHP44IfoGWk4+5vVCyKaVS5i7t/yNFK
ZXcFLjJKOQdDIWcySF+vSg2eMkotUn6366XxwTaZc/ABYQsx96aip3F9zv+0m2XfNKbAvGhXgkBb
GfRA1OgEv1xgVg3MsuXN1NPSJJiSALm8+W6lywYrrFQEGuaVj1Xt3r9znJzSf0CUA883+PW0r7hf
NBUw1/OYFELrteZNnZk3TxRWjPfRWZ/A45wsB2p9yzHWFcDUyRH/RT3fZTKgiLr1NbdZE4iQpGAI
2qsrDdzhnAKQcEbFfDRPqD2EZHCWvHG8p7yF4aw3KIci0xOy3RlhkkobLay9qfDYxU9KZ0KvW8+x
jeqQK5x+83OQqP5JeaevDj/sFeXlrPU87LhlLtme8EwPgV+S4ChS+DqHa1YUq1F79Wb62BdqVdCd
m/1XZjYy+PDV1BMoROm0QZZF6GJYhbAzOYbjLBVmdA+egfnjt1rHPRfKGxGibEeHokkm5uO7BbwM
R7rPT+auXv0NLlAR4zR/9B3J/TRIGLTWoDGVDviOx2uBUVw43TJ9cTQuJALRvv5sC9RffVbFcmqj
HzleSwjqScVphFoDhfuuyixIoNk8g1o53jcQkwRqtPT8GhvFAdEm3ccDfK+2vD2ITSQTRkda0rcz
devdrf3WCIGGXd7aXDCzal1BJdqWh1mso+h+pdjJrH3iZndzJkqEyCJ5E/oXWfmvbyKWA8WvJrPU
SRbeJLeg0uGECrZ2lUYa6dsoLMGEFP0j4PFM245j6Vondug9lzpiIBB4TPPBVcF2cVq4+YrpHIXH
Br6VsjkDGU5+Mp+kTSdK1PB9ggVucxN83jXjUmzGF8Jk2YDE9ndvn6OVdUq6Hk/iApyxE9gDCNVR
Yd7vqzT68b6k45tyGBmPwi4Izh2j1K1s5TngB1HlQGeah0aa9GZWCGSi0KX1Ewyj2ChSqV9EHuLi
gI5TesFfK4XK95ndl+Iij6/yCjnmXgaYwK5MXayR+7+klwu+3rvEV0SuJVmU5JAJvsSrwvjsKcTF
GmIf8fhNhJ8cABdSmYjFtDta6kHLllubDdZM/FPjJeDLwgyovZvAnRzO59actFg4LpUtjcnlNujU
QnptpJagx2uJfO00TmJea6oYDKVxmEvx1INlAWF/EAGP0U/slHDCWcdPykHrm4qCsw185GYvZv0s
Dh6VSbNW5/FIBE6awz1r6D5IFFQD+285xtx7vNoo46NZ4HsecNd+yIfCIcWFfjKDallFYiu8wxJF
Hgc67hihZoePmF08wIt7ARcIlqdTq8yYw3muZgyBuwEVX+7rjaB86xFvDNTwYBx+cjjtsYRV9/lq
5TTm0CMiF6zQvZsx8ulDHVubqrEBpvEYd22beVU48n0gup6HVrLduXGyhYpx2FLaLbpDO/n0VDgW
tRpjb3Hqe3VpzOJMeF6rSVOP6UJjhUcG2Zqy6Y5/3+motNA2T5+84MBFA9zwWQpnvCrIJntduP0b
qORkUfltS2R6Kkx0x+EOcY3vw9YTGz6kUwtCXURysgVqytyYAdZd0GFrTqz2NF5fG1cGVXjxWM6V
XauxMArypWmEvHbGu6I/Iyaq9D17BpckRiPRba3f89GpB9oVH5q24swJHf/6fszM95v9EsP9Gafc
AnxRfl3zLyz5yHjJOV298uMkms64Fom1L2IAU39qh570bLvjsQymaK58+0wp1fXgw02BPl+y4CcS
3sSRmjjJiQp+Z53uqVQpU7kt8V1sa8i+W5Jc6W8tQterh/2kRYFV1/iVuMRWxVCpagTw75dWWJ82
p48nX5kW6vaSQkphVRBEjlKz1dc4C3tls2gCVHz2bXMMf/DEoEphBzHrWxmsYfIA3+xntUuv2Iww
CG7hC+aYtGXuiTuWGIPp6m4VeanXnLeA8D/qrt2vr5I+hH+S7GKvLQ25iZXl+cjuHMrteT6mGJYh
aqfo98B+zI3jnzTYg1mDWDstA/WpprCCxiBo4sacA5TCdvlzZX0PEFz8Z5tScfTRjslQ0nnGfInY
qlR52BsrYArWGKJldCuga6GazBzzPYKYAOemCxKzUoIGhwAuNf+ELGJPNWAQ/eFREHUK75m3iAWX
CNK3lRizob1z0nAxTwogo/oXASaGeTPGJsf+hCKV2NsrkxkyRCQ3VY/M9vFL3+jUppDXzIghwKLD
PlcTAHst0c0m5tS16zQ/QbuL9fZmO2d6cbiVDiiXuQDjzI1NGk0/Xo3o0bCUFZdera4HlPBaMYZh
oLfOmIFTTNoOJAV/RxrtSMabbxfmHRO0u7Sddz37Mu6EvB8DCUHACMffCeU6IISOjWO1tY3enNhI
8AkC4LnP8MCTBTJF5MB/5vtwmpyouOfQYTIhAeh+i0huFGXUIGQPNOGLZKRgmVEkxnhQeEjhc1sV
ZlURYnkAtVlLSqbDwYK2xTy5yvENDcQaklNUrzv+q13ioiSlYZweU5RQ5vCiISW8GqqVFXVeiJXz
J8iyeHxc+VRyiKZWsjg/8J7voyMD7NDsgU5NUp+zZlbHXlxuhdtIb6Xx2z+tGkMRzth29hR7HPfn
ufI8JdUnR+c1qMI/zuslcqewMLP9U3tb3h0FMhojfWDJ4t3RG2zWQhpgrgy1IqRzfR08+xhjV/Me
8FTHJk6PYkCYENJ0DdtimlhUHyzP6cteLRP58bR7HqV0Re18hhE/QshqA0WBsNyJNkUHdfwVITIX
CTFfRNFufiaV89xFqX5pwPJkEXGRmliE8kJV2ffGN2kvTIHkQPTMGluZA3ywjz8bFj0eYH1kSq0F
vUQACLs2h/pNAnuSGX2VWNByfvx5OFpQ5JZtQA7uK3AOf5h+U/pTgrPtC7UpciPVpe1ZCCEqnWGW
Vy4saB4n5eft91pH8biaelKbQyKNerkQR78ydmCXd27xULg8hixLwzsWdMUnYInUEjEQ84JMmfuI
rTiWVVPRjdgjVony++CrpZweUDWelWeI82ka3m5cYoN8ZFfppjymVAsDeL+mF0kh1rQI5OovVENn
s5LyPHkDE8fJB2UQMm2ILYPDmn7kYUJiUj9p0UXhmTfCQBJI197rcZUILM2vNLgJ3C7mSbyC4t/W
+sA7T4CBVHOStN+PXMK2M6zXUzSrgcUPs1kV3Cyu23DQNRmpF9AcM0oV+P8cK7D703uzeg0criUa
Xa/fT3e6O4bY8u/1U7HXoFAG0DWwFRYYF4Cmq09tfxbWfx0sYgMBF7Zuw2r93HbCnj6FJitl0GAS
vj25obyvm7jkxK0vsKsnvnIjSgJi4TtITKVods2BeeY7mE0HDNqC6dnm/VW4J0BzYHHH1fThvr/S
DKzGa3Zvlp5B0BXIJcM6Y5qQYQbvyJdWiDxvvwKHzG5ONNq7Sri3Qk8Bqu5Yf6O0DJHVWzDCD6uZ
w/1ZQ2Ai2no7QAWeoTkcB3ACe0DfKJOS3zwgjsNzhN7ww4r7WSMMJ9/wWmS4aWJZictAEaTHjNSV
+m3zxvoXEu8C4OmMAq5XBdQsLT9ZBA3gZThqHTE4UUM2mY9Uvg9NfZ5Q+8DPsIKNk114bxZ18r5L
uYOBO6XmiBEwVarMAO0uxEl2Lz0ojWjzJrnpWvdUTa/iSUPVTGsoqUahJLqOr5ImlR34CbD0sPGr
w733sUoTYDYockIMpGQ66l0u/O3zB18pyanvJQgU5QRn1GsUdjRREpx+PYDmFlHrqyl/6pIQybAn
akrb+N5SKIaoQAlbiOrAZOCWpFVFogfprwS9WXCA25pnRNz5wlvrFFMJ/m/+2cAlbHebvoNiz5TR
z5qThV40d4KEkmCn/F26wEbElxQsUm0dBlb84vgRn4Cpaxwliivbh9xLHsGq5f1UNLi/H5MmI683
3jbC+akMPKHkLsJPckd5eqKAIwk9guntrf7p6OJr2RRfymTj3r1N7Xp8PBj+sIU5knSLYwZdCpAm
X1pkKfXezLmkmPy2ggH6aZITTYAJvMnrUEd6LwvxKWNCdp/xCB+Wf7bUS6ix4IIWcwbjJVMC/Dsn
HyJMt2ks785kROiIgbzyvj7S/2wZ2HD0sdxT7PRrsBb4IsphZmr5nquGKMqnJbHkuggXG/g8TZep
dHSQ1anH7GJHjLXZtwfAlKy2vrSUbbcZylKki9Xmf9DNcJuzr2E5r5PMqMves+lZe235+lJkiY0V
zMRgZ7DHoEaf63nvLFsuwk1uaX6a5JZsMIZT2xzBHtWKiOZ43EBOg4Amtt+KqkkDs+KnvAFmfklA
j/hCfn9aPWq95alkt+5jUgB8litRstcYUgFUG+0i3V3FLZ6ZfvpCc0MbRo1Mi51W9y7f///oT1lq
rRX5b0iaBnLQs+/ZprEyiOD24o+IBquZZMJ+UvzIXU7ECOKyMCX4NLGDOMdBB4WZZZRQoMzNy09d
8/ZegIPFbfGTkWHy9hvil46RWiW2FtRiBHp9evcxrLBhtGIrGjjuU7YoR1Ep8J45WmNAzNz+REGr
ySPNgqdapiy1jzuAFBRNZJqrGsEXxudo8i2VMe5LOVCPeToPZ0e65Sp1bKZC9VbNmId5kqu3dlFi
PJy9POypOUDIyB4HA3nQw+45S6b6T7jfYEo2yQ1fxPtNO8tGccX+9qm4A+rzbr5BVNXFeCzaH0QG
aWXwFRz1OIzi59Wy1MiP4mFbM0omY5gLnBf1pnES8zUeUtiu4uGyVG9BR66CelfTBnz3uApkkjWG
V2Nn/ZDdMBwTgaCPRa2h5sDe9KaKpqnfEoi3zRAYeYZsjkgGiRshIyMqGpNGtrUrBWPdmAQMZNm0
08etcty+qY0WPEB6zB/SmVtMqtgfneQECLKG1UZtphKFdpstbVbRX3GAdQzPGdMN6/1evJsX3lov
7NDelh7+3l+cYExi+QuWuU+xl6JdxPKV1hN7th/zFps7YCe+j3qDcaIRVJssaKbZHjB15bnaMgc1
oAKvJpd0G7d+M38otBT7C2BSaXXuanMOsH1ihAMShtw7mqMsMS93AUxTSnv8er59/7nfHtDhWr+T
Fr5teaoUA5SZNWLLG4lSzO+z+zsIt46V9wxNeKzz4D86fDlNtifl0Jz1vq2IYpSoO8W1q1x48ERf
F2tEovf1UknK2ARB1RBTBfDgmWCy2TybSsCMCT7JCteTZpsbf0IBBh3dEOVxvo+bVmEK9FUuQvhO
eXj9t4nMPhfMlkDP16lc+MtE3EWw8j6TdRY5ipx5ukXm8uoM7iYuZe1JRJn7W2BJaZVRwABRToKS
ldBjFjlW58wVr7lsYEPv2zP7ARA37zrBmP8LbfDXifbLrxb278fjYtdUdvYjS/ktyXIEhnumwBDu
OeCrfpLQi6ZLUXIbqE7FXcWNAoJvTJp7R0XhOf2fZUYtBguGPgHwYsEAj6lf8jWwpckg5EidLaJB
HmdMXlYZjEPhTodb6vXiMo4DmRDSVVjRGlfeXg3JZxQWgexPVKhz4jZyLDc5fwktr2wrktkvXLmc
b85XpKTx4hMzS++B9CFFYv9D/dpzHNSZh444jsIUBKUcf0IYSLm8ww5rYjMynalWwJfxfkLm+rYY
M89t8t2FPVlQyTJ7ko7xmRBVBdZzlE2DAgONnXYNr590XgjyLDXiRyAjxW4T3s9qV+njSfqRUk6q
/yWOICOqDV7fryHqrmfk6nLD4aDd3GN6tIsVjApwdAc8/Ib9mo+rr2pQXQ7mjcbY+f+qky5HWRye
bqJcu8fJhwdPc+c/RHJcaL1a5XZo/yjEJIJ5kIsYjj693gFsrnh9qlF6pUcgCs1Cei8uWHFP8blO
Uj8vqbdZHMbla9tvFNRdbJ8SphReWau5YPR7yhLel+pzm/zTueqZlLT4PSCDckTJVR11Bo7HuxJF
aNxJkWEYZti846ivMppAw8OpqLB74uHet1/Ds8cQHbztWMh+BOXT1Kv5nc94Ptad/aYhiJK3s2Dp
uCXtESkmI9aSkQPrt3fo2yOODsDyD5FUEOJG2Kt7MkqzRHU8Cwhh9QgihEeGwuPUCxUaV8YzcJFo
blzvaXpe4QCrSQmz8qJKJA1yjM3eJ3/cYFhnm+gRAHqtcX0kZ2SyM0JfgWn+tF+f+Jvm9wI+8alj
z0NC1TL3NMZTURZeK5MNtRLINuWuh7T+H5uzZ7/NJXx6sUB1DNaOu50dGpnzu1RFErQF1BPEYD/r
dObjhoWN0Nx0S7q2BhpuZEHgJWJL2nviH/XJKahInmWjoC7t3w7XzhgcFSv9D79W8X+FX4o4AhsM
t3vb8ynh8UVkwsbSjmmekFAlK1Cg91AE4ymIH4KPJOoZH4b7Hl9v3HYCdhy8C4oKKJKNiKUa65b+
CQmHU50H5IZiv5VXV/VeMWyD339ilch38s7ygKnmk0NvyC8YGlMFmYoneuXB80JbVlNtfr+QzVAr
38S7yEIETJryzdRdGhbsM8YQ81VSQQanPkMH3pih7Zye+VyJ2NvucT5IuafXpdhBzdUhI2tJ5U8g
ydlTFjkmMW/39CycOSr0lFrKrNzmy1r9z/bKn339mTZO/4A72C1FcPRwkMBojfqVJWQm2pMyPbsh
rTEedaY6jBb6GBhA5p5u7YGR+knvR5AawINaa2BkFgSKTNPfm2hQga2qIV5ahg05H6qjqjmEHBpY
rL6XA2D7XLt6Q0xMC71QgM90sex8j3RrWPgMk8aJZarCKVQL8Lihw7RJXDTeA2wI9ZtMwQRjiJXf
h2Pb38OjwX3kwqlAitl1YBGhSwwZIR36hThxmk8iyZ4ONABQlYY5b43lVyOCaMA+P/daqlGAiqQl
xgaHA6QR3Aw/dSr3P6WIEDC+81KF4w6fZaVr8gIfVsdAse40RnNvJ7qoiX+xi8VK1ApWnIntQ2so
5kai5kbV+8q8LRg6HlrLt3KxEi2VC8EuSboMwP2io7aD+DhqX4i4QQj5BMTHi5SH2zkya8qImTvd
K+aI9pLtzOF66svnYUVULduu3zYR2VVb18loN11MFDhHrR/0mzVD5SyOSoTGnvUv1POKzUfKi0LC
glbuUUlEy9dQo+4Z9SBxLDiU+VNqZgvdk8PqqupWxEd9rC/TRFGM2BBncISftYSBnqWajzetyMMV
IKkVkL5m03Yp+a1rtvh0PzU7JFTclfnfymZVV/TzQUucyOz1u/d/ryK6hYdDUczUFGirJcdbKTqR
QOafTnCUlBqiMkx7+xiIzFg8XfYdoaCwY2BODM8/m2lDH91fDYsVii463FNOppL4chhQF42qAGIF
VO4aajfCPyxgJZbk9m01+Blefl01njrVvOMyx7LhGmaBmokjNzOK+F6RFU7i1dITBpzO5ZX5n9nm
wbN6kzwgGKQLnCSsNf085BqT+Kn/LQyFRYRRqhvghJ4TRyIsj6TJiNmBvAfFPMpRb69vVCAkyx4m
IQRyOvw/xKttaAzYVEybfBk5H4OjdVrfZl6PVMx6qWIfE74Z85dk4IPAPoXXtUvZZFXwKS6bLpsU
2Dc6a18SN/zK9OXFqxPyrBENdvvprr6vWqZhs9k4vc5zB3PhQSsC7SAEFJVaLuq0UPs1YspqABKD
XtB81mopGegOiKNniOgsuzQOi7FNx8c/Ea6+9cPJlUbAp85tKldqBrB+v7qgkumJOLYzMg0oFUQi
NbNEQiNkJ0OCrpTBwLgPebfsuVfBKL5QDc2qEviDXivHjBICvmSkQDwdYk5lOSbmcAaj2G9omT6H
mAiHMQT2KZVJse+H8Fz0WffMIApDtRkCRQHUJ8i5rdHlrKBeXWqnwES+eGcamJNPg85ttgNcJRWz
dCVIwVFk+4iV2xpMu842Ug5TAZs4N/lDTMl9Mb0WAOzjMZHA8ZrKgW7/Vu9BKDm7CSeuYyWMKwQB
r9VTyvGDcZOgLUApXm0QLB9hMYn5GD5J72teMfMu6hkpsEfPYMvfbpHt9rFv5KMIGxNMx6g9NRNk
QUnj3AARvntnhJaPjXkczIWwQ+HOc+tkOJYLBAsTa1k0F0jhTVQpfWfoiQc4BVoVdQWg6hDaz61Z
PTSIUAj47ufY+VjZKgHV9A+0e46/BQHldjn7+E+253Kxg+PEkLs6hZw7Q2pEx6oSCWmHgh3a2Z3n
Ci0Bjk3ENB/X2goQcspjomPondXnxZGs2iIi3vhZXA1YDKizqJQNAfAW8PnOBE9iBYdIDZoeY+iT
e81Hkvyh5ke4sK2dBEc+hOuIMxnVqwpKOfPyA9FHk3cWbRqLPwU9keIjjmaqB9w8xlT2V2Db7EFd
REP4C8uMLlof+5yvqVfpsBrarKxhkDvExAVVLhVVez3U5quzckgDi2QIw+tnYI0QfOPanjjXXidY
csnu/WmRjFdxEGWKeL4bm7p0kiJAbn+HAba9urhAGcV1oBVNPE85LSkhmSncvTkdfh+huosIhFDS
gOh8KL2vF0vp/hQx6lDfphpK0JB/K92YDFSo9DdseHxul6TzJI4JW98xNaX3U0ZdauofWi2tX6Rl
KSp0X5b/H4FJCHIt+eef2pkUh3cb4hKUlaAh6XYCwIsCezUBMFabE6XTwCr5Tk1s0v/kD/NfZveF
j5mS8sEjHj3lkOkhLfuaVWRxnTC/5UK8f4ngcqsjBKnrEUK/jeaemR2h8MGCFCY/Iugm4w3FzdnH
VDdDryRE1tb9Sro36VvIH1PucUarqWBE0Wxl96dirUSaqcY0Ig4DOLBEkdk2eA5Q2xjqPAFSLt3B
+Hx7G1mwfiDBaLK/QyNrH91QP+Yn4YYJmIQ7plmff+SPoBeutqi7In3d2Y9VP0q74vOB2EZ6SrgG
mwwbl/4KJlAWOjV/uTcUSWDBEfWhM3winMDRtRx9PXjLf5ra+bsO0Px828ZdiV9/bTWfj7xPC5j2
10VQI95swMug/KwNZqmB6EQQuChyjvAp8xnkgH5fF1luDKxhXiU3Ix7plwzkkHgaLQYRWU0108KV
3e4pS3X/5tqaMCpzMqHkg3PhbqqPcv3ZI8+Xxb+QymoL2Flh9f59+XTaR7hCRCyGiCcwSsX1IcGL
K/cCjHpLr1p0Oh/bZTlbtElyezaZmuxhwSl7SgDdVBDLE8ERVE4ni1Z2Y1r96/Ik+1v8XbNqdDbq
kIhdozL6wE5CUb3gQjn1eqAjhM8aQn9qca5SfoT5onh9GiOtz/jl9OZ6lcdG7WBx/imhXM4Q3gqA
8u/HGZlT1tvodpqp19oMZQzTB6KLuIg8yapiK6qrjPgjRLkUvZpHjrnn9sQ+sk2a5py2PG5sxRL6
5wJAo5ym2VPXxSIdkaI3sqUOFoEI03oEYZoIyTZZGGeB6eSa/1Jktilz8KEWGsIYq4azy4E9ZXaX
zWN8mG30AXe1wO5y6vvBiQd+2o2GTue2MBkZ0mJhlgX2xKKNJclnUtBhsJ8kcD3hQB+wW7FyOPtx
C+L+ebz8RelyFIHh0Shh8GuGWhe74NMxNa0zDBp40ppewo7J7B051IEvRvSBSlYy646IcceRx5IT
SFMYszy3N3zpHA0Ik622hdOdrMPP2yiBAiQHbqueJwzsG4JQ6W9bDI4jUuz1dmgImA+XZTfJWPdK
MJYLweOMfvwRQJJLbsK8qaqKHuDpLn7ESEy1gbuWXNeA/hjTTNZEjxD2qRBneTd1qp7ICV+fIrK9
xWS4xDsf138Bm0kaeh7F3BCpH3CeHqU2IaVE5Ck52gygQdp4d6dPPcjfF0Ng0wyI2yHUqOwPedzn
J6utTWtluvfcaLwYY4n9bOXqPACHspf5eZDFOWihpZX9bvTEOM7PxieEjbpG/1lNlNZRVWlKVi+6
NUkiZO3G6DAnWm0FR/Gl6HOvqsvZXqODD8JARBrv1Su9M240ubi4LKG/RR3R+T2oTSbaVf+ypDSp
NeMkKdrDGk7+61c6q+CphIaND99nEI8jGydAhaaVuV1Au2Qojj/+N5sU7ec4cclDjpgvLk4aShc/
B+zEYG2cVLSBibqIK6zvRyrKmJRsWYAsoxX6kl6vtzQH/WyFs386W+tUktFXgh7IWJ+LX/UjnKdQ
crDN0FcoONeDzTxu4dDwK5zad/f0u2muo2xpddy83PYM6Z5+2u+lUc/XgXVTqKd7D2p2xQWeCkbW
zx5cnt/dtgtyxryZMT1oQ1dOYwCy6lCYrTRbYmJLLBzny6X+7zxtu/+XfeXEksWW7S56bfm5aWYR
JCRRTfGfUUuxQ3OlbAEGEWEM+3txOZ7u11V+RAQRLi3NyGsCgisb2oQ0kW52OvEdci6Zs5ZzjxRV
Rhwd6dJyJyIUBeMli0zh7+q+fKqUI4ZSRs2wZNjgo9k7pSlHvCPFIiiBuT+1Th+bq6kqqGdefKDv
jzRuT+xOk4UJde9wDy1mhIAU6HOMnPxdzLpzKZgG9IEyb6/zjsoxY9YTE9lVRfvrJnVTaBKW9vHt
n3cTOYhZw4njik0zoaUkXmFCI1HFX7hi7D36tdSMWP7s+sBO8sUJTwgHY3diviF46Q2N8xz5ZkZL
Q1soJXacwttPdupipvQrjJ3SYRnN3bque6/Hjk9gA0o9buLrQlFE5UD9zs+1b24Dx/zCs2bRowXD
buCyvmC+KVDnHxhNFo5PBu9vVw82tMf7OXpZeMLtCzb2pqQE7Q1V1qqKBFAlZosjOBSpdHSUvUAV
+AaEInn8dJNnDNK2OGbI9aZncAGURjjLtwiYUVitrjwHgzXnGauq5Fh0+AHBZ3I/gb6B/7CI14uk
kCOFEJofXYedg6yAPZQCTXc2e+cdQ8WjY9gsfjTkOohl734cZAFnehyr4l5tIo103JYT1GvQT26M
XDdw9Er38jZ1kDUKOt2DHbBSfO9jfrAszBdsMQ9zWMUIRKWNpgc2xTF/JJ5gAfy9uATCm8psW5uP
jYyQCuf9QPw4f4un3cao2ZQAq2yg6tcMtcePn7DeSK/FeX5SzIRKdYdvaIMohvy9D/cosIHi4ue0
2drE9pHaGc7D/xvXTc7dSGZf9ByJ2U+rDUDbvXVYIYkJjAzsBwv9ZYc5WLAasyiWr1tzuAWPTU/c
BvAjrUa2zdl0soZmocMSoJKm89G2qRXk7jKq+oUpX48lQYYRudCrtUm9jQDVCpWNUYXgGvtTAipL
FQ3ltnCiodCLVd5LdgUV6zDt3rdTg6P0trmgZlr826vJUnACfWZcvLDDN12MV5TAcs6kOxquopll
1VdrGV+yqLPjOtxUfp+i+5RFsjQe4VzcaevUTqkjSBWzkcwoV+AmPgFycTZLbcZTuPWqrE4iT9Tp
nHp7HiMhuUMVq6VxmNcyaeTqI08x6hR4qn151Ek6vWR3XkzG1ohlfEOv/+lX1Afy2BxbQeIVCFsC
iFwJNqdCDzkPRok1PVCnmjjqfykp9vD+Py/K2Xo5yU4Q0Dm+PneucvUJ7ooKx4HB8WNQL+pjJrwv
RGcl9ZsMIGfCnZblonq4rirnxVSDOADBcrn3+3ROca97bfCSuskNNLkN8HCuKFqgW2zhP+M1O9mo
raCG04jq1m2sTqpHKzg3EXv02/7EHK9Y5rHdxn4GnI7UtLqk0z354/pKUYE1AqtyqaOo8rLS7hhm
wYH2fA21EBkwPXVByKxO+A+b5/fRlTSAQqPWbPIjqrZz6wK9erQgUTWcbRIde7v6F1jyhfxiUqFb
W1l+c7Skd2Sf6beTp71fvohwXXUsMEvv79weU3XYPAaF0G1ylBmGm2Zk0+6ucsOkXpr4RMMXlatE
TUs/3dnKF39GYXjgJvDZv45Hw9yNqB3/wLQ2d71DcjazPnMJiZpwqWheSpDfiypnYqSQHKqiLqaV
PNqdr02R9e8qRT9yZtZTZ0yeUOnX4PRJYM0KFdiFdvqXqh5mmyavE7D4j/MFJxA91ps4ECDCHEgj
8sDmLE187E3yxEYl/MunwyBGn+wQlDdCE3c3vB7RoKRRfv6lAgoF41vnzH6QlmLkUbDMPai5dOPd
ZRbvi8x9IfXem9Im6aqYoSya7bA9goImS9twsNJE+hQZXOYRJJ25V40Say43eJTjhIH8nkDaQKni
NhszD99jRUyLDi/zvGsBdIBPfDYjyyPQz7a0wO+Kk1mKT4NNZEd6JtdKyVvNRZlC6gmO/JzImW9C
LXGvxzROhVomaRdE/acFErqTXQj5FAoVtOcfPp5vxiEGMFU7qMIFFOmNMo15jp+mOyqpAPZSwk2q
+SdcVaPRWPL52LjJw3GatEqK/nIkXYMdd5CmhqJSFzQk1rogiXtk13JGYkj0DuNdPpLGc+1jW8yY
DDjFRAGibKmwu/qLtmYGTRtho6bw3xQa9/aWR1iOJeYvI//688MzNkoidoZSS/vidAMOYIvhCTxZ
HqveHomrPnm3vFPA+6ZYeiRJV6DHKm535PzDryaNSm9VoPn3egbvOzrPStbxDRJJADixiXl+a+Fi
VcqktBlL3gNvKW+u3e4yjbr8IPmOXafGejUVoVCbqgFzmXIstz2N5rTnRjlJ/r1IpuTcACSbl5+W
i3K9a68/OoD99bb10OTDnj/qjIEZkH8Zhb2jUWWjjXLqVpAn25RJfjKWrek3EZpME/VWEapmxg8m
vds/k9O5LDM0mEHhTjvTC+q0o6WnLOUTKivlKqFHVpwMDyKZoqSLhRCxjtFaykgpfKAuTYCiW4A5
2H1b+0HinxqLvspuaCe1THYW8a+AYtjWqzUx6VFiEDn61d7Ls+n1W94l0vKzuM+zqd/FtD+sO+pT
mD4xYfqju5e4iPGmWsjWwmeLLOgZJwzqeMvLOBglnhqIYHgO8cj+10CZW4yTUC0wnQStJYydx1Bx
Kpi1t+ehyfO0vMNu1oRYpZaZN8xDErokJBIUbC95pt0sQuaO0u7ZTn6KGJW8XKuOyk826CDSrvmL
QNyb5mqAKzy4wAxtccHL5ui/yofg21RvL0voMPD/FPZGe6UKZ92Erdd5RszdNDu6N091Q+yB9HBK
WJSiV43liWPaI82u/YGMqh7Vb9sFDxBCF+neMj5v+kkXSbU0nKSw0ULsMDFYmctHaYk76jRNupsg
CjO+f8NzQ8mM5Yzb+VP5BYDVRdjARO0HB2hBlZJnd6XcAazYd6XVC9Qx46tpDc6nU15LX3yGc80m
v/5NZcoAHLdZ/YA8Il7JMpFLsXrSamC3M2BmYlmhfiD2BlhCr68mUCU8+uqIB5oakGI6a3pnGMFL
jMBI/qWBvjLlq0dQS8zodqrIsdWdtd87CmQ1WofC93MhXbjGAF65Sqv7miu/JZJPS5jpgenl5AR0
KcnPyhOrE61cCCug6OyxqoYlqpGxi05vVq8uWLtttxZqs9uHFC9cHHFqfqJTuf38DFYCSkeBlaUh
7+Zt9D8xNEtziFXjLfoCO9/DyiIwb9ppiK+n4qhe4vg3p/i19c3oafFnJ0b5iNcIbkjlxd9nl/9M
DvIYhwcm8yfKc0+cEtbnEdUUzMozjJaYMh97igcnzGJIni+PR00qjDXsaMLEoLyzY8fA++SD+zyy
JzXTBK1oSgpbt093GVLKOMP7Kx59FW5RbmhJ5KhT1EGhOQChoaDTUJAgjLdR/Y7DVZXvH+AoXcI4
EPAZ83Xdt3Cws5ql0K7R/vWL3f/VHe51N8WLZ1Yfrv6vohDPYffc2JflNdpB/Wcl1XTYKrtVQIH3
ZzJk08eOp1KSeICWkUf2PbsoqmRHCfLL/bEXu6MpFACwyVvajk92SV+doEtyAW1WOzINxwYdmkEx
8aAm4K4AP5NCfFT5sGdyJEH73Kjtyr0HDYn9UxZXBRbVe8DRU6RHJ62MBBLFGOaYjgEUPCiHF+jR
2ZAtUVHVvBwheczcD8eAtnQVFBbwZrkiC/BubR188phfgPdYqYUKn5jZ9aw0Tf42RbZr1oZagXgA
OMdmTfkWJnSk4GzZ2KWCA1TZ/vZVVaqNobLdK+40XwLguNzVQ00YNUElOEH775JO/3Dl1CdMsHLP
RB8BdLi+xbppzYEOltP94XDIOTWD15pCp3Sy1p2ORZ95UawZ+SlY/wA47qOfDo3KqYuilGnTBe07
zArAvqgokahC4eXPit5cuq/fhrnBPDLn+kd3cBtc1F5n6DbKgQwdfoQ+6tMdQjiqJpgQ0KamCp4l
1qGZjLOhiP+zMbBY465a1AbdkwoGQgwgQ/8E4dGJGCZ76qiJpFazTCuSXslDBpAz1KTdu8gi2SCu
K2dZ1JXBVDSnONdvU+sStluoHRBeKZ7varVVSzaA1dlLG+8Rgx+g7Y/fk3FuyYurXiQhO0J6kOlS
m26y37octzGsL/s7CaLKZ1JFBGJzUq4e48RJwKFjc/HKcn9MwnmG4pM5vUJovrh80AFgIeF09RDp
QaYgwWNXTYCiBN6IMUYDiAYbXrXgmVNluIXfFnuKIcI8vNcdB6qbK2h6X3tMzVJC8e0d9QjKzgVv
wU5dwZ50GmfeIF/KmoQ7BB1JxaiKMlE6Aq/rbEwdaaCCdZCA/8VC4lNB2jcbGazc68oxiEopnU9e
Ad9DPj2A3xoHIpzTTxjWb8mG5U3JmpudgfGQuYmaB6yoCDmpkbudJvL+NgDbipK319uAkMu4Qp6l
iIS6+ksmd4TOAVYx9UpxpA/bbjAZ5O+Dx5Wx5DZDWYF1S9+DG1niHULtK4kEtPBLuYvnlLluUd06
YAnyYadN9rq/MEBC+/glm61Sb0E79cqWydRYhKtVSkPBpp1E2vDWcji2CZRMm5rXGU+bcsdhsVaJ
lCRA3LQV787Ab4lswPWRn+oAR/5tR+p3btRMSLGwW8d1ah+Z7M5/HW7+d/c1FwJinV68beXyKe8h
TF/DDNq+Y2IHrmM5XzDvh4V56zw6r2qsj3ABqxHbbcNbjLfi5Xh69XkLftXcalhFw3p14VV9Bosm
7JTAB8suPd1SyVni9EPpr71HbJAptLLrCevlHqSGpPFb0XY+7mAmAEkVxTncwzcqeDDCqgNINFBg
vokMuIRQU3LSC2J+OZgVO7+iDXFqeVvXX8Jkgc3MGvsmFvMtRVxjyfH98w8ydHw1wLZjEgrEhtbB
7etcmcqiy7f/UADST66SdnFyBRcFNTaCzc3YOGHvk3Lopi8hA1OmoVZ2ykP8zRIbfOHCfhqohGX6
3i5uT5oEjNt92ie+gtCeYzd+/yt0NSylCTkPFvocgs+pfV/h5kb6eiW/br3ZSsWO0XUdyo6OTuY8
nJc/xF1gEYyoi9eOdMtGUTIGYZytrA0aKg6y221vxylSkjJwnFdjlkJczT7to3gwCZXR7dnrhXEl
YAKktDjhUHj1nV68EtiyjUFYhnTBi7VhRg3F9jYQR9qjZHwUIESycS10cVTdMjrpUA4H7W3ejqjH
sWQMOpvDIe5F5me8o9zopNRFC7bmHMoIg2V74YEJro4sq3epXBIhepVFrtEqa9iIXqlUHpW+GqKc
1jzoiWp08KIMEHjozlewYHg9EtJ7qcLJL/Ay5u++r7bnZHDLKf+pJ+lVjeQtqhWHrBnoILRiIJdv
XeeJ+57e4x5NvOILmMfHMh3OEDRFodc90BUNSJkPMBYs/2MGFGm8AyWFhF/wAJFk/sPDol+sDHcp
JDCrf125GpdOGFAUhLo0BBNevbG0iq4kPdCDZkHqadbhKki87ePLIeips3Mktt7k5R+om6t4rmmZ
TWi4CW6HjVZsr7LMrHhQJIzLXX8LXKJtaGaHaiSucI/D39jh1bbNHmrnYD0uLmlQf5qMVlqPRtYu
O1+4wh3b4PiVBVNeT3Lp/9QarsNStmqujpFz5G69S+rOA8H73ptedGNW7CGl9kY5fyi9p5un6Eyk
8P9hmIY/eXxzE6Y3SMLAUWRVBSaR+Q3ydWxDH0WAyjYlc7XAy4VGesTno/dTtzQ5sGprJG7vyrkh
UWG1g9KjolZ2DxnzL8fO7NO1/NFEVzJIMWoHFUrxdAQEmWJuMMap8yFNGuQoN/4/pt9PMKDfUeRP
TfiK4Ph2BiGzCMCYFdB7vIxJOpcRTt92hJFMMUcNSvWV33+bT4V8r9hEDlIyy8Q+Vwa+14thBKjE
n658R9aIjKJqEOwq4SbGdQeLjlRciY4JY6dBiPF80QZ8XFx/BOqE7tp6tcPF/IJyBS1z9FjV5Hvy
7laNhOFs1eK8eFHbs7rPWyS9ib8dUBnAk3xgGYdVjWkQiLAZCukEHUgIvWiALyKmR6o0HYdyMlgi
vqReBMuiZsp3/9xYIQNBpLfIm2qBHnd+EXac0Lav7t82GizdwgKzBP0GTjONnG+HR04PrBDws6TO
dYhh037jsB9vMBV+g2qAZsHFH+0n3FTSpno1XF4H13xYmP3GUuCixwP8Y08MYzUC6IwhLpuYFNYm
g1xJNs4LPvZoJfNrvAGXW0uWzsJRfFKGFd6qex4W7pi/MsjNlNymChznUP78LxMxYid+VmcSTs12
BDDW5pRNz4605JS/fRrYhlOUgi2OFzpRJLbw/mef20uwvaXeeS31XHO71Yh9nIQrbwK8ossbwfhB
LTIgYJ50YXsGV3sSq6x4e2jva6fYG+mSyKuc9yHNtZX0CkXCoUFbE8P5StLpRn9dTn7G1NoR7c2/
YI0EMUwjKk5YNYZJG8KU/YXzMeaA+MBd4tcxYEcA2xKRrdPxQ78QRjTnSnxf8exxlInXBuCxxqyh
C4S2xNhMFSkC3OsH53oB4l9K7EWH3j9bliaBK+j3IaRlUkla4AlN+1DjTUOEwjV0Xc6lGvlexeMC
GwKj3lI5tAKcdp6wKVAiy36gogoJ3qa0pvMayuCpA11WABH4eTwEJ4m/J56NlIztITny0VIVcAjO
t/xAEsYlNTqKaHq7GHeetDtRsuGC1ql9EU440WtwHmXKrnYi/3GDql3YTOPqQhQqdQtLFS3HEgWB
YkHGJB/NNqU67IIjY90dRn1xKULHNVv+rZdyIisqhlWtku2kFSVQ6NkMRp1uTcu+NF6s2sZm6098
Lgu6Ti+sFbjsJ4bUiO8uL7nIZ/cH78VucZ5HdW4LmBNJzSt0OgrmlLHJ0nlfAfPYVsES8Qz59l9h
U5p2eyeoB7mK1I8SWZxFxcGSEkDNYj9yWk+cEFJZI7SZqaXJzuR8oQZPz7RB13Rqm2FIpqn6FAMe
Q2SdBo0CxkCi5BiZJKTQnWs1mvv0p+jgnpzEG7VQtKsPaS5TAIopRp2tckbU1d32DavRTPEyl+4y
cvBHejGbOxbyyAOekTJfmRm+PSpE0WNqgmrTtMTflk+AB+uvDumYtDkwB01rXqxvGIflb8Z2MUDN
JI2MYKo9jxI48RAupv/DY1ZyxprfhBlyC9O4f6WIZMydG9T/6iw/iqAGYbjUrB+eJZ7WxgG+F62v
S4OjnnqiciRbjS7aRdbr3Rhb8NWhlVR2hLdnh40DzJ3PECp2cx4xMxNljuQ3aE1xecdjXYJSVNvM
SFnX3vtubNhy1dTiFVsBnTyINe0OYJnkZgpl/pFQvAuvD/jod7u9T3f25flReArdl7oqU8sx8yYa
jX8tcNFNjd41xuMz7jEXnPa0IjENo5qjqlXj2gGS1in4/e7oJS+p6xtseHy41FJzsGmogGziczU7
mn3JD6Qia53LLIK5iLeyUncU1zNDPbwBkn9qrBbvlJ+tXqWxbvn0bklunTsGW7LUqvCYPGf1i99w
jcUXLYVE48upcsfhbpY7Q+2xj+DLQ9IcWy4++rgQihnTsxcFGBIixzjmdUnjlf+dM03beg52g83j
6flrZm9xqdQ1squSEpnERKuWRNlzL9czqaSpao8K6k0LWVTL5TKecKbcQMckhtTxb1IJYXVPJ2sw
Hv0ROLwZxfGWUiaGl7VRsg3ltcWG7n1L4ZPVIu/Yx7PO8YOwpoO8zXF8u3aetDgoHgKzylGj7zIW
1LXymXrmlmowy+GEsYYTpiPjH15k3orBX1FYRy//FTZfUdAQoH73AD7TmrBBW1nNCbA/Ng7jkyPi
bT84Q5nAdDMu7h7AkvuscfNX0KNCxhhyJ9CJDi2MVcM8e2MH+ayIZbxnQ8lqupQAtsTn3p9Rn+8C
ge7mUjoHedajlutSLt5dL0GNZP928lune1EK0d04PTRfdyvxNIDSwaT67/EuFkLhJTOnzk1EtfZh
adJ/a9/IDjZiiY3qiSTWBHsQ06RUnu3l+btP/TxTeOWLihbDIma/rvsbqiboj2tK0rnjjIOX2E1G
AHT3zE2ETDkzCeNYSqzsjdetU8KCRa8VDZ+m78EMOzKkZ6gXlBRkc10PXnBdO8VcVOH0qpAnKoZK
s3sQVCZnb/2z8B2GDTjWY0U5HqhQ9drwTqgU9Wwmx1Jp79EPLMavNbOjsyHB1n9UsNfs0MymDpMw
CtXWZdI/ry3rE+Gi8wkB7ncAGAsgbke/zt5g0qmGW5FUZx1jr4AJk652Tk1GtA/zVnLnQanTOZDT
eQ4ZoCsaaYt6tiXwXkJM8Mk9lukzCzqr+TWfFn5Oxl+FwCAfoHp6QDzuy6eG0akHATqmSZ/YNXJm
8BMJt9e5BMB2PQT33qnqG5ujmTp+Opqh7cGCVLffZOwPW5CBVhdeK631YIlPBOBCtSaAwFJVROa4
CnRWSjIZhiG6bGQcYqY7jwYEb6+b2SidlL8EXwBAAKfPe9NcRU+vluo08LZQYDWGFQ6NHuIYlkcq
VbMUDF6/+Wlrt/1dBTQ3xQltnP3gZiUxPvpBolNvAXhlELo5JULhEnh6b+OhYeCrDkuA5Ixv5G5j
VsbU8xKMWPfGayuOxxSL3k5CCl+MmKcRZi6LB+8yZkQUM/VWkreKT5E8aiiuz0azCYErPR/BxoVZ
Pdp2VJ29GS6N0KNxCHfYeaJ78HzGlGzEjrWqQ4wd61A4ikAEuSw8DXVuF3GJjLwCflMNBeNSzr8c
hDe5+gXqiyx2GCfBkZNFGw/sXCY1zAz0ntkXSDMC0n5KQJSovcxR7YNzna3BgLw3IGX37TnPz7un
lxY8VkZ11jwsnnk/qucWuSuVN2ZXi+hkNDDkCH7RxTUyN3twjuiFB7WGP/GlHO1B39+VeOI7R3zJ
pD1ja2xefFNRb2OKrj0Z0HXVP3mAAWdQ+StaqmaqSv3c8w7D94CVLvpiz1ipGoKXfQR4kD2T0lXq
zUWMxz803c6af9IdD4rgayI9rwrFPP7Pgjbvzfhpg6XjPESo/o0Gw/+8dXxhlZtZTNUeQbJlW2ra
dSD3rwfNvdaNgogDfhkkq8dw9IFwnj5GWsU9R2ZAaeFc40Xx4XBkIQKcN0/rm1+fcBTNjhkcSl3V
oH8Xo9w7/1Yfn7dj9dZ5/YhKDFF0gofCd2RURY1cDRfNDNWElHL81u1fLLSFKM8gTA6x4yGoHVxn
VXYkqxojwmEQo5n5UTBYNhp1W6C+XS+/MSBdvu9GgFAfZUw9kkI2bBtjDfDcpxHHkKiON5YMFMqW
OAhWP/VLjS9WD0vbOXGQe3cPHx9hHipQ8r70957f2NPPIBhTm3ix2lQy71V6KgTtK4Uo2MP3Eraa
OJbqdYM9m4HAYLbOYriSFAC8p3xdzEejkMBsoSizPeg61IRj7B2IYJHCyI5IAfzvIxKT8yFO+M2Y
dxMnKPTeCvQxg5tNsw6zDlNtzTmDU7vsE6KPoXEyHO43ef8d0V7/nbCp8X1sF67RXctrJ10QD1ZO
ZHsVAMcUKE9OS7wj187Z3IrKAYIjwGnONK6GHwtFq63T5A5rsIpJ4s3KAHANHuuwIjLuPnMIWpvn
lVFkwoiDzDEyHOXbzGWpLuQ7Ohgfz/wAMh0LFBOI8DbiSrFr8rY5en2Nald2TbaEIff1Dx1alXH0
fCuJRitLqnG8tQMukN18sId7RWD/xxmDXJzmtbyjIay3/Yx4v2yqzbfMbpEuNeJ+r7S0244ctvDT
uUvT6C34RW7JHMjuzJyUT59rb+2CtPal75ENwAb9z4kgROJceysSdtnA/FvLCp+ZheXcQhI3tzRQ
5zW8KJcz04uBIhEdZ7AnUG9TlzeIlVk0gam8r0hFTs1MSdFQzSh+QrXckrTHQT09yuybl2s6in1L
uZCMz80TEJHuxQ7wnMnecKDTvVspIGLPnxNL0xQrBU4d3AmTAV4ZBAetCxYjOJdXMb0XT+m82ZFK
PSnkCk2tsBCDTj74t1ppB2zq+5JEtUyN2/4GBdhpmByMr54g4EBlhC4zyaYn21H2C7mVcfpNVwyl
jKAN+hnhaAkMaJ6ESqaJ/EUJ9XKd5XXddFj4vljNNr4c+AoTZ4hv9Gtu6lVa5hCAoeT5n9hIKrUM
5tKWtkubJ4lI9rGwYINO197bPWrld9NvDdUF+/Kz5CyDK65JnOt1cFmRrEUP8HFC0JgM5kMM8gqx
qB6bN9cG9MtwfTT3Wp3dQGQKp8gwiOgoGf6JlLnwaictwpUI+NVCkc/fX3L1BGUKOP/Xx+l6RPx6
drAqIJo+T75E6211BhlxQ3yehdB0jm25VIDM0IQ9Lz/Ha9xeZ8RgyGLO3kpfPzGZ+S3rd8Bp6DpI
nb2z/+1z21cn930woupRWEEkto1kb5ep2Rm9JN8zU2pOQs0iX4ZEMOAfsd2dHn+a6QFeHBUxF9Br
UrnBzMV9Odn0lwBH2lt2BUe3CQRcj/501ipa9Kmw66JmMkmHoG4IW/NalSRjcXv9HQeAZisWINSs
SaKqULGoClSXD1HC50QktGMjnrSGjypBFz0ug0Sh8VwN69EzPTyxUb1H1UKxzyfpSVoz6dAehRGY
u/5XLkEqC6uVtPQ+TnP3eKHNBJM/FZ1Kf7LV1706wGF/EmcMA6QenjO1kqUV9+Cm62bu6NdRxMFq
m0rS94qgsfcuNPkQ3qY2904wCK2UN6CiB7IaiJ38AWpO+Fd1PXkOrxmfoHopV2w6gcPZeIDOw/QB
fm6XRwqiW4E/bbOzgdq9S4/w6hPR52OEHk66VlkHRMo5z3LQR3b+lYvJPxW0cGejqE6HSwf7Q+gF
NSJ9S2vpwj7sto+p8oVHorrV4WR6Z5XNKZc9m1vJrP+GY5CS/XFq3oGoUiJ6sVj/B8hKuxy7I2yh
9gQDDdJ/4nAY1Ue5QMRcaGDzP1pxsWyh0GOUr7gORL9DPgRl8VIsO3au07ciX+pe5iPAle/uMPZJ
Cfnqs3pGX1LyKdEPpEeu9svmKQAHpInRiOvPDsD/byY55sl+VvXejYlhWtnxqlFQOheDe0k+MV6R
c7w6S03bXVGB35jDGJceqnyVdmcizKW2UeTfyr8AeiimUxsjS3S0LHNnYLpU2SNNEBylALCj9Bmj
a0BU5BOuWomlW5tLI90297V9/rd2p1TdhGAb4PpDpJSzboAAgTETY8CcMY2afaWb8jyNK2TQFj7a
fba9thKBvVoQEuVPMeRmM+Tb/GDRfHDa+UH8vFXpWufu6Qqc152z39CbZsscK+c9NLCDorwLRhXO
hIzwVmzG1U66eAImlN6pX8bBcvZih0fn/HEoDmJgwintjPH/4HkE4Yblhm9iEeAY2CuLMWhT55JW
Wv5gGOL86umwRUn6zYnMe2QOdlvaYN/RQgETbi4Teo+iNFguKXDeMcIuhS98bHolfQ44eQ/triOG
Yvzd+6cOUF4Diw98DZ0mBrJn5FoQ/Y8kXRcOO9zEg6M5+Ve9JstmrfDZl+9bxq1jWVQE+4JXm3nZ
aVKlnsGQ5v4I82KtTHH/Jl46u4CCDFEEUG12OIq8yrW5Vke8ZFiehbGD3BcYehAWlh6thSbBJT4H
n0fbfkXo+xDBWD/8rhGOPciu09N2Yp09qGnLAPvLLAvgSRZNBdTToOmkM7aoBWQMWEqI5x9MJ0Xy
/JIOZthoCBiIjYaBtxkPvqhH6ilKc+OfxwT089SuylQ9fQJkOw5BvwgDVwnEILjKCJ2pmkg+veOL
oMgQAhnh/hFJQJq1Sui9YALXZmvrmQChVx4MG8qqQXqWxNjhgqzezZfY+KsSPvSxtPlfkVk4sVKl
7eNCgG2N7rylyzZRzDXxAigBBaLeT7WnjwERcVQRu20Qttgh6DfYrrRPKoOZDgKL8+fvKeJiXB09
uh1EnJiwyfolGo1JH+vNdkWa3YihGj+2vLe8FOU3MQh/3dC6mILsHtQft5ArcrizX4TbcaeSZPCD
gDM/TpiDSZ6UWZC2v6nOCat1phUazMi7L2VFI4SQIBTLnccsRF1sGClKj/+5Hv9/cfi/1aJCSvoC
XPmAUgz4JOpY/H6e4AI3t5PGLpUQuVIMAW9tgttMsVl/cZQqo5KX5yoPWPT4TZJKKVEN/WfwzRg4
g8z6LakVtqUsyJ9TmZ0Y96aoDqcPxRUHWAJOSVAq/uMYwQrxBvqxpDdYcWO97x7dsI9YOo2XXIVi
tUz2cpL9T0q9me/bu1MJ+BQPK0F9eCUyO/Pc8YiIdfMYgUodmqnRkz31hqwjlIp33rS1zsAWrlto
/yBePr3qqwPlr1yZAKD77C9k1vUJr5L3WJcuAzI63+XRJE0/6CqCXG0dojsMJIH9J0laJJ7D2D5Y
W76d4eZi4oKA+w59grf5m4NH4bZDamRNS38J0FdLMACwcS16z+4ihE6e9PXpoAIjOQhNIZPEE+Um
/SfoOihll9FkwvIhHNiZoQxeTzwvZI6WoGiPS56ag9P/XrPGQVuLRqwWAbszF/r8nam4ocPwZmgK
TmkS5b0W6sKY7GmLn6kAIRlg/GjBn2S+9yWgbKHb/yWlzdVU5EjfeOi3SVa2EuRVI9Obi4Rfxg7b
OvcyCR2YlGp3oYLpj94WNe1up0eO75Q6b3kK1fmEvIVShZo99BkNb8Y3/hbI5Ldgbe2GO/59u90f
AgG/UksDpFOjr7lPf92jZ6mWJhH/4ZFPtU7jbX2ttqm4VGGoacl7UTmMs84Mwe2wY8SjpJM+OuFf
UHTw5TFiILgHo1l/czugIxOOsSDJzB8g6eZEOVSfkFf7liHrRawEH/PBiG2owNGmnvif+uiQlrOx
HgzqbpwXQXR1VrUqTGBht3QqMbj6FBDGvMNEznhG0f9cSGi59IFYXa5RqpB14WHYOxmSH80uc0qv
qVwfNJJGMbo6MPEpFLe5epBn6qSDmKulCi8BMwNWbcCRnipBhry91gpAolCMhv6huuhyjdwxgLnp
krykDWch9SJ1SlRWEz7DzGbti7RQD4ke+DVaF7+xj5CEE5ei7TW2EfAHAILWCGZEEh2Ct+R038iq
JUTLN2A+7RPNkFE3wmvTIvzemDb4AV6xC/CEvTVPMTPozSyDB6THCbc3Zk3ziplcFWymOckuft25
d9rtBZmKUfsnQ3+n2VnqdWimAkaCLTF/VivUHF5z4GeKpERy5X5/+IFaQoydE8hoE8od9fPrpOCO
NCprEJodZF5L2fJHTBG8D1Hbm0EqgMm+JasFzszmKBiJBLJDwyYoqhvEl9zSSm5B/dINo6l7RqBK
Ej1w4RZnR4pn3F2XFuUzh/qGk1xhEyNUrxqRUrE0A7N2Ly5QRsbo/ziTNz/gixudY8iKsT6uPGfd
WuEHp3mQfUPKm614gIXlS+1SA0ovnKwWmrGOpwNOp3Ofp6EVk9PvpzzvoOwR4euTvTG1bMiszi4e
YvEcai/djUJL8Et8SwNW9osTrWvDQ7tYMHyZ8ryfyGBlkuNG9z3SyL7w9lQzbgDSgXzunhtI7o3n
0XhV1Qxoii6m8cHB99bdFHhyfUINLWNkrwY/yJVvq99N3Gmypj9Umr/+loX92vKuu+IcOMku7zaO
WPf8NMN+ihCvOfH/Lk05HPO237HoCP5scBa0gTTZ5Wl0nnnj9zZwaoJdRESAXaxS7NqdMrfuAZgc
O6+E2Zfz7De6ba02wq8lNwGxZXviET6Zlr9oY4EralAb14Objp8cMQruQ7VmKhG8L5gMpiw8TiV1
cPvwhAUO+DkVnsUI4X50yiqtEz9vZ46UmIiNGy75zSd/tLtg8ycpACMy61p/A86lFWZgxaFHxFIs
n2xJ6MzCw10V6T9mCMZRqqoM6amhKH3AiWaqUsv3wZk0Dvyy55t9ffcRO/jvvq0GHETnK7JWUskw
4BSLNhsSC+b0IyNR9Yixjnu7NaPsk8AWI/Hy8HELqoWtIJggqOlDdajTDa+ArMIdyyp0R2MaPRzJ
Yrh6S4R90UdcaQGCdlarYvXAHz1ztGASiYcRu2E3RfImk/C1MUMWQX/gFYW5AVVflHxKto5mghQX
tjf/LT1Zo+mkppv5khr+WxjPeLijFe6UkyA0D/fh/9BofQQGeGBuvp85vFtDPhzEVDg8KrAyOLkP
sSLkWCZPcak910GaNUzKYH8D+Shwr9emLq4JT1vkMKcOuAPIyhSF7Z6C6BULWyyZ9V5nJD9NnrfG
iykyy+pGsJWzNUu4SgmfT5n15gsGM7A6rlkMLPSt6GBEEiaelcsmIewEwAt9LXNwWrDgVvoPVAz2
kqbLZ2xCukygrSildYIWonOJWGit4XmxVLip32XisOkPaTVZd0wQA/3fmWXSireMJb1CCmIMj055
Tkg1uSBBdhuEjuCRD9r3t5u9/SDKz8/e4kk2RKyHdCLO3CYelLo35ZkeZogsCour0ihI+fsfOkZx
2F2UnX20RlFhB5ihoMkcm8ubW9zzJbYh+sFMNo7ogJf9ZbIobZ/ssKf+gfTL5znO2ouSkbMF6hyy
lnSqTb0OVtz2Vhx5VLNCuDg0RHRlKQGxymI+47Us97RLsuIQfuOMJSn578bgr1GNPJfxn1vtdy93
PY+IL8M9vHhfk98JW7HhxwwdK8xcHIx6vqcFoPfXrT7pKCR2Nt3c0RTrASVL0phPiAwlLWdcMspd
fCY+Q11n50cq6R7VV1FVRdaVq6phTAq381/2KGgvi8Wg6UeMkLgiUdIsYUs3PT9KA+/NNoUKXqhr
QTAc64+OsiamgeLJiNPkCVKOHCpHuH8UjeNfqrn5tUvbDa5szkK1GPBkvvHJ0TNzv1vGOSXTqQW3
gWM5+n2sx74tbsl9YPcKTnpyd5seMKU7LKqBmq5R65b1S1FQUaQzHNLd9MZTX8AOsVsfoP6LxLX2
jLHGWmzRqEWDRhTpaUwFFOLYy1+1hGdBHhDpLXK1bg8iWNuk/Uw2Lbd1wsgCM4NZEPd3Rj46f7t/
hNcAy0VggneZM090laTwZnDFh7RcgscKEuiG5zz5r1I+q6kvDXtdcnXXW/PITjUWGVhs8LI7ZXt7
wzv7UTLBM67z/LNjNelmfaipnqCPnAVe0puiAk+KMwDMVWLRkMQ/P83p3Mno5iJRvBVujTzsVcje
4sBFfAZHeqmyczQXpELfA2tHUgT8kPPD7x5YJevbAZkgSJK4Tlk+9P4u2dFq5Y4h3/9ujKDxPpE8
+rPxz0P9VtQzUGn0/K6OPnFbrDCAJPAknKY1iDhXFkhn4dDaaSUxHcNQBt0r/LsGcLPLWBsTx74D
+L6WMrTr65iNndasvh4mrPxZk2F4mkAZ/yUq8Op29yAxHGJC6anZ4oeGdIOIlHMF2nFv4ROvpyJk
1y+0w4dlBCtiue8oFEqXFffRZNh5IxLXiLCPfQT3ELokfx2sVLSue7aHuC2Fiwo6lzTzmiJLMCP1
i48bhyGyDsRBwKftbJI1npci++WIneAiQJu1QT1PBIO7qUfu86F3cDCeCiVPgQGfa+zTe5SZNG+S
aWi2V0zdKjb2pYYP/pkQvXaElKr/yOeT5sxh3K4QqoWG+TOJ7pWPj+QHPVVkavthNue/92t+QpJh
4C4SXml6/e/y6pG/jVL1VCWfaAKS9Q9IZveW/0HTiusQGf60Y//oBlIW2brjeX2UcaiLOD6m/Her
eRt/LAVWrPJvYc6YFjlLSuf6O1cEx+sfsYcua9fyVqeqWCCsLZ4hUBDJ/A4AB8ZiApj+cPHKluS6
NFYQY1DYIiRxIH/O8XRO25bodvihwqclqQXeFAAmOuhel0J+kT+1j9bLHulBXyKz4hH/Nibrp4N4
sNhQhyxd8IvjhyjIuaAUB27RutDBg9DNJ0WQ8rxxrVOwWi0n9AmO9lMrFwnCh2q90FVX1Pbmp1W5
sv7uxscg75fdKS9IpXZRkvTJQjewokGk6+kztjTGHduOIpeeNwa3de2z9m15yX3YbYagRB7sjlJP
NB+ImfESL2r2tgas26T4rigFNOadEFmDo+46ox79gIHQi9bzhUT/hk6KpBnWenjST5bD06HKH6mz
AA9TIqOCasRj3MFoeLM7r4vkksZRUarflveWWjdr2ByA773mTlXG1SbAMO3UHEEGzk58PkLwG+Js
gkcqrc9zSJjz2mtyCgho9f+WWsJ+4Fele9c9zSzelzbMVsntUpqqVS608k8Pwk4LP17Z53vN4l6B
FwxEf41oS2phH8J1+8g6QWsdoFMMYwG+7Z9mYA3LvI5u8JNx/vLMx6499l6MPgRScUpvD34+RcLz
An6x2QgrRazH4Dt3pVM6m07CDWFAJA/cEc9eAbH4EeK9R8OXqPjigIpSd4CVS3yMdOs6qBMsYILy
elRyFeWW4yaBzjzdhrOlMfGrJt3ics0ut4KGzQbRDxOCyFiOEh6Qwe/tTS1jyv0uOYNTpPHbHSF5
kUlIREQANcAzaIMe+ZUshtc88HQVK4sRPgYlCTVwR16R14EW7ZYL7DXAj0V6Wq5DPOkvytuWWFjd
v89mq9R1PSFECQ2d3VPcuFrhwDykv2hrMb3dFuhAyv+NF16Nb9OfxBBsKqDG63lGbk7MyuxIcop/
Xvzk9sg3KvVawbEKDdg/G+/jj4N5bsNka+KcjxdYUUZKLC9J5Pfwv7alujrtgqdr8soET0OnsuUv
s2n3q9ogi7pplZOKWQC5AU5tm7+X7y7gppdDEmQWO562x3d2jO+JM24bae1/ESvgca0TARPaiIIw
33CKQwqyqJbp1970z4IKklFBRMmOjZz+u+SqoCHqngvPz9VL3QdAO+Xr9jnRAbgru5oaG0bjf9GK
mwKNglglzvUPmtKM00rRBtZ1zHvvbsvy5VtEMYJ6Fay+ERK33KHqIHqsq2EapXYjmbELcU7lk9vg
6f/GOGbnI5u/oslLsFIfoedvvjAGLM81LTmHYYUfi9o0RTfbq1c/1Y3PtLKPE4pGTGeOsGUHpaQ+
DPlGDeo5KMD0dUWeZSIfm6NeWux5QwCiUBXGneUllutVL33c04rJim0t3Dme8RHDFnaTvRES0FRX
CEvfZ/17LcOt9Vo0lj9p831+dUxruaNKfwcHpBCjPcGQrHkYo1+W+1rbWrSYRAlcAZJTxxqBoWPC
fsiGkt3KAv4dUYYB7yhqgXEfFO2iQJlbhNC5sZOZrB8iFA0u6QCdnbUfMGwTOLHxD4sp24iVOY0N
WnIMhCVHHtw2kRh5hII7iMV1O41mDrzn2BOmsu3h+UOxNWwqOOVotwrbCPqAAXQ9PDCzRE2lXnFU
kis60lRTArwmdbE6/3PTgUuuG8X/cxy7FO118Y0sZpNDPhTdlYZfNOZ+VJbugkdKnWSowcyXMKEj
dERgpDcjxT/URwtmqzTjT1l52kb9aioJsWmJc5K7etINynXykPCdIXxk1Okj08fUKxC6qh90wkIO
xVGVdE9Qu1WXsDWkVprbrThxDOgPZ2ikz9LkUfcVVBQbap/UFy3hwoVelfW6S5T2+jNJneXbfq+O
+TEEWTOdEhDD2BvoWFXoNdDLSBQ2nj9dT8MIXCPfWNgtuc+jTk5gMxSEuWnCTtYv42yDpllqNQT3
pCexmY2tM9mLWAjdbhBcMChAQsX1UZwZVXLd0Cu8jBEAxBWHcvOpQjdsUJ4o7JsF/CvjfZvHPVwC
HGurOyoNKY9TG5fNT12hZY8zi3ecdiAs98lk1aqJLv2m1W2pGpMAlMkE6PyWQGV6lWSpLJxyPnYX
LRyP2qGx6TJTojM3jJ3LkxWD+bZyEeXp6RTDhEPAO1ffJD9S2pRXF1HaX4kYFU1nFNlG7rcyjNsx
FpfJBozclsteHBC7KtttFFEMavwAruroDWsBJRhf8KwstgQts0J4s4E6tV8SQ51aRA+R3H7+QEk9
G/RA/DZwBhijYfoy7xIfvhgj0VSV74btuXSdpEikOD2gS3DZQSJAn0QwxAr3mbOALGgNC/YN+8tF
PhSZ3uIgZS+yl4/CFAQnQ8guGxssZceLWOBJKgkhgI7vERmoSp7puJvBUr4n44Fv3KQA74nn6Pxj
v8v3kPvpDolXvJ8d2c4n9A1HpOtcKW1ugnERvpTsylk//EYEnxj6vgVcFSZ0nNQ7wSRRd1UVRmJi
O+3jaXx88G+8ENPFnLmT4pszkM34FIrdpc3BL2VsJjP/NUVErP0gkVaPTqh+4Wi+4MnhrFoEkjHN
V7nPlB5kp8aVDntxlUbp0ZWnVj7C039tGGxE5b9o0UZU9ALApJX1Yl9Y5zzAuQutaPvJ43k1imUj
d9x+A78U9Sc4WFKiQrszlAMcH6DmP8Kj7KPPHfVpqaqQ0EOUrI2SYUxTzJu3PfMJ5GzH1gDmuCeO
7fuxU1KINLB5JValHc/XiJuFDYjslgEE54IPY6FCmrlWp+HT26KX0hNO82c2XDWdyjugMVWMIKPN
J0ktqZEbs6MiP1JHqqmnzsNJU8drBMT/WnaG3uffMBfBQulM84iFHASOgctaLQUDcZMoJVgVBmgv
ekJ+CsOzA3xtKVoVDN1LrzIRRKxR4iSits3rcKR2fG7U3laDclrSXoTH51+CGt1myf7YLdzr9GXV
uMHFfNv5EVhN5RfBj0BQeAGL3WWkkGhA2tjTkkMqk9MG/vnvwzuahntMKdbo6Fuxx4w/Mhfv6kI/
kf5jag/Yj+m0V23tB5xYtoGuLyabFOz9KEyYf0gNFmZdOdWS6mIfGs9gNfibsB5ph4WDjFRY4v/t
pgGrCYTEc7DweUCLJ7fdV7cN9Ome9jveixFkru9KeL6nGjXIe0mhe7alKe8mafdeYDfZUqbWsJko
iwDuyTaXvs3d+Y5Wed84sXFRxDzk/O2lO8YCxaT1o6Gw4DK8B8llitocX/z1iZrgIhVvJFNpEIPR
x6JmNPVmhjooqUbnliV5YvCQhW2jXuvReKIt8hjcybjp5Nj+6U2OMkO1vVBHogPts4ndkDQhoJD6
9OF0YG7Nt5TWYtEH9oVdYFas0PPTf3619s/eDN7Y+fl/RqsCKDnc4RGo+cuNIKVgNVIj5JJa1oMO
d7ic7iXxpdVQyT+BF1xYtRo0gja2FoovzOBxloXJLiQNxNX0MtpleM3Cu+2WR+FkRCMHt4p2lttf
ixoEvUVLS+BHVlEMJdRImjizDHMeoIrGJwmLpzFqQqh6U2YlYtXOu+TCviL3Pn4fOKy69gFXaoAI
AIuhY9PYOSoFj0mWcA8kO0+2ogyE3EVAYs5TCMHXVNkK+5cyvdObTXu1BZAnknbNT8NtfSXgqRpf
XVax2KOaBH6JdCieoTSpz7+sgQ27yQmIjtR0qqutND6yyzrTuyd2urSd3qNJgaIVku0YW6xzJ+Fk
TY/i+p+RzTvhhrE6FVZSEPwZYtnHhO0ooTmmKkcwCp3TWtQzSdzRvcVNyD+4+3q8XXOvj7b/SXtq
fNEUFqv40cMye0JOAF31wiuyKuROp48K4y7Y8s9c5cd1HncG8Iifh/p1+xiLZ6K56k3+CDmFX7Pf
QaeA/5PBhrsM84TqDOE9RechvqJcKyKEbuu08tW0hoCixelFunsbovcMXrMBtdEJqR9tJLEcowi2
Zc2LFAnnVgmftGMKy/FWJE5ayoHTO9jLCF28/FMX3VG8iu/W+EHefl7X7qFj7/bLWFlGn8JrvG8x
RK106TIFFZ0ORtOw3+jq+KLaEq8Msp9IOdc0u//tF2pAT7Fex39h/zbCiZr432aReAqaE0b7CFa1
PkM+oc6z338W3ahAYu+UqLjb1Yy0BOPAfB03XpiKL7m42gf8OvytjXRFDbGz5WMs2MrSFUWa8vso
k32v14Wve6w9mlEMSENh6lijf0h/s2qZNUhZ1sPe9h7u8OTBTbsnedinUs0xIvVtV0/3gWtyHKZw
DBLStNVObTR5LEpZQgpxnN7gykTh4zAV791sjw+u3a0JTmxaDkW0dQ9SYMLtHxxLpOh9fm3wf4Xa
pKw5jdnQWFuAc1Uo0D/Z9TV3MjNV7rtamwjA7OEd5IaqpW25Fq+4jAJOp2UnwMvXA9dDJXVoQT1j
XixU2X1dPikuCzEWUHHfjx1P7jKIwShgz7hdptVeGNp5bI4twiFPVWEE4YPdMTPk/iTcxUUUmIeF
3si1eXz96kXa0EPnrG6MLbwzh4/t8SRDxt6nDC6zoFM0TfsAOg+deab3TJ2i/Kxnss4MqxVf4sU/
xFMRNld5tLLpdck7bsqKHbc6pSX9UOuImVJ1aLC5kbbI4gjgynTu1Mr3rpYNsvX674SfqPpX92mt
mOodojLL4sETtxCbA8NjHBRAxb9ESaylX9r0UVA1PcXIYSWnmAVisBVXgevdXrWnB9TCmpfaNbe5
FXc5PIoMfk/hSrFuT5mAPSbiZYSHOZ2rNwrMh/8jopCCxdLXvSlWrJs3uUc3nPlIICiBaHbIaT+T
Ju9JoGBTenX9sysypDiCN4Z9VxzwULIysEiN/NvpbcVviuY1hI9hOTwEc4PMa46O7elQia+oXuvH
Z+FaF8I8vVFXzW/q612oap2y0+wiEMc4F5zhRLLqNpIhgsIHUhjwz/Hmy2UMj9zfhzONXgZFRqLI
1qWzn/6/ZxywVj5NYqWhTDNZLgugoiRZyUIOqU8dshGfWud8It30ueB+LbvpMo60JqEHBcFRIM5K
uUj4AgAVsIIntUT6zOvvPtksVykZUovCgB+AsXVul50aAhuLTfjLvMWm3+BXxHyzLNjJFF+SPFp0
wAmJaALMZIrBIj1P6KwXmI9sdQW9zoiYftc+s2XIcLuCEe3FDgOuqbyrMDjgN59lq2jxoPBNS7Zk
j5gvPYC3FqeSN/UEL8XP7Rffkt1nV9hSxpndwsT3a8fdwHqwmYQfH5+kmrUB4DMihDc6TM6ZlH3F
jEC6DtAT7zFcdhS07aPeJTBo4RfJ2nhGMhBoHGA30ubphMV0GWrrSvPzDWq3bFjX4U4xKof61pR8
Je04IJJ1zGLvkc8LlExdbq7RWtWT+Osc4CJnUg6tCRt39xj3gr3Q068ddpaPlBWZDxMM1qseSPcu
7DVZSgSKjXyB8JbF0bFwG5JEMuXLfpbkCWLsx7B4B88sKEawcKz0rNLbv1B3h9VvQ1Lfe9kuEnpB
GeKyqHU/ZZ/tiqMCrjPRqvRE5ZVPai/YToS35X4tjnShi3Fw/SnhcVDS5D5e2LdFYCHSz7nnAxjO
JmzaWwZ7Wgs6kuETx/jcn1vsHCp0zznWKWvuJ8FrLH3Armrf+gE4rXjvmH+gQledGxood3Gl5y/4
DgP7qJ//k6jGQIdIQK70VLmr7mDUV/zxK2/4mvLM2tVrLD6lhiP1cj+aeHLv5Mi7vf9u5dOWrMlk
n+yHJ606oNxhtrmIgCJAzgpWKjy77z/QSJ/6izxfZ6OV7pCYx8uK5eOSlYIR0Q0xG4bhrYMqx1pl
hIDOVlaZnZUy+ZCR7vdoobl6K2Oz1vP4c35qqiyXcG+WjITjuH1tuzZn2VXCWNHYxFqMUpaqO/8h
HEsYf2CjLS8DVOHriTcJkUlq06xf9xkU/xCfPuZ6D8mJ4khnFJMPNnCl3y+Gts6wV8PELFZCSlfc
9gAUFCdQVH7B6cetjCdpCMAJUdUyhDkdIpmWgh132FHx8IZwtTlnVz2sgjfNUkHeKpK0Iqp5hKrJ
uZtNZ5nbQz0GLbWe3Bw4M/nyRo7S51aATWd39A38fIbt7O+rQdZ8txH2gbM/kKdDwHSjpLqq5elw
wKGdmEFVkTdcdIjb6nL5FnYzTPLMySX56lJ1yKddOgjjfA/Vff4rqvfpXob0i/UHs/xJNBUk0bvV
82KEZ7I3gMgva4p7Nof0XVdbsDWGra4AipP/qjDvJVmZZr62cLL7diKvVMj3Dwt8MQLC5Tn40UpS
WncLaZyuSWnUwm3URJg6qc+tbiDe0EncIcdSYkS2XKIxmYjGZEX7NnRVBx21kjBeB0hVvf2bT80b
fzNqurrYnCZT82eza0VN8CGlf7b2SpKOBLv1Z1Ji3h4eh7mJ6fyQIbR2eLrQ8TsmKPOIQpW8pl8v
G4krTyOBidUmPas4KC1z5OV0fYFcwtLSKon9V5hIIaFKuqgkkqahEAqze6UrdFISZ21fDOWotmP0
xoU9uRdQ8x88Y+PCYTrhIWkSfiXx/6IX4Ts5iiGYx1Qv/mGn4kKc5EA0XgTgHvfWa639+fHNSnnu
GIBKTpL2kxU9hB1RXAoSuIoCd0f8azWw3aZBa/dFdmzNnGvN7nSfsDT0fF0y89wx3k8dJ4jxFU05
lkyJFULcMh0kfgpLcAvskk+td8U1rrocSEb+bBpgznKcR3C6nJGxXMS21OnnsYxwUQO+ketFj1e+
Vwm5j1z7JaVSl0plmT5uyQfxrieO0xJ8huLS687+fEfyOp6UhNDEit4+oKHFNpo0PrL//0lOxrfV
AdwuLHTansIW4YFT0IL91xb1fgkHAvp5mk+s/RgCaXM/9FETT6H72Y8IEFrlpVRLCF8G0UoLJjlc
FhMhgohvhDtnzTvSKT5M6Gwjq11wEdCGpaNSg3O1NQZm/Di2n/r5fV+EMuW/O+TkVbwi0jcSENKo
Xler+5D/MHoWgKTFqVUWr6pYnsuRfi8W472r2A1S7zIiPOiEcgyzHz6/I26u9sFMllQODB1nc/uH
mKuVwKNbY49QUg46vTlzOpnQqOL0nDNS0oB/KNvPL+vJNqjce8PVBxl77JYibGJtj/jehp7wQCcc
IZXoYnTTNDgPls62ZtzUf9jYe3jMHLmeZcdUiHkud09zdz0qveeATXl6lz/ewT23u6Y2ZVB/w5QI
oKeWDLQ/Hy7okN/Ne6BUDh+TtkUS/W+85vVJQq0GBNWZeId/frlEsWtFuJiyBBaE7xF1RYHuXBjt
6TsDQs2kJGYFztlhdKOfHv2qBFbaCP1TP9H6DcdCwy7iUQrdA4M+ZQKL5tN9GQ8XTwfsXiP5zA+5
wp9XHmfRNE4J5nMIdqYxabAXdO5aQoXlEutY+1HGSwNv6i8mNvlCjiAWpzJz9HbgyizwRdj9124p
u+/n6IqTNOumegFWHPZmcyvaB+Xrk0tnBpzkdbXzc6tTqvKCmC9chtgnZSNEhweaSH4ef6ch5M0j
9/gg17e7R1d6TkTanhf58wt98Hqg/ypWuZZr8zlSP+C7wYham/aJ5cUQJL8LPWmO6D2AZc9Xt/qg
X5kkNr96ZHpGS8g0lWmeEfD+slMpzprZ1zWjiM6E3gsak28PA7mG8USpepvlGgDGw72KrNsORYZe
iAZsjjxkjRlPsFOy6x2eGQdvKYacWL0h1WCL4noHOiv9jNksxEwJ9KBI8ucn6jU4ImuPr0kgIl7/
0prNOwx0ehoipWU7pQMUu6MI9wERXYJJu8QoWTXhFZ2/N87irslK397F0UQpQNb/1lbbLfqRoQF0
qvjRnmsXmLbeaGkji2koFsVE/za0TdJCm9AnFayH9GqUayPvvxzIaqnWAj+ThaDtzelIwEapgOX5
4yCLYkprZTHPh02Ombnrdt9VEbwsGC7LTpnr2vzpYG0HP3is8ogsMkysQViOYAeDi2eUMMIbHFG5
XRqSX+gWtCIficNmkxsPokB9y/O+folahCUTw+FFFFlCqQHrS6cFx1MUEmxY1Ibjb46AOmUfhEgG
sW24T9R5MjVmzxdBYa4zGrNPqa7vWI+VnvrqVFqYYy+uXt6OdPIfOb2EEGiXaKiQ/ctmFYmAtfxN
b717CKg7/e4R0beZxXl6CP4jFQhb9VJI1PrJPTqXiggBTUdGPs4K5L4ooR4E5vtQwe7PC3qeVZ8o
feyXZs2Te2WZONxw0I0KAdnnNPS9+zMM460J/9hiDDCDBkF/ih31Xh/ViVlhUeFaWJiOd61EkzXL
2yVkhtAYthgc0Xg5FDmSjJHQl40JCT/2PoveGLXc8Eaawaq6xyJfPW6VuXXN5VavUrDWkJ9uL/YD
TwAGxiSVNs5RjfNKJ8DE9If0C4KvJm0sPa5GC+rqaYo28CFOdAT0tV9m9glgCG9SJeeooF2azGoR
vUoL0osvcfxJ0cSpEO8SvJXzyfoDXg5vvQ6bz6elS7ypC5vHantY0GeKZXRcqIVz6rC0iXL7k0Nu
s8vx/z6/5K2LjmttZnYwA8HM4TGMRPKq0Nup6g09Sqbb3Yuv1E1t4XIt7i4HVuPRpCAK+IPUTu+6
RuGHeHl8vpJU+XO9KEXXwx0s3Xm8KJS7+mSGHtHUXDsnoMWYJRAWHoiiNwE/35nSzb5pzq4bfEPu
rBZpKmjvYnuJJj3/iMZDWULlQyR5SNgzzZLv5wFKOi0sd7gQJG6HnWkbcTNLDo+F4Zy4MyoelVGv
RcCCtQQyt1i6bQsA9UPHVfLFNIimb2tzaFurJ78ooTI7P7lsKQ7eWJSG6GVO9dpl/JaC3AZ5g+vx
/hGqln3+W1QHpyvUMVM0R8PwKgMVV3xyJ4fDyxW4MJsNDtKo3S7qyFZQrMh6mH5QL7uLnalLpxJ6
wVeELiVV3R66eCJn6So/iLePPe8EFFW4/0cFFxcbfsAr/GOzu4Vw23MA71nayixym9p8QgR92Y/K
4yuYUcQvvs6Ksa1K2+RzxeAQyL7XWn9UXBcKh3ObjiKzObHP7EXN+MGdRXP6WtyoIB9n/GDmfdwp
yusH6sE8o8XNwtuHdedH6eoDkpfN6FNMvPjm0MH04AL5uI6xmBhHP2eQOF5uq9iJbSKLRbj8Lcpi
VNOEvwBr5zc31C6lkcdDgm007Tbjwsr4tNIpS0Tg0qaeLFt3//tW1sv8b52CyTSAsKdjqRwJamXq
MDDDxDROgHIN4Kh+0mEDrKwmfG6P5JnnwNm34i340o6QK86gor6hetUi8ePs6DRw3epvdE2Ft/8X
xY4w0FDTZAWsjutOOj/O8K5tsD+AS2jA0niIUabeKoXFqyMs8Qf7Fzu3BYspYF2RnUAKhr2hnHjr
h/9dGlTc8ZKc0BU1ur0Wm2NG86KWA83gzBwmFUzFtxE3NMV9qK6RDV+QH8zsCD3Cht5CBiLZNAJu
UaGw5U4k7BHo9lgQ53/mAn9CyyvxwYlgc1zUxbqYO+tovMq7jTJNGn5FMDt5MkT/8rnFEIhPfiXW
sn1mC7ENQJTIpojd111Ytd7QEAn7sK5ulsae1jQzEmB2oYj2yTZNWjIj9JTlzMFB8hRPEZH3FqXt
rwYmb2s8DUtEMQcClXTz109LG9ZTPjb6j7mzn0riwSpzCwQmb9744wdNYJ8z2pUGljIJzeXA4L+R
5zdzDDfTLoJKMZxHyyIANmUifzVhCBQw03Konnvy6QbXT5LSsoUfrrlL5ha2j4nNqcc8mjOdmS0S
r+8GFLja4+DiH5AQYy5UhTLAAPQDHDqBw1ciLRB/xGhmxzVtw3mU6BNd6Jqd1GipFzW+G8ImmiWi
ekX8DArAztYIM7fGZLno7REo5mdretlQ0nDGX3BGl+ukJoxyocGsr7Fh78wKGkR/hfnfKP95JTW8
MPv+qCZisjtCegJkaSBQMersblYf1Kfeh3e3ImxCuaSbgvApt714cbyBVCFKgTgBabmaJK0cs9uc
vROIC6WG0eABjg7h+LKccY4in3cnuSzEgXPH/kCXyuEmsC9Fsg/lDyhQo5SAbc7S+6TFS/59WeB5
w6sRh3SYR5QWk/cWzrqWeK6SgfVsQZBXvgtbZ2O/HKoyVAQA1PA9dRSil258LwaTJ1Frtr2Gec3I
mUXWdZAsMMnXidTULqsyxHWTfF7CxKxI55sS7buJLOvefdNGv+OJfbl7cECONGXFh/JI78QV9VK0
s0R9aUS2gM1ewqn81a91/CpDsfOvXZp1ku7KItB/P0SWGhUDM+XOdMSYQQVNbvdC5LPY/zctwsl8
//09lms2t5oozbuZwJTxG6H5synFFuDa/zW3V24krJSSOjAPZvUsJeqL3AVjiRZN4CDpiGu8dGqf
mdJQfJrOP7L+dHYVWCJkLRHlzCkihMnVCC7OeV76VU5snxbdhimNWzYcEyP0dre7OE7hjcusF4Ix
lw6/74fJqb28prsnRAoRsbqHnQfuW5w9dKsK2J3h5bvlnQKXnqIITkphusZetoKJbumIgqZopDoA
3+slxgDqouytqFcrS7JV/eIsDEKlTDCEVTQgUL05+c66zIvrZn/O7Sh3WpFlyp24BYg355hWsouM
9K+1D6mFgd8PyssG/vJC0f0LDsRxtT7LHEydFjhB7Olcm2mhLpJVxIisInhvPuQ0rCm/u6cJGwts
wrIrZEtM1/yCyqWNqbhZFea7nIgs5+KyocPEHoZMYZZVvRGRiWJsuhgSt6plIK3kKUsM2tiiW0mp
vgv0sd1O8sCmY1HPRHoWBnzZnnjQNGTXenkeWrKam8YYt7/jb7OzgGMhcntRF1ladnRxznxJs7G3
xsiCUyp1RTYTpNeydEz3UlXsE6XjCBtCwDssqMQ+y62OV9FdCLGNmniOXr/eCh6aDqm+FtPiAN86
LLsQWxylrXNedZeuH9k64ZwTrQ5jMihshdSaZwhOTV2nK5MpoUywzP7UYuMZP/1KyLNcvv46MKaz
WQIoD4gZyuK+Q8O8CJmSmH8EsqYgmEgWIVYaPIbbLHCtZY63CVb8W7vbm+zKBpF2E33bTQb5pVtA
UzDRLD6a0wwHvqCSaMFdKoC8M9ut06F2xWEwwiw23XXqmMq47wfj+ClC7Ayl63eNnHSwstFsVcjA
aPHPVTHzb3CMAp4MUbiXd6CrTGuJITcO1hsE1trR37JzVngjPyitXpxQ6YbrHv0awqJgRNFAu9p5
zcX3sMXzW4Ur5Vpnf9+Hdp/EdvxuNRPl6ZhxhkGBaWiYNSSAfcfEnB9mCqdSRRR5e/v9o75ykPpo
xUAqNeAhjnRMNcLQV1g1+ODjp6iiNeo0sqMq1/u1x2g9DeZnm7pCRJTJlF+8jghaw2cXqpWFslgq
PV0t3VYDhSwCs9hG94K6f/dnNP9uL2L9Hi0MUD5pn+Nroa2hP/eT2DNSbD+AOb11EQ9QtLvknNsJ
Q4Yv6KtvG936067+zvlCP9jUfQzpQoKuJ1Wqm/aR5vNRn+2t81rhahm1Y562LETTxcZAC9H710ws
X41zDCbe1CumtwsK+/BFVMkrpCYvhanx6T+F+6o8TuQ+T1Ig4EhZvJ1ct4tDwcUzq/ejVGi3rJhU
bmdi1zHdM9FhX6bqedoDMiCMzLI93I9XJyAHsLDD8dqCFZW72pcQNLTQiNm3MOMGjCTzMUxx+Tx2
DAfzFGG+SJ+1VEzmsmgMtMbGAxkceVeiVAfbPk+B9cB004W4MzFjXK0I8f2i/EDVK7Omib9IAPWt
6Y9r7UXB2vmtohLk967cMEyjpjpRRvz55vZKHjE/0If0PauvQb422US3rSQPCXd3bxYq6/cavZCK
g1lx++yOTGA11vwrslrBpxmoHKqGx93WcyJvmKMXzKelVyU0zr0rqehj6JHo3DVBuI5iB2nMLEfX
cqzruByl4uVelwP+hGfCkjrRTqpf1oEHCYG0jG42g3ceOs+Nx6KvGNysclF0wXdxzKnxCdFhwLIP
UUwcFW2HGQylRaLDHRNNgVjQq6t0vBw7Iaj83YlCBvFI5fsqgTqhPt5/MISUIxXtWjY/NtYHEnCt
FovZ/D9cta9ZlAcZTY7H37Q7uwGgJvQ3B4kUEApEQoIzj40MRqCLGHkHwBv/eiFOYf5j45M9eI4O
Rfga4M4UwgZXaFSbPsJXE6u49hOSRUfo6N3zhrGRPKyiyWJwX3ewlZMWzXyis/MOfdT0bMjFZIRA
ADvifylRu8yXwQw7Rb+aBY42AQGCN9cyap7D81CuDsC/nKhdQQ7SzOHQREbsMsPIUrWaw4CUCNjo
Ka/JXOa5p8HJyVDHDgZ+szoWyctTsBir7VnUjP3zWEQCqWu67ALW8qnE3FUYlv2p4BFqm6hvGk4x
juNL92tZoEc12dJ6CfWznRs+YC4uyeyxU3f/C5uwM1FZKZkl5Cqun7qAWul6huieWHWnPgZGJCqP
RpvLngyQAfqXqXPRjW+bTv2N6tHn6hIv3PfFFiS6VlKE85lef72ROJibcDkw+W8TkpM5YT6+84jr
m4nzxincPj3g/MAVvofaXSeYB8fOJ+qm4a0n0emdtOy9EInCQxTodtSX86M2+/HH+i1WGXU8db+m
NlnySfb4b70OD/G3hNe0MUPqRE4fDVykEdKFkLAsuHUpbnFhoplNBGKGjL1LaVbjPyX2SmyJuJjp
oPWq2UCzrshb1+jWZyXa2s/7ltIWAhaq1mkt6goyMCFO/LHcvmbc3BxjKliEMQ/R0/OSVPvC93rZ
OceXCYJ/Sn4DsMfmyP7s3jRuwnyR+PychHDNxvl01LrSf7l6Q8xE7ZayxXmYTYZr8f8aEcbwm5m1
BZcsbm9GJHVS7tUfHtNs4aNHHJNlOdM22/cU5U/F8nIc+BLIIl5Ot3IRxaZL7A+74ysOEtvh8CbU
a/l9nEQyKmKSmZjJgmS2CH+Qz4cnVMExlUrp2lHxLDHYZgk8I1rEZCzM3ak6Wc+AAXUL04OO43TJ
+lJLBEU7Y9Jcx9UsmpYcl3+usFtYo0kAysuhMMJ1sWPCzgy576Z+2Tz7fY0SJzw3ZPr16xGPTQIJ
y1QzBaI31dEdFmlP+gXsaotKKtOhCbjEGRlqbanGmybYKQnbBC5aKIBHnpsgZX33tG51Ep5j9YVE
VCFOmIDyH5H7fksULJIxvrBthwuXe5dyJDLRYdJriCEc9utOJUsMpQxmtYbUmmU2XisDBd3l95wL
WDyWLP+s9OsEvE7hiQ3gOm1ix6vETXxi0b0OOiAPHQCIi/Aul5IPpjjn95ppRo5LLR9o5gRetPSz
Zp7Wlm4XeNuK0h+e22/1phnwCkmQ2N8m0A/zVv+Y+sOUTceymmfy2qbhbiiOrJ9EtrNCxtd9DbbG
X9o5bryrc52FXm6QItzrCk8jUTfMa8f8pBTsLnnpXDPT6Hgtu0SbMs+hnSwoNAJsR4DrOry1CsEi
C7/xIJ/KHnYmNPOVGYKpRJsCXRhiEtgpOq1kLvGysjT4c9c+LB7R6FZyPqED5vrdIEqvizGmKAwn
YPFUTbPGx4nrZTymWQ6bKF83FcW15jhUfwAxU5+/Y2H0fhxSC0a9aHZB7IpKUIVufN9UPTNN7ieW
i3HWAFNkzWFnTwXExM+Q2+FRAPq5oYpUZofhDK1MPjI4yDt1dt6sr2XL/GdlohkiTSX3dDPkBNoP
0nZnTqpHWmchLbb5fqoy/VPiMn0uwgRl+ShB/qLWzeqqJL0GiDHkwAJvMWX4Zr20KhKjNUwe+Dhq
5nXgMK4zysS14HPTcOc9O+EHseWFpKQ3CTDGCz1INvBf+7l/XeLYvjZ1FiN5sRvTsxdD+Xv/Sxk0
2ZoQIR2g6KLTGXj+jiyETCP2kXHjXuRUqBplMlm4fNzUjoT9dsE/EhD0q4iTCrAMQB+A/cIwIo9E
/hpvqU71pvEU3uxavIpcRjO8aoXWvmPpf0oQwG/z4kJnHN7NHT1r+ej3q9zfarzQRB2QcyzAz8FI
xpsenA7IDQzZslHd2VqZJweqzCShBKhRIvikg3M3+IrtBjrRuQqA0BzbtQ/yDLn029P276yz2fTI
I7lhxhfaJAjdOufTPOMhuNkpnQo7dEzE0jcfWgUgKQiCA7Zq7ASOfqoKICKFL7MxJ4v/PPqBOZzF
0lkBoE3zINop+n8Nekk6ItSZjGKCFx+u1HW0OaVAq250k4AwNzjh13EyByxcz/FlMYSLN6WEmvTJ
SwJ1++P/rr7x4u/mLx3J2ViFF2jA1pBkhY1YRfm8sNJgaFds6/xQd9GSvw49mz913DYQ2QKd+sk6
JkA3rXZn9bFcx6vOUSHjYhFIoGw7BwnKAoCKj2J/0fYBfDipqaS6F17ZGbWfgEDPHmr5L8NZck6W
8nJdEuUJ6y5/ZtUB2+JmNcR3VeK0+xJSU3upYEuxobLGc7M0ISn1Cmz4rsKgy3xFMoi1aDcD1sfO
r/ZGbfsVLVCDpCN+WbY3QiVITAwoNiHL80eK1Zd8XRWzhdR4j/ngNr5NBmFwSY2ytf3SP6UFDlsr
5n1Ym5WOX5rfD91gnQ3YbVqApAyuHQz/kdk/HhNzVJUvP5OZgjjNlCtQiXp8HyJMOjH/vvU2NNzu
Hf9/pdETLIjc3LlCqUhHY95Uw8IS6EQWGV1KFk+2s7GJsET81hZiLnGvhPnzLOnrQKelVtEJuau0
OxPKz6vOWZ2+9r3Qi5IBg2XmL7hRG/2O2MWzS1iQp6oMGrKFtYk2RwhamcF6Hylsrm+srkCTQZaC
DZRCyQ/W92f9kIcRCN5dVet7QxfSsUcNzeZD83O00CANCt9DUyI3Erx2V5So8zvNLYdYkfR7NWd3
tUKNTKgHbnVCCQM9PA8TC2UzzCqTdJB+ociCR9KrnPCflxSdvn7eJG46qc7ioSfaMH2sUAY7eM9t
1hkJeuOGv5EjTxSEgJPwQGsX9QmE5QKiX+GVtVY6zJU2yFHoZL2oeb9CQCwGH4fyH4t7akfFx4na
fnAa3dq17e4FhACKU7PzzieWH51/H65EiuTm0M67IwdjMRX/UYBFM4X5ODVU/EnPhRZSczZixizE
LZVzRV8/v1lXpgB41cfwsh7aCiLfpTygJNLRuTZRP6THM9y5XCJlvEpYf2y9w6r7d84aU6Ezpa0m
ri9KNzCNA9wmhwrbDrYMUHQ6c3duzsIrLX2q6SBobWVnsOwnYB20bCSvQougdb+CApOYNEEOb+g2
+6tRRDabChtG/LSzniWj3fr0iEeeKaMOmRIorojyC1mbUpyiQn8BI9co9xeBZKp0Hj491z12Ijhk
DijWmwM/4ibUVEJpLqsH6QYsx0A3RmG1Z95mxrLRKNfebFFoSm3O437rg8nPx6X96TiJEwMH64S5
sRUC1cgrPOV5BOahnd+vlhxvu8Ah2mfl2xu2xii5m2FWax7tP0P/qgJv6Vpz1m8+g03Otft6wS4x
NUaZm4J31/g/vt1edg1cFO9brpAKA2vZKTpFtCJG2VniA0EY+zk6ZrzUmsVyJ5BtEPwEY9xM2RLl
x198w8mV2d3pNVe4hIPlCRRT7Hti+JNGj0f8BHmL10CPSjST93QlC6D7zfuTcpwUMEOBHMid9By6
8pbrZEoykEFh8mFlrfjnwDXPXWNDNUR5QrLI5HZtCOT2xvQoOr/Ep98GRTiliqhWAEqDfrhuGRpq
VEus3WjAppjfCHzZRwgDRLRHnB3NTVgmwUmu6qop7yJf5Tke2eMrStsb5WwUp41sNMfG3ZtSR/Xh
nqn5BNE0p4KQM0aQ6pWfie+amnkRjw87FcW+Rx4IvD3Jh3w+Qq5LyqG1O398BD9TiVGvHRYyIHpf
6pCUHuOucYbRnpacdV75u2GvP8TlSrhAklrY7NmgmdLiMdduob5u/K3jsOPuLwVyB1cXRrEj5CfJ
VeRS2O8uxqV/9ijO0nlbdwdJPNFRBCGwcpY3sZ+qov9BxN2664SG9dmHb1zZCitduiwi7eRvn/bk
JbET7rCOy+EqXpyS9wgyj4+nQZF8RthLTX2iXnoCdLMo6s8K7SDWzHLKJPaukzhHr5sPd1xJPO7X
s4CIbakFKpsOcDrxUWtr5Ms502fpNUOdaIb14Psrq3uTotEE8Xn+dykf8RVfEfJFEGk8/ggH9zTC
3vrbxRWTfeb72wuB0SDSoJeFV1hxHWUWzY1QGFPcOZVYcA78iCJTuiwKZ2uLM6THz8+Es/k4bC0U
surRKEPgUbXANhCzzyeyYYai3C1X8Osg03ygWWKjlVa+AhaybD0SiYBpNIoig/U2fKgQ8mUKL4R+
I1a4JYIwwQc6hoj3pREjk5Ae52yjk7CQGA6pkzRl7McBH43Q6hYPIaPmOyMP1bTsHMgccqTIWrlC
n8wc2/W8gmyxxZE611cQfe6FFjA4sku5GuPiwBgBZcWux7dfbYbFOewfG1zhkdRgSJdvu/9irEKO
n+UjgQefP0aRDFL9R9WGYIzwz86QF76kBN81piOSVs8vLEFZ0zVsjTbE/pBdPIhNmUAN87iQmyf8
OYW4G9tBCwlgsiZqyEXgDea7pFfH8R3R9YdDzWh/Ld9DYA9VPBVlOyMa4unCJCffHEuYZPHSgESr
R6mhnn5O17llyYB7Eymg1KEP8og1PL+feClBroFRPVqu1o/gSVgUYbJTve/xijRImk9Ngs5olpOd
zQoJiNbztmeUII6QEBf6fiFQ02sxKLG2qp0VHJt3HeXyez9Oow19AwuE40qwtj42xURikRqy1evD
Ldkdo0X49IyABBiDOu/pqahkmP81JWDT5GNC6MHsc66uuRwc/IrzRVfcqkyQB3q6hQoGZbhRrlaY
9fjcDmu/D6t4VicC8dxN9Tguy16zJMd/+aInsfCZN35aqaVIzAHQPDVBpB2XnXmZAaLdD/PZkUoy
+qoqAqfrvi/6rVGCcF76mSdcWHKav0E1RZxhieznUpzFhLevdRsnFGolq2S9INaTZRl66WAr/Cns
epvotveB4puwOEixpQceyjUnIk4sE9vdW61xApOTKMz3YD+6EuTfMcfpJ/tbFsrXdiAUC7K2+3CA
EUleK/XQztM0LVe3lSYmIFrz2NnhP6LG4+n4gK+EJwleNZoa29zdC899nB3z1vzo5Lrq4H0jth4v
Icx/YqL9JzuRBhObIGgZQBsi0WtOBv+ytOJnEY5gKruua4xRVARYFwoKMDBLii7yIki5QxnokFH4
HAwz94u+UZhD7k65Pffmyh5kF2nWOQZyZcMe21tBeeh//3ZR3izbDkeB+BOU/f7GTmUnNWsf85jn
Es4gmnAStDQC0jhLAAYQ1u+X8JE1aVF8PXTTQFeX1EOYvTh7/7OCi6TbPgvAsT4EE4mSHJrXwKQT
ckKHUXOcKVhQDIVdlCPwWms4Qog4z44mIHW/DPCZQMdddXzBpcThHDKQFq3jDNZBFH9YnBGGbSql
00+ewDx3it5EsLnhkQ/Yjl8B82cdZpFC/E2WZfp66mitodeajEDOFhDXLKHnZLbDrmGr4CLhCv75
nImChAwU9bL9sq2pICiC6+Q8pvm/LJgwKYOeSyLa2iagWjMFiw8EkWRC5mP4svqL4aoWk57Ct/af
+i0fEkrXbXqRRRp5wb1hg2C11t1w1izVvvBWiXCqwrR4PdFEIxkANX1AEchKMAWQBlA1s6rXv61D
CAogPrp6GQqnJxlkW5+NBThjdKCxcXJ6yI2F07v16YBD2pj6YDXSpHreHLmlcD/k6MqR2T+0ptYu
OQMfiqvsJravlI3bPyb2HmT9DlPvadjwq/VnHWf6mZcRtrlp1lvJaXRdi8V8VtttKxH+3jaayLGy
Jv9ml2r019m1m7OjH/ZexI5DNV/p9A13bhMsTfaH6MQu0RJQBSl50AiVhwdCWmqlDJ+lK783ES88
W606R3vqCY9QqAQKUldipazYRpzuwvCOLWQdHnZJ+OoNurvsx4agK9vW7Ax9TJ8nRwRv+/mG0fQ0
cY1DOdkfpi4dLDfdOTkTOtB0np9RAzGzvhU57syvdTaIFDD5LAEXlMfmbTlAi4QJULBFvAJmy/Rz
1cZfhzbanyapeoVb+HzurmyqbG/sGTePjXQ2OOQ/PfYGl09FAaOqrqThl4RzR+emeP1YdALeNsfG
QSp4srG6DdRGqNQIqryGIO1gve34qVkrtrw9BCl9yDBUtVlQQV/kLcozsDN6F8Zapm3Sea1/nkNq
WQa8Go6dlWplUUPi7QZfQ7uFBfSgVfVmwGEpQeel56C5LkLTWXYQwYvrunMtw3tSuAImQCS1NVAh
SmTTLtagr+zZmAR6auCNASa77xVjUxGDbAl4vKsCNaBue/ihTO5sz8uS59MR1sUxXVzbHYtMDLJb
IZFNBIL5eUXdS3/kUqhb1TdVRW9BLdk5aUkpyrVudPxJ7ZJy244cavSWtIJTOJ9G6VUhlp5oB8pp
gORpFU9N7euIPgOPquRiSKOU8pUAnyoK6izekA92QKgUezde2c7eVfyTnzrjiaxH7Eqa9iHsWCQr
W//YOq3M3UOouj0oag5x3k7C9YyZLu+ZbS81KMQFboOfQp5OqZd+yZyMcXtqmXWua224pnKLEwbf
eqoH7FE8izc7Jagtl9xL2H9jbQEx7ni7woiqKik1xZOdUH9uGfQDKzcQRBAUDStr+LXt5yBbpMZG
WkqKtMZGhlzoZgg/CHdfT4aBstgmh0w7qv5tnIIVjoLpjN1MCIfYWaQtBe4aDpYezQjeKIwjc8gY
FXYYpnblF3wyT1kzcaQkHM3FahG+oQMqwjSaS8x07aKegqeozmS2cGSie68UnDu1pKe9CEFYb9+e
nZ0X229gKNy6JxL4T4/ST5xPff00W2r8G4/Lq0HGJcafvQWoTN+DIvhrHkEPk6DDjlylwt5pU/kR
M5a6XIaPiZk6MgUptGxP4sVHh5T1I41IgbnCDgGqlz9ugW/jiG1lk/bVqvtVzvx9GNY4WoPpBTpq
IxgoTN8AbJU16MG8kkqIGJlzMxNH7AS/E8y/1BDgN4nSTvTRb21iBFePG6mn3nV2dQeBLLA9Dy5f
fmK5cJyBG+Q44jfiKsM2PQw6IkOB1hVfOgtdL2CvxyIbhx9YzQ/uY7vRc/cXtp7nwTCML71Y6wSg
hgYMsZBw0Be9ddDDFGilX9bT8aynslAAmFmXSnGYPaYw009m1NYdZwunIHuvpRimD3cPow+k3ECa
jMBZSc/iyqDhP9K0Ekc+l4eRNhbO/3jsK+TKiVW5aJli2iJ/Gd7jDmhqJN+H3GIOiwscWFykr/dx
6iEUrvQTpsg35frvVDUnr8nAZ57xyy81Iz3rWpkwbDM+FSNyoMg7drca78eq6U4sm7KJ3K4Ox+il
4e4n3KRKE6u2v7/QuwvGUBV7Fn68OdaqTsE8YhnfFKKe+jE8kxbbiR050suR/3DnkU8FGcRlkcBd
hN7fsbT6RSh69Cqq0fB8bBUmhgYIkLV2ndSaHWEGw5gOTMK3Xurn4R6UjZsYrrjh9lMw5rrchION
qd31c5ftFk/llSiGPwhCuLU4QIVldkOFJYhArpMPxPKsl8aES0f7/ATPFI6Lw4XkCJRJDvNpF0z5
RirF94zsUkOshbdb23NhTD4Eu0r5ZzX96h9wTDYFMCCecGZK1hpzyv7FzlbARGwKDh2vaLkLQnv1
l2ZLtzYGAPqx59ypj0iNnAZrYn9MDmo6i2FT2hFKKwvFwNYGrPkvQZuH+X4/rbx/Jx6RHSULGP1a
IyDLQAqQE1OR10W7hOh07Rs9JJBLCji+o8hyZufLbyJWrSgXZhpHHSfWPxGRKAYBEzBhZp621id5
P6yeDfdkGAj7U/CqV1rtLsXRtP9jiwi6W1V4LZTKsRmvb3/CwlDkgC79FOrpOGiCHF65UrAo4Bj0
ljhfP6p2aDO0BDU6aSL90wKrhNJ3lMf4OVu5/k67neQemba6jVxoiSYgSlsr3CnOigp8s/hl6DmR
9gKPVWGLy8iVg2ags0r+wzG4TQF62ODIg/w/+kNJAFF/kMX9tBd5xQiUz03dSh2XSgZVa+e4TLzt
PZsBU+Eq1X5EVkCIE1/lY39+mO1BJFupZ7RyBqu6Hy1TBtxzEWN71QT8c26WKNe/9Uz0JpP1qQcX
H9rhUL/nW/nvrYnOV5wGqtg2HP+45l00qE0I+gAwfZrm6E1UKz3lrEvdXYZLHpKtBCrZ2Vbjk2LE
dgdLDjWTVZlZ/X6Sf2hpLsjRadedTcJNfhYB45RBFUY5kFufsJnBhk54jTcbZdVmf7ixzk2U/HZX
p7vYSdrjh0Aeji5a8uKMthu76ddtT/Y25y0gSRP87T72kiNexfhXGGFpyek10+qqkrIALEcBd0gX
1do5xgM8KiC+tt8zILDkUj8PsUs/a7yvQ9FhdJQ3ISud6iZAjtKUSWxRWrLLj9UtUZY1bk7yxVpc
oxl4kj+iiktzeFR18ZEOlTgW2Xiavv4mGzD8Ea+L4nwbMG/tYdnsDmj5FZy0pQmZDdE035U8dWWn
53dpNgrMYSXrniLwh5/6GNdokY/zhg8cylMt7ZgOgzucyD7F4EA1o3LLquS81TM5FaBtKmf5GsWX
YKakDUCYrq53t4HYOeowWdub+VjlXQhWWREvKhtg7aBrnoos75kioHXYwAZ1PBTJ9ge8WE1YCRS9
jJcQ+g8WLIfaLuFT+g2WKnXUoMqLhUCw0HFyTG9/hPQY0Z29n1X3jQJxc5umeZ4Wwd4GXkOMKReN
axpz8IGdIA36AB+3EB6DCBbhaYIxoLmoLmzpDCp8BruzDMrGbA6Y23zagyr+S+P3WVdJi1g8ADAa
EtNZg6fuOBWktJLiPZRg/xjtppWI5z0fd3mKokgik/DvXcRBG024jL3Duu9KzwRdKAXREldQoElj
2wXVa5WtJ8HrN2yK5uns98gB0IHvoPPC7yhr+qIfWUEIv+sEXdgCVGwBlaghuUDKSuAj/QX6k/U1
Kl2divgixRf84F9C+ruTxRkgtQ83Sj0XBmoC2hzJAb4aFMfXSUJ7qnpabkR631026jnE+qJ4UAci
TH4zrGsaStm9nLb0Hl87AmGzv09aTD6ddBoXGqTKi53kw3hbDniA2Bar96DrvQ6PYPR2zG8rDWHW
QWVxCNMWTxz1Eje5DIPa/VcrxUDbgkaDEHW3VPXVzlwk5P0gX/1auZj2TWsWRZ1G5x8XzFDUsMWG
MoagdU0yKMpFIguNIyWtjDJdATNdBFLwVUGiIALbtL+2wl9uXacP1/8F/RRwhqvnpAQnkEV/y2fX
7Wl57OFlniUhVlTTGACgJN7SA5nr1DFm/jD3UlqFpLMsG/UC4oYo8u0FJ/VP5ulMDYeq/9e/k/Im
TCUawMaU1rErU+0GSX3E3U5+TjRcZmc23JXdpyR9zA057PJvE389Glurmii+llqYJxlmN8MFfJXW
qRYfSYckQmbM6NdQvbRr6Qem92GQzf/DO+BhM56sm2ZqWU9Mgv+3vB5eQyT7wwEmMCdixGL9SGyg
lREZo/36GBP4jJalWV1CtwEqm7ar2Q9jHfLdgdlZWGyHewichkfIgIS5YCGBSUKlkLFCQY+PRuyT
1DZFaNP5LUiRU+pSqGHyCrLGtT1NazS1eGQSQtE1c6KYPyJpS1HuY7Wfv2rgWxTExEyihZbHWBMm
mVE/Gr2imS9GM2ID+HmyXPcS23V3OGLp4RazwNM3jH/zZB3oDzMEq9C9q/ezk7wpziBj9+PLiHzc
P656ILLQRlDpb1C4p6pRP42Mt1DoryLvnBMbzKoSZJNZxjVt311TbISq43mAp/wgqjJCMxzi6VcK
lSnC3EjwECdevLduAbkWeQ82ZPpYj27R2/G+nNaS1z+eWxVjkYUeLtTlTLTr3Abf0T3//V6yCbqN
zVKkG3qEdj2Zc6I/ODtoca/e2mNI+T/snRDymtWDG+wSgO/6zsrOrOSEMGx+Bysnec4pG4znfuPu
JsnntfwvHeoo9oBA1hTsSvE2VgehDL6KecfCWl3HSvDEQBjcw6+lKqGmtajzqpfqoywFwcVFyZAa
nr6Cdu6TYyntXdei0bhtUH28efpsx6j/eHOb1j8Cp9AXvqBvdu5jCL31bczSbf6q7vyXO2kmVWMd
8CKyAAxFw/dudYWcgK6a+F8+EUZUaQjSuS3KLLHXNds31rl5kgXpOuL9yQPwY48OJlesMsGxclfm
6K8oQ1w1cVskkzK6ULawnuYKIWq6xBUHEOgh5YbvQ1rpniaa9OqmXo0Is9NgjnixzE+ZYO+sGhZF
AVKjHxmTBWOMuJjY/8GFdERtDgRYm7gS7Jm2yeOLsakeist+ZTeY/2sv0J2g82X6FXr1UgkhLU/h
EGd3lneBMEMQIgM2tpEK0CDGL7v9Sa596/CPLisGMprIwZw5WtAIdOdhewMJ9raMzKpFtpiU31PO
Y0dVXb8ffsE0+Qnko8XHnTgIuc6dMTWehmYMjT9clJ1chSF0CO98qmX2DQlnad8PuzCvJUXDeboe
xFTY8AIe0iDdgH91Q5DMPY4GJBnZId+4vmZM/evYjGb7n5XKXk/a70gXDhMjUetbAj2V1tfr1Nw2
xBWcCH/8bIFhH/qwgs4i+/yMOyyZ0fX2KzZ7iPRefhIQMTQutz4oBJSqZcSjpf+C9BwI7pipqPd8
Cz7MXfxR2T1G7r7W35HEcUzpwtxWhpbvLOlSGY+4WS3wu24lT5naN9b30YGb8V5tffEZ9a8lqpVE
ALxb8ZwL51cn2olnzs1y6+YMg1p8jBRU9zQr9vsdFiNkfNagVJQoJIDRMCN5oi1nBXD7OyhF+pYx
wDkrnGtLGSDtRBKumZO0RPLp7TfE5JNS870ls4XZHoiOPZUYcIR4C6HC1puyN8o6qyyF5MSceVIU
oL5TxM2NTu+p/X2ajF/ifYPu1VP4AFFhVE2QDgwYa8yJvC9HclKG8IS6NQq+KRYEXgbRGK+VfR2r
bl0tXGrWfdNYERGBTk8uXMZkhZuNXVyIElzyQo42o7hFfLTf0WPy6QOUD8WuE3lKGH5HTqyX1YO8
7V5WxqBNvI0J7gdsjVGM7zy5hogiu/Sk9odTQ5xrn0RjyNivL5EayS/+9R+UzxszDG1Ovv2ayatF
AyGy+BIA1pySXF9O/xY5h7Qjks5/ITF7hbJFuK3rOA0rPHKcze1NyEI9oXsAtyQhE6LGfNAW4WA6
Ds07Bj+vp22ZS29JsO0gJQWZS+Qy3fqN4rDfBAnP/uTl+vZ+o+g/EKf1oe5aMpBPjOsu19u0kHYG
IkfGx29qlRSOsDBshtZ1BW4BfJo9llH89e2DKqEI/pU6uiX86hLx3MrTIBM6Ks3eLtuoggRCol77
eqo5ksv6wbUawqu8B0rQ2jgYFlUAkjUg4gBRLZ+iXWj+yrLeU0u2BJFc/Dnhk8BeFpbs17MWNQz2
15FuFtcqArkQthRv876/3IuwJYE2t/0LwNAWshfpPD4qM06a3MgV5zsCMFriMFHDNe4hU/3Dngm+
gqBNEm9c0ViswAglTbjaiZKk5e+hOkcTr/x155FwIoNHwJjnv/BFS0J0z33M4suAroSQEc5Cac8e
CQwknwITuUluSLRhi5THmt3hWX3J5QghO9WM+F+HAp9c2SHPsuIOLiNl3VWKA6nX+QlTv3XNmvDb
gjYdv9rW2tH7RN5CYvj1VV+M9ee4l3zmitHsJRPLAcn4PEbPCGjOINPaF6p6sLjiuBJgP6D+w6y2
gSHq4f4dBcdMmgICsGjLbqcBbC4uH9f3kHZVxpre4+cbu3OcQtqm5/h9zIrE0eLmSmIKBB07IZ6G
eOmiQZy3ATKy9Y/0JEUgm4nb6aUbf2v7CTNu3q+OaI3gRoxJQrKy4oPI2FsJVBSZTNa24l6zKOBT
URSUs8pNzxrcT/EJ//qbkH0EK4t1sj2lShoR1kQsFRQQEKKzJ0q/KhndpBOA3CrDRNPVtfdDgfBr
9nmuHVTFZJYEbk1zuXc8902ky36+duoSa8w9LWDXZLW8WtUPhG6LB8kzXjEk3ge+vodhFpKM4YVX
FQ2rIv1RCQHAokFF2PQosDDqm7Gv/SY1onZXu4eOS1zoqtBdMOa3ldrJegH7ft6Ufgs+XA9Zgz+o
gDOdXlNY90zOmiSR6SHntrHouYhBlD7kaaK7UmvZupoULch7ndQvvQh8jt/rVqJ5SHihTsuno4Sd
7eN9oAbbqyYZEAn3pAYw0NbIGpZ07JX5dYs72AQhoPmu3j/ti8Vddj7roilgmh7kT53zxy2XfDX+
NQv/OMy7VPdrwQgyjmMN4lP6VgZg+WCTyAg6XeWms4LZ3mRAp/IObl1zrgYUwmrcOo/Nr8ictPh8
pcfYn19jnNvwCYXeeBhEbsSpD3AEw2fwUXyBhHb/w4pBxBFBDmDAXok9UacHvWOxQEFtoEH1fmhS
GxYXpY0KU6t5BysWQePCKEJpygco7HRR4UYECNVnYVn0eFFLmW2I7uJlGxzbgI5HbhoonAqJFR2I
2ltdD3DY2vwMOtOvdrE03cBLEAaIB/23ch49XNvQmmCpjLpSWTJurhGkdm0nrIqdmr30teKHVwbW
M8jf5/2yHiMUjG0pHGUS/9zm6u5ofXvpSuOEoz4iuLRUjoOxtRIchZAqyg/xzbVMsj+nbu1VZ06U
yNGELRZ2qNVvZ3N5A9UkAem1OQDsvQO+B+lFFuaH/xIw0ne/AfMzAfd33kQAleMlNZV4z++P3tFB
PHFxY8B5RpEOhFsQ35gnuC4DyOfmQapIAO75VVln1c+PbA6xEAtJgp6neIe425OdF84v57STsDzC
a+8Nleo7KojO7S0GI3O+zxBMmESkr75P17qVPEHffjP/SKey3a5nENUFNPluBHN5yxTYv2bR8oxX
xPQLxXHiaRgtHddbeqvQBihy1Cijg4qVuhsc9+NCQFqxIvsUzOKsUmjuJWm8oEhOLQS4HD1qewq4
VVYMkf78MSgLtV9HoS6e/lZvX14X15itqclKLFIVZ7mgVOCZKf+earLB6yX4HD3R7akq6AIsUr23
IoUJbzs3RM55yUOT/v2lmo/0B8XYQr0Ztu7l4UyhY13rjzmbMII+mVhSBZGBE6OJI9v3K0ebcQrM
NRtWySsrxDttEFRKckY+sJu68FO8/qEfOvmdW6iCJcy9MDfj9boAak16MO8DuL+wXjfVD4WGt4sa
FzAVVQ8/8nt+n+B+C9LVg2FG6I7ajBJ+J4WlZDlVydF6kI+LVFgnWkSeFsr9FADzv6l2R370soWD
dH8nsDBn0GBTeoNTc7GWzqXyqmYFRgCs42v6sy8WpjXntMmNiS9cbycGaVATGGbN0bDwwZlpDhCs
6sJv9/sjlTQXEcwythMu3a59IRlsWdTUvFnK3MAZi9+9+tL+UJvRVV9jxXL/Dfz00Pvw3VekveVz
wzjeZVUpuPVoOPvBdp1A9Vfj9iuzGrOmd9YlNlAkYHCajk0AM/AVhOy25RT2AFr+oI4/rr7ZZkSz
/piRLubv8FPbicLG0sN75VA+VYNPfefzTt+T2C4kkeDkjhPYzXjkwX21o+lIcd/LmLH+u+zTAFlm
ysImmnovtpdOroH943JM+w7893awQrsAh82LhkqgGgbPbNBHsP163tvuwbdUtqKFtg2zydHcz/8o
Kg8jC7rqTUvEgWnOEnxAiYebs++FLB50aakMuvQ9RAhHL2YecN6v3VO6Pe1R4BfcQs2gCP+zdQS2
Dfy/8hTjE3HDgo9guFzq2gKwwKbEec6mVDM5xiklYx8dCdADRY6wL/P2oroR5R/nixkzhvhkYSQi
cuihgUuRoKBcb9srahhd2uENXYkktn1gHl58tlh+5jkOLih8DHYi9aDnU4TwRlqF//9K4WdDGaEv
00kL+btVyrEPG6Wh640E2w+8Qzn1NKlpOpMK61JL9OCbbf9BUymgyw+rd5PNfIMNxmppbx73xgvv
E/pvcZOhisYeRE95QXF4BNBkzcW0ezfmHz4u4M9Py4Q12lJDNdDPAhXOTQe56lIFnqG4D/CcEW5V
FAAua9vNUO+522R5FA9lczRudQpGSbwSRd5nfFeOPpPz9yyugVqYdWVycvv7Iv7Ge50103S7VCTS
2QSwCim6e3WYzBzX3/7MJNUULbXhpuQr0Vbm9+PsoFw4EHYz0IqeOKdquUZvbbT1Ge5qpTl+cru4
dHagYZ831wnW4Z8/gyOpl4fgS/huhjZBPxd7CYAFYVnxQemg4K6zVLhYy07t3KH7Yzb5fKWOJXgu
gg3Y+OlSBvWfd9IFlP7bQZ9AqCrxpCQW4oQ5zrGuJb0iL10a22zoCucCYoylBM5iOE+brTtyMAwh
JUSGULKpYVChPwwRZhI0sqhO0hYyyq4kaih0yXduZut3MEtE5Akkh/jst442hcux0yO8DkDN97Mj
yP9oruVtUB4uTkWnFJiXCZzG6dQmMUALaOWTq5rTIshimIquCxQsusEjQaJwosjytXO4azEkesHw
LHPrPb7O0CXlQ02s+SVSz/w7H+zLHzxNZNB8/msrvZwr4zArV4zZ/5GRH87nT7uEpUVy+TU+Vnw1
q9+eYZy3rtyZyzAAw7RyvAXI/uzlog18ZWNGiQxfNDTpX5l+dsfwHV4GujFl97pKWkmKD5I3zFFb
ab4H+DejZ6OcvkBXvlhQZfk5Q7TBSg84ZJC7CZf7nMZuwvR5T7fHfUhBXpJ632c5De7fbxFoPFsR
TMWAsIDzD3ftX5s5VYR80SqGsEbeO/WDWZsIU9HsaVzbFSWPXkrdgEBF5zP2H++glBZTIf9sAqVZ
JkZvJkCG2FyHAZ79SHY8B2ipXa4kWphhfNGiQF6Q8r4Z/iDWiHEbsr+E2zmC773bQkUCAwpI2aRN
nN0n5MFX2LWdSIUxMRh5LPYeWacM6WsoTtG2SUe4L1CqIKc+cfpBjnc3dZX162VREXVLVjX3tvoJ
/wq5bHU+/YFhJIc7w+LgcetK6PpoXrcOHFpG+85CaULLYh/tsv4GEr0ev/4Dezuz9QhN58HLB015
Cy3K82HyXieozQSB2j+YRPEuvc4H232FAUcw/+QPMOr2ZX045x1OzRcqOQv/xYGAKGKAI6cJ7qi6
fLs8ZP+R/zmzMCL9RToM5FA6yQG1O99d9otOAtI1/NNI/Egh34NBEip13oQQUmmtPqyASXNdVdH6
N7MLiOBC7rVrp7YG8kyfjG+kylXAHJdQkN1WxFLwzwAG8t6zerKROYj3cZfgHSAYfbjD+Yzu/UKq
HN4lAOJ6EJ9fRYxbTviJHCF/P3/rtUS+q27bXAhZEkjCL7ILUTZ7Mav1MD883HeWI50U7/M38K6F
IdZ2DKaIz6jrHasNQAvPhXmvjd61bKIQMRrYxQRut6QpMuq7GT3zyqU0rYutK1Z5o4PE58DV0ubw
7v3R1bYAj7vfVPzYfOqEoYYKNTSeUtYtE7BmOUDhn2NYB7iRQ5ccAeGhdhc2wZEyJjFF0aMw1q+x
vI1ELwK2Tjt7hkXkkDvDG2icKCNUMPG4go18Gml5MOv0NKiWadjmjqRMYyNvzFZOVsVMv7HzTEob
oBm9HOQDDLaJNnNm84J+uRPGbor4u7FCqWrfuA5SvtdZBTuKRYDjNb4XE8DTpCGBP95FLGdkFjc2
Limz25RCa9peXkEETneIrtLHZfznAmmme1HrzhbSn5/wSu2LN9BOGHT/oXHvJCeT9QCAr+zf1ia/
6O6e20Y9Q0h1XWeJ5Jqxzh4j8LcBUKltMtgw6cmdoA9fWoyI734eIUUswzB2zhLY2RC2W1FhJxiH
+0SCyOsPIqKPpfZKK7HEZdE9kG3gGdbSu2aoiv7lUlshCzhDmULjLsHkB8ObhLQo3gz8muyhxuog
CHrHXb1td86Cb1l5oeNNqHtMTFzGHKAz+rM/9kwlMai8kSslTMaWgyfY1KHF+h230HF1NNGZ6gd1
saad6+LxWwPOu599kICFprr8F7+IW7gHtskqgXjxMFSY7rEVXTmklMpWBsFW6GtpQmzp6ecb1R5y
It0kD39BwsePHtNmr0G/KacwZ/iLomTwGAaI8o6OFzG+v5dG+lMTuXCC/pk2Dr0RGKBDwcL58hyp
hAQ3HNXNzaj0spFlkESMEq9jnYanVJCYgQulkQkt22YYAfQSUouwK7GaBMLVdMRPzrLdQval8nsi
fxUvA0WQSQHuZgIO4vXIEnRrnTUe/l0Gi+VwWZAT4pOlghyd3peBvkI2TUVosg42bjMHFALJMEeZ
IqLqojZk3kzOeYzIpD136sot32wo2s9zdpsAjjpr/c/euJNPRJ23DGbZ4+cJqrQ5p/fRMT1uOJcZ
vcYZx8B5ocqdbgnHxujHxSfLLhfeRADe1BsrMjGYsTzIflmtCi0BAiFfycFdnnmOmCI20ogzNDQV
4FS+wUHIlqDqRC4TqSlw/gxQ0eW9q5JrFiFW5MK2wxIkvYl8YxBarWZF54h5DFWSZ3X+Guh0GvJd
ZiAzOO9hLCq3eQ/aCqpe4sxb3NLzx179SVJK5OCq+LRS+EiDU12MgezmBMF5GqvrAEmlI16fKOKj
rfU22qRs1dmv+kPzyCg5iQUKJ/3fLrqEHW6nlCUg8b+pk4sHQLAJ+5PARdAewXBLePlTbwmnPCJs
+aBwD3fYA42CYE5QEt69ObBocqWPwhGMDoIU9rYc9Pz664ygq6zy0tePIg9gUiqmsCIjHAqGsIla
hFlufCS9ABkqv6BPQRMpVUeeLoVMOl7NFz3bXZ5cMAwpKg8D6w81k3R4g/fw2WFTQtJYZGKVqPGi
DilbsRvPy44iRqylBaHd9Tp77TlLO46Hm1U7OjZy2WdGKuAzzX0qWjCb4XMzOwhAaylmtzZHaLK4
swGoXP6hWEdxK81SbtGJ1v2tVO+0yut3DQReg1ZktKt436b2yQsFlF/NxythU0WLL7EfAQhcqxPO
T4Wtdl61WX5gw/yJY8JYTSmiEvYIRL9BBhsehy3Zo1+yBkt6l2IW+t3lJ4TntqdBiilbfj4ZpZ3o
i/TVczDEIRyenfpwqwUXu/PnTg1L+KTnj9JEZP6ZP10Gefd366mQbPSkyg0qNCebBS/AX8rh4IoE
fkjsrr6WX/o5rs0HOtSKl2lZf/tWmvQ4E4iRIEBcouOfmQZcbwwJNXntbuVTeKbUAKJI0eOkcnlh
A3VOhMoiEFp5N/Rz9Sy93/ZCJHVdP2e+2Z6YNpRyJV6D/HCXLKFRK4JgVLm2L2jhtSOubzbSqdqo
PZ+q78YtjN5ymAEp3ZloG5sd/MwQIM3yqkE+FGmppDvw+ArD2GyCRGDdWcpLJn5QBKHsUD7auZGW
LO6ACI+2LdM+kLeNo8jJZgyo9V15uWI9K+uVTKUFmKT9K3NZGc+wTLs32gzNRrYKmcKU6kyCTuQa
C4juzm/ry1CHRL2wZNBSKxAz5GNjc1N7iDPDEa5Yw++3nHUh4en9S/KgI+LZQMq4E9V3ooE1TgoZ
0BctomlayqmXpGouQB7TMcWMF39w7xkbWm5Jg2HW3TkzO3vGBO0WTXnJ9aD9ThGRSnHnadKvv4Vc
w+3p5KnXm4SlgCj1KTZEspeIwgR2aTcxNK2OMP9tsz3kvsGIEhD6Cf4sjP7qdreEc5fohu8S+Fvk
osVIkz3rM46lKMaKIOoNdgb2Vq3JArjJ2PpghPugiRANc20pS30D7hagamawAJC23tlgXFSvBSUn
HIhoDeKuKiEj3VO6ShFHxHmpNQ1sJJuitTUDidVt0yd605pOeOUZVEeD9tNkJscveBSYq3o/ZAhC
8WGDOeMzql6wniPH4g1NdQJPkFLBV/MMx05d2h0O5kEi/iYERX2AaLyGfkISW3u7jsPVpigF9HCi
HGa4Vc+WtteQ0vQ/yZJZIljUb7M1tT7H/y5wHXoLDP6eVi1+C+yMzoN4ewp97NlFkCRofDqAAwOI
S7lbdkHsRAxB+ZLrNKhaWXXGFfq8TJPfzTQGMf3mfKIRh3uqD8ObRACam4jTa6Dh4J3qHaxk6zgm
4wgaIKHckgo0ZXIPjBXimwyaNDIJ52oimYhL2dIPPVleVKaIYCugXXlIUUASHFiOS69+ogQr2Cfi
gq4/Bx6BNP2vHLmc1w5aLBpepQtKRMxXAGnnNs2WWbeHaNHO/H7/FYexjp8AT5njrFo6bhh4yRze
pPnzouQkg2AIyR4mQxKDiIJmPv/FzRjvr+4Djtbo2qjqdc4YosZYOBPPn6qU5t2a9jbjwRRGoSoT
gvpSm6KGGEJ2jbzYviNxNMvLj2LDA0iTbXNb8kQ40Vb6vzc23kiMbfPc0IfhFcILATRxCKz5ouh+
BOjsaw/lU597LjUdiTu9Y+Tz7urylBYAha0oi39j4itPjlz0hIatiZsbE3rffzImEokwlVV++l2G
elPC+BSdk7l+51SIDJf6uCXaDN84snZDYihU9AbredpuOlYzAHOWSkjvS9T9+iR9gWGHh6k+JIWS
n6p/B67P5SqrYJBxaVZNAliJVrPWq+XUdW/UbCNOxArb5ZJWuSIjmc9uk8dGuNaePj8h0zL7s+Of
wQ89gRS2hbhW8Y3KFh+XGOgnaXOcZxwFKaH+3MZW5s5E2IVfpK3DJK1s9AEPT2BuJ5fIWRr6doWU
CqkLb9TlbpHxwg0MonoZ+OxmljHnU2gml4Xz3fsjh/3I1ldOwsWi1sk2fBP2wzC9x9OalL9Oh2FH
ZWkF5GdL54ieTFZXrqL4/lf0zZwrA71Wl5OjKEXLKJq0ReNI6vv4+tnPNW3iGAvJmnZO3G6jKuQt
RSXNs3pdxsfxr+6v0JjuPb1UZG1NkRJqBEVRMau6Y5ab0aCWCnEki+fu7LzoQcxTM4TlTmcyccGN
i3gxfiqKJjp1JPmc90tJUo+Meztd/FOgkz2XLFqe1pI3Bqtu+4Zw9Zdgg+3habusWwUqRmA0ixx8
tZJlmmfdm2FjAz6jSnWAxaBXPoQ7tBXlScFAk3cRYLMpD7LK3I0mRaipVyK34Md18K2uFLtTEGy0
5sbTLPS4DskD4k5roeIMtQKvgC/KDXHDTdJEiC4kHd5aN5gAm1/ScZ1rfeE6e6TQa9/88wco0KBi
L/r5YAyCgze7XsGOhfB+HyVMibG2lvOWRy+z0Sy+Rrgc0LVqJzhc5hB8gjHOtC27yhmAyPHB2Q45
LZN2RE4eyW20/vSyCyu+ESJFC6g0yk0IP0Dio5pdMVaQwYlbOgSDRw5APpXOb9Vf+q3QD0rO2+dB
AfsaiDYWVz3+iUlj/D7fNIFN3aUhQwEjNO3peu9ou/jT/F9iq0quXv0IIV5pM8jE5ZJMt9VnpJ0I
0lUIyOH+jgLkzu0u58EHahU9lynFBbxWiWzFJn80bUFfsYly7eJUMHyBwoBOlqiC+UP1nHl4t3OM
BqTrfcOCro8P+54cnYMBvm4a5HKCV/hepq2Png5o+smEtNuG4Ktp996TLqN85ewod1zPJTw2mRWf
hIDiwqNBbhyb34Kfh2vEoXWsPlk0oTMGhpuxhyHu+I6QpnF+1QjlxgjQXmQZ9xcwLUgGsMTJE3kc
0qjtB9hlV/0n+evx423uFG9PQRKdT52j67e8k4TXxe43e2u8W74Xf4g/GlcGNyFjv5QcU7VqIG4A
LUg+p7oK8Td45xRYWnNjVvDSHKrn3gFom6Asw4+37T72Y+Tfb910CwaOmzoVawWFFCaDbzZxmGIW
8LlJC8icJWVERMhoUmiVDRVtc0YeOaBELASMof4fKTRPBJTMz1J8jH2iuk6tEATJ9s3VB00Qnofx
IjJgNZfCP9n9dxe7W+rOsDyFOJtEk/JfaldCBsUfxNhzzNr3u2o6czmMFhGI3A9G/53rbBlu6GwE
37ZLQ799MVPL0AQLBRMaSIbfNu/ryvuHBLnMBN1j55AdQe1o3Jre4qMiJt9eaB8ROdUOUODbjnN0
FZ46sUiQ5PixKG9QA12BQQMmYH5ECiRDlhl9FNZJCBkrL8W73M1HRFXNoAujXqIw5b1kY7YrVx6p
8i58kqOs3l2zTqz+jCPYhi760V3YzwwiuV3hwRrrS7csyKghgxParEKh7EnrXTYtms2waVfShq9q
029krNGwpx/wLv35S2+2PEZQSKTcBhw/Ec4ZTST3ghfLodA5IEQeoYs/nFmsgrqaycS2iqM9liwD
iTzevSa5KS2y02JovQWx5AN3E8hm1+X7x+DSEf+AZzL3FTry1BEkbphzDmPLoBffnKIDYHFFFCbQ
mETTohWCwXYIefGT79wCLvKwVPfhFBlHB2XzqB1vZJYBGnh8mx/ppR1uTAWr7qc7wwh2LvLf24O8
qyHaP52biUJHX+EIPy+NN7UjORdp+29q1TIrWLdkW/CPiOgIttEphjY9+Ypdc112RBUEVbzBn6j1
+RuY9cUHwQQyb9SzGSjkDtsleBxM9rdEh8kiMGjCgSkL8etolnB5i/EEnslsC40tugRU6+XlIqH+
nqtOQMLNGaI9amez4NvPiy3T2ZpGS7iq85bRzyLzFmUS0vRhKzhKvS52SGVpLH6itwF/MnhkTku4
07IQE6FXafo8MrAKALR/loMcixJCE6sRM/9RwlTWsh5yuRftEvarGNYzf+oVM1ZbgDCBRE1VtGzI
0ZceMH0J3r4A3fKRN0z12IhVHTpCVEz4mTTkX/BCKE+WWNCxlm46Ab4w/xiT34CsnK1jEtWaLxu0
3OadaVDcNVdnZNcAl0ApFqiWWnoVDVrmBrROmraajTdQsJEcHvcchSo0MKYeP1N02WRD05U94IKK
VZJwUOnBb2Opkd2Ad88uRtkCVOwY+iiNzrccgRYd4+/Ki6K+QdRLB+m0t249tuODvFIdJD8nswLG
5KWkWKOw2lbgF1OCZCqPLDmbiGQmGVmRlw00ZoQx/a96Z/5rUOwSEnj9ozfCqnWijrx762FkYI3r
8j+xb4U4jVWnM9QHebGeMH9b6INpqkbl7aCb+L6UM/ftWHy3o+Y7+G2GsUbvazbiN7yYmKxiClFP
7fON2OR+AvARoCmjjEZTSWUn+MT9k8CGCCc4ktbwjCP47jUugWQ56D+DsgUJoKyGBeAW+W93QwLq
Zcmb0um03wUw7tMj5Mee2k77aqie5vuW4Lk+yWy1RgeRoq3SSFp2Zt2kIkK78wSuxmLOJIaPNt8Z
nPy6nbXqJi8MW5O38vCGrBWMDh2NCkFANkYJhBEqmXmWpDHiDoDPTRnCIKsg2mESTaJFHWFk/PAB
dfCQiwvrva8tn9yfik9thkCWu4/Fmx9X1huOv34/OqD4thZtflbfXJH/ee11VMp+FD+PG64Q4ox9
rv76ZxSlKlHgc02Ty1zCK6SwT/aaccWsv6V86zddYDAIi42dzloJXUx7uara9bjiBhJ15CsCUezL
LwBSroC2i0TBPWnOi2iuA1QvDBFi3BVotqY4CB09EkskOlJmiYDJPT2ob+QzIexOT5ZsrxbJrr4y
k/F7xXTPNQllgEetf4gxb3qvbvoP7mW+WyQVC2+aldjPWWp6AYJsHDtuXSlpPCMa2F1oj/GjQeOA
9z8NGJv9ehMWQezsKJZyrVpsy/utX4lxGLMnhcYa/NUDFFop/voXKWXkgGtiooStYfd/iR+QeYnX
1TjRgouv9c7clC/WmshLQPhLg7LBQIjo8cE7s25G1Attz/UZvQzurAQaJ3itpzcmNVjJ5kZrsje2
lVxjkzAv7TpNz4GkIgBKLsJY78rh0hIwvYCpMEOi8ICxRmeUMLvJ0dpNZijQXMS3KPj0jyrwnJ/q
H9213U391NJPLEpoC00pZrHryFEu7YJ3Rq3+hUCRLpC0dOHUUFFBW00JDZQJSpa4L2K/0UNdkwGp
fP+ddwITxAF9buRl9gohWt24Ex55c//fEdFgdDr2zsKh19vg04/+r1Tk3RavE9ACpOkTupnmZTp1
zG3dmOr0tsCKn9P43zIKu683u7+KHRmf6ZIuPzCrO2rKP7WlO+ww28l/QjVwiRClesyw6GNxsPQ/
cKqXv+ZfYddGySteKjvbB3q+keX9ymDR9VvlHnH49xp/avH4DOTxdTXjH1R7ANegwvfTYKJPl4JZ
6rVdLgpgGiGaD01FTIAJYdr7YFXBfFJ5J+Unys3uSvapa3qEh/QooOPIyagTqKK8i5Sz6iGAI+SZ
zgIvVsf4kiG4sDgvdcfrD8o9gao7DfZygak0k8L0NLhM/JCS8SF2hEtA49UYsOIf1tAtvP5LqTbq
icKMt0R7VZqbkF3rpaGWlnYkbJH5ABxVdA4jIwBGiPm0yNs/fh4VwpVZnmQGuRJYD3jPPtRKTitf
vQ2ehbD5z8/xw00L1oJDO/+LflcCmupQR5jGQU3vseF+2tCb5Hh5Vh1RNwa8XYmD5v8pAbajAmyP
GjuWW8IbwpLBrjvIpxk61h1hV3cy8X8cFU1Im+w0D/FYkM3CJK6x5OvqHA3Lt5NqaW5W12O45IBj
uCbdKEjWATgh0n3Z6d72AlYRrzd46B9aIvPICYQ+gBpIoGRQTRGy8H8zr+XVC8ej6WDJtdue3TAZ
wMmAUXYdFTKIl/zGtnc5u+t1oLhLBfYPuLdL2xwAR8iHi4+Ev6JXTQHci7+Hl//KAxtNac+vlpv/
PBJiO5y+d9ZVyEb+7+RHhHC2XkwIKTGHfmFGgFrGBk0aggJWSu0vY5b4j3zItQGld9Nqq/35R8ay
GR4mKKVmsNfDfuNB9Dz3S2BsFRiRU5kRcAFR+cDk0wP9OIJKhJltJUwUbrfGSkiDkp3urtLXv1lr
2TgYMGIEGqeyxGMC8IoGQiHArMM0gNsVBJEd0uPgsvEKQ2xi9Wyrfjziq5j+H3jbHpv2XunrJPns
x8iHVpsAd/fedmcXRprAOADNcWgVk9+X0H6EMCfmIeZHb2IKgiX9VBdtVrqH5fXCytMEyAD9WpYO
0vFLoJOCubv+xp4WzUHKp/SXOx/C8T354zFZC7iOhdxNMp6YYMlDluxqKw6tYfKAk1/5ybZT8dsV
+/HzNLxCBKCUT16pTdCJRBX9NH5PfYs/m4XVop5NqQUBDOtaaYIvzbh1s8PPSS9vEHdHSCy4Xnb2
v1lnGodpQaZLdfiURwDpLlamTqnuwk9BF7W3HUMW1A+gB00Z+sjU1W9qvobATZJx6LSjo75XeRi3
yZsd+H03ORVH5rZfz93MtHALhYgA3eZKeNdeYsA+hdE+oSG+ePcdFBNwsnAk0tVnAVxhZNG69Fhy
7MMIrXc2rFepvd3QEMBX9p6KC0OVC5pNr+AFYpB/Rnj7y96cA97dCeZgNz2hgSKR7rnIOw/cqo4I
y3hjfP3aQe4oz6IWmfgGvKMRAfBYq/FzaF8r+aQqvaQIPd6NzpeHPk91umUxeOPs28iCTFhQYP2g
dkZLVAe0ddzoVKg0ML3FrPimcy+/sukrZWEFLZcyY23vJG8iTWVAt8mdTJo1ubqMAA+OKrp86zck
xVG3N0gQUwd/0c+AZmsv4uQpP9XuWcdK4MHY0NPPN9ceG1B6VG1Acu/xqv6niaijbLz7mee4iia+
cUcx+2r759kAZ1LgX5d4v74vOYPI+pwTkK35Rhe34dQdCddY2AbAn66sHsaEhL2aZb9YwsyfoVAh
8pssESdJDywY7aCb5z/UtiGFan+4ZSqKw9YxgwhB52ZPmOfG5Wuq1nyBP0i4w/sTu3Bqh8yTssw4
ls+BRdTKhBnbe1ywgaH8qXdqsI8vP1nsmqBviqF5nr9UsofAu4CXaMnLXhQforAqc9o6fEZH0xsD
IzfFYLOWgjsLNgPTbLM2/lTLs40Z0/c/579zQRtZc0weF6TWR3VAD96cAR/2E/MxP9RR83zmD9+M
kdL82CFHDQetDjJepg3WL8XQKolJqE9eBP6aLUBO4u3WAGa2eNJHIudSCktF1l4oyMRj39TLBimH
f7273YUOjKPzojUc3EaLfXhxj2jnRIOGxT/uNPeB6yCu1ttg0/UChjjFMw25GMrM8vsRpyOPTtG0
jiRRii4OlEp8dzO3FZWJZsINKca6WH/Xa5+e+ZLt48Gl/NMZppp9Yl2g3O3HnHq0P/ZgFGwYctGr
fZet/+tx5Yb9NsIMeWvnsTgwselMLuQrz6amT9utK4U68OsYKXDTtuw2JoOomC+igvQ8EBb2e7fX
RARL5aTF+e4rj6tABKoNKxapQL3NBtzggK4pQalAk2CHysgWqjGUnUGSKShH3zMcUu5gctP8hvUD
ba74fbJ0ijXhwt4ZXiZaKBarM1Zy6CFEDzuB/znxpZEQbE7qxRdqVdTgSmm/CForoGqUVPOrGfnR
5EMr/wsB4OfjSgea9OHwT8X5fAihYRMFJXZYYNYJgUoapYZYKRf4+ZlZu8nr6uEHZvbIwvQVK05q
26KL+BBsQQiT7i3wcl+IFeDCcIpIkH5rRQ4YEsucSF0nuKqGhwObmr67gfLD7uO6mNEJQWAhgKdo
ac9qAlQiT6pr4Bf2/lbubrFOlMpmIUIO5owWCN76NoVG6ocKfU6ek3OHjd8++1l8gR+Xc7ztkXxj
TwW4L8VmNOJ3Q1VpIOytBjr3ZIyGrjXsOOSdFHOnrbjTL9fGKUQ19koYYsiT4mChcFwNjI3C0/39
VanmyeWTYF1A1KsvyPCmaSdZKhCaQ5hH02hlxG0ZZWb/vwKnpSoIkI7UEGQwQnEpsl/3z7CQl9j6
dGVrCXZcs+3RE9utzXoGZ9ic72wL/X8IdJnSWNaQGz9dkymJrsb5FWSYKWW+t2gyXEUW0GYP0elj
/TW5Un3u8C2R8evfGsXBnWSjuLW0irIvDqrsBviJZBoX2Be5xD6mYI3YiHAfWILlpgWaiU+5XYCk
4oBkH04hmSuY1QKzu5KA7efl/5/6nygJKbczWJamssb5kciNb4NEwsPDEspWMP5xdnSLplwIrBd/
zKTIgcPBp5dAGnUtBXSvvHueza+xrxR+papgsvhUSLbCCoRA9Him/P0wpaDxj3XOTBE2FNYNfKph
N6ELCNGP4UhVz0xXWcyNz04drgiJsLlzYwQMTbUt6qwWeib/iAgVStDEYo0iyVwQxu2y73eEeT80
ddFMWQZn1dYqpwJsNq/sFVrlPSWPycVJrZ4lTZGp4kYTHLWEZRbwlmLQUeLV+andNK89zCsKjV3v
AB/tgBtTiC4EUXo5Sn0zOmOaQ5R6X2wESUdLuw6/rpB/eIEdvapORRBUGvwW1IZpGwWYm75LduA7
C97sKsUEF6trAMxWwt7d2bTHkVpVqTAD3ma1bZUjqs23iBWT2Z/yDZSTzE3nBLotfs4YAeBwyvLk
/TeoPAfeuRdsIaHPx8nRHe9XZogpVvn3UXEcVGSDW/7yrDH6b+fYJXVzK7SM5y3u8OcWwMKAqkYW
03cFLZ3xIk9g13r2p4tYGPQo5EDWqg0q385flp7+uUX4TozWiBpVWKLdm/JM0tJ3JN2T4DTycj5U
18eNYkbIpue1QSTRilQESBS2R19kC/MmvmmHdElxVt4lfc3Fz98ebYZtVrJCJVotEo73PV/jv8vw
a+JjFi64VFMgqa6oJSg/jIl1XDZZ3POeqjSDE+zDi/Pxlt2VEBVgB72Xyn4jIXL4lg/SUJJ+VdgL
B33PKE2PreQetN7TT2Mug5mZB0jxmJrLs7skCJxrsK9bCLug55HukJmg+T21u8JATWNi2pQzBYzL
sHF0m6IL15PiolzLfwYgbjfWkNKFDv/YY/xOS4En1yvJt8e6qzV0k53y1gBq2WGiOFgg5W0+/6Im
30SqaxaRl6qfMiSh5IC3DwqDtE64xtE9nYZzHEh8z4+g4Na6EEItRVHOvcaWSPrVtCyepFF2WbzJ
UNKbAqkeLVhJLanSpZpBgLF+MyLkElxKfAee3rf7JqSTt0+e6EN58rZIaJuvbKPGKxd4+PRztCZs
pSWkJbbJWSNmb9Kqe0Oo3DfnS4lzVpXWMHBEDYkIecr4YrvWs7ZSDNv6i1PS05mYS3hlv/0yJO1i
0TUz05+vRS3D5v8n21gSLFgUvGAOJF7JFhdWPDNvuD7gZPHYD5OMcwu8A8mAEkqFOBvDJiVcDnTO
8xp8gsnsETcJ6YBKqW6t/WTPnhVEkKsQI8wMZF4xS9E4Egv366G6874D0ug4I7WcRvygOxrZA7xB
eFmxISepKbLNqFGJjhayXUS+D8t1q4NMiQyT5qJaNAUQjPxVMOFTnP5NiTse8/u9VwQqNgYzpIvJ
FnXfAij5LwQY4Pj1/PVrkBS3ntSJAQbRNeVHuMA8h282PjY3Gu7pDvJqFwmc7tghkSnrY2TKCtDk
SQcO7fbHJu2mn7AcWZXuv8cf3HC6Dba7Y4eNOhVGkmBm4yxNuOx/tzkd8kHLb5Z+MgTKhTif69yo
sREyPtr4HZWkiUzmU2Tk/Btx4ELOw7UeCUUnk2ZHG24/uhMGalo0bNAi2rPCbmojqz4A83FulLtg
c9wOh4fCb86e+mg0e440+zRLteTmGDkZKLTeYpRrfmx0TstP+1RAJbwjcnUHLUWN/OWhlNY7u79f
TpsYHrs7ou0GBAXtAQi4klCNJwUgN+/oswj4ouJeOtWcdx8YJ+EOTlWC4GfFR0qv1ELXsmRTR+zs
sgbWOGe0hpioNwAsvKaW3w96W2/n+f465lMrNsA4VPRjZGTOKmeFk4CwIVZLTjk21TzSwLAd/koq
GQhCX1+MVeXjWBPN8z3tTdatoh4NDThbsgfVGBKhyPkkVqsa5qms8B7nONuA0r8Ike2oQIJJncZK
BNB/g7IMb0Buysi71ee368v5wBqrQ71+gTz0mvRgDk2jUhN7Y1+X/Z6rM6t2gKYyL1lzWwbu+0n9
aOA7PcSVHo/kimL913ZdwKUATTfsALpysHQzVCPlBTddm6gd480I/TmJ0ZYvcGp+d9y/WpRa7jFY
vld6dXp5nEzmlz2HS7c5Im4LY9ju5rx52CZIgF5OAr45Lh3SETq+yDXRZvFpnvQ05sf/FjPcd9gn
9X8mcAO2JMajzSr1mdYoS0ORfwKatnqRuKdGHPf5OdQQSdPC4BsibTpcO7u7rSOnvgo4xPvm9rVm
VyjQ0eSp7a5lbAIiaIZTSdCu0yZG0XA6N0KZdoGRGPYm4IClrro/fFCKBQ2FlF+nI2CitznMONmV
daK1eHj18+GYtJkoQzPV+GmxP4HbNkeadjAAgAHZzgU/C1HlgQCzBqDaLTZSUDfKvgazMutEIJl8
lIBlz1Jm3j6eKHte24ra2GeFBYCvfnIpNN4ZHKiHRe8P18XgML5nlIkWWePbuIhP0iXzEKi5fewg
goB0W/7ET/wO4IvQ+OIfAxGXovhuORAY7Lj0HwbtPfGE0DwBFyJfb9CQ5yLqX2hyKRu0WtZlY9cL
6CGDjpmFksKRWbROXEAjikBIAvcciYiAp3jOH0F8eCwBvCmPvw4M333QnFA96VU5kJoloDPtQQl+
8QCDmi4pjynLqh3qznFNOCV8nr8zJNw0USN5dn2npXmq1+wlAhr+GuvwmvwDlUW9v4c8Ok4LuYc+
uA8KvKm2gnf1WlMkOgbIdAG9FTuIpsQkK2TiMWMYLvvFeCJ9Fvfx4pL6uTor9Cfh45Paw2VrsuS5
ueR62H/zJCAng6XbBmHkxHAqXEXmruGVHAlZR9tQpWyrR+uqjhhMEYntoy+Rh89Z0EhN+xdF0JvS
f3y9CQ3E5xi9TmX2eCNDMDjrlPNssf+xvvnwgIXylwRLp6lqoz1n8Qg3ajw+DL60FsrxHN/M55oA
hPPjyofJJTBPdW8W5CHwIrFFc8h2pDPA23XwsKPJlf5wrsY2X2+5Il0Bg+M/hgPUz1RMPGlu6Cbm
NbRO91qrhglZwtNcXEdTtE26/HfbjHH5BXN8OupLOLNiCZWgsuyTM+ZC1a2wzlLoDfBu5PZnuv7I
33QCflM4ydbWav9S4N37gyn1wqIZARb6Z5UWTtuBBHNd9e1tPL+xgpshDwQWvzqSzGgM+Rg7aNkm
KbvpdKalFn7TXMrfV2dWWtFkZfiDdGe1I4TOorOmqMXcy5aOYXGcjibOLDvvqBL9ujd4kFW195wn
LDsZLBiYnalkwgJvmcP8FWBWDG3PUFm3YV1HHdNCBnRj004gljtO8f8+2F8qOXoFEesZgVSdxLX0
DjelZbVd7H4raTcXPHduiRjHzsyXnI/sjv3dTULSVGcj3p0QLiaAgTOfsV7//e+T2Ie/fOFc3Lvd
jZK2kEmiVTM7VB+xh0UkOuUWz0Yio+3VcIacNJIb0DL83QNhSotnyQ+t3RyzlZukZkf9EzsnvKAk
DUzSzoBQ7+BpesKn9wxcG8ESIj0Fx3oqmvmWIoA5x3lar6/7koyjP6O0RoAndNcaAm3uqONXBf8g
ov2VK77hXftirzFspg1ViMVAc86FDMSzdkEqa0OJUAjBSRBFqxjH7X1G3xWLd4cOfQLM5VnfYEJf
A4/IbxWdeUX4W+HXFmzDfvU5jMHF9/ga7+2fYqOpVDQ0+M9+cCRVMmtF6j5IU+j3jbUw+/Iwu9UH
lrX4Athzlw4jXP9xfeY0+Slz8pgV34nngLVUwPLXSNI0PsaZpzAyady1Yp2uOZfVzfzx+QS9YB69
rdchecDGxHSNRlhQkfAXWh851BmXFUo1I4m37YUlgw2sGI22uk8nXrE7mwXsZXjouGAMB2A+6/Kz
rGdKX15ZKWhqvRNerPX+U/FKrf5NVJidBYr7dxZeNEKPSOkMx5/Tgt3PGxfyXKtphbWoT5H/Ni5T
Y5T85odrru1kiUjPZAWQPSRNUb3qrZMbIZiyQtOcimMgThZhnvO3rzT0C0X/EdEmVQqvFsRPZqSt
+LV5p3DNemTSKgyR19yNK4BB7zDKN9NPKgZTyy2yW4boue7XTrDzRU8SJ4z1OPLlBuLtF+qRbkbX
U0OdAeh2QIng/XSfynZJQT4r40Rdix5Ne3NkxZmLc1YwFras084OG28d5uHSrs4LQA0kYTkiv6Ot
wno3OO/Egs9NTMWNkBqjl6jqHGMC82JvB5EQgia03fHWjpiKiAC/9nHhNzl0c6YuSjT/eXjQO59z
E+7HEu2MFxDLLgP/8jvvGsBszc68+4LZNvcNYEgFyzfXyxcd8P02SgWmzlF4yDI5sC4Eq2aqtg2c
Ccurwcqr3u8hbrHza18tyOcoMjWrnQ8UQL38SxxDRIHPQWd6WG5wGMxkUAouKB0dSvD99jKQxDRw
/zv1ceO6gveZx2rWqGYIwILRFF6exY8/ay4GNy1Z+ky/xNKqC635dKtM1ABDbM5l01oTzcDhU2XF
x3dnuHWHbjlvEgHFR3rLiLiS+lHz6yjDK1G/PzbvmzYeurAj+6/aC+8SdvOm/5JIij7yH7VQMlPq
KRdxp/AUetDX/qcgZmihhj0NYLBX0HX63cI3b5ZkYCFMAcAfrCT1R9f/yl69PM0lekzGckKdflqS
Gjgnv9iw66jDyDnhdu7O7bJjVbDmUW/7HEcHT2UgC7XM7Ijg9VD0fVJ7Awlo+VpIisFxDq4vMbiF
ODlVh8cz/P+UKsx7lP1qt1oW6d7K7cEgvaFdsgDJjdHSMBbJ/uZB7aNXm8Et4+kH/TwGvz/tOXeU
Tvj9eWJmpSVoqQz4NxDa+Gg3mx3d4nM/WtSGHFhYsDo21yvu50o1iS/9nS2ZrRLuHGlbJk2btKqO
y/djdE1WeM5gLDCopRy90/KT3OKcAzMUAabWyZ+20vcGeVhqFjZnQ01+7A+RIkZ4nJQxW9Og7qBT
QOVJFp95BcFDMs89CVk4uN5YdxuSSi7yu435s56OzKm9GSsTvf6/UjV2R9vefnyyJAuc3Jw/9twY
YF+3XoTmg2ooud8qsRvyIxg8sPqTneK/yjd/+kMen3u2KDrjM5ED8cyHTY8hmLbiwj+nHVUTTiIS
S3hrmyQuEhUgudnYiFbHRwxeuBr0BogFjg6VIwZYDhWASDv7azzplxanTelN8dpGuBiLPy7MwNtC
gjEcdPXRoClu1aaCoVhjSujlbTO51mMoerbmj59GMhOQNvj4xLw8safEzN5kn97WYneLrYvDKjNY
X299CEEkGOMcXFMzv5mj7/h/6oIr0cYrwsguMTfahTUgptAy29daBTQKm5C72dzuLo9GBK89DKnN
kiFvyGkVX8VMjTgPZPsHmsj84OwzZ4HnF/XhQ+QylcOU1GoxYaCR1D2jWe+dpnyTfkoU4mXeUft4
ImEq+45z1r5coXWzsIifljzP9T/Nn2B2TqBHS90Q28Yjk9Etr8mLXMC5cQffhsFAc/446uwBIR1g
gMZ3ZdDYtj1yFJTXHi78mJUhQfz4bHnnoEPylzlVcUXec+qdktf5EdMJ4JWO4bxEcnMdMTyI+97n
5j4GTiKlDbgcgzJ3k7MavloGtTlvRYJGDOjSmTvlqO1aMCcNGcQrBGFRVn5BKskyxKFWx95SmuJv
S+CBSkT3UynR3KmJx0z1MFpyio1+P8wWtWlsuqjWksyEffx4E+uVXZEzBUjTfTXb8UHrOqr3meO+
7hLYKAFdd4CuFDPi7oIUjeB+dv/6B+c6qJA8GgAdasPIQyzc9eV3xB2O3Xu2+zDFwaZXNKrUx+sA
a2D8lcRbw7cxjnXe/bhgezIKL/T3SdTUnJ+pafLzPiTnsDlO6Qv46KrvHNFC/qYmL1JaF617Mx93
4dvIgUsfnSrMtkwpDHedY6TnhVPz8hyvqvHNVfboTpdhiGYN2eQ4CF2RG6dV3T8MmIiHoBcb6KG0
i4sPUc+tnhJYFBGX8LurSpcoSPP5MS6SrrYsL4WN6lpVt6a9hH5qqmHIHdjph38PoLRORe4Okvr2
Qwu+dqiczC0YIWmRTSPnVPrhHq3AcxkDG24Sf45lxvQ4Qb4/Wfu5SYLZnF/62A6qMRGtTf1rMdR8
HfCKBcxudEuuJu7UWuWljRwotWWDPOVwTysUf6DfDkavYHwgKcbRTZ9iNumULoo/Q0DNwq3sh07K
BxTeeNVFmiopVm5iy4Mh7Kxph7xkghG7KxNVZ1W8u0usRWdKNqXIAI6Zb4ZXC1aOToi5uSnyOHPH
QfMsbpF256J8ZjafSKEZzpsgvvgWkuHUJWq0AmVVYl1Kum6j6l2KC5SCMIuVEeS5a9tD5Wk9PPrA
0dL+xUNVlhdrqF3iK1WABNjaTOVxuQ33DfqcPR5LAoX5MSTIv7GxAkZg2p/kf1Opgd6cFSN+h2Et
SERkB+A4P+EqU4U+YwLqX0CNpLQL2VE4O7P8opuXR/VS1guu2VqqZpOqG32pn6FAlApRg6ZsJOYe
EDnFMdPswplMwpUNcMwprO9kwLfD3vlyU8tL5qBiZTaUhBAc2cb9VQ0E3y5uzi9JgbueKi/XM1cW
BptQiapRCmbmstE9rx5JXEXLaknGeFUmjFNL8ByI/pIQWHJXb/3QglZkPplQrAHJVq3UJut9eF+R
r6e0GbdtEjVP3ILe3JyGBZQKnzfNhabvBLWqnubw4Zq93SMm47usR7XKaE8yGTp/YXx2z6ba9OHG
MxGQ1QtI/kpKOe1r/shIZJGL+2aaLHj6aiYBNAP7hzRbbMLhLr6o77kRTltLLzyEgkB/mrLLz3bf
6ZiLggvjLhBhR+Pj6q89ynG0RZuPR3Tx2TSak7a47rC/DAPSCAJWJynt6L7nD/daoL8owjoHVxem
CrZWQ30osZmEG7B8ywDqsvze7hQjFPSlhd8FheVZZJlTEuLqmXjAg5YQkfaUxwVb6DEtMf9ORKbi
/goOA9CCFCN181mtZqjg1NjdJVre8k708l9Yyp5rr9+quv3w0win7oDPRkoYTMHDqTo8iQsXfpIW
XeOIoM/QsAEph7PHP6awH7+n1sLxdEDWlrm04NdM6oNuDClNJqSvikzgxr6jGEXCtn4GYJYH6lVw
LO3BvVZ70BjmIH09rZ12ik1OlEsVCPOhcO+0LgrUjlU4cLNAoqm3RHkCcZ7m5fxkj68iF250shfo
YcV6qKenhK/S75o8HbYovD43feZHXZFK62mbTrHRaDsB6jeYGiScCSfmT8oHN2Xi1KePSC8NwhzU
y6HmSc+Sb36Y/fLSUxXFlPBoQkH01s1mHaD0coAqqiZPWJ29IDrQNrXlEQd9kW8N7TlDBdLrRMZ2
JkAldrN1gATTZIC9XLh//R0w7/bA2Q7iRo/u4KkQohN0HFfbzxnR7cj+j4CqtBy+EFfXo27gwVi1
tLi8hrWwUUlSOtIZBGtyWXYAWNhiXTaGkxkmt5usbPxAncW9tbqdLdpbNb6ykgUAadst6KaG0+o9
QD6A9wzMlZkX11yVrbxc+oCXKWr7YPhSNzXXSSi8Z+bkxzGT54oCcVBSlkgWZI0WhEqb5by5BDvm
SIVJriFePNhySlkhcwghLRAEVn8yIrrTgN1ZWnHKLk0IiCTYqTeN6G6WdnfiawwO3hpZsqtpEjWg
4yVB/0T4lOr67+1IDdeoHmROEszQ8hBgdPqzRvMl/ZmGk8UpQwf3G66a/+4wQqi9IrEHL2WnkSKK
kdhwbfOBRKL/ktTivu08tIUGdXgj7GHfxHhVmT7mQT4K9KRGNDydrhaXabsuoNZXJHy6xRAK2txy
hVd/9IHZHodq38YQ2JdRV2aHb0Uab4QTmOwEJMu56Y3db/ffcRSP64bZiDn+4+zUzPSeQLg28cBa
fT8ZbEeNXKUh47rVphQOH3+GBljWHbyIduI39QQVTrb8qpMKfaJphGhXEv6s5L6JxCRvpm+j6XDA
02H8/txHujejgQJfxQeOb5TfRjBhTYHvwxs83NB5rqduK/PWJOQ6sB2LDpogqQIIQPesC/y4Jxcu
Wnyuq+6dkdyiWGfAHn0AcPkOhm1V0vw1EcepMiGvewOsWlaWXaff3vt315lBmi/NpuhfLjdIzaU4
rUnV7N8/GQ5m12MQzFiUQUtSQeX2ZAJA2IVXtVM2kvKTDWkppXHuGWAQNqpSFtla9EfgulY+lXgg
Slh8IS6Kfiz+/gC9XjHpVq1sadfTS7Kk5wWrM2gw34KStW93Jf72Xr6BdR8m7frcue5Ln0s97Vmc
oP6fVFhsPqiSkqVFzR8EB4xz6TmZObigrQ4c6zl34I/WrmmFUHCrhxFd1PStltErabiN9djT1DqU
+Vc3xnw82wq4+z1tKB89S9SrvXaR8FaUVMJmFj5d6sCNo7AOu0rRcULpit7YdlpuQcnCq1LDLeIA
PgO3zW7+LF+0kWcXPjIiWbf3CWLUjtLsJqfvcBm1TFBFIDLAhDGYcvYuR4hVFzbNSwxyJWYvmek2
uli1ODODbkuMqmSoe+iqgmPPAbsxXPIelNxDvzLdv7voYtNMfUEw/kLSs1uIeydGw9abUnPRSndV
7u1lAwrTMt5QO1mA9DCyuw0AmZWry1zcU38aC2rS3/Ibycs4oyMXZooaSwLNht8V/8Xxh7J3SMPg
nIcVa83KiY0YhEtad/IVuu84K5Akf+r95+iRm8S2qtuKpscd9Pmbh41X4e1LQ+Bvxqr01jlBCyEi
zuKPKrPi70HSplOei1Xhkvnqw4SgsB6Y0cEedV+Aj0CLoqaEOw/yW47ChamT9XntM3eLpR0yS3+w
yqQsvIakpJQxnH6v1tQsW/wcVAWr/hYBIgl7fA5l/ZWxZsb+NTx24HHsy5AGQaEfu1b4GKSHU/it
+cM0blHgT9i+29AEukzaZTyZrrK3UiBwWpeEReXd3QD2LDUuAPYK7qkE8Vm+A9pImkW2dWCouY8T
AiXSxOy/mIFZXoe/FeZu/EgWEic+MLfVRLxc5GIbUtXLLKMgUvG2bs9HL2+2ZnMF90XFzCJ8LTEy
KMqXW51ecxGjx3qPJg9rHfqmJIKuPQCB2MQ/5+bQqOicX57KDh+9j/sE5hpUKqHCNlzs+ODzLBiz
F8yvUzW8M+VxwI0nHMqFCtkvE60VMWBj5ZpHX2FCtgqNOMlFK1LO6ylkHZmSDwxo2yuqggdYGj8Y
2NeUkaap0TqTZTnjDaNV8tH0AOX1lUVrnNYOlaxfH+sFVmeI3ShyYsJUMGrAG8ctU+Qz8BtpSzQn
B2vEjNoXWufncRWXbkJ7zy4rw0L+b1Rqe53HXJvnQmkLlZ8xyo+6fl5RqtvS0cXRmxiXfHwpxQXG
eoY65WYdT9cfJalROe1U4uCYbuCZ/dPkmSwhlqZTdYkMASn0PWNCQJIJv1XPF1bcxP1277kw3vSC
jaPU4A4ZFpSYGmcGsgLuZszDlHyO4OTaCPjcGKKDyIC3y4FOd3OWwgdLsTexGRFfjTZLA4Yf+ZEt
/FwMgAAI0E2MeQS9Ujz9bNt9M5qxFivkWMc6iBAeai29PlH9G2kZrUv8b7Gp4GuR4UVv4w0Ui8nY
nBcOEzeG+vPR0Ye02md6xg46ukZiMBWwGpNY+Y4Oqd1tynkoOJXp6gPu4IFWixS6mZK1clKOd3Pb
vjiBITII87H4Qs3lNdsgM76hOUJR/RXdNKZh1m/8srDmuw0CbAIiahMvuDsFzWMcFq5664dCYjq4
a0DJ8wzxl//92ISAaAxqaTDE9HorAja79pT2fTCBlC6LKEqiFZ/E+VpaspvSecXOP9FTWdymXtV3
CZnNUGFnxY3XoWTdXDNrhCxfaJl8J6Gjd1YKjrbLXe/LtOrLOcOINWE7pnrIj2D10RnWOwGvmUN4
BzXuPHlEkBbTbHZcg6O6GeRvzKFI0nDouQOxvMUsBrGHnN18BlOkaDsINEFKAWDjJ+8BVHAY7Cpa
IcIe2sn2cCvxoKFXb92mtejW0NZsFesHqanHV9IscMWIqTIXZBMfj98anPDf/KCb5xajkyRWaZgH
lNFRt6ZeWXOu2mf6OML+nHTz9nDosQyTRs3UYohol1jq1piNMClvuhMVGq59K1PJ7ZTopbBQV7MA
pMsNXkMMvaiT0/2HzqxVBl2nSCvlHp4BwiBTRnDRdXjrxi8NPly7zWwxDD6Qadx6Da3o6m11Drlz
61rblXGJ9IEPPHoPmvnkWwkf1pX84Q+y8qz7RRnDyzmiMMwEThSXiEcOjxOaKbbiuCZ22y/wK4Zv
pDXF0SEJ11xjgODG4U+3DeNuU9rz0G1D1boHLRTuq/pRPnFPBhK8pUcTNyiF8swh8qy5SuprwMhE
fgp0H2GEcQ7Sif/rhA6XbMGMgYkM8PxVpS9Kniarl17BJmZFEhf792kbgucpkOzZFJzCEFnAupsI
/TAO0qLpiPC9UQjc/D9MPm97lxSxJVZrE2IFx1tSFPr5zGTDoy0+oArtlMEO57Gc8KVNVqIUGbcF
oLTd8t64gaLus3hGxWv9vl5TrI6XpiyGCwsvP8g0pDe438Bb5dN8KvAb2DErkYSmGDniEnBEj1QD
YzH9A5T45l25A2mghoP44yTx5zxvUK1cXTUumZdC81bB5+Nqpagh55O+SyRwoHoPtyU9TadxZSs9
L33eQjWNidtSZrVpWH+PwhZW+3zwc7i91loY7frYmWe30qeKeOyiyR8LW5OEYvSlDE+sNOKDyrzf
YMkgLzzb3eAKt7S5p1e09dpq3zBorLxjo9+sx9WMDqR9lFm4Y8KTFiLKKHn+UA9osRYMVaizj/WA
1jqoV5F7oc5lgBbiAww3vVz8+cN0RdavlRxCNnrJXVQgMCN1ORiv5Hnwcp+ua0MkokQqXykKD6IC
hQ8KIVBUiglPNtp5iGSfRNSuSttk3VEosnA88+KZ8O5wy+NyVollZcej51Da841bYe6zNebI2/zZ
nPlCZSetk7bYL4PA+rIHOvMRBriCAr9558gFTK5G4DKQDbajy0dg0zE9xniupGvAfqhQOJiJB5PZ
MqwSsnWzDV7YqXLgWSIyC3dposFdGNo6ur/twbW4jkyCdJLY3BHdAVlozZt9ld3r0K9SozaGfwKd
pyvZJ+RALRCpulTAGAtx38359UHJQILvo2vIevQs9uJ2DkUK9UJsebLkFfPwiR5SL0/uZE+GGa/Q
BnAT1YSPZ3OGM2vEMYl0I3QJ3O+26ZRtrr24MGfAhgg0DNvQfDqOTiykEqDOXlUA+2IR0U4e2Xny
LFEmDEReci+3f9txXOi7vV/mFSolDARP8bcW3iS1oYHUj4tGlA5lH9sUA79whPSPVZKGt3GfF8+A
DcuIN0cJjYVk1OXVVK/DNrmhP2ealh7FCva9YhwbAH857Wwt6i1L4qO0s8JKgyOpRfBldqB2cIAO
0zd7qW5EKXOTKdEarmjskZjlOZq7JFklJ0pR0GLlBnxrpVGobMu3WvHsvewXN80oTPnAqixVJneq
MQ/IawPe2UWhZl+svE991xA5ht2Z3Rkb3OkaRqXNm8uHllNVo11/2CkVy4QuOz/KuG8Xkcljs8o0
ICJQvcQzgRayGwplHd4S5eLGP6d8fVaz/jdDVGV6wMS/9jlntCrNw9J8JgUrGY0mebODuqNOu2Ri
awuwoh80dott/Rg+3p85P+0swUjZVkoWBEJEHrbxTE82nJwRDsy8MenJdMIj8GKnQfSb6Sv7mtkU
1FlHSTky8ygWR0O2RjDCG2NpzCfyMXEtaUEzu52E38Ga/cvy2VY7J3zoLGE9FoHLe780Vvs1P4H6
8cY2lUQodAw8NALIpNbuzrJD0kgDu/Gdqj61WNEv290s7GysIqzZ73GutbBE4bq+JETDT7Dix+oC
FXX8ENtfVyOJj+ppE0rymvzkgHh51rBF9LUgSnkcrBdkZreKRPiWSkRVYtplnwR/mTRM/cHUralM
8JB3yEt1c59DGhCc/RAWLfmz4oo9E2lFlUwecuDgHe/wg8MYhAd4iWYQez/8ShXIyyTLZffpNasM
pSJ+7EXl8NyJ6Ix5I2cc69JuTcMLjwCnyfHb4sT3NPEwT7PwwjDOyQ5ttoRarwYBxYi5tFNm5h6g
P+V40ey1wNl6xQoI04pK4526WAi+f89fC92UZAJDhvlKqm0Y3w2e4YZn8FLjGIBOeiutkztXHf8w
+DojV65RnqOeqARCQurqOsWx7AG7f1x2OT6HuSDOD26aX7U/BIuSinThUOMey0G8PoKDtR6IZQgA
MCkjgaepJOi9YN8ix65AEq8O8NMTKwZjNcqDBKY2kw02hLhPnja3Zi8FTiFLyU/s4B4D30qbC9nB
nV0xazmASIgzE1n4DSv9a/vhuO8kTjsUt4j8pjjUovvM9aPI7RYMMcrn6nOf1Cod12QpkGMFFwO6
+g/WFBRrr4J9yv0KkHOt+fus607ZrdRGuxQyUmo+8o9ih5CrqIg8q0VyhruF/LIlJYB8/YeSX1Wt
8ex3xh/B6VXtu7rKyWeHyzX8GSNLHvSmIbuLhZq8ihYdSfVFfIfr1yOi+8PkSK/x4wZ9fhjhU6/V
FGfpvv2qH8eD8H2tnc2fe+c37IAEDTXtOr8zTByKTQfx8e7nzFhN5NmUmLJjA1RsA5/Fe7EsnEN2
WghobZ3FbGZb6mw9csqn4IlbFSw2RZNxUV3QNdi0p3ZeDdeFZtxIfalJrf/ylnEJ8InI3cs65ps/
Q7Q8kiGRsK4CxFYbeGxU0Q36DIPR+TH3AV5Kgejm1WCnXN24HyRUkar0+aUlnCIKXMverWcqfyC8
dLnlVR40fNvd/b1dJOUcSqFexk5h2YVxit+o/o9bQMpcpr/17+wc7+2mw4dFQvl9UZIACdfg7owT
RC/8M2kkXTZlSfQvjPDlUlqSJnxOpvhJ02FOQBrUYpKFywdwBB7JunMeyuGycDQ3wuud15dlGbWX
YIjVDgebRco6BcB28LaVKBMwWqbMS5dk5o5mQnW23057Px8srd9V9zCXCP+ha0/ILMd52Z2xOgKs
Zvlus3bCEcuHMZbXUpeEQcqdwh74gOFP0o+SrhWHWiLwqd7OQ9DOb92G1R0wxQRt85Ql/4+bHoqs
85BS4lBrMussmtdAamFg88yoEXLc2yNhDg3+Qr3cSCluH3TOj/MKt5/CMJSrY0DhBw4BRf1cSsq5
da+MReWxsocHF/EnENc+Sjbq7xBBaiH18Boyvbge+MV+eBeLVX1+PkC6ghboVns29YMbZf8Pz7zP
6Hba9/ifIMQoScFaqi9L7pL/Y/mNVRZcMbK7062S2yWRJjaXa5es52zwWi2ZrTigDW78ie4/mqaF
V6R273kEB7vKDuWcToukNAKXLB0VRKf0vreIiuqpTBBF7xcCopF7sg3wF/GRP0IzTz99x1E5DHEE
sn3zQ0x2DnO8WGqySq6t3Da6LBhNdmtZX0oYoorsV1GARxNoMTIh5C0L/kcPmWqgIDK9hGlxiKEQ
0rmr8c0Ldyk/ez8n06ISMlMunPT3z5e4P0v8QsKgpij8IKrC+IoXmFD9J+xpIVxmKV5D6ymjy7oY
sAIbfWWeFgMEFM68GCv5fjtJlJYBwiwWaiqyVtj8aS4hy2njik37N9pvNNYBwKxqCN6KRL9e6MWI
guJ2MChbQn4cz3Y5E54C8dVw7a9lyQtbqs8TNgeeOcKVmN+iD7ORnP4kQqmfnskf4bOHZTwAqmUR
2B0z7j+NtxTZa3SlrkLcTr1pgn2GmuELTa5l4QuJqM2n+Y9ViOpUGqoZTKGHhqjg05tOwivZsjSc
HoRpxE4PA15vvoShytJ6PNv/4xy/7QoKO/63vWzEGxKvn2CsCvhIGj+1CDA5wizTfNcMyU0bdzPN
IwFHOvZcIkTNm6NrX87Rx7EK14ZeLPf1lJWhpsLOpyqRSzDzxxiUhO/sXpMyqjZk/9YOolS+USND
TsDiQxtmW7qDsTVd4pP1bGkNxDXZqS9zEjlTR8ZOTb1oGyYk8Z/bW8Je0aR3vueHN6kcHnb405IK
AkhcS8u32NCTDl1BTyK8VEtMqPxL+DOVhFPyL4qMd1Kt9B0JmMZlLypqdGocZ6L8z67gLH3NHkd8
hDOzURu6C2OhKdlnXS1aZg6O8d0zOABp8De7/NOXx8hgogBdaIz9jvn6s9QH7u0RNrWxbhP+zfQH
xn4+ticqjIRVOt7e+qEsV4KJfM6p7khk/7H5DtOJ+il/d/dRBAihmNq4LlXM1g//tgZ/NYrS5d7K
NhYU5ZEnt2p0MBRTCEjNw9MdoCBDU+hGo7vXkOW2lVKxJvbqMozohuqE/I9QMouPcAYk7H+fmkLP
QK8mKH4iwPznLbglzQ+ywh3eoMOWAGTM5naSGrmxG+syDbfQNzhinej1YOmKV/vQHGms1ua4m4Zf
O62VhIqgWCNFTagpS0iyNrimCj6gz4qldKpaNxxtoZjEYhZBT+bNgR+iHh+pqCE0BaPgCgk+19oR
y8EVU2CCuJu6uO9pJKSOQmuVC9rcYdm1ZQtApAQLyfl/wkhKEB2eos76KdQOvohzihiXiPIfmFVV
mqgvohV6iwkEPDA5zcZb0ijHcZ9UmIiSXDRGnyXsACAO38FokpEJEtC1KQp45B3wchBqXqEpLujc
B8Cegm+WPn6BiLf1o0pJpF/22qbV49h0buc6ESa2ewetUbTVaDlqnWzj0uRRzW4quTgJ4npSpol9
9zDkyJG0Anl9Pc788w0gU7HWPJUNvrptlvC48zM6H5GJXrXuOf/3AQQvPmgdNyosrE65LmhWykz9
s67MiJrjKBQ4Hz0BGXmgNhaSuEdpIMmi/s3Njs6fowzdUMsSkyzKNpz7cvJJBUpdI/kOerBvIweV
qYtoZSReNCYuFhP7EGI4rPJEut2ggyGFK3+P+LDjh4sL2Gewt3J2APs9afQF2GhsN3a4ehLpfv/i
w2n0EuThPyBDvFu7gJJU3+w1WZV1PAwfngad6r0B4N+pvBNgKCESDf7zwuoNt7QFrSafU+EbowpB
WsrnD2VfOOR2MhF3PL4qrTpMTQJ8WFSgqjMSI5fz3H5LXeUBPCBgCJH7sIakGwA793vFLirums6x
rRPQfcp+yjMfH1jR+SAOQOVf0n+Kg9jpGycrH16T4ALIX8jpgSIvrQGHdv1v/jeEFZDKIKjDSoYk
m2mvC70vO5SXmzvPGv0HygYaA6WS+WTqSDyIPdtKKOHdoH7ruEnb4zqRnXkdW2tFGRGCV04vBpKc
kvkvXQ408MB/uBCg7z9sJ/Jg/QvJnCWwAYlP1k6UlObJi3LopndaomsF3lIfvUsJCILOh78ueAXu
KNR+PmdJF6n0mxxwdb2Jj4G5dLTioK3OvKGoRljSxXP7YgxvfyBe/LFTmq//WJ63qkvu0jYhiiRU
+JrM6hV7MSCey0SUNc7P6lvDHGKa7Me4WQfd0u3lhFdMNwpPxS8W77rcPkXytWV/5bsqKuq07r73
Xrh75IzaTqCWLfOffvt1wypicgMWEt4hF2qiF15568fhbq8xcM/0zP08qmnrbO/i2zGMusD+VvjU
t4mw2w1eIifWctMK8WT1kw//1ncRIEOUGShK1LCKVPaszfHfJxdLkKBh91s4/Q1ipd7Ma4oYs/BN
N8wLoyj1BqGFxNGhejJtiQ8H6Sl3L16aHNsnxDnJJViiqgPdzIGtzwwwqED5J936y5Gbobue7yHp
cW/BMbm3ATsZ9BdHJrTG5ANexwddPChjLSKLL6n1FOW4gdLkxuIf1FYe6sHTTUrFpJKOe1sltgLz
RSPqFRDaro60MbsNW8xyF/VBfAANANrSnS2rdMUJjeP1qNM9AcuvRItWjKMAFsI4YlxzdOCwNxfn
43GcVSV/2ADbyCYilUmx2s3l4yyKqH6UbAOyzSR1m4Ot8ucIkLtT1SjLBdoEHRXGDLwLvvl2YNDT
YFC3+olehHNWe5FaHbklipYtR7P3PxZ/5eUoAoVYZq7sAcO7eWmnRSuWEqPMPZ6+4/xlF/xc8JEY
qzKsHiMw2QXyXl8wxKChWYUJiZA/8Le+YeAL6rvXDSCrvIOOv+FlMQGN3JB6+Hig72puA6nDqi12
qR8k73rnry/VAnqp/icE3kz93pfi2hCugU95Jy4pYxMiNFdVwb4PruXw/NDrUOWoF6HayNg/Lkpj
myFq3O6tucCvL4U/nYeR1PHjVb/0p2v01LS1w0j2/Zdczk6SIWYmEMIE0mdtbIjygUaPFf5G3+wT
yK1H7pzO8x99FnuIXw0SUvqmkth85FOdgLnjzhRjXzEvY2v9Z+RH5HB5MLSsPR9lyWHOd77viXt0
9b3vgrfIbpkcFpC/e77gQrA3SvERj1g8TjO/RAxn+n0dw2FDYlCQexbryhU21EviaJ6Y4ouYURsj
pVrigL7rwampcDR0GSe9ueAmEbzYTROrV/gyYTOHrq5sKOfYkCi8goF5d5M2ApdgWJ0xrSQkzGqV
t+TdD90C+h1NTSvC2cZxqPKmW3EyMDO6WlsgDCznddom/LStFZglSpefD/l8Lw93sHeARUR2ZSMG
idEbQ13XdzE1ilIL+/NpItc6Jq6LaIp1chV4yJwSOet6Oc5l4RiYJx07TPrcpxY67w9eT7i+DUy5
1Uq30D0BTKX6XE8Ibk+25PkasGXg9grcIEOY1NVDNU8WxysaimpyYF5tYVfri19PAb8AwmjjvLiO
9W3sJMdbRzI7ezc0jqROeKYwUU5CXGQuBKTJVH9GgynQiGpAMcuxXLluM0AMJqc/em5RJRUXsqyV
Jjnh3XBaLef5jG1eNDue1dzKXBJ1W2C6aR+exuy3zP4kOMNFcqf/3kOQUw2HS5+11ofl42clANmL
4pShQeT1Fh5a49Jno3jIAKImJom9U1TAbN9CQlWH7VxC13PdqlSRugkERjWfR3J+cmP1ED7tIfG4
MNjfy15lLln4COysrua1Bvu20NVkhInD7/ujBA5Jfr4FytmUl4xQzFqmGpmCPTVunS9wGR9hNY5K
ImFer0U0j0iWyyOKid6QNedHpAOwY8xb99fg5hzuuV/HO0hKVpa4OUC61wMuAiGjvOkVor8WRy5l
LMVVipQ8/oGRGTW42EDGv3b9B4Yhfquey6obvSvmHagtBexyCfjTU/A/D7mu9tcQQ4KbZq4M2aOO
xwyTL5n2Qy8OJGDOK9ZJ6lVSEFf+a858NizzDFctRTl5p1DNEvD3Byq4ScuW2RKc1r2vOWuznuoJ
N5/SNGY2HuH2Xu/8LDWkEXkuuGDsnQz9nC6g7t8kRt8mOVKXWsAKqubL3b/zYu9wc94lQ9WkZSLb
B6qFBNNHSRPZSsKKABF5sPTxjfHYgRBASba+mDv6hgfFvzEC5PSlgJ3BcErPE/xOrb+5OH/zv/Bd
7se9k0e2DEFJyyPfeAx87qUVeoWA9j7iPa/uKBVc76HFlCo89hggmd2yZgrgi4cLHaYkIjq/3wTH
BI8xXGSX8O0arNuVRUntQNl9HC8UR8hqXQqGpPsLMOJ1IZQbvIZU7nRX3Lm5kL6YLN9VlNCqdCbT
TyFDSnBoGO0lcHmZlYEdNVkrBsh3cllUE4TLI4igoFYGiZc4RVLiORjDMQs4Oq/kYYFbPgfmz0NJ
0BsX/v1WzWKwfQhCD+K6kt7iu6/QvIz+0/BgBgiK05onM9aJfEdaG3HOFyoCjOrWXoGn8omW+P2d
RJTGJeoXWSm7cy4EhBXCCJQnVBz4mWJoP0vlQDGBZbd6bjbMpHHXThNdXkl+YHEzEUz7Ynkicxka
j8q5UNnOq8Ie5dW+qsotqncvEEA7IeI576iiegxF9ag/sGKmpwya+tjR/0WeFidgxjh3mikrkKKf
0lqafDT0syt1NQJd6gqj9zvISOo6JVOjDh7dwtbzY02RSgVNJGXLH3p1KdzsytRUN6fXj6ycXIon
SdN/OWLO2q1z9yz1KYHIIiaYDOjfpslKPLOlqQUPDZ0SbzF2pczKySQwvEvPceSMD0pYkeE+nhJF
INFkZvjQK7wfZA84X5jT0FDgakOjhvieONY1GT8lLwQ2AJyUHvr+rtXc7p3wf2ErSgWNNt/Y+uwH
jj15+hq5Cn2q8L1bc7/AuTRUgUsD4Iy3J+QsQf7v6l5QotEYHTDZ8L3kg31Z5IoriBbVCcR7ZJGI
T+kOFkU+RJPt7+qFe51Wdn6XDpAEaYCv/YjppwXVIlsDjvtyvsVrVK8JgnhbJZ7+Ym+AOr7SJso6
J6MB+BxnpTZpB7zkLO0B04EPKJ5cDRN9+s3Cn4M2AaUVlp2h8kcsastc23jA9V2OLe+NJ9bQfVs5
ktEW2UH0GqC0nO6EVG8ix3TUZhAypBrrlPUxfkwSIpTBbe8MPYKHF7pUmjKcX5OYuBygYKDZ1vsV
qAw4TXWQcaXFvGC1i/wtNbCvWFczNKp30WSkbHF/Duqukj41zuH/ur0Aq/y9d2IQcRA7XhZGgQNN
aIRUNHs3ihmC6yAMQ9LHse40Ac10e5diqiJymY4pGz4hA0KZkjFtbxr0tmBQU9IgEDryaInkRFZi
R0RJSeWgPrAYdI4e66FR33ictujow6zL2M+HAkmDnyNF4D4Gt4jP9PY5P4aEWS/72aPjxT+JjOpD
4xmSVq2EFWMuy3xAhqneYW6OgPVX60bjstSCA2ocu4KRfFftCd32gQR3hzo++WQEZG3kDAQHHQxj
sI8wex0NWvyU06Z52v9sQFXLiTOHqGvSF+QEfppc3+WLR4pufiTVkZ1O2Q/boHKr597lkz12Xn/r
Pow2dongv7CvZABMafdWv+N8vxiu35+GwAnA6LyW3DcvoejO6mjvBXByND931zAqDulYHDxxmZ3l
qD1FOfCZu7eGN6vjTQ9BgcM61BLfoO90sPO0IzxSJ7EjWV1heJu6iIVPPkiFRTq8J3tk2z9C77dm
9pHihCNKEFOzUP1zU2g95fe5Lw+HMU6ufS1vm7+UoPHKZI11x2Eq0/C8mLdzZ40ZxZjUHX8P4Yvs
1wbmWIhwKznqUB7ONjNJBqYSVw7r64ML7qXb+ARWVFidH1qKqljxz/hzpxrEdh3HlCFs/oTmFZTd
VshBlhh7mHbx39IBgKzjqgBo1/OeYGRUhCrsg2eVxtG7OnovwkZijpfXGwmAp/AU1btyV3pXXZ9S
5jUgMMxXDXooyJVmJ5jvts8ZY+klOx4dk5S2FecY6qD9nbLOcAbCXNlhRvvXzSkD8BCYXtxuj0vh
TUcg+iNOjbwhMaNPYevFSuG3i7BlJJ/fvyfaUfC9/6aE2YJdXNeRl72CYtAQu4ltpXR9zVIKpK6R
OEwEhDyHXnKxwnrt7oH/COTP3VXZIuGx75HsgWHNxUT7n9VkUjc9EwmSNM1hnAB7/7YLNNFka6Ag
Fb9Oaqo+qe9zIWXGQ7n8r1XLdcaw1TtaxVLVzoFdnu50Kljw6REj/LRCfQsUfDbWCoORrGXqGk9B
fiCfWfzjatyCmuepDb3RFffUGMZZ8ZJ4hlbuW1Lf3y4lp5viKpRoWeuW3JixSyG0RfUkWTKv72vi
K8KL+SLqsj0HdfgvYvugGrD2Tnb5/ntPcBX5PphCwd7w+yul2ELXHAwuS8oC5D/IdSpcaSlHhZjw
OMTrQHpf/BomNo5Aay4QxKECB9+7b9QJ62Yo/AN9MRO5BjsDYg2WjLOG9dTn3N6E2r/exmtHPqqf
DcoSvWLSU4QHhzlH4YFtxSwb4wN685cyATjXt9MBbnzi6qM1OOpFkwEEdKPasbop9qCQ5XObb0sb
IPeDMtT7/KpyUz7/RubvoTcuJPalGeON14eySQq2kmTQmXvta5fTRfSuKDV587INn5guENwFXh6m
1l9JsfLZCd2lJPYqmpuZQd717kMaM7cG077Zieio0B60S6DejyscRqCj+GdA2EeQVBu197Xx6Br3
s6Hu/EZngEIE7Cv82fVS/Qt7mXrofg08EM9ew5yboetPiPfj+pyWKKXB8FujtSErwPrGQne5HkWv
wzLJVVonG7Z3PI8fNwP7P7t/oC9LsIwbL+4j+1Z4D3djCmW35xeTbmK4Vlv0c9j5G4lr2tJwORKZ
YEKS+5q9Ult6bsUZ6Khf1bF/oMwioGZZimKv1IS5FB0usPbV+XjqVam33ewt/AiAF2fvOTnC2hX4
Y/20GLvu9PvGW0nUCvXYetEMDsNcR3r7o8OqKjJByFwWgutAOOYDSmfZC4bZdzxaMKhzW4kegVpA
F8STywzlCJpdbh9XVggMqEEflw/ovtVUdwN7vaWMgsH6BPopMI/sl83hhQhKsCat3/okJpapK9jW
Kg4PyV7njUfoZrAaiqZqVpxliGBB8JukWLctkJqYguMu6quC1OXG9H+wMGWLZHzaX+xIsb4oEChf
NpnVK1yiGPXS2xsS2iOWImTeJjSub7052HgxOM3Lz4rO39ZE/GVwvIbHZ8Yc4TciMJOZvuhNC3sw
zFIpj871mjbxyProd0y3WO3J2etChNqcm4cGYIXXN3VjQmEmFfsDT/cw9YruoHwTt26lSfbord1t
61eYFna1Py+ERqJE2GIHUa8bXAmf9HXBws1+t5Yg4850fY7WDj2XYMZPZyTTcCvdVGxRFHfX0KM2
vhw0r3LxX1ILZ1OTaqb/o8KTqGe93lbCY6OBFBdfpRkvWSz48iS9VwrbDWoy4doi4RAVDaYtRoMp
2mZel6mZGSsKTU9qn275exwuUKpU2LMHA0jeermffUNjaiSLwOaszVvmvno2b4Rl4KwG/iHSAswP
urhACA8UBRzSdtMZ73f5b2xb1iU9owtXdn7KH6vewdwZEiyPrnabSDKEkIFnGyjWDuT0PFRtxHTy
8WQ2BSGYnqjSx6A0c+CD86pfQaZ27H0BVAMXykRP3vsUWg/Rb+CpnSyCII2Da6hl4bMlyDoiEho4
5DHNNpQDTf9jJh/a+i/jet/oxJ+8g7CsIBKCC+d6JEHG/9YfmM34fREknf9E209mctHuXjynZdl4
HBUUyNDP8xetTc6ZCHi/oyLZpTtSsK9TcQAoDSZMeI0KfN/7+BB1ZtimhYFI7E+W3f/BXGEu0Kq3
M6nS5Oh3WdIIsQ4ezTqm+yrnAYlPMPc+xWicMmVtPD3dwTfV+MwTkO9MDaQ3xj7Iina/uj54cWm/
YQfjIFHGU4Tbt0NTdEQiAh8125hYiIkl5srZXZMgyA+v+U01rTxXTKD3P2E6xLOIDnqMI927eFNP
rFh0vB0J6XbT1H7CMMtnxygf/V0vofTLYiV9qTIgZdx0ECSHwrZ4pRhDwsMDyGnfMDVwpoDosLXr
slZWkSoCtYnXzgwRzSkXLqJYCjEng9+D1cdOvO3+8CC8VyCdL7ozqh+NiF8yxcnUnFjE4olH2jxh
omjdMzMAt51bQ19rddq09t5esovEGGbzcCBa2QH/1BJ0wJwDrtDZiiftP6ZaVBQuseKJYspbB69J
ryepOM1dp/na0KeroZsQdcWASai+pxlJ4YZGILk3iETiH8O3mJkVONBkUGDJCoNSzgqvEkrcq6Dd
uMe/u99fIgGX17YIZpCYi97x/YX8LgTcqlv/xeY3cuQj0pqMnWkznmzi1Camyxhxz7d3LasWM6tT
pBlUEtYG4j6+Qp5mjF7mbMrszWVktklRLby7ypjNTkx8hzHtKGSkLFfblsivfESrTU06E+a0QsMe
dlBJW4YR50EBvX/x5JonCslwMdCnIcjpEm7E5o9OmVR5nNCcG+mC5LjroebSHZG41LUe1fMBsiTo
+odLuMIcXKiC8LmZ2rbOjMWewb2FWje3INvwXr7TtygY1PBGz7XzY/TIzaSte0LoMiwE7yr7JsQD
8Xy4iJwdiMn8NIB+89pn1hUN0rQ01EFeF3/KPM88zZheD92bGElBjOfhSMUwoX0GLOEgwOyAUWQk
2ZB0hIxNhiXco5ZizNSmvZ8TldX6/nuOWrwDVzh6Mi/0DPXSpYx/i53HeogWAk5Mk4hqTNB7pFn1
dRHSOWUH6x8LC1vxh2uF9pvQcm6ieM1c2GZZ1W2hlxGfoQCJ5xkjHCMEnNUhJJUsAFYI8cCjD2nS
cA5ahrKTEMa2eh5dhMRm5bS6DjYUyorGf/zrceS0ivTC/D74NicFt0sq4FNFxdvp5E6+FmUxiyG1
CZIkSuZOnWQ4+5ftaNrlEwO907APGxqDGDrelO3jeBrVZCkfP2YAVym+ur8FOpgCLjqQsADb6YGS
WhjlMVVJUCGo3vX9XGPmDkxMyR+1/KZfeg/z6NUG9BQVvNvG+yEx5yS4pSNwocwXi5vWxzwVmIGo
sRtUi+VilGvjOxeBzDHOkCXRXALT4vpdKFvtoUw3G8nBg1iLb68e5Lwbq1WMm05FtE9KwxQOnd7m
uDNJTjgiME9gPV/cjMZPRHVzwCfe/3TNy8SxnaPNqoQRhwsNS99+Kkin9N6+mpvcKBBuUy1SFWK3
zeOun+5UuGoo7mGCYYJFsJpmzdOc8QWZ2CIMLrNoP5F5QUeei/TPCwTDMdHJDiy7VXyC/1AEaWT2
VV4IFhw17/Kjr5k46uFVO87mwZ74uRy0QL/DBsxXEjS7BVEUQ+L3FtqJov+MeVVuy/7Ubz0XKIYk
JldRajHuMfJudRCORAdy4PpfX1s8fkgJT0PBF59WkVKktJ4G4NTug8IvqB87GdCYif7ujRoBz+9J
n5CfbGFSMlI/jICB81QNPfvUOlZazqu2aTUZQsLgmjJmvcEWaNw2vWqRsdcBj42I5s10LIvBteWv
d8wSRcFclB/UOaTzLcXc5dQwZ3O2sNQ8/hgEwInZabqjDczmCz5ZHzbe7R1ZeYQ2Murd3i5qcH2i
GeswlFKhKYvz1M8SQF2a2dJ1MFRtmMroEcVCh96s2OHclFoiTTbg+RTSMp4EE72REbhQ2fnDDukw
uTQGUhZO8KTmcxrkyXaF8Mda+WWdI9R7DQfOGV8IHuP/Li79u/QRV+AMDd1oGz9E9KIbNN5sPvnY
3MxphmLxpn2kjTxnzqN5CAU6GKDL8Fd8rB2iabr561a5V5gHdpFJuwggZ3kb7j60z9Dcah20VdmM
VJRRvCLohrZQOXp9bSsOJmhJZwevQ1AoRNFGtkBRzQtQhWuYRUeRIWvpbbQAs+WZShIZ9DTTWZtD
cZfqdOZvmxjFTHt0e5hA3k9B0sumNdP76zFyLpTUA19myFH5znRiFlEURh/NwOgfnKjwKnutCZG/
qxN+BI6V/HSIs26PMOXEk/JqE7rMKcMetNbl+va/fH/Fbl66kaCdDLDWiyTih0HXqsfSdCSFhjyk
RxqRTLYB7Z9MRUO9D+gFLRhE71l690edVS7sYoQhWtZpKT9jjBgyAtW26T5/ICw76wMSi8jF7yIH
BSSNKZl85BNehd8OU6sJID9JJkc2+1nlrHenomf6eZ/eMvy3Hb0z9htUUUBgcS0sk/C7UMH7e4Ze
VTnWfP6QDkItH/Nztj6nNiGh6rhRynkWJKYS9wzvLJvzavKDfNxXFv/2Y1GkYl96mxgBxGBbFFqz
yMeHL6JoZDXHOZ5BC2w1PyjdOxVAFx1eN40JVZvx3PztVbSnnpU4VAVG3HBxNuBn8n4KnAuZ+h7C
lDAyWI+V854oU12hMul1Pb9KpADNgXTkEF7Q+3eSKmRi2Ko49aAohFGoJ1vHYK1jHgfj/KmCCud2
H4PGy8HtjKCVIfeNcakXWk7GesEWmY+yWXNJztVXvYAJErODVBGiE4At9Cw56HiAxwzTfnIT3Br7
2DDnhYlgw55HRzXNaTAgx2nV8V93WjtGrpSEgKKtc8/OhttU8EBXG5mdNbVCG5wUAJ5p8idfJcRP
OBJ+izrMVJFqb9RO0OfvMd77qmE04N41c1HZ5NUNtEW3F8/K4tzyEvVq+diJfB9lmP2+4qVhCqXS
0WtjEaruWUyJKpP37M2Q9VKbaidQWj5J0U97nR9NI9+twRFyhMQ3YYmIoFMjXxW34D3ygsP7CJVN
QqJsLnQ4FuXQeDWTD2bCwV+mrgyvvW/u/SS54Ju6B52/r3q6GraIe+M8fOMimBb87fWWw4dWnbEx
6slqDvuZ5fTrHYsc4BK8M2C3P7fH0flfUrsVBS7RrRhNzDIWi5UBZjJRUe8E9TbCIZRKOl5mI4sx
rSmeqBuHC/0e5G+V1jELI1ZD6dD6pTZ+C7Wb7aN720v+F0yNAI6kuuqzyy4JAy4BSVieuCabTFSL
oWikktNqkA9IJ8Ezpvbp4gyNJRkZ7Os/811pt0ddszB0I1h0YNehHlItSZnTF9akMg981xBHWO1p
cCq+NKk1wiB+9FaP9Tlz0NlBnkKzv8/IIoKIywJuNbK94e6hBEFv2xsMAmmdvrmkYKbXLYdoqXqI
qjU21OLO184XzL9VKqF0xkXc2vCElNu1/VYGJnDgqo+j4A6zg6yyIWNgl5e89AZRH7GeZ66fJVJs
h5JJS4tK7D0zERryA6+ACb6EZFXX26Am23MoA8aMHgIXS6XnKHAsUOH+RuUYUhvWN4Qa84Q20AzI
h4EQt1JHUEGAJE9+pL8ooOkJb18C8SQXHiJ/O7TwzfD6jMUU9iByDu6nesBJfs7eloWFsdym1nHb
iMCI/6DDdEt+RHAqyMato9S6LgdaLwWIINzp0HuRyUCdg5Sv146bOkNvKmGOGTy3ZXr0PhjPJmKP
STeq6htRwlAu+3Br0odO2YOej7qyzY6Vy5ib+70IvApmJxwkm8kYYaOd7wWFG+a7p8AIwZbZUUPp
JOlawLsqFUfMpPzfn+xalyIjld3NYtn487jWrEm+pv481cTp1GbTZY8J2k49Ac6loE+xeLz3ez6S
B9D0C4ar33s58f7HCvBmS8qAfvHJfpQdXRx+0nQ14DeIZ/HiXTDzWWfR08ap4fnTKyTHliupUZcR
CtPLIfbTbNkjPeTRzAlNNiqDUXQ9d0/1sgBWXzieN864Yb3x22mSstMlLwcoEuWkd7CKBGCjykAA
XRktUf7i1HTmEzjoQqk=
`protect end_protected
