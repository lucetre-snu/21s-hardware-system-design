`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7OtZBpltt/h9CD5IsJBmAQ+bQJxazkQVbRBjNJ7LWO+cgudo/XA7alKhPL+qAE8nYmt8n/nhFV7
1FHJnU9EmQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o0V8lbvMs2u7Pr48iEK+soyjigqgrrzx5HsGK4k7Ph8gI81XWNRtIljFPpaeGwucYu/H+gPVGgh4
LxNZUBJhgeC8kZr5P0UJ497gR4WHGLQSo0hvtVYHYDlrxnVk2S/+il/2gMAwvI5YF/lKiRUCJMb0
2mL6cpx+2git922rE9I=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hIqrLT0Q92Qul/GeORaSvJHHAIqLk6EmPwtSD3Sw8K7TFMN/pzvjFhA6g78oxGwtYju17YRUOAPP
BxWjMZac0YPGSx1A1AySaj/jWf8/sND51mJS4hxixMPKgd+iJln4gROFDpToYNAZ0eBhqGsKoRPf
Exo4YtwLGOksTW6jkb5XyScrMy9eg1uc2W3HXgQfQg9hr9gpWWe4xqhKUCFXFb9eiIDe3eaUQ22t
Qgz9S0YooH+uhgkKhXgOsKoG8s8RO9q+oyyLd0ANkoAdDySOy1H2+qKDhuJHoo8oHgkWp+t8x1nO
sbVK5ZibMfLbKeRbGwFkFsj+EKfWfOy4ck2AmA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O+omGGx7WVLIBeJijOGvFCJZ1IO2vxCm1x3fAW3H6+gw883MkRTmRZO0ddVzk3pvzQaBPeJUDRsY
1XbF7OM1C/khYSkVv9TjyhihrgNNT2rgkTkWtfQNoOMnsmtYkK2fHBBMyNXzHPZRBh+2VgTZHxjv
olfJ+wvlLAdf8BqZKWo1gutmRCut9sBqwVpKtMbEKFGRBnt2pETIJcWkewW45hEmUxoPlXpgWrRg
sESpeoKuutTTWJor2paEV2RoktNIWs/+x82raY47L1AIZ3uy3vEVemolA7/fyBhQXHdXuWEXntN5
bzesBXIrWmoZpCMSf+IISz8dywoKgC/dpdCKGQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pc9IPtPXrLLm2VmqSrmdhsB2/sqloTepqxhS9rXzXINDRuCWOADiBYd/5aw6fJ/PtHP6hvfQmgPM
pe5Rbb9vXhfZlTdZe6IYAV6ajOneMnpE0SRKlyLpgkbpQbwWF8Ta9x699vjybNfWF62AYBS3D7DQ
b0t7dD7uNK3C2oBkpBFbB3y/rTrUlQxN4AZtlp8BUDmTdKIOwvLfH64R9omltAgRoa9eT5fKR+NB
hJulrR0XnMdnz4MTDv9F/TNStcRrNIf5MM0b3o9Lm2heOPvkpoBOr22fj5c2jTQHuYFT3gyiU8GP
rFykj34Hi9/EcnhfJs9E3mtp1Tszf4e89AyXHw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rp2qWT1ngiwszVInFfAgNDsqirvFBRH0fhGMVLdTcJjuZF6cagj0r5deSp/lHSGQXbQ6hn2NE/pT
sVS4xwCY2B03TkdpZqI4G+dZXB8686b5iwRUQ7S4WwcHb3WXRb4Df1OHJ6dgH8h0dIOxvwXXNlqh
PKzd3cQ77q4ZzFc8bvI=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JmHrUUSZT8PLNYfmwBtqUH6qJ1p97BdaA2q40RVMw79ZG2/5JMAd6P3xNNzdIISzZU+jzu0NYPxL
Z/zfPbolJrCwAck6UGljZ/OOpPHLUDGkBAu8BIP536kFNfmsl2/w8PHTByudSnwDI/YKiNqfsxGP
M6Sq3+TkXml3dJEoLhHWDNi1mL1f4wADZ5vEh09j4ryxXNWZ0T1vCwLDq6JQfC0fF5S+fWguWeoy
y4GDwuB3WNo6v4nkxnIBm5jk34GhklMVorbQQ90znGRfAejdTRlBiH1jH/CASbqnXiNzj4+1wJ6K
83Kv1+Hi6TU2vQtu3O5wYTXjTMpJrASuG6iNvA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
Ir8Fj948lg5AH5dwlwFpcKnX/0RxFZzmQFfNFhV8IHe0equTtPTrkZWJdiG+Ahwi0gGEHXzzZwtz
l6iltspJ3Tk/iV2eD9xxmB/2QMU9ALQg+yGDHHseHcVpMEbtwEzQJKhiIzhEYc8lw59DDJmF9SRM
vxJoLwm1049/brrzS84kKAvOoBSoYUZHbs3DP/TOlsnMRLckBJUtmdy/Vz+ktDvaLIX9ygjAK93u
dRAAQdlrfFgdr7AeE9NskwzAqdmnvKby4D5CKzMLGziLebv/+X/AC++a9XLjQA25rDPkoh05acKj
W5mku7yAvOEusNtaUehG/sgEfiiaiRkC5nhTSfBf7O6+1Lqjx2Rhxu4wfySbsJSyKMh6mHLkVWx0
PUhGSH+otz0QubgXEJkvKO0dQXA2cJwMo06BW92GuUu7Bv17SKkN44uoqkuHptUu62ajWZhUBv4D
OC4ypnUscYJlYRtwyPhZOsOhHElXXnwzPCIUZxyqstrevsArcnK1GxBLXtuNXA7DmmwR42FLPIi/
OyYmyzJbypw+c3m2S1r45dKBlLbVjl3J1yDd/z9eYRRQQe0grhzZnDsZXB4Xehz15snMZd+jmeC5
+v81AMJwBUa/JrNo7SRsOjFsriuPyrQ3+l45SIOeqyISV9gT4fGb/IwZRs5AhmC1dspkyIJ3kaX0
dIltoxR3eRIqinUw4mQAl7VzjH/764gbTF2paSdY9fj0bt8s4GNdGoENhpiVg4k7ukpJMyQp07ye
5bOUjC1jtKXj2Sk+XqlMtYzkW90Vl4LqbfvNpT7qYKoJkhvYMPbrI8RvQ4ZFLoitB8vOkFemmfNe
hcmCeD3wHj4U71vLCgpIM2LZ/m5zYxsdq51hDfT6KxQTxEq/IZX2mRaF2qhcDZR6XHp1FYd0LtID
3345w81vRJWOnrxqKpjekrdYGh929JcJgQzKJ1oTlfwMiMsg72f5QLpeZArhKTAVOM4VcQJeMTNE
oSE+rEH+n4QjIIgcbaFWbNQqo3jYhWLQpPBaYoOKcx85RQuqlD2RH7tfl8tuNHC7wlc/R4fjuaSy
UTRfZ/tNVtenWCtdwOTRugHXqZ7DgD3z6tlyjMbsM64LVVKrmA5SW4eOK/M5gtTtrfUNOLxeD4RR
Bq8hKcaNXL5c6IydtzvTPwHdkpEjA3tb8r4TX5/f3TWDG+F8P7GQqKA/B3S+DoFyVSOLS7eTY8cn
u99PcBI5njC0jyB/hrkhcJ6e7+yZ2PnP88G5hK/aGr10x83iUD7+ZUyy4DAB5nyYDLLxhKs7/SLj
ClV33znHoUp++BjVNnwPsFaSWuW2GmHsuw8dcsUZ8fZhueRH3M08ang5d6ikJR+N3ZvTgHrK0G6a
Gm7S66kHhJFHXcdzRtzbDTYIRMaMIGFnnFx1qlnCMIBMYLhNRepYu71s2yQON0fZD1VI85NF9anO
jPX1zn9iswZlXdhrlTVv6oMJn34x3bzGUxTmRQg/w4mT010qvIvI38Y+jcU0WUnSyoWcDK/GeZQE
/owxJxMkEtwN2zIlpf5jOwqPs57+RKPKi2AdNTVExEhE13F5uajX0CW/uM4SN8fqJlg0IHgD5Kpx
I6LaTALJnS8GG5Il2qn67bt/FmcIq76w5of2nFjUylYNlsh80qeY6RIjTE6Cv5y04kwwx9O6dgiw
DJbTCicyoGfSRZzeweoJ0m4Bp0eswENpaj6WkeQ/jc5YLURs9oJ+X7PKw7c8DCkhuyNtoBSpSVKr
8nBzz4d7TMZulHGp+Z/9s74aJRhrxJKJijwg90WEhJI2h5PtgDdduhuzjSkPXb+Lv+Y2zJg75yEt
jpozw9V2AuH8dywDFQkY26yXehh02WFXS3GqH0iWNBi+SnXzAjaKE+/Z/uhW5tgt3yqt/oyKa026
Jdoi4//HehLJtM3ATm+pBOAU+rQYqZuJWhnz7xUYBiJfLBFLS+bnM4MqbhdzMNfdBvMCZOOqo4LR
Cs6RlN7Hs7IKuPWB0Rcaa/uYU1PJ+sHSI6xGqaDqe7aaWbXDM19Htb5asmvwpC9f1fK01EVVhWj7
KPWZTf/fQkt0YNoK3sqqt4Z4BSjHvROWKwlRMwlsIw4Veo3DS20wcTbF/QdYe1fgtskyYHteP5EF
eCUFzdROQb5sCJFMwyBjnI8ekTk2TRmkfMXBJ+ANz9y37xToE7aMMEM/qs2+oSUHD4tdYNcQNduC
yTA/lg+KHkrrv6U7ROdrrW5bMnjB3p71urJs2q/AJghnL8kKa7FsCtr07g63b9dnCP1b2rCaKE8B
nE2xSQbSB/r0gWCMDveotRRfrVAEPEmkOmvn4LV3hWNXJK8pHD0fuJJfOkY2Ryls/r7XuSQUUokH
erS5uAFP0BtBbFC9e7Fe9bOjbTfZwdiCW9j99EMvfK8qAfgqRm/dXLI1AgZJ2s5x69GZy3Zfid1b
yMYoFxsqyjRBSfakQVsl7PLuS58LFQAdiBxomc0Qq+Lxcf9HfqUFH8fRaRL2TecBYWlGoAp6NYD9
ZaVp/22GU4gecxELiMO0xseRpkzCs7HVu+0MFdHShuHTrwh5z4loRTrVC+STmmMW+oX55hjHfb3N
JepEiaeuUCd+O0j1bsKYuzu9Z2PBpfuDave/JV4EXsZbp9z++OlnfbcMI0c1kggPkpSBtwgqI9Mz
vVRuwNWpfnIDyqhjZTucHynO48ZysOcERXYrrg2HHZbxE3WpTreOJnS1JWO4TgxDSfwNbAYZlsCS
wUVfCY3/YEQUDKrSDq6Rh6t5oT1EKRDZ7SAW8BelC8UO2zh3YpYMc3tyEZYxdzfdGxuI0WeCNjWS
6r0t7GqN7iEhuz5kns6rHTIvuRt/benmWry5jmxxaJq+k+j/QMUO3DIBJRcLOpHFF9I/mZA/a9jG
thSgYAO2Lz3qwbzOmnGGeNwOFA60kQnadYvOi4xefn/r/WPaU13J2enGFqTFVimI2R+AxHWgfjU2
m3CaOgFRdrvxmOHg6nQ+HOLqFl2dP940PmXihs5spjXZBZ8cPB9hzzMelfEH55+lv+HquJ7CD03J
DNzKP74eqlBctKBWohxXWEO9zIDj5rYDZUhQTT94bHHg+eCVMtZ1SGQmMGdw/wGs30FqHwN7ZkSF
HDgkdExXAbOc2rEBPjhjK+E7x3DyhdoW6zVKn56qYQknADgZ9I+mSLv61oH241qLFSOBjUkePZFR
mg0En6eyxzJBeKZwaKE8ivaPND93VuWOdKBNhG3WvjNQ4/j1rRvSWmrojGWyDDTiK7dX0AaJJTQH
4R2YOcOCvKrrtnzYsResK6s0cTxLGGEK8ZWhZJQRnDlOSEa8dYIUHMuiFFl5GgbzWKNUhVJAAXcm
0mmdO8wpO7qTmv0lrFoi3gaFk4FN/2tMNI9CHiaMmBGpj6tIRCiL7TPtoEerP2PNy7wVWSUQ9lZ7
A5EH+eT4/7W+tFNH/UW5qVhn4CnY0696cUuC4fiqlFBQfuhZXB777zEBTo+QkWtC1YEyCbTtqRzZ
9FnB0+Xs9StSSxr/5b5/HfYuxycq68TRrdXMtiOJyHpTTkWreK8aZ7yuMvncoMbcvQrB64arsTbu
6OyFpDZfPN3z5dvper7fOrKsI1iqvEHBxuNwmFfSGUmszhq2zbBRY3bfVUcfT4dj9eaHeVH+2gSl
sg6u4doD9x71yqh8zE6UgHNKaH7VKHvwyyNAPhkzirJZ9hlPejBhenAUN80OM0kZskF8kXFcG+L1
B526V8btr2T+JOj1Kuu6z3Q6qNso+Zab101FORJ8smFPCkLwzlTE+V3k4i58+1nP/nu1QjJQWRBi
OaV8n96yUMpSVRr5qpN5eHcxwg64Kz2CSlcYvhbDaYVA10HQYTypZyJRhFSW/kyCSOc45m7lJcpf
g7qFv55MRv7qIUOoHg1qBs5sVNNFXba2o7Nsrxe6mLo60dCZ4yZchQomXQy5yopFDCYY2TBLB1Xg
ux2IeMR6Db9sy+OhyFa9pzp1mE1xDQG/jlWarS1tG7G9XAmFim47XNeHoaFTIM45Ze9sGBs9p8WL
Zh73DB22zs+fMll+xqmfj+Q4Hq0MCyIbVCdNzY+hzb8PV+2HavFYnYJduop7x48Kf9h5Tmqee80X
LLNifzXONQaq8FHkdfYhPlHhUL3fDAAioOIekznf1OsNoQgGivAHIJlmYHOTeQg9JM6MiIstbrPn
mCLX5/bw45AgY6aflkEqwUMMtqVrJmcyM8Eg+gvHnr5GoFA6pQ/F5GW99BN4To2bbgz9UdtWmZvK
+q6np9cWv/GYVLRKbvgeBAlcfmLQzSWUswvRV4G+ORdiPhG64vvfE+bggva7Ez7uvGHwmjSRff6E
5HgC5l2Ha4taMOqQ3tkwI4HFkgaDvqGKYDKcOKnLD5LJ4Q2EHhTwvp1ZyBrI4/SCVYHCYG5j39dS
+qR61CLrVQMBBumTdoPSXI97WA0VmBJvFpK9ndjwfr4NdnvvknwsLcU9jswYt2UT6YwSo8D003O4
fytfFRnn89AWt+BGavDpvFDafh/NP0/hJo0CuS/DBES4yUYidC3jBUqo3XUfmt6uxvX/zKfHCQSV
8n7/OPJaMWkxdTLmPT1PxLz+CVxJXQ05kfdBQ3VZHI+U0OSZ1R4OPpSxxsiAgRoHJT87BgYTNyO2
RB9Q3H2rAVVQYMolDd2LMKqgsmto9z1hAfboulDaDwnkyOEyQYXxB39pLlO8QUmP9Qwm+yaP9ilz
7ngAIoSS+3NeDlyqzD78NRs2SWEDY8NP/xdTdFBPKjT5aqnDj6rRdRl22y6qF8nLZyWlBMuXQeUE
9wlGHKJnNf1c83ZPtsHmUo+1W50ZXZnGQvvmkyrFHHPZvtRxmfdPsPn32OXiEQbOEOwC04FQS1cj
SI7TT7dEwwi7r9H1QxPPt8CfRE7hHHcOYB2jheEpwLMmjztbpcHaR4i3rCuGYpLq0sOkqrEkkAIA
ymuEHnTecBuI2S1uYNnAGfaCKxx4kcZhSvM0M03N15AxJVs8uVVWh2xOX2JQJgaE2f+H4HS0uzeB
pgTad7n+p38Hu/Ki3nvn4KiIrkbbw3Fj1C78E87rXDUpuz7AeDgjS+DDxRYKQspk/nB88+HNCr23
tfjOkx1rt2jxCEPKyXKPjdaxr7STO6+q3IwT+u11iB5bUj24qbNyRRjli/+arCpOoqI+P/IcWg+M
xAz7BPhWk6OrbrSbe0brcUmRhdxXFI4L4138s+Rt+SEEek3ssTh/pXHSeR4eeXcLW/oICHaLOBVJ
MBxRUo1P6Sqsows42lqq2NZIVHgpg0yIWsNvmUkakyoyhjBLO0NsdYqYeudgLlZVziGLCVnvoIs4
p7rMelLuq/SnpRwdrIQgZli/4iILPhGOl6uKrTBsKk4a3WVXaLtOsPVrsCZB1OWK1z0ChI6lJ3WB
tQ7tIn55B7h65ZEFuQjNIX+RvUixZARadqomtZiC/Dhrji9enIMahMuUXu3BGMl0y9i2VY6fia4x
CpzxSq2Cj9migmvysoMDGBeS1RKSlQ/wCf7EXQRhG9p0ShTepvkxn2ouDnXvsImxJRUI9SctGnPF
25pleQry/sRnEcQ+PCIsRlbru2kRpYzAWxMb839c+08QN8BwTKTw+KXUKLTy8Ylotsz94QL7WiZW
V6EtqTLDh1HbmvaG0XpU1c9veRNMV4VEAssVjOQPslw6AxgM+n/Qx+s6YTY21HN9QkYEhhPJ6jDn
unKkG0IwZ4N7nlPhrYMpO9EVeBcRiLXHxhKSWXmHBdeGvpRrOx2Tx9NUDzhbJaut9EzvlQCXfCKs
oaUbjs5fRKD2qBcsXojmWwS7RnG9vE1PE3UO2QRm0v4ruOu2/a9ImUPiKU79XE7RebI+ROMulhm1
fN29eXpudg5gLYPLEFSpT3nHSctA93fYhMu9Z7xNfW7tKBTYeDGxyAzOeBGj0sd4dkRF++LHVc4t
SNmKR/dH6jWcX9EAOeX74yiVNjMKS2ePNC9d6bQX9VH/od+TGzDCiJH4Sa3d6lTrXxl6GOy310b2
rSAewDne8P9JGLp3VypBYNnw7MgEEaj2MZxjHB9Jv3KQWQYafba12Ly6vqJEhTbEdWp3Jm4A+h2o
YTdSwBUDE1VRtoGpCHjagpT0FqY3NgkP8RSMt0tJqW0ZTHwWQBmowfpY6KqUs8YAd5+aEIIjmgj7
EukxfSuPTeJJjveTJB2k4dSX4ipuTgCJXe7wVKcCDxj8WViMJ3TomWd6gd6/FcPdz8g0aDcb1JJD
dpnKkaBA7ZZH71SyG5oyX1+g1qTk0UlOVbYm3f5BdEF7V3Nbit25Rk5FH1AGZj2ZgIP1OJgbtw1B
Cfg7az7wCzl2XHOzen9cZkXAf3OAQGCuwzL/v9DG5PyG0W9ECiX8Ew0SO9x2ppNVvQUH0eHDKJkC
NdCb8oVPgvSDCi1BvrX3X4cqjjxIYNvgetfimlTCASD7Zj6xcTFKHUDM1DhscOxNtTPbRIxJqOBB
7xvPAzrxnp7SmKVVhTgvdzgLaFu9CKKWcJBFTbrWhavnevfxE/jlRAuAGBUbx4iapL0Hdmm1vNSQ
73PiQmeaD+0m2BULWsJVtc3dTTIN0hT3WYvQHS8n/5cNGeUA+63dxzWYesivhEmDXWKPe/fu0AAP
dAYzeb7aHn7TRzSNXMGLMMnplBGls2T8VHVt1Av1w9HlSbDF87DVo9FAaixbci3sPVZFFM52Fgu4
GH+f/59XwMl4E9VZLwoMUE5pHJlwP4JTrVnpzATt7m3N12Zf4NQTD8dFYhqJAV9rB28t3F3td8SK
tjqr2V9gE2n6L5iH2h2i9fy2BFjyNESywImfjPDCzoYiYM6FoQsfd71m7zmMfWxgW48wcUqG0/hX
DPwuJ6mCendPS9tete90ipcuIVb9ikXAyaq74Ts7pOrhko1xnxItfBw7CCQQdP81cu934Bvt1QYP
5bKnWWwo11Eh0n/zR2C9Wek/OE2zzdXd/xs5G4HZ557uyGYX+vqDASZrXjYQ13Qz78CfunHxAKKR
hqxyrkR/vSL/Rj3Jy1temvDuQHlZSPFyGW9a9pbsI96+YyzxmkEUnBdh1ZGes5RLGNm97hJN3Y8G
A43RFIWgmcUJwn6Oh8WIP+j1PplvLEIF3XEXcmOvtTwpPWX2ukJ7AIyvQHp1kI4SK4P3ymtxG37s
CyJVaeDf11g+iQ5ogv0inr4W5wqLRbXjV9mVztUTrjvmaPc6BCYIc85clrte3chDT2NnF6RVHcNa
Nw8VmOShh408ffR1W+4900Aal05CdaY7t3URepwp381wcFOK1t7BaUajdcinU9xz2copzBCA0g+s
w+Ji4JFbWCZ/BL5D55emDsAj5I2X71DieLQyVHsdveloZoA8kDk+i4M6J/KC7FG1cK8oneBqsGbp
eS7KlyrDk+KNg20wf+/c0GZBKhupDfZmiV2c9vsIA+5soTPUGl1l7GeYO9edQCzGutpZLBQ1vQ4n
o/laZDwcIur8uMlQNzabEIqzv6ShNQuk7sH/G70l2G9QGQGakXW8FZvOavY56A+vs7Op1vQKvwc8
AHySTTpMlZ1cf1rv2wpOkOCc08mOJ6S7y7arlwWvcFbLJNfs+rZKQc2TnHf5VORXQvVqDnfeeXro
eKR3sVfkkqH1r4iiRjo9EC3ZImuxXqDlXjuyTdB+6MfWdeJOuMzKcaeY+vOI95TxVJ9ufYgefF0W
4eW2S+SE/u5PZK/Hhwm2xmo94+iZ8VnVpi7aWThp5cuUbypXHe0Ag8T78uIRgTbQ0eAQp/Eq+Umn
JBOmXbTRWlGB8a+9behPu0Xp0PKW7Odsl5LQwcuNeNc7mQ98ZNJrHcZ7Wp5pVg3sPyvvCu2+tFru
ZroHZRVo8hSALiDqgeb+yrY2TEZQhsr8UOjPJgBhVsHo9OcqLZFkoUZOq799/rQfEqCIqqyKAnM8
8ixm17Bl9q+jh8yqZCSmn7Go1HAvYCAvHUNK88sUf9at4kbbok7ylkzy+1lHbLfBJpse4bVoyW/z
3y8wQG8gSz4fdAkT2sKZHJpVKpoUuKpYEwqqDIgBczfiKwZ89G24Uh6qY9g3sio5TPHr5bnxvEua
/7IPKZnKfW6kiOoA559nMGSuZV3/srtU8WX2C/JPsJykALTaDe2yzfnU0UlyVTbNJ5YPvoFMNsHC
9FTE2qioJgn6zm6BtVOeTJXAEsLEn864U+y7s1qio7FwCFn4fF3iBFs7C7ncwPxsQJHnX0ANRDzM
on4rahM+U+pBboHJJqfaTOZYx6K8aAnHzxNAEOPbi6w9dUUPJTBG4Ru89SQgj9yLAYOqK5TlNCw3
8kzXjoAlr3TH93CDkoCF7aa2oIFu8ypknQMzo49PEYPti1NYieCjK+vg9dc+vNuqsLTFtPD+XLvk
SsdcHwPQMapsifpv8T79h+TP/8MagSpZJ40D0PWRQ5YVt8rIc5uzL9vWyRMUUwQh13UeMUswXTdc
gWM7WLehwZpmfaR7BueljqB2N0bktcTl0mcO8dZhza/dOYVa2RltvIK2n2Th6bx2xHL+woNjjGfx
M+zyrTdFnrL9YKiy1aVG8ocDQysEduXkvDl4A9EDRsGT5Z0hH9qpjewShFUVwq3CGi5tC2DpjGc2
umKL8DHEOHqewB6emzh8GOU5SWLknkLfdH+z2scBL85MKoNMFvXKQP/DXs+4eH37+ALOeIld6cah
6wTdaa5R6hKkFR+mi3IsdYAuXuNJkjlLmw7PBt+/ZrOhM0yXdZadAy3sZSfinEsivEyeHJQ1Hc0c
atxIPKj2Z9vtvy/CL+spL6DUoCMcoE1yC0Ki4wbBknhJJ+cKWF/DAzbI1fEmMluO4CUjYpwyi+oR
DTM9KUcyMSDd7rA7gMY2iqdd9D5645UlPd0vdHpO5ciTp7NuB8sAsOyn7+8kXL4k0LoRWb5kbJMI
piPIzE2/FPe93Xeol4CcGgxgJSEcFks6J5QHpUFr7sja4IMN9rE4zN9VCnQ4P/KaNYSOK5NfNhvz
NuXFXRWE0+tESDqYO9vE1VCh5500zG7ayUMAGxZWtWDtweQXj8E8tw8PWq/1I8iga3lFBvHbJqS4
7MTNTuAnkflvtwTCz3MTViwfnctOMApK9AfCY4r96aKOXSQSrKNf3u1pirMeShdI1+GO6a2hn6Cq
KrA8PtMiao3UK0EJ05cPW9C2EhbtAghPQgG+ayZgd3n5DbTvdIqUkZxWhtju6IDmE3Mbe18zJxrK
RX8i+zPsOyh4FIJdSMYK+PdsaJ+GuEyhsZV80Q1ZZpvVPHPfaDeFweKuDr+IljH1DyoJt5gRCV54
s8flPnZuZ+Syo+qYnWtWLEPXs3rtUDV8TTthg5QFxSf2JmxHhUee+2MTX2ZgezTlMvQAV9+wErH1
aqKUKPXCGlhLIKMFArIaXCm5m5b35u32zp3/d3q7b+k//Jl8vrooDvF8UigxePN3QlhbfAdGxd8j
kXSMh40E6haFm00Hqi5NhRcIkwBjCKWocqLcuLzDj0UXXF1T4K9RX13jITzhweXfcHQwsLiG/+Oy
aSfdYPclFuOhonjgnKySCjXBcWUuQ8IzaFcURM4D0egzUDy7mMwfOf47FpTccW59Ktq9fkfB0Qs3
6D9DCtFWRaL4fDH2Vc2VGIVPCm/rGaylf1lYx78vvSB2WQ4SFBdR8NA+XUPyAnd0or1KR50RHuhj
U4puw5puxr9pdU/PFK9fFs70iJ3Z8on615i15OLio71l/VDqkMwBmvHmB8yM0JGMAZdGQavTBlal
p2x9t0AynG8azLcHJP7frilPWkjJsP4JQftlFDXWMDoL43RUYQIGA+NN/vqTQITSVHFDHCuYx97P
f0zzMxbuIEFWZ/zQS+rM8YZIBgjy93TStZ1ZeZS6CORRrM4UaYJ/0bre0MwsmAbL9rAuG5rPnAl4
T3HNjIDZc9doX/03vdCgQj+AmkyboXqfKArO3JidyWI6Y0riUdx9ZwAjgjM12++FrUkzv1q9ggGR
qT0nK0hTQ1+M1a0aMae45VIDPAAN22Ycu8CMF3TvUEC6c9P3tB3sX9x8bxJ2CGMSEHUIhNT0N8FT
XKnuz4kcvP7rDO9tRs2NKLNBhm0qP7rK8xVS6N85Ur9SOHRKleQU1WdqMYYyHaTprxjal7okLXBm
cb4cuzmvWVwKRdaLzq/Hh0AbgYFWLzVu6vjAyHBmeodUMSq4wH/T544In1detTvxsI/NdCpQeoFQ
Ct690pv1ylLMa+/LY3nOzlXKthcR6sF9ngl7RYlBvUJ3pN00zyqt97Wu266TCsxHBJOg/UUvQh1A
LpBT7ewRAs8DVf/DxR71qI941tyTLC2W6HN6ZfqPOORKDtjRWn02bwQTTL+R0WCP/tPK4fMaVzkw
2A5R6gQtNfEqcYXVMe5HWOeeJ7lH5mncWQP8iDtsWlnSaEj4ehujCc2bQztE8nyMAZb+o8eIk9Uv
o/6vIO1z90gjXe6lMnZhXm3y7N/q5BVSuGQppjAgbc0XVAUt1OM8Rn8tSOzny6Il2PG1sAKp5AoH
YVVgEQrfe46ftV5GSyEDzyDJbsbsmr38z8UK/F1uiuTclCRvjP2xaN3qjMPl1I1UW3LKbSWfomnk
Qkpjz3tia8d1w10DbFbr2jEXviWWa5Vjd0PSLtFVkYWn0I0dijuAYI8ObQJTN3NSMmD+3O283eR8
H6ZwY/4O/T0WpLaEYIBNI9UaycllhiqtxQqNPEKAVTGZvbTXJKRZKFpk07RSWAiyMzQbTJ9jCCKI
EPNceINwiPr6WoeOX7/BFKvjlNUmVTuWxzyShKwyAHwgoFfnle/fJhz9y4aTIQKhY4viF3qQ4ZEd
hgHhtLzwqNvNDy0Qshtp8JmNx3z0XmSBjay3PUTAtiC2Zu6qpp6xIEnHGB8TNnJ/CeUUSPSgp6dt
4IUlrwkH0SQ7aAMwZinyIuausJx+Y+tgxMvuc1umUjMKBjOyPS1QBC7WKKHgiCppm7ZZ95Ol1Vw8
4UAfs4d90da4Z1e6RB/7V/vl4+wAinJYXvj3+HBdP8s5xqHSg3mMmca8xXw6dqASjjKxifJtACb4
Uy8P9tbxpxcFmSejsmYoz9KYK/mHY2z5F6p0mSdlC1EvrEG4YWuGq2QtIPblwZLRCj1WGK/RsmY+
nYjJAltzDEbyDs7GH7lZbutb46dJPFqBTDt6T2rRl5X1pMmy2WJOQSEPs5fTaannzBgyEYNuOQAQ
Al1pimhKhP9Uv2wqSN7pM7eTz1uRFpj5y3QgqRSONe4c/RkedWgVDLdpMCAIlSK2MLhe1dWsO0Vm
HkEeAyZa96RpkMXXtkR40Fp04lCKe+m06jEA3b9PEKzaPjFxINBZYpC0SWgrvtdao+T1ESr6Lsap
vgH7WUmJAZunj+WRW4HGotRPLA4eBPHHuJcKF2kELhdUygny15cU+UDrDlgQqbXXh2duy/s2PmFL
cqDbaNo6N44Y4r8B216BW7VeElA59xqBcbTUcF8zDfjsoPMZyHeKeTfdAEaRYnY02u6SyXCZ2RBG
aswPJ3D4RkehuLOajAYv9swnJpN1eBrK1UGDwgHUd7XyCd4H2tcWo+loIF1TbP/XYAv+iB/yrHAu
24J7u1QzdqS4j8r+pXpB5c0xP49CTk8eb9snjuTUz+wXXmVJ38/LM06r3gVAvUEgUxCckv3Z5cnN
Thkaoth5ixgyNWpD38JK5ojQko5ZsH1umxgQY5AhTDQU/vDI0p9wmlUbIGo1tA1hKnBeHmP5iQGx
blxm20GsVNPVd/+XOwHQwVZ/nLg4cRduP9HNB/6nmHBNAGJgm1n0/l5f3c0WCNyRbhSCGLfvGEi/
IkGulVjJ0cuzhWDcZF6sTdP+UqLfxcGCFCkfTHOHwRtaq3zLe61cUUiiNDlHav0Ii1JR4mCa4Uxo
044VmcQS7L/6cvd4ARzBR44FeaaanWvDWq4hNiDkCYYV8i+1qDpYXKR9UFYHj8+YsUiqhasF98b1
cbQCjbskKgB5uSBY9BMWaAaUd5np21ltA/rAOCGdGFQejbeX3ohFo5LIYC2HmgG6MUfklS60yd1P
zxD5O0t8pUETd4VNkoHvn7m2wWZzfmukt01Yxe+qKQEqaHslrlVsgFKZSLgZAIuihtSwKzblPMDZ
aQQ/VHlapgXpXJoOXWyZA9LqLZ66ncLfz12Y0+PUFtbd0ZZ2CoC8iICUmLYcB9SHmsWGkxb13X4V
3/OVF47x405A1HjfSV2/wnSM17bQMkJC/Zd2883QuN47vF8GhLyu3QrF5M4p++tKj28MrsftEBlq
WNirbHU4QcHbZh4S7Zthg6HvZcNT13VGRQ/8xaJ2uXiVMq0y/J56AgEcQ4RwJzmLP8L2DRcL3ckO
PxfLN0JSysdLWC52r30C0wq8C98TZPzJlTMBQ7FUa//vVz7KQgNNooyvT3AHn+ILzpKxK4dulx+Y
fWYLB2HiAJ3CRKIRv0urL5Ju7A6Kjp5hiDOUFYBoyB63sdR0XcHa7a6ozA30ufOJARF9QO3xdKtF
mQ3teh/dFvuoc46CMfxj0ZV6IT5A67WgxPgjWvk/7850sZhC6a5SUqsLpj84AeWSRE2yv2UzGzvI
eKYfAzcOEB2ZfYwsaMsVoWR64CVBrnMuSma7JO+OseSHxTTTwnR5HE/LpeWxevxZt+NzSbXLrEux
/2wHgX1ZKqgMB5Ak7dsp4igOH45/AqCZx+E2y0b10JnOk0U6Bo4rZDo3piPwymmg95z3pmlfOrhf
uhrD64WFIWaaDhxMIFJZNwMQEYCqGPccc52sviwQLtwAspVbcKYiYu7Ex3atBoPyfOpcqCzohVlZ
PTWd/r1imMuumVo56LjhrAtDaTegaGMh5efAYHvdSxCFhMJaAmwuNWclycCxf7q3qEj/CF4Zsqf5
+flhfOAIJ2wCnDmxMpguyEA3Q5csqc3uPVWVu+CobRaj6R+hSUs+vLMvDkF3Y57hgKxSeXVtvFDa
h3sWj+K2kA7BL3UQ6PWcWoydoCegB0HlMUzjMk9zcCXZN7MYyxnvszpbFlppboRPXoqqoAn7seGJ
dNvWeZVudtxQ8RyAqfd/UhTOUyfSfF4psYYUYpwPbP6Q/KxBdjeNNnqm/glmO4Sv1kkYuHIVCWEE
r5AUkFO/CsKzG3QTxjwDaQv5j2T9EaWGKk06V8G0mnfPzi2IPj9TgdGvIaP6ghVpzGxlA0o3Lycu
gda9HD1BNc8qiGuiIOyHmRW8jcjk4NjRw3grGH6SukC1oVsX9nYwOaR+AD3JQ0twsk1O01uHf/FG
KEndot8Q5ylhQ0sAO6KJ7BnQFbANIdyvSOPrFi7gtn9uvYr6ri6TvxsJN/adlcbeXgUt4iGRtb1w
yc0gaJCS2RzLWOPQiklnnSWxewVDNJ5w8yVfvCgj8/QUKlGRATCXvTTjPX7S2sQxgKWFVxS4OjfU
0tggHDJUMgUjnB0C7e2hvmlJImMaE5zsoKGJMIg8j6NBSnxbHCEG7tHIxgFO3FUhiMMdY/Nt5Jcc
BQgXUWkyRgmVhdyMh7tNm7/V3Sji8acDGA0CmEvkqiALHkId9HtGFFpNVGxPMdosvZ23izWMBVQ5
481ASkOmkt6xldtD5l2dgyOctYHGzBI8yCD+LtKzb3pThKhrJMTJ6vAIJzl9vtEshwTGVKJNqVxu
4/xnbG5N2p18bFhCYPPGZz0MR8FQq/ai3HVfnnk+7LmkL4AWTX8uzTliKtW5w1Y9FYBGdvtv7R9u
isLTx76ARQlEHxWYZw6i7Pggws6sGsmViyXPG/G3PC1ZLx2ilfCadmQsxcNLCT3pWIQgrqlOwCsf
GF9tQNJ0FO1VlLnwV6jOEJfCzq3vSYRTShyQkhh8MVHYeKBkaq+yPZeu4buPpBV3JULJ7EXKzGco
HTEv+CvEoEAOy0WxpLRDzHZdWisM8pe8Qeg/u8X5o8XzeuDEmY8oKGyOFp72DEl1DnfLCRsf/maD
78SequhLX9/c7oEUYL5cdjFGf1+hp4fUHXn5ehZnoerRh6yy9O9DhdgwwYvBzKXajwD4OOj1xbpq
J4SqEkDdWZktGwoCTmCBGB38qXSvPB8UV59MaLTayNavfqoPCtWdpS7fYBgsSef7+Vwf77Ioi50h
xzRub/0P6pGjtw48FCI5fWIJUF9B5shPz5xDbYlBVDYpyaisDOexRMIK9e3AyBhchaR4bRT9Dg4w
9CxmDi/fSsB4gRdtslMcigzD6EiqzDkprGAVp8ci6mfS5r5ioWBkH8DcYEUG5Bt3hD3YEMIT1TBl
NZhk3uKvFnk8ajW75JS9PoBoDFQIYtmBQOPtwPYqk2pcrjIi6fy0LcPtldmQbwg8hpHtz/L8dxjf
1llTYHXRxfTyLd21+/dbQlmI5l384DFi0Dv5e19XMne1ziZ6WU6D/hEEa1pWQsDa0dZfMZb3nZV5
DqwXHx50nixLBfEFhKlr7OwlTWGvAbdq13TqFz68ptpdHNOBaVa6l0WtJrq4qfXfjlki+3n9CbTs
a1DLGkYSOMDeHQOXY8+AzhUX66DcXpoOMee3O+VlMszr0muJY3w1aYYrdcTT79F+eJzie7/zKP5S
i6f13Jg2v8Nd1ARG7Wtq19in7tejGU2203gYvh2LsfXKMTl8ouXn/8f8thX4FnhK3KFPRBEmchcR
zhbLamvY/iOuZftfILEY5MIQQBKqJIuRSi4V7HI1MG4aYff1qFei4/SIlMSc3HnYWcuLfSGI+tQo
SrvQhptJM3KRP4U/BeAwYTbaX44P9kIHvUarKmobBUSpP0V+vX3x0qpKzd8CznXPW6LaWcR8IJ0T
GSydgpixFzCcFgY2fVTZmO4xM78vkvmqNInZy3b4BYbKfFc+TPC1Y4aT2Bp68pHmh4eVy+4hvdd7
iw5GvPUIz8vuXdAg1/I4VWyBjY1dpF0I05Rcp5/gdU26mzolU28BLXoPQh8kmLud3mF6sEvR8MuE
CSWIHqc+Nrkr9OkKrWK4ka2z0YklSyTezKY5fk79nt0R9+oWjc9OP5bzjB0m7XduMS98wEIzNd9y
8lFDldYt7MPB+Pcj5E4ugcNmlydJgWK+dWZcFLKbVU7j3fYkgRIRXOuVQr/KBywqxRbA8BgMyzq0
j+wJ6EHbDyZb44VXSUcB6wcQWo6T7JsDg69i+Wifzg5JlCt6LHmMii7Fsqg/ruBXiWKlXVPxwRlw
XugPLijKZEPo9+Zt8iy4q8tJMOYeY9oTIJURftyOfXqkveTRHZmhsqn1/qcPFbOZgSA4Xo0PLxFD
FFkuQj+B/s7fC4gV5I8mIU5yMJUEROWbmO/rMredEJqSYb/hSclyC/osvbMSK1Rw1DUxMDEcq4Ut
wKKl0aeAz1z9jzKcgqRYsor3CXt4PEfmfkESWJCvuyIY2yf9t/ntPp4LBHzvS/v2VfMpHi5TqBgY
frSm50De6+yOBl6nE8kbmDj8Ba/rGcTYda19S1YkNQRU2awcGTN8mI0Jf6dr8Syagebunvd3tc5/
NdJ4vLGll35blY5yNxQ869oZkaAkirw1dMIndBoeT6HQy5s7L/JGmmyOkR6G/GfxaxNkp9R7bOC8
9sYxUzH3v8xEZlV/bdSW88iqcUzuOOZbgDb9nNh0uMLqA0PjfYuy+tWfv5ecMVai9cmxsEm2BHYX
2AjL1vkCJyFsEt41+mDV44waYl+ULJg3tT9kfco6OKX3Z101FCL4841lF2UkbKG0vgS8fEZ27taF
0sbNIwdnZNu4UfNLbIsWD26yvncW/gRkSVOcJlb6H74mYJz7X0dcq3at7ifd+Dxk+lhgUI57FG6v
7i+MCNhu9ofLa30Y+JngLeZfDOQXL4pyVnc1GWEAlVrUjhatUDMcjm8425/tyyyfh4fabLZCd7DV
UObxhq6ipV6Xv95dJ48RDBLC19OKAL8lp0RinyRM0pgl+xUtRbjioj2rep/5qa7FTBtq+gLPriz3
ZWNkcom1o7sKudN4DjiPrRnD9SH0LGgxrTe59M8FHKe68kUcXuJ/beafALgeCH7KN+GyHPowAaO2
NzLD1O4gcK/rsAFgsWjZJ86NMrEl2IVzXhqL490ZeZacsDhcgXDuJQf5L9Bp8jzyDoyFKmKflA7f
ZMROiJum88thqh9Dr0ChKcMshly/yQj1hy9mzURqCyQjYv+aYstnFPRAN7wFg/ummswUtFRoDn/+
+FjpzM0tU9jRVHe+/qynLVw3qB1oVVCaz1H9lWvHspZ5NXkk5qkFz6dUd9mFVxGXdk7aj2Ixqsqd
9M0+gUjw2a33OQJZoy0cWudkjWpLOgyWtRZDRIqcYcwlcWakgvAMuJ8SomCDwH+SczXcabzkp528
RC9ivKI7QDmWJtukyRIihWhxJvTQipLbeQGKkDxJ5YOyYdhWfChpf7oM/RZ81TlcZ6ml03kV6c2o
n6UGX1n8g2sajbdxD+yA8JSAL+3VIDdKXNpcr+mv70Xw8XjpXRIA2XG1uM0oCN+1xzJm3BZui46v
1+49fV2/jPIMRiXOMJ+kEdrDX7m8f1xLc2fZ3Ee/pVOiubeTViZuUz95PTbFGvcRga2O4f+cMjdB
5f88aiq98GJicE3GXKaiBIomNnMweh9uaJ4l8+U7AvW5z63OY80aD2WoaE2iVi7WviXMLTLY2JfS
WoQonn7jPsctmhz4KBBCPEtjzx+s/HA6pyF3wW0v8ewu+6EG0l8m1ArIYDzOaD88a1MZMPE2BbAJ
g8JPw784YjCNycSVwYJkobyLCtFE1rMtKq/J3aaUQjWeJHspYevlGOlsx2ArnhmnTt+PVn5a2B3G
7zrHxFZ1fCvp4SSwhmi8E8h/mI1+jC7SEDH5vM+vz617aN3DgGXTbWTbBuJ7VSrSdsZL8WUQzqnE
nWvB4wos7G4TPuNZ6EfzzcM2lk3K1+o85eMEqCdM7rVwJLn81KqF9rw2M+s3n/YIZCxHCjAXUcjg
0FBDBH1NAsPTejstwXiJLbQZUoXPIm6JO6asYWOmVABbo+sgBK2XvmwtbAnSQvMYolfeR6IuGKiG
X2fAPJrhOnjkRAn6RuM2elt5IJzz0FiyV3aQ8Y/VLU47GyC9TNOyZ3ZTOdFYx9LKnbJ0JFNzj5nG
wFG8zWFH68ex1AyUSTFpf6GG7YUXdBUYJI3QexL3GTL1txzJalGfA/IMGQ6W/w2FkENY1TskOQHT
jpOBSUwLSCrMFyfwuzHkbDAMcjpxwgvPx/Xc7bxZYC9TLIjWblYPgNTpXBeH0BX40T+vRZE926Q5
GOrtohhgNCu8ZpMIHrslQRLb4Hq/FpauKBcfS3LvcSxGfJSXJ0cvvc141NHPNzov9/CqdpLGORDj
I6Lx2608RcfgJiufL/Hu8yXFEG393fpomvJkginqQ03hFMrzWd5vdYXbZ5dOA3G/IYqiQrWgU6CG
SlHAkLRUhPYRhP36AV6D0CNRHt5msqKtCegsQMif+VvJRyS8M0AqCaBN+Ws1o627X+N6xgXLc/g0
EAex3uL3nTWdODRPSn0eXlAdOXzQTV0DE6U+tbkwmiEDK86TbSg4ETOmD6fDVWl4e0LI+ZlXFy84
ddWfrpRmGSEBpw9CBokyoNGJvaIwgkTT6cb+dT5a3QgWLJ6YIDLFAAoooqbocG3SxkzYvFkSZfIu
/LuGKYLwRAfcQe7zSb5LotQYmTyp3Bwmw7Sl4YIBltmrbWISnIYHAVf4AlA+8kl0JpFsRunP9iNd
gYb3rzJwEb4lTjZ01tgrx8v514pbTumSWmGyrDyYmBOe13Hle/1iYDje97fg7mSzUxVAjKe89s/c
ALp2cHo5jpBwa49xWhWa3uu7pISQypRk+oy3NxJ1SDS2J4JuCLjrzrWoW7vxBw5lVtcMueQ2qzJG
oQ7gbQ8dN5/NV3WyB+zwX+wmJQzvvxD3RaW7RlGIRkM2QktAEi4Zk0c/FMT4YRI863lUybvBZgBb
J+Sky408y44XrYFTCzWW5c9/T2Mi98Uqtg07bjMZP9gTcf7T3TcLzj1J4XLVGsEKB14EfIfbf1Vt
XPYIAnLOOWfzvQShZi7zpAOrwuNPY0HI2Re01RZEYzht1MydodzWZj9wo6tZYI4LsrgtLZpwWyLa
huwbdOp+ihqHKfOaYSct2V1KU/P9xWUnyBTKKIaBuRlOYIc1p2ngvr9yJTClZ3My2VekfSaKuP6l
3F2iu3BWdiY1avdSTd+9oFk1GWC9R7TWUtvBagnkVMwawxfgxycHsWsUPl6MI+Mror3d60k8+xc9
sPLe3CGyXnJcxl/SZ3pcZzqOklgeHKEbHElhzD4qg878YW3SJLE9rxMWb3d6q0GJU7J7NlnmpG9N
BcTAi/rvFDsulzytkNXAbIBiWXpAdNyOafoC00QAOyfvxZZY4DkQYKfBZrt51Su+QWcO1FVYvl7p
ryJWTd2AMoCp4H2kmI7rGGJuf3/aX6omG4xSqZKwxUimGYkhn25lwA3VN8JHYG6us3RRO/e4RvWx
uftFHNzWd2+6RSpk9TBFuaCPW6FOgI6llwK60OvWhXQmNsogGm3EYACBkfCynwfxWdIkXgycxBZ6
c5SNCt9XNGo8L2nZcHpOFQ48mQ0p2U0dPy8ASh4ncBhfyulEk5FLGbdbvAy0KWug3coBvmsafIhm
mEgrOwoP4J3jYQ0P4t0BRCEgfYOHBJYLqBhWEy3o+/+Rz8ZjBeTRhueSHLiaVzr4FahbIoJD95kr
DO6Yr4009aFAovxbFnjlZ2I/Ifgvz/2QxerQWcIRm0QVh2SjlQWkaEdi+jw8PIC1NFqJFebyYjjH
aaBYfPcZG39fJvwa0ulteJfns4A+oEeHQaxoo8p73vpEndUH02RgmQ4QmNZKHu0fVs2a2IjAVuKL
zQQsV+BJ62QyREgubyQkkJVIzRmExtfUMOZRcvnIHppqcYVNN2FbkK4wvIJZwqNjMZT8UPI+7N5z
SZHE/Xpi70holaS3PmwWwK6nMg8AY0FCb+FyQ8e1CTB9USBJym5RQGJ+1f4V29oE35pzon3XIdly
lk7YAh8e5j4KTPsTzPZhTQBa5l5k/+qHM+yOtybmM8ZIMy4FfdWNpmrFXo7YFNJsLSPHg2WWfjmY
aVHeQE8m5CUQWmW0Iq++TKhdVKe1HKS1/VkVSLZmR4JEMNmWWt/dgLaAN7eKr03ezfhGcRexaCPx
V7ywrutwSZZtVkiMlDz3Is4wUTQftHTK1KZWMWAfNOYOCK5e5wUcKkt23pr5yqRBw972h7gF1jgN
2PlgN/cY4X7gBwptgxIrChyPvqBnDuXIcQtV8X/q2dDxEf+pelQeVw8KTpTjDIIxVPieIoy+OscW
RZF9uTTT8zn82spQad3q/sp0zguLpCrHoDex+tXf34Xjyte3ROARre/EpKsNPgHN7rwPJ2L7dcgC
0PTaXAUyagdX/LCmmbnBwgR/5dM3CrlUSS34AJFL7ljlFLJmur4395xyX5cdVm+4di3q9dAUx8DG
/hHF0caKYdPgAuyUcDnXDAf340oaoMHf8SX/gl+oIAyD7U4OGeuLBgF1sXxSsVYXzI776lJl2rFj
bffGvylYTNkGkJbZJbDzZzKrywVLfg6lmDOS/AGH0PZ49K6Br3PJ9CAAO4AOvdvVwDEnNRbDR8G+
E1M7uDFxxnCKh+WnOqtwWVXzByYuulhv2ijpHk8NJkWfBBkRi6iCIOMkn254nQ+jQ/XBdmXITt5Y
edu0+mF9ldpswJUUHrHMwEMbl+ErBqY43scONV8RBfywcs3twJKJrZVoKrm1b7GQKNLFdyet28Oj
CIpOz7GzFmBJujZlAyABfN789HYy05Em44ZkiEDKHBBhde9ubrKDT4HUG8XfgYeb/BCuzx6xRvuI
Mf1cUSa3JxqzFgda+6INNy3cpEYSEEQWF3TL1yTwSRREedw6/zqeWeoyXMIGxcMt1EGijGO8fWpk
6z2RaTXYzI/G3Uh7uTJFXUVc2VzOROONFnz28QMStxKs8vdEQyIZSbalK1lPYrqcoqR6eJOKfVIC
h4rNN75x9QKbJOvG8fDseVjgqvqva5vDdKjrMYM317tomz4xAqt9voiKKenEV/HIHQRPVaNuk7OU
AT5uiD7/l++FNLvgnZs5t62bT1ohQ156mTYTozqZL+fbSnFYjfevzfGiNbxOPm9jhFK/s8TAJnin
COZjoObmJgSKYNFHdVY6kjvcQZLoaK9V6OfidQRDZ+nwPYpNBF/am2Va8budkIKXJE+rWQuYhvtX
xqjpAL+VvQnGCDTR/PHVcJhr+lwZKiw+q8Mof7a4CoSYkeiZJmjz6h2dt6wBMeDzweNL3AVRa8Ou
vSM05gTeni2Xm+6o8vosndv0D/K4qgYUiLiVO+9uLgc3MM8PAsaI/ph+Fcu7fpNHD14ZhtT8OwBG
ns9/7K8VZoJosZHINvAEhE2CgueZeyy8DycRZrKK9R+Dg2rNkplhO3qJhYVBmBySS/HU+b1RqK/k
+WKZCm1YiCDRTzhmEGfKDS6IbMTv8+82oFt9GaUKWL/EwRXCJSbSCDmYC7fzVc+Pb5sD35VolTLo
oSIKDHlD+KfBkzJnSds5Ph/EvGzRb3eIjdFfYzyrNwTc4QzZ0Q2gtXvcyNfza60Jt8wf6WCH2tUI
2C9AvI5rEN6xeC9p+sRE5KiDH05klnKNnq5+5z3SEgSAi1ukGoZmS0iRY28apo3T3gDeyFnfMb9A
Q3d+SRAhBQRtUFXrZPkA8A6VewufonZqGhht5iAz7MHcKOk5Ghm3CMOAGw9s+Mcp2AWMq/mRo/CY
Ql9/wuckgH7BUrcFxc8BXa5OAa3wwdFzMZbpuPNo+GcgX7PENVPhDen3qtxVDSgMhpfQHf5ADG8n
LpHHZn/N3w2AnJMc7YRzPNNt9FHWT1aLCzHKFsQsnaEakXWV4R78CCY62IKvCLcHMXtbRPAE+wtE
RhBkpLUU1j2ZahnZB8vtAkUhe4LrVRznI8SaOcKu0vnh5Mjaw741J/1PQ3qNgMQ/YEDw4WFN8dnS
GOgJ8vbFdxepH+7kzMIkLUvHM2sE3UciAR7egUz0eMnIBbmrsOWJDGVPvd+lvZchtV4nbhkuyEP7
lu2Fq7wQMNNBsqpiNUbxWlQh49m/RamqnjkRRHu4rs2RXAcUd/Z5Vmgqyg3m37uZI02BscPFkT3p
w9e+mm0PSVm7P10dpXz21WZcSibHGPK/Qpf4YBRaW4zrBMO24+UeoqlNNrMhsGOKHyaia9wmngal
7IkE5kpsvd4Tmeit4aV0QOw0AjggHFGhOutv3wFKxYKUt6AROoDpb8mN1VYfAfZXY0mGi5j1HXta
yoVSNLJU2FWoZvpVcFggFySKKIa+JWqHyUuRa9zBn/4tMkJ+uXWWnMhQa5NVIy+aXSRSnCYxjfuN
nUsl/iZFQ+DdGdt1qqpNb8aAEmwIb3GyNV+02tN07hF5LlRRIg92RWA2diW08C4H+Rw7XQzGho3o
QfOwn/qZ1l1G3tOHbpRt+hu7rAdGOhnGAl0tbvDANPlpnIdQCZK8SZW+Z4Z0hiAHYKtDkuVTBfdE
GOC6rhkj6C2JPhDvw9sqrnUWuWQ4KvVXoSez2Ja8jjprGIXU5t/AeEU6tfvwBIi5MkQyJtU+9yGD
Glx22BmjlFqy4xpMAjz3ZBGHD9j1wjJLNi+oYf70aIw8035Kbg0IWUqIr97zppZLEzP76+pZFRw1
Hc20aOxlvb806xkqiD3J9ns8VoxXc0d3HMDHyBTrJjCZG+1pn1/w2N4rlFZeJrN2Ww4Xru+GZsko
nrXi6nniNdCGmwWVdjWJOLw5mUULxINvqDfMxouHwjF9xK2/qs1nrJHyggZ2SwjD4D//k0UtMbVI
NGR1uV+eejE+GZib0SM1+zj313VtMd6n295V4BLgPgcBgfYbmGaoA2BrnD+2OQfedzlc9haAsxf3
GTttWFRfmlEB0gm+y91kas+1/zAfMRRxr0mXU9F5dvekLzSD8+ACJRebWXzsvTTh1QEfXKz4coTh
9ZkNVyzlX+JSaDQ08q0NL2TbL46QbeozeKvjse7io9DsXg5zfNqVgjjPRLVKXWI16Fq8/O3Tvafs
BBwLgnFvWvx79pUGxuOodbIf0H5b1lGGGfGQUDHtArfIHpcBcdUZCV+7it8JHkUkFVyMGn+eeQxm
dmWivSXnY2u1a5F6OeIqVYMiy3nQzd6fOqNYWw9PUrvVpftNS5KSQ9s1rQ+a2o8BHFcG9wjK8zlR
mg79Z2xRgiD2UHheGw1PjXizyvNK0kL+UBXGzPMjpBKxwQA0AU3UBsZPIf9v+0NwjyxwM8+7bJDB
ytEDyAqAXIHjjY1iguAnx7zGwMynOjL8v1h3ie9nYMUzsiGzYxOJjpvihZN5hR0Cc5edDBcwLxd+
rdECeYfAFlQaiiuv/uSmNFu0aU69GVedr7xUPxvW9LfvHZFYmVnhg8sA6EkKmMqVw5HpM6G3zIKf
EKP7mQSgFk1u05KKGdKJF7UCCDmYllhNwbOZUg2hdr9I6yIyLWBAPiNMAuLQ2KeKKT5npO3r7ebN
vjemRF+4hnAqjPjsSQ2HYROZ85XFf6p190HER1gaYm5Gicx8Z8y3fzE+m7ybS4yXjPxLNj/OfH7z
o+aPxYoA+D+xTvKhFQ37/vtCQhrljpX+ttOqxpz0sUQYclDf1XTp3VBmTmro9q3wl5juKjBzFnZa
7FiBA2X1RZkYJHQWGbIJEbS2J70gufIMl3EOn3/WgJsuyO66JxkKr6E9AUGwGaW0tsWRg2BJZWFk
cFrb7dRQhDu/KQ7r8XtvEANEiEVxyFSfzxq58MM1u/toKj007P0sO0AEBluK8S2gad8zgk8V1+9R
iom6HEmzAwjdbCU/r5TN8CsXozH+NHQAf9v3EmbfMxgwKBwczkeqA21Pkq2H1qnd8TGEarYohKij
f1zvM77RcInoVYnJ7hXHPHSzbxnZBwf2EAoeozEt4B1oYDRku/FQwi56yWBcis9YS8FNb5FJx1Vh
grmKLR9UI7omB3bVuhh69tq4sh6J/CSUX4Hj34WqcKlGKf37SWpoAerjVoF8ohwiGruW4+cw6zBr
R20HVUxUJfd4CKJ0HQ+o1EkNeyqsi9Ve1rkGr/MnmBdzagVOPZytauDN3kNJR7hqOzGPYie/mitO
tg+FPzaW8/QZVjETd6VeM5QMkzvhledlugzhM1FYiVa3BCvk8/UUYr90/z2Xx9Py9ASbI72rLSSP
jK+hXM9AZTLaAT5Ap0nNxeyyZtwmLjmPc9No9wVoHelgftavOdygNhhIqlmCD1SP3LJO1wQqU74r
NbpYXgDg2zN8kx21f7jmosVV7PWbCInOFEiCOscCyCpey1aWPYGA97z4L1SQXhDwaPBX1Ad75d2K
ZuoaetIZRaoS8VrtW3NtanwvlblANTZvVoDrIxQ1dBLc+R+M69sJOYg+ZnOsybak0WfMYOgzFjUn
UDzW3h/JE2o88tfbXahOsz5T813AVLl4ocZ6yCZF6gDdS+7tl1ZQnQi6HIilZlgFAx4kSqBs8Pi1
mW0xg3+Df59ADq5qiO7E+jB02nXiM8AIS00r+D4bIxR2J6Q7B8QxrYMG+TXa/KXjl8yTqz83nSJI
HiLeNoiTRWcfQvmuugsG2oURzq7qlJPyGms6MGtwVPqmqQos4yEsAbsL1fuBHmIJl+Py3zCuGzIx
HnColPYWo0GPKoCNy6knwba98AeDfWsCCOKOj3AA76zJLDFnINxU1gawrks3+Qt878YVDjFIDJ52
0o/w9DP8f31MkalvqICwGr0fNIN5fCBEcUNgQIF/IpTzR50jizUDM2NnqVnzgFOVnfdhm/Ds6KrB
1w5Ucf7pae6h4G6eg/0fQcyX8o0Zpc9GhEIQ0m/diew51/RdgI40ALYnMTPWmQDoG61n8a6kV4An
SDBz6CT0vwcqavtM6ZN6HATRztSRDNGU6LeA6RbD7J/X+K6mKp5MvZM/IPTYeRJZwVzvPMb2pUsu
bWvJbhPCyBB4ms+q5hWGJ+2FtKQRH8+atgIxhqQo16+cOTUHWkVi3gzYPucR3ONREuqCMDFZvzrG
Lp8CmNfwwPVHimQxosL4IKUX/O/c8/fpU0p7k+sNFIHxadJ+gh0LmBkvpMz/xd7hZos+udLM2TPy
w7EIw4z/hY+RNdGIZp+gF+ryTdsdMOvewBn/Jc8ffh7CtudP4jpM9LqiDMYeqqjU8Jkwil8nWQnR
vYahrHQ2VqK4qayLXl/n/dhdQ/pEaupc56BVDRfYswIMaQb33XTkows9qgSjQ0E524azAX96rBe5
eVR92Cs1TyjcBr6dyxg8lfgsP3HSo3eB6zDi+fGDoQUA2wKP/k0j2YxIgmx2uCKlrivC7qshXbeq
T1YT/yhZQdI7L7JfjXkb/oxUvBw68Ec/j7lB7femNPJdFIuP7tye2pq3H3zpBYjTW46u+nS+B+Ol
K4nldsOnEFUVzFVPp/VbAB185qD4WL4yHUuoyogWnczkCQa6eNrJmWqhCE7NW5/0NEqPuK4LdHL5
60uprf2ijxvLxjsDOJ2GQQmKNEfEqYt062QJBsj49Tq8UrlZw4ARq8WPXVTGfOxcg6cN7npCgDfM
1Ub4PO4o1+WmN0W+Ggb1wejn5Y/p0RsrIY6RE7OQ42GDQkxu/ifEuV1rmS1Ahd3MdrhRbJ+kYkAY
af7DsAlUJ3+cgFHrDU1BeFUdbclP/aztQJKR7cVaQrGifnv3M3CL5fpiNS2X7CupNjfe3UBLMUde
anetiIpMH1fHZjo/b7GRVbTFGOERvj+4A8z53L6wsoWZZ2iMeDqCi4OkgFURWRTnB9oiLD1B+13E
B22Au6pCwawdiAFsSyYiKr9gTnPZXEh3HIpe7QeIK0Zm7FWuCX/0a5CrJrwL2ft3kwzgsxrQNstV
wPIlh5RKsT21Un23PCZ/9vhetGMBvKpJ27IMD6n9F0XjnYCc6ESGcWKpOeBhh8h4CxGhkBcZba/4
uL3E7iOBghgOdjisHUbuePL6lMaU22toU08l+LBxkHBZK55WwszL804ez0ONJpsYRPVri1EwE7HN
LHUsxiSd5APlSTq+onidZJtv5JQbGEE5MEYJuDsXbC5P3+11OiwipvwWZ6IzVBWRZh50WtuRRZhe
E3FErAcw5FxiRkNHbrqddAgkF1xcjYJEIxbHeYvsfl5lJ33kp6PjfivhVZWq2f0NlLSWHzU89rbt
wp+f72+wuxwJsC2ZS7/ZQdoD/mnwPYFsVPFu8bbBodmK10KKoY5LOnccRZB661ImsEmMa/bJ0gT7
dW2owk8fcVUW/8U8x2/OIxZUS4prYKxtPdsyFDeBmcSN+Zs1GfB0QPfh0nbGfOOnglyXcc7vR5eh
UnaD1jvsP9gfmNo6TyRtyD6159xOHie4fLk7xYNsZVXt8yelYYadjx7LmkzV/B9ZKkIMKm5bhxG+
b5O/nJLhwN31kM67VxFKWuc+sLb9u10Mvi0OHZMhJ77qmyohR+meqgbhISlviTxhgi/pyZEZqeAR
RcNJhiDcSQxTmh8tcF4zd3yR3WyQE3AZHB6tMU6JKQhk4h5Ea0vq8ZyJO0tHZbYsL6xTy5n3Sl4Z
iDQdtc2BQWrMBJUAHjddxwHX4p2qywbCQQN8rmiXfsqlSkV7S4tkmruZ5mgdDfloFf18Ty9HHPHl
ZFUEe4ZBQfat/VdXyBDbA1xLonE11NtDdyoIGW9wpVOZa944TPQjNZ+m71fHPATjJP3+88UW9Tit
V/V/bRUULITq4jE9KZkAx6xYyiYZGT9ezGVH4AUBskoahcjNOkK5cVfK204MrBpbgkCz9HhXKZRz
orSGwgvCJYM/4r1tlEuY2XEHikvh5HOgGqCmtYtDLsZpEBKt/rmrs/dPsO1P9dSbr8++72XkXOR4
oLoBddgUr958iLji11zq6478NiEaqI1dpHXN9bzHZuxyWraoi7mdsp1gOh/QgjrEnNfQLJr5Ap6d
c7cGDIroZyhcLh9/f0aG2auT/2GEwsAPQpxZ/k/9BhCiQJNuZpS6QgtTcToJTPxxls4JA9O1R+Rz
24riTRyWQLNVZKF+yA15zsAtvYIvWKDNmHcbl3SVVUyKH0zwOH6poaype1OLecYGG/GFn+vosnhZ
YhscU0JdQ8V/bY7tFPt8EEpyQHWFIFSVkkxX0sH/dYsW8HTXhPv/kc9Jg1/V04NP8FQd4H450kxw
usyvB3TE5Pd7kLZGGCTrApcimK2Q72APFkGyNl+CJ/eEkXxqGHyjmCBd8dzCIcH8h1mY2wsOThOz
ky3nJ4OYqSrQGF91jdY/U7zo2qHSDRdZyPPzYq1eGuNU4HCjcioH48tnpAm55q2QXYaRrSgnaT+N
/HH4pDnUyEjhmcw/jxNl+uLaQOxE+VqNhUKalFKQ8JhUmQvfw6Yv+xNb4HRIACifWcMHZL4mhYXB
l5gz5AjMRv/41fICRuzO887qEmNcvcE/h6Ks6SM38qY2MhFzTEqLJ3xPapAO199xxvwwp0hhfAvm
XDpvyOBF0/ouOUtiDSo4eBYCM3g8M1xkweNJhr0IN2xeEdXOd5R2FxlyqqzSuGxubMPmjwrXo8UF
5KoJ89gEq/0Vjs38KiykON7tyxKZgbDRDjzIrYMtHyDHAF/nlLIBn97adJvuBuemV5lH/1NU7uLw
2+G3kdzVSXNiJhNVeMDeOlHEc4VR0LzqywXrPL4SJK1sGL/ooQss69VsgK+SxZWcA/3A9myxKq/J
SNLH5zNN5ueSxS9HQjh/eF4LsKd8w7U0oifJECBVsplxJUAyoXfzXAjKcUetzhpcEnBkd4gull2g
hzh5atmnF+p3j3dgueEUoQvb+xs2fjtTw8F4nnRS34XK+PWnO8VGxQYu3cDvt8iYRmMy09kUb0+o
n4dZviuF4rlFAT+dTy/V9UkAQ/jGuxMm0b0tsDTpuPZxpqbvk9ryANs4KACPJBdtbaPGiy/3IGFd
eSK+BG88pg==
`protect end_protected
