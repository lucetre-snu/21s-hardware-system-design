`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UX6PGj3SsvCyCs6e4WTW/JyW6bO0ab9htopBE1fpgzTJaJckW1Q7oPDnbjgu//RZcJa11E+3OMah
l1NA8Q1Omw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rTNLM41zRn2jlQ7+LnYfCHUhUy2hjnJkVIwrVepRRi4ivTmVgYw6JZPqwMwWiHFpud1djXcpBCOl
7Iu8ATp95e92ukyl//KHCHvSAsQjWuYtwlO9e4UWLK927gG2lyV7ifM4GOZ63yIIdpEqOugLzbKE
TuK2vaI3HEaIvXPaFCI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NBZjFovwJ6Ud4AurKWrTfGaTSetfP60XoKCw6c1otuyw7Bt+uy/Wb0uNhWyV+Uc/FjdyZxHYPrq6
wvv59PFvdZQctZ6H16nvIBY7p6cF+vvvFPaVElH19FvZ9VhrZLLt1p78FJVXMPBt/n9U8/TwsvOh
as42T2GBFzwMWkIF/kmL4N+KnxDYiy/VD+fsk31IuRy4ilDRrITpfmKHw1iZPs456Q5t/JDNW59P
cvTJNapo3YC8XIY2dpq6lSsNTLlL0nkbyufC+kTIDhhhu5MszatagsUYBFW1lvIzGxRZQyf+pujk
D/nFXMNtxXzgmAxgrmb6he2M+RIK7WOGJIConA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FACL7SADPYaVcXp3i2t3xUzgHH+p99cDppaqGEP/aoAmWVER6VAzsdGol2xqIrPgnRKVT6AUgciG
bAPPalrwX1bJeXv5pB+8NJyk0vmOpePdZg8puhNKSguexS4UmrNARBjOkoyPNd22WzazwhV3eUN8
IeDsnvCPEjxgdIxR6V/yIluavd3TmB/JlcEqxj5rbn8KJeSEIEuVJuj1g3O5evgTaYIUh9nVsu1c
UCsNhbJxLJxaIvhDJcmYTu/liJ27BUGAd5vTLve+sgv+N4DisxFBdly1JQha92/JsmDVIhhYWlRN
aJF22OFr6Lrec2f2GxpLH0CyTuTmELTjnVD7eA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YVRBPFUFI1nTGao2WdWdHYr94pFLkHltHipy/MwLeW0wURzG16qFlys6O/D8eQ+2KRpDxWqUVmNZ
TliqNJ0logq5y8O+sYWUnNVGK4AO6nMVjgQGneyAIk9RTw18Qow+jLSG6UpcXIQ9gS2uuFecxyc7
77ryH4/SZyMQfkL/JY4=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbR4iEroecb/C4aS3sn2HvpeKitXtP9LkAc1a4kbianUqI6UBYgStnqXOJNGzI980S70aIBSdQBG
wein0qVBSe78rz+ESN889uk0DzRjV49jDvZ2zZY5QPnkRxc3mDuAXa0Qc2RatOHyOwHydZLCklll
XqdRG+5HklDgosgTRryGyReNDiW4Q6g89IAocFDapWgEn4vYiuQF+no9+Y2MGuwlI/p1uITPGyF9
jKWeQUsz7562Oph3YgxmWJZEUTh2MuLeIPsk1rQS9xlw8FloFxLKR/0ZzqkB7NeNFTMXEkZ9a3/Y
/CqtYZmex3OePoiK8WrQ/Bq7xhQ8Qmy0TztDUQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f+jEpcDQBsSK8Q/3lvmrwbGoumBmz5PwW61HVL0Izp+3fFJwcv0eIWmyUP+ix5TxxmB7LtnpXMoe
TAxcrOK6ozpJrqvM6hZl3Tvp3T1GrTgn/iSCD10N9dPKVrC7fUk0DTBDhUeyqTbWlXzIy8ABhs+H
CUK/UiA1D0qI3b4eDepd1YkzbMwkMPpzrSPlCBoxCKCMbzbCwVDE4r4KPSK7FkczWRGbQGIFMN5O
snv+oELS2ZUq7Zu6sHfBshTC8R5wu4v+OpE+qZVYjwC7YjftfzqDtfFYY/oMEq4Vi686d+3GGFl+
gZyhR/mxNviMdhUr5LPtpffXBm4SF/pAmppLgg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fjUcRM3U2iE8xCUymVhRo20elwNzAeA5+pzpqvDcgTODIcWo6PPJMkf2NAY3O8D48MShQ+9vWurz
LBwkZ2OPwobE5AlVOWprg8MMOdTnI0a0cpkAnOS8M2K3aj/XfwhUS8kO1ZZoonTP9xove7krs6v4
QnIPw1681myg14qLdpHYU5eSfsXGrqqWjRWpCK0qxOgbJlkXI39XHJoKAlrrAgJ4Es3ez2x1/nAz
0hN47Dsjx+TPUd1xPpjZLH2qsuqoVw+cJDBPPxR1QrsPy/vxELU8VlWthX/2Gxvt0eKmZStFPtxF
pSWgxInJVoTyk48sNy3UoLFzJX1GIPLEEmJzHA==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WaCnqI58LQKNeNnpRG19de53PVUJkaVUs6+PXM6O6SoAYNniwtDNsnL9fE2sGwVme2r1xzdSTQQM
6k+4eaLeXhIOYq169zjhAhp54WtgtKgIfRYoKj6Mneekx16BHzWK9rhiHpNiJQsOJpiXvyEjg6Qg
PeUSbw20kL4R1X8LYRjleN+wRtNgcTE1wk1iSrFUbqhd7ctvOn4UDR0vk0pA8AQrjqwNmsrylTiE
8oElUf8lwqFZkQ3QteH1K4F7P9CTQRp/pAS5gbpYFUrRqpRCKdqSnfxcNAsLRIXHyFKtXiunRDoz
zyKeKoO84O10/534J0I9BvdvlfjDRHzf0WRc1Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98368)
`protect data_block
UWlmhOdpAfVh+y1ncz7A5PG/HnISFQ98wQxgH7CkEiLlPqyqDEWLbaPS7q3IFLm9+H9ds1l+Mkc2
iV+3uXSq0SqPmDnBDh75Sn0l0ByIlJj3WcbI/buoDmg6bcKPa+tCFeyZavsOd+H4Xycb4VKYpDUU
97YM6qLO6GseZIxAtpEtrtzBGQExnSmAG65VaBohuSBEQ2PcVLl6v9I9S/UO72Htn++WNVQ7e58X
dDUAxXr+OUAJVdfKgnFtQULgg7ZsmuYgaNBUkRiyiNFHJKR3ZLbDgu8++/qFTHEIO8nzfPggBshY
lseacBvKryCWCKt7w0BAyxmzsX5LCCtkOojnv/h9Tb1RtTWFx77KlaW9WXNfAn3rZGB8JN5UQvEO
/bLDaYsOPKejLpfX1XuNOmzfPVkm7qOF3oHQI/KIinS9iMCSIUzR8Bt4UXR8utOYa4ukorM04sy7
zctBYSHEpSD1n3htXaL4+M4a40oHLwA4rSmjzB8R1GLa27CqU7vVtHxvD0mdU6YQqOCE3UYQqwwq
Ca0xhmFg1ivorZtT8/97vbnDmWkXNhH7qrHUNbKiO0KVDQ3fQOEvLAC4nr5lzSjYphHtvNuva/BK
WAAlJ+PhSQjii52TexT9nK0CAW20UO9/u5HhJT4IV2F4vMJzzV0+FOikNYFnC5CrMAirGMB9EnKJ
wk5eB0qQnV5eaOoFzgQ1AofeH1TBU5v3jBoQ9RF6mt9RGHlActyI68oNJUJLgGx+OZrIMIZvqooe
yi9ucCFAn4AnbQEoyHQS6oun3OC6L+UpmaTjn+5KqpjZeM1WpgDWFHKeHufuIhpwq6O03AU5PwpF
RrvQK33JrkYMLrvQ9LZZSBR2x+WDPz9cQPA1X5SMbWx0/RXzdOVDe24JzS8UvtRyWupVzWayenYh
ijZYrOioQrN3lgfb76zBh13TTlwhuwxD7cJc5EDcP+H2FygmbmyOwwvEaupB1tYvyzgrJ7y9HhJY
7icOMIIW2Vu1gk1r8AZzPskCh57PM/il/ydS3FuNLmiHayFP3ULc5UXkQNEje0OUNw3lpUk2Qp4y
jYiB8E6Cmjlos8bmYzlTxzL/I70Bn55GHCk8kog1O/nl/i2eGDaP+BKyIZnXN+zavBCGh/GeQ3Ui
DUkDrKVHe/tn9U8O6Hy2R/32fNUsT2ZELl3KASW0t9UTs4qvK93IAJ0eK9V1X0L+OLMML9jHqKQU
WP7TLjbc5U1Q1q9MSfn7TpbypIDb8X4HuTpvmTyphPnMD8sQQIv/RFQU5YI4eAgsEaGt7Vzdt5BF
MbnlSZz0fWq4icRLOQ+G8cja3yb2eUPWZcg0F/vLDAkbq91UdcToOtxhibfr8qD0Yol1eeMyyH+J
V/SRaqPvQKY/38Lle61jSLDdd5RC3WqMsl1sZH2Q84M7RQUoIRL0jv+pWkN0hbZyrKCIDcBCLScP
rkXvEgqRIAqhj24qHpFswNujlyR29SIq0BfZFEhq1+nLDMGFNo+Xyu3g+7FxLONvy0ilWwYuu8WO
A7rOPqNBVG3dftraYpltBtwEIXfSE/sbN5L8hWnfJ2dAJrN/924A8/tRtFJ2r1c9gAVTq8dvDSXn
E68d/hbwQhBSHuMUuQjdiEjViNTHsraJzWT/WiVVXFJCdMP7lQnzjsY0VInLZTjI+8ZnVovOeY6J
l4PhzhoBkJsszzZ8ylkCCFQeKJ3aNGBv3epQWl9G3fw1JqtyT6WGDY8R/nNYcacCrvZlWUoLm/jT
oDVFYINqeHyGH0/EXXC3Fq1L0yTKWnoxBDHC/YmwReKEbutzPoSaC6xNWgt9QMbsJwT/snrEscMd
d2zDt5Ph2KymASfwUiKo1HLQJIWuweD3owNAR0hXTzbzkGQgianZuqQhdzMa1fR7joyJGHw85Zsp
038MkvqPRTucZQpRbw6gxi4q0LruhNLjinzKS6FcAPHpoFxaPMaHhZxtcllHD2Fzr0sJ9sp50tXz
acF3XiXpFZGcAsnMAnI2ebe9l6mcH8p0wr3969KqWlJnWx1Lfcyrcfw7eT+mszf2RIKdpCvpy5uy
Enxcx20KUKMdrzLdbwK3xeUzM+ISHEfe51+HbNEyM+4yAUsb4p5ZUTS9UpCtgikSlRUNkAMmG8Bw
rMww5VlT2PZ5uC/e9ZSmpzJHVhT1EBBtDhOK2860DLqgIPiCgMhrI/mce7Atae92WxYeqYZSEDoe
gmrlAmMvQviSRjSeN1oILdGOdjX7UpZp6/Vqd79WL7KusRxA1XRm9ZAzXeaINYQbtyFr5lYYcmsA
qc+3T5V9FMF3k2uPDuWbh4hCc1A1eU8srISBh68zt/LRTm064et1hVbwamUMTz50hX8lAlSFaGtt
+GMEMwjVOairOC6nS9jzbO2hMTApaFkvivlT8v7ztvwIlPNXO7pZXSwoyOC7FgRJHz//nhNDuIfe
9nyvxGuHExg0NTnvxWgaX3atZNKoKWMO1D95MKYzidI8x1xOTD3G9AUVzXVrp36TRhgtz9K/Nerg
kiW2QFkCBh+3NServbyDGZXzXa2u6kFnGbkMMfYL4i+DOfILc+9fKqNyXKzvWRns1EHP7UyN8atz
541KppVI9M8xGmvIT4oH7OIwmKyIEN4E+8Osu2ApgzkzKJzIZd0N5pRGt7NhipR0TuZ3RQOUJls5
6+43+7ne93ChLU9iMmcEn0BWJhp7osmwnspnwS+xikb6fhKwtWaohlIjJu87s7uSTuCoNbKzKH3o
jR+n/e8/pS1eyjk0hmaivjPsDJpyxutHqsCzZ2Hr/EhzIbVV96k1Hu1gnCDPAzKfoUvYwZbGN05F
LpKFFPyn2hEMcGpKLS7CNQSWF/CAMaiQFbmpNdTZtF6d9ixcjxBW0g2upK7A4tS/3DnogUPpDjyX
XI5L/qhKg9y/eGYvvgqbQ0ewBhFsjw7ufH3YwdOGCSw9wkNP+wq+ueOFMIWH+rMn/iQgF0PgfgfE
CazTO9Sr47z/xunK0WMZP9eVViPYcUOj0x1JXxI6A9nHgiT+++v9ZhnQm/6UzVGNWBDX7Yt6t9xD
vaIawEHDtql8jyztFiODdWGGtHEEpPSrxJUB970s2IP7Kp3rum0I66S7Qw1PFVUxtXxMG68VlC5o
gH06kLYg+N+coiBH1tXZieQ5wDL5eIcx4DLuuVQmS2HC4A0UNqEcjIV99oMn0F3bFcoJ4sPscym6
DNpKcjRkfRt+OBc8GJfATkQpttmrfAMYVW/M5B4EDFjunKTVOjqYqwC+w9VF29g17vxonj7RIqM9
fD17Xbnz69nI0cJTmaHFPGAIiD1NWNP+Ek4yxZCbAX/UFul8pU+3G5IUitB3joZ5/v4ErbkEcr8i
E7/oWOfFXcrAEHv+OxteEPH8ngH9Hk0FlcNzcXjhYuk4/pop1OXffqXoN6ywRRuXKTW0coR5lHMF
ltnfy3wTC5PP0iJT75XN9xH/dMZcL9vcM4fzi7gLvlCRu1+RXnPNLnd6EAD1nMlb63EA+EY2x6Zu
4Oh4FwyttkgVlMtU/S937/D14u8OwGvG4RddZ77HvrRvlSvWls0JV8dOZcO2dloaRy69XpBsD8bK
1YjBz2FLKr8jhOOZlB5mGn+jX4tTTIz2DsbRP1LbiQyQxCBFqId/3n7X2aQHdpxiArzM5R07AkQL
5XTFehP1mv0sXPSP9zlvzrV/A4ANrdOCXH0iy7QDFezirwHWG2+KqBqs015lbPVDI5IwB7j1xuWg
PHmFI8NNpGcTs9JS8OMEU8uEb9M/+L0XuOPAuQf+Km5VkHtIR77aA/RWrAM0F01G7Fw/PsnL/J74
D/Gj2OiqYshe6x+Irf9AHj2fj0T35Hcy3o7TUX2s96M4C1b5sMieV9rH5l4cf+Tvyuk5TlaYirCM
Ul7MlBMOVTtmTFgmDmzaI4CrkVNa52oq/z4K65qf42Ni22ppwxl7W3FbnpJeRlyNRJG5dSZ8TM7S
9PFDwAcHrnMMccRRnqpNTNIokTd+9E7jOAib7/kRahpe89dCFs1s98msJg7xzeNZgl/zopNQEhVL
Q7fj6zWSt6+Ft2bQJMiJ7H9OSfB/TPaRBAmIV78GtRmwvu1u1kvn3EXxFn/W59qRf38TdQCQcgtE
xzVsEcQQTLMGB1AkDyNmcolwmJpf+ePuExp1y+GqGnTc7UiOz/FeSIwwC52d5faMrGOJCmhlWuIq
qp+YlQmCQ8cI2I5AncOOEM5e2YzbJndJbeAVUIqVEYYT+ji6MsMJnJ/jTV4LPUBa8Q74KK7nlJz8
aQf7Il7RDv+VvLlhgtm3N+VvA1/vHPinEjEhRWNoCnrqMsxZszuKeWxT8vyWCBRDKNacEmNsdBJa
kg3BqCSzigIJ/SHSslzbnNwi3JS+rcoQfiZ3IEf8B4zIycXsFox6kj4KThwZvESya0KZ4LiyWUc4
SGYRINRzEH3n2zCCzyd5pCto+6NdM8ufwidD9PrpbTIaATZwUN8OKCNIs7IPUGIO4Eob2prxXwzz
uIt//O4p6qY2jppgp0H5XczFWQzw7AxoLnsiRCgYhwxrNii4+anlCfxHxKuZhNPLd5hh85zYBDeM
ax5Z+BZsWoG3WY4+Q2LjwakLEFkWzpgcsaKhil29HRBnjNdaCMeFhwymVNGxw4hu8g90ZffmbvHa
tQm6wKTVoVfNpJHDn2z3GpXUj7dDjU4X8E6WLZhXF5iL3QF5GLWYaTgC54XoNwMXn/MXXTzcqueD
mGVatcPPzVuZwOR8osA9Yr3fjfl2sCpDK0hqVtVM8inLSJJE2gtY9GDJZESEhy/cAIZBWM4Ho4+A
GtpBUQAnkO/gFDiCSSGPt5bNFnF4HeurJZCQge3ND0OqAW1h6WpCULMjeX9zslWRF2dhZ+Ydm7+3
kqOD22HPE8/KiYdYPZGs3xWp1/3myLGMVWz7z5MbKnFYvduq3KViOyPYAfIzj619Zh4wYYhrFhYw
FvSz9jL9MagRpEA148biZHXGvtHq97AIVwCfdFScd8ne/TkqbGrdhJr3Fry8qj5SXkUpeX0QFw3X
wS+19pqwKJmbPV4c4kOtp64W4Bi53c4NZpmgHg6RGYLNiamDZJ25iplWwZRXNjxp8viqcZ8lYFGi
8Z4ke+jh/XKk7KWX+SCwwAy2O46QkjT7O04zdSP3+BGka6n3c0tON6uiox7JnCn5UZ+7T/EBjY+h
vlDcVgQaY4b7qh8gr8pFiYEh1YpVKa8z5ixcrdqrEnuaOU8DRtT8b3++oFM+NqllLmNslXqMtHSF
l6Cr/J2MWsUfVk2JKnxCuI6fAEnIyKalBE6vbQePsY/lZN9YyZac4+DPxizlrH/LGfqTvppaAmm0
rf90HOQf3ynyzJ2SsrHc07JIrXR6xpqhUUx5lZlbr1DiuoNx86M3OaB8ec4pBPvvONSp02YeGxOB
D29SCL+eiKnVTcV3oJ9dqpBODGkXJS9uAbBfErctH5UTOroHlFBISXPZtKj2iB1EFdvfB5LUwrdS
1o6oLjYUmsp456EjTLF8nFNyEJZ8chbLVXP/8xoKGCoiPgE0HW5zxSeUHuVDNZHN8gnHL1SUj7bC
f4ru1Ftvnb4UXK2yfU+sW5ikoq9EkMKNI0bD0GrEAnf9qE7O9E07PQtb6jTduOyUO9Tm1uBBkVM8
nhB6Jwr13bl61efN0HkxD4xavh8hnyY/UwxFzZV4kTd6YXinZF01pV4zlmEbIQqqlYzmZFkZ4Tz5
ZHkyuaUBImq0umeWqvcKSEP0vg1HVL6fGVXM82nTGXz9h6oHbpApNR6WytsynUJKXNyGxO0yhfsR
jYoI17U0URC8tlZq0k8tH6x6+PNkKH4N/50YqAIiiBCYuNNx2aXuY+cm/wV3oGwocVE9HUlK4tDe
FscGsXFD7wT4vMtxpV1ZK56OfIvC817YgoMKYQ9nErqLER5ZfS08ggGrtq7Ar4aQWfbzAyNYX6G0
sPQZdHFgpH50rPx28q6TxtNdO/vkLAzTdTWfG0wIDBRz9TAAwIlRRGQGNqq3GktFtlnbsCSoMRs5
3m5Vn8xu6ojODi+tJAVZtfI3n4HsAWMw4T6O1vjJHysTJ5Do9ZovyjAcYryCeY5415vYhXAzVp4s
87wtJp64O7dyV3On0YfZKWx6axyFdCwxHfpRspzv/C5O8lA1AEFzws0fQNXSzun6WQniYw76Q9LZ
Lvrrl1TxgytGJDTEvb4G4ik/dl+7mwz1nNIcBbu5F+/kqSroXL8Bl23/rOmvn4qvEzNMPJDcoL1W
LYXxiPn6IUithKVQb7CWH4VY3WZC3yPIdSw3cO8UfWMXlUbxi28kNqu4cwMpa1lFoOS0N/7aaWfv
obHDvgMm+2sYNHV1NZEp65TEHbQNNcP+KIaKLNAXAXGvfi97Pd8dMPQx8u2XHA2olS4R+YUHP8Ob
v/wWVii2A+VjVQSjMRhWFFiYuCGuLSUqPWfgJoIyzRU5DSpU1NPfSr5nkIselDc9Cq+ejpd5JSJH
y6rXnVJ6P8uDCzHavd95wNK4upCP2RILre1FOCCDBGQtOBwXT9qjjZf3jo3MJgbrEPPwRqz+33OT
VHLZccQd7lHw5XJn79ot+Ur75tapSpUf0s2Uh6TM0Us+yLj0jZuja8W9s5vta61xu2bXXqQz6Xq6
FtEsZ2gtM1ZdPesNrRDT5wLk6MOQ3+5Gn/hyvuldLkDlBapnwyO83OI87RGR73TXt3ZF2fqBecH4
yDzfVFuc9S2Lzw8XcNEqqnM2G86+v7vAabPykkeqkZS8yeKBZafu7L4RweY3YTxsqL/ywJ3+o4aw
Mya46xB/bIU2yW/a0B3sc6B5bak9O2wf0ElvCTbVDguC3rKzn+kI3YJPz2FXdKvXoVWr4jV24bwE
rGOVlraYl+2S0IQ0TRLwQ8WvwT2eFEAQGcwCX0uT0OmEqjC1Gv9LzkkjHqoV79Uvlkkfr1pzo5La
jMbQkyPhgWG9xnKbRUovNRrnDMVKEhklAhhl+U7gK9E7UdR9csdlXCLCIuRGr2o7Ot9Zn00XzU9n
9XEPWg1CiOxkvkgSATTB0AwLeOu3z0429nRChwyk68RPIz0ghA94LCQi5Rimrv/HXY2MPQxQ5rKu
47MqKHMapA7TklNKOWLjdCHH5VNkK7qNM5tnD0Pigjmz+rThpfmN9WlbZp9g3SHBnYzFmoAChbBK
J1ArR46f3ihmkTYHSk8zOHof6fpoMGVU9N1skrZWTuVkSjWp3D4IktnITF7ubN16pWPFO3MyqvoQ
idz5knMfaZAlFIdsYHhICI6nATpXIGYkmT4j3UzTjlsIWGGb9LEgWOL2vSgk4b8nrD+l64PaKGQl
kVy8kmajP0ITcbPAW+VgAGj066l7sIPhSckqM21Ja/GgxnxSf5UZ4CMHF9KxT87ylS5cvN49M7AJ
u5f10EAbWFbkHzxy+NE8nxHjezEf/9MW4GbeXHTabcOFdTG+SlW0kJ3RguC7UEd2FOOo6prlhzdO
+NSqkvhc0DYRZ44OskELwxLfYdGWk4a3JVCxlAw8ToFcqgf7hZ6/sUZtrX0/tYSbyAc8xnNcKWbE
AvcpITWZYkqC/MVi/AzVn3hOvdQeRJA+Tcc5bu2GvroPWvX0NmCiuHLq2NDj3gzUW+HAgCGHgigq
plzIdEtdQiqouypsPzosVxuZ8z7G5BIzlA6ePl3ZflZbvMnNI/lrkV/eNsVj/ex8qF7Ldow03/wO
4zKW+2SyUJD3qWQuuFcBL6/afpIzttrzsItQWORN/SDbDZJDKbdyx+inDdNpEwObFXU281QixxGk
+dKryf/KOUxiE/WUcTfso5QJDrbmwaN8W2adbAxTdzlfy+eO0eTvOPDCqEWJmRDnENN6Rtzn1cxp
u3n7xoIeNlHKnMzh++q85sFlrYiFvA0kdAX97kAcrUM1T80Lqkf2iVTvhsOpBGQEMeaVmXonlv+F
dmmdaa/RL3DSEkiJ8ZrE54Ea2kRlIUeIwQQGfGh43fBz+uroIWo9BtTokJylRo1bBHm5ZrsBldXK
mapKLxARUxEcdIEZtg1FVII9bRwE7ikQmlee0ZISJEw52nPS+JvOFmkOm1nn5KBXiOgM+O2JV45c
WQ+PPCS6ww5wXuKrOZskciwgiMv+anN3MFHoRb1KMzMgJpQ0vqKjENe5zuPRrkRC4rohijHSP6ZG
X/D7Twq3ns/98wYWnjooYz2/DD1/ZxFGwXTC0zyzx/G6any+3e56L1W2kuHmOAsbJSddqI7i83WY
BrxgPacy1Ip6sIj1mgH0s1nRgyvLAsDxtzdIztYKvqPeze2657UCE9eytmX68/HAKr7NkNx/9Dtf
y86zhFg3r0xGTpCkkll/74eRtTO6qnblWWsAUWMj7dD+SZMZeNjX3VZSNsLjYu+iZ1v4kN0aZWrr
sbnlNYSRJ/2sLujQE+QtMoWxC0uFEZbEZraQa1Yjcreb3ssKhmPIw0nm0SDhsXpH3nZHFFMouXhG
W7PkzBUR4Xy/NVujL+yd87McccAY2IiVpBLaKTVGvfItGjEHcSyJQ4cJX8i11t6UdePxsHFYZLFi
jaZUcYZ/xxJunRSMjkdjy1efxCiWO1YF8HPRMGCKAZ8/eKDD4JYSHyVc/pQXFBKHY0/rakFcAvhq
cj1bsqAESQ4GyUm/lgADi+cW+KamXe93ND6HjOMjq9rn9YB6ZDZMWmXLco+4y+y3xEZjo/E60M94
NbGS82jzcjqxXPFTedpn1qI7susqz9e8D5aRLpRzP30H9lV9Fb0sqX9Rro3iYbLegUixS+ay6Xji
Qo8WultxdjliMMPmlOFeReOvDfX9BTGEl6wVaSI3tV/mJ/eNcof2RCO11reaAN/bgr9fasn18bqh
YMJ+fdroEh7uo+fYn0moAE2DPpeaojIpQabwhTlfljgAjds8ncGvH9pNJkMb/IvOPW74rhgmRN7S
PWNsc6z5sqs3nPgblXT/Rt+haQTmdwP8WWXwLSuJhs5Jkh7D1Rl/VeQfktgWOjXyvLUFI2odwtkM
2PE0o+soZ7qSayC4lRBAI4KWL/2N93XgW4cu6HEdcyRhCwxItmndnV/aSSb15VoMCvpmh43o74L7
8rInOkPJ0VD9YCFG8pitujsgXiLHfay1x3ppxBdAuaoNJr/PsO6JG3spK8DWgkHV4B3BQdYfpD/6
oVDRujRxbzMAzkXNDdsTjmvTl01J2i9YWgU0/QQKA+cmR5Rcrfxzv+jI74vRYRjcXB5FFmKUpAG4
EkNsM0wnS4w2uYn9F6vFvgf7ygmwEXjgzkFRO4rSflrwaShQwdBoG4CgwgfdnhhmTA2Ibzc2eSHA
bM/Xd2q8x5mMdLbX52NuQEMZ659gZbXlutuWDrHwHOLmpfDVJGnoywZGunnMK5wgiPLf5yHNWneJ
6pjstyGgJ0sEZ6vuAc9Dt051nNMEvCRAwZK8OGnmSjQcoC0dZv0U4Fp+tjuLV2yuWBlAtwu9atpe
PfqrZHKP4kH4V6Ctly0xNu3B+r3b39FpUksoQ6QzIiSmqtIHb6mXz/dVSSB6eY89egyPNaogytpD
867p4eqL9iDpSzVzfOptxvSCrBwQ2DhQGdVDINcSTMbnfaiWVF1L2i4cS5nBJdSoBzAfYBcNdNJ2
EVz74nPgJ2Hfhw27Ig6/93GrARTnmbM1bPXGGxIfoTV44lUKm2hsMpZKVgBqLl7J3N1hPxHYFdP5
TKcfUtcCV9XESJOdpnKAqnkc6OYDP/4rCd1xV1TwSbS2jqQlzTUp3WImytPI1u1WT37bHSwPX3Ss
SZaXsQhBFa6O1IxdzMu8xKOeo+1CZC04oQXXiEhdHFIlG/XlMtAwmy4O9lpB0qOpdS9GzXA40mQT
3mKbZCbQn96/Ufav1w8Oqq6Bh2gFDcCRooGBkV8umU8AUlE787J8PKHIjglRdWeTv2FZvAzEodat
zNrRWI6WcxjsBNcjY+7/hqGF7NVRx5dS5u0bYTPhjOinWdAgIExTwvVGYwnVSU1XlZdpzqCYFOMG
YcIklEPz6ULUampOL3vzxZIJWbGACyfHn43zZN4TFQt+b22/jcC4dtBkTV9WoRq/ZPRg+zMMzyqA
ozWRLtYIZZslumhWfV9tfOmrcibEblnMl8NOvME6y8N3wJiFj1Dp6K8HpyzC0qmL/WfVreX0PY54
B9RaDNitFNC+qvQUi7MT1ESwFm/UrlZRVp4mBUBLR6fh+cuM8xDqBjeQmZf3+HuBByE19JLx3Vb/
kRReNLVw67IlqVg5eOYKPORTidSU+ah4t6KX8/dbN4wTkJy/TUDVeaVabIP3q5sIS+kSU+PS/QiI
Uj+w74yRG/Z5fFKUih4RjjP3ISWLDahTTJLjIfTQHEIH5D4UfON4KJmsgEXXxacoqIm1cTl2wFR6
36emPvXQEZfzraCD6j88mSjXTkJRKfBbq7kXJpqRPKG6Xlrp9f8sJ+axQ7QHw9jEGaZ0IuzOBc5x
Gy01+ZoKMcf5rXTuCyXzyNfeI17R2mknnKjxPAoa19lKy9wARSsJodiqexQPRF9gqAvnVsscStPN
cD1//l0wgZPwJDSrA3hKmViNUaehyXlYejCBN56DIjQUEWuU0Jr8WNIH84Gnx1kIruL4LunZJQtF
k7gGSW3BQ6SoF9hNbraonViDETznqtbFDB6/I89udM+mqnWFJyIawE5TMA7bD1h4UzGf0El1UQa0
qGddQ09F/Q9BiKXk4rWfOYbGuf7zhaZSYPp5Zpx2MlH9/HmVLxInsOPV/1iTDCg1XPtgFjpRiz2F
jTszDzbOxx7FPqxFoYvRsy3UlZZ+3Ee6by3VtrsJCdbp9jsmKw9wfwz7H6GU50KJ92/Cgp8jQdk0
1Km5xFhPiMatmiGRUgHqgZoLiraV5KtCnSOMqtyaPTWUnoNdxATELqUual/ZoGaUBnEvn06eCEWK
pw9qAlfCeX2A7YXHgMpLN3J4SKSjjaSl0Hi6HT6gGLbKR/m2Zm5fMt3cNhlyI36nHoBtHubY5ZI7
ETlUVth7QeD/wqzQLCndfiLBrS2G3HS6Tdvsb3/h1Sb6UyttmEeqgHZxFgZtt4uFOOQ6dWqxwpL4
rzYGxDq54hgmIJBk6tG2zDyqtukGYM/SwlTwGcNNrGUgHNv8Wy+DMOUws2zYvoT8KtTwd07hee61
YhDHFq1CphCl3V6u8/MAMrnm/cYCOhcQGlio96eRMtrL/+9X3uHzWF5xz9m1Ro1OI0X65RLLGPkF
kGgp2o0OUnG8jt/BusPfXi30ROHwJhslZFfXJpIYXDx+AA0NmXP6AL8j3vj2GOECYT8CadAQIDFL
CQ5ewk3kTJoIH8/tSFi7nhDV0M8KzY5OnbjiMM/nMgPZwDwvudRNQEk4G8q9Fc6I3OD1J+YdVLJv
ohuQi5aWthQrhWlpM+/bEY01POvjGxfmgMNVxVf5MtvjA9WCmr0PmrOD52tOpk4Rjkj4NcgXWggy
2ezUeUbRIyXluNxcjWYUwfuWRnTDAtpGzKycqO8rbp53OD2ymiGyelH0pU8OWWOMHsleSKiRebCh
RWhxb4yCTJ4/9DiGn6oFQKRpJXr3YW5UfYojXY+stoU29CFc5HJGjf/fzWYDX8gSpmVITGhrcN2a
sm2YpPMNJFzzJ73UHgSkrrWbcNL4p8WCWxfT9l0nJttP5DiZVVRSGvPwkm20uzBjn59NObuKtR4h
nkGBLAgOmOI9Dp8ZkHIQD/vhHAGyDXifC/Iak/sgsJJ8nB6U3W9EFTMhamJ24plG9UIVpEzjIfXc
BwaIlXbyul9vbTCsbiUFZ2FJ1x18ay62DQ/RssN/+9FgM3zGQffdNwMYugfWRuvoCCJViuSUH45b
bEOe1yAJ4xQJkkSncPyMYWFExnXv+vAFDRoqVA2Zw7JxzPrf5WTwCB0n24CUw6OyKr+jZBlZxDtA
eYtLap01X3Foklr+LOSQ5FnME78rqmE9urS16bVN6u4U0AGdXsu1++kWfCnPfJwvyMBWLYZgKj45
UxmilHaVEltgjsy0mIZ+yf/v8LktXQ+adI0U+ITDaB/yOQBozu274Tj30T29uHmoZFLuECxD3M9h
Ld3vs5Z9S+kB7SdBYKTvmoUZaPXaAbYaOKaenvAFtCZK1nVbGpOwYJmhd5dM1vfUsQRw2GozQvZc
8GG0CwWS1I1xgCsfGV3OYAqPXs0ujNr5B9hvMUyuvjJt3p/At9cE92we2S/pHE7K8+kQqD9JfLLr
EHsA8EVTNjj/q7uzwUOmV57+iGq9TqJljR/G00NGDOrGUuOO9ZV8ecpE63vWxtYzV9qfEgB7a8ce
Gz19R2xtAQaIPMVOAxJUdDlK6MczbEvR+BcZwZmxBRMPfCIqv3IesLrhK8aLs2CR+SwMNzZD9tTl
43LhtGrxgZAiFDQzifItzDw9FcBJfRco6TaRWh58IKfTxPkwJTeJyRHggiHII8zpVMMfr28bFbug
qeq7aO+vTzuUb+xzPOna8vLyg6XPStDqxhpUTUh3uwokOplQW9W5n/K+5bQhyCr0xPQM+1FHjp3c
4aHVDIESedifspW/gjSv26X72jdK9ZDcnU2IA+9/nB0g39mQPbBcs7GOx1y50EzNdyN35eCB0Q7A
HrSGKDsg4X9nRCr43mV7K8LWKKeQGLebILcasaTlI0DmSPik9NZeJtfzzzuGJ4JrN66zhsWOjk36
2l43mkPVZsvoCps2UIfN/bABAnQsF8HjlrqalPph+GQH6+5SC2PANskNmONHP8YkAC4q5EOhrzoj
Eq9orHZ8939drUMBxMX35eeBN7MmZKgb4yTVJhvwQKq/Kmal1Y3PaTXM0jSJwKbeuEY3BPynkuKN
LFNzD2Uex72X+UP231S037XrCehPzwl8E13VFoKYBxIZJ60scrEnxsww/+aFjcREI4/076uIAM9G
wa9c6Ae30pulUthNREg197YcH6QmY/v9zas5rXU3Tmc2g1lZUx6Aj20JfElW+8S+dWS0SAvVg7FX
1NdTPBd8hP6wGLrM1GO/wwNjW4al8Q70y3Hv+5+dlANA2zTU4f/MCOkOFkuPJPM4deANmnT0RgGG
Wh/Pox/2gbhXEVedosGpVBVC7T2JseCgbkRpWOV7oCILAB0hdM3IKSGp+OFNWr2jJ2ozzjMUsOTh
GPohRqxW9oD1knO0H1g8PkXZ48/Vqr3IwUZBSj36L1UV/7Nmy0BeR/M7pifvC9PXjQnbACEEE232
SocuTN2i5ACWVPhKysOG0R/vsDE2YVHXdlbptG4CTaxrdtBNhORpXyHcef1MUf+rtB7lSXCP4nUd
h69UHlot9omIhYt7aTIFqgUt/QYoZM1xcli4RrmlzeQdd4uSLWNePuGt1eFvMPLWKZmMm9svmfwm
62V8bTCBQe8AzygrVhYdkxrPLC5S9tDqoY2jAmBT0UZfeZOgqnY/NpgQJUZAh3MlV8D3SxD0lyZF
FRsp/NZxlytBjJaKllKU/VQIuNh7FjxHDR6AjE/10WoBYsThn+XUoouvqQOAnxsDAfNYl5K3lS74
HKeDtZrUTynmiUiuIAoU//EKIMkZqMdzJMp4oGa9kHvEBRbyP7zbF2ruc5a5Y5I22o8TG9VHxggM
/1oxyfNzYtUtc0D99lE+9JTlLBS96fqyyY3Vm4UG7E4+7agTezlC4TgjUPJzS0bmDKOBS2HgZKYT
mahuhvbWEVo9R1H2QjMqdfiLiGv1V7u0+YW6Gn+e1ox/5MLkyDlV5O+8QclLTUO+/EuDhjDpm/Ex
Dg2pL6xh3rgxs7WZI2JCs8Kjuja9dIdlhybGijbtYX7VR2c2KgZesu96E63PiHug5myWBuXlrYUD
mmKGCzGBrFvl8S3HkeW6UJ52mn5A3TsQHXPq+o+m8p+6exJCRN3QKFdM7rg8r1Yj1WIwwrqLlQiV
EPIk37rB3W6La8sQO7GPrLWpq3mM2vTRg9bRyJOo2xdCWmaJdWtra+JMEFPyiMl3YLDBsZl+Mwh+
Yj5yHUrvffI7Yxg5gUChosRBd5C67iV69V3UvJPZNg5zCJastR9IvPhB3+QyF5M9SwN2o3vSDnUr
p/nr93WGMhupxkQJhaRrsOHk0G+bqGVJ0+ZgPz7s2GIXDF8S3b5TUEeS+LT9p+6h9BxGPM9Ns+qf
FpFEV+WND2OW73ehwHsPC/83tabC442M3iinKwOIWIvSlYENrK2gxHH/nbvUqS/a4mZDcPgdDzGp
lGJ543sef2F2fhnCvHITNnmZ2uQmtCSCjrUf2YgATQzL/b3b4yXqOhoxsD9qDmGEfof87CJ+oLHn
isubWrbR7H3fjYDCwAYX3hVo4qEQrDYnwogsdAoRXmVPrCD+/DwFwwDwPqxUPwqc6parcKba3Ul+
XAqzFnuogz3sr61ati3RgQ4KHdoUD6mah4hpq5e25CkNkM9I+VpbDRvFpl+Q5W67IkabRYpf7fKS
g7Ppf/X6J04qh7lBrIpSow38wVfd6CSg0pk9lBtoSg97b5aiA8RLk+TmMX9kiOBFpuPi4Ogfu++Y
lnqriejGjM/6gSgaAHet4cnj6bu1dEmGzBssFrAHvNlRZ6Xtw+JV+cp6GdB6G9fAznYYc5wfWiQn
hMWF2X2hqvesO03rS3+rYR0mk8+Y6NB1P7ml7TCxLNf42CTlGvnAdNNS7f17k2uMzU+apTaBwhAG
C4irGH6JgxGPqNUNR6CPP92oWgljQoXUvVsRv6WUn46QTMCdHwop8SM4JVfi5bDrvxgo/L6WKshu
QSO2QccLCsn2KAG5KJEIFv1BcZCN9+2CZTceIMG6JIjcTEmkzRyebkdiIqGkbzlukU4tZFCISBw0
B7UxmE7spQjT/+zYlQ3dXQOtNW9dfM27N4TwEwU77/fyZhlRUqj3nPw7bQ8YmQdRhqp4Vbcusl/P
k4ZGSweBLEzjt3XWvtBODomFnhDh2WE6/Nmg2LLuW6gGCoT5ZAf7Wd7liTznS2ZnrR6RiBXmRk4q
Iw3YLmtCJ/diCq2h5bWXuh/GgsTOJ4xXHFBGIXzJ+FI9Z/KowfIG8KXt3ggwMQUDPlJlN8MaZ+zX
TE085H0qXI9iYI3Xi3cpVVnJ9YaYtbkyPPRkjm5c293E1gJXCa/LABTymTn1tEicMo562VQAzktH
iJRbB68NoWw+NSGNgCmP++1/gkpNUvXHOF2DRr7A6asaD90f7B6LLLJphWkWlOIGcCVanMi5vQ3i
EBlCTblBsC33jOJ2Uv6imyHlhv9p461A76/Rndz7maiYIjz6AD+qdFxqHGnkZ63399FJ+ebTFYhb
NVaojkcRdFkhwwdct6TK1LDygPH1R6QcXCnA0P0TPjqcgVuklj1a9XeFaWEDFGqPtW0RrT7ljOUO
9oUIQsUvzgvK3/PyyF9dieCmJ2o5eb8vOV60s0XkLvSvI5MeJi5HoOAeU25lNT8kMQfrC3T4xYdB
BmN2wE91IYJvVslzyu4PFfRMcAsz29KL39vYVP1Ey1BZOeeC7HJMadC/RMOnGNY1S8/3ZBIgFD5k
j72CBX4EvcM/5azC8UJlIBXwaZ43bX2fAW0PLB2+FglIpk2znBYxsJbLqSwWpSrnldalFSeAuXeO
SsOGNuvKLlGfpMZVhYQXKvHEas1styeIw7bb+mo7uqasg0LY0gLlmzL1lrzDPXn6nhwEr0+48AhQ
qJg91SgrqZ9ZDL+kE2IKiM/C6q6dy/H4SyWBdMTMfVUN3hhzYoGu4dj7iQb0qq+U6lPCZ9kpaRR+
vJ6+y4DjTm6RSYYtVNBo1Mp3Gj4qQuQITE2FUg2HzJYrx4/CM8jwOpBw4Zpda2x9ZJfYQriBV7/J
C11uV4Dxpox183H9SgstDqwu6fhc2RY/h7nb7vQLO3p4l2TmGbiGYvEAzrCtJ4BV02eNB+5BsvfS
U1/MR3G94jY8ukiHHY/BmUCMoa3FJa129nwvU50zDHFmqOcFipPTivwGdaqQuqTgIGVlNnGLz2tn
WnC35z66OJIGtcV92WYovhuOBUzWUb1oapU4VCAs8pDeOUyjEcV6m6lcRqzSxsQaO1uwa1b4U2Ab
FAHCEv/crLk8iOifhZMB+BjCl88KAU/GXY5WDmPTPgUMTeJnppFg6Q3Toizk7pRvK1OT/bIxcF9a
tXwHGMHAweoEEGhXfMKEmXbaeD0Q72eadjXApdl6rvITktEn2/LS6csw5Ew/zAccfwhautlMVYdy
W84EUCyMv/Par+UUir344LPFu7HBA1GR6AlXrk+x9ZmrqsmrtQb5sGTWSG5K9qqEIL5z46D/A7ot
CJ2LSRmj8kbOg9Ey0/xOfFfSy4tB+uBd5iMZZRFjsrw3XkWABvUYy+IrLwQaGxBs/ab+bbWpG4hr
M5ORb6R9Pzedk7F9Or4IJYcP53ssqcY4p4ekYa2toVovWOcpjHuIqHhSVBfrLOS5yVlZCDlClXYj
5z19wL34K7kKdQyJkjwZ1Wg6orCwe96XvWqsF0uSxCWJK2i63JXkYBCGXICHyUg18PxqFQPcP39x
sOdFPim4lvVS7yBr7KaBk0leUA6t3BZEjjan+e2HkC1pln1mimPgI+DfxIAAkD5aeAfkDLHk1JFr
MUYHTNKV75gozIwt0vM1DZx1jes7m8uigr44tKu+FurmxPVhhjDbEpJTu81B9/AGAFmrjJsB8sa9
iP+Kn60ixiL3KwCO6gVoSDUjxGEaQxaDpUVTPzbrSWTcAdvUD5m4i1m0dBQvHiSrYdpxr/GLxnuW
gb1jkAeoYyhuJSGeIqUdhXN/aXIZWtNioU0gCUpRewxL9K/iwBBnQ8L5IOVkK6BQsXmFP7Kf6pll
HXsnczSrn60+QYCW8XAgLnvd3UklUPxpXg41pj0jruDGG+IHn9Hyn4udTQRFbcrnE3T6pZH6m8OS
MDAEzVbNBmPOv/FlIZt0UPIpplIfUPTOBKtyoNkOs74bb/HfSpkdYqNuFAj4BhJWkIqSB9v5yCHC
AiWIHse2hl/CwNk66OmaxBVqBfHLUtfc19fVYiKY0HIDVQMAG5TxQ/D1J4ifOs/jHnVQJe/yQl5w
JTrWyp3Oi/QFl8+FY69ksWZ8cLB7+mFwz9ogmSz+jY1urWxgUhKoIWAMDnx382kwGq/J4tLQ8z9D
ut7aS9k//CJM4g5Fy6rv1OgjFlPpCqeb7b/xWAXwG9HW0CgpaIDxbvqHsX5MyIMRyEBheyFpAwuL
p+lXUD+mfzG4EJ2Bx2mXfRtutaFup2DEF17Jiax1ON/64D0WoX8QX35FioCsjHCS6iRgcmFAxiTf
bqS4IfW9iTGWcUTKnfw7Fd3QPy1wvijG5T9HxzbkZwb8pjdJsmNaZ36uVlV2tr6K+W9A3EvB8dBZ
l4IkGBNDqWvDcC2l74l2q5Vp8DXvwZPYaCoGONUBGN3aqWJBmi8IaWGcl73QVAJzD6VUb/1KBkQz
a4SEust43IP5U3hxwarfj1zw8WmkuR2wqAQQ1RI2T7QTGwe2LxAhBcEYmhyMpvc7vCf8KYYm89bA
P06RV+52aa5ICqHktOxnknncWSV7+igauvZarvdvgzNhxv6QDTe2iK3X3QwvP1O4//iSIiri3R78
KKPV+crMYwrKF2Ct33sJrRTBNkHhma6wwwXtB2bfqs9W8eX1RLLMPWmvVYG0qHMh5m5XgT1xAb+B
q8XTAUCesTG5Q5L1L1wi4GN5VWB0xuETvv8A3k1+wJIbmNp+Yn+xrn+A34mijPdQbyreqaQShnzs
vfD991+X0SJvwZvLu8D0sVl+G8bdXomcS+zH5yBYMii9x0Vo5zNOMLGyWNDXVgwmo/dSWOx/IIy2
K77DTZ0vNX9Ga/XmwOJni5PwM+5IBltn5g0P/2bca44v0ll4hOzQ5wd/Y11fLqFfZKjfyf5R+2/4
8Z5WD6ESTOCJJiKPGSVBy++BW4qr+IwQYLXR6m0ddFIeuuqA/LMh1wFxl/M0z/q/XygUm9LOSwMP
ZVq4cj3db2scf/4EQHCL2rMMVO485D/2HcDKmFB/wCz/ABpWyQjlNn0xnQQQZFQoSWsv2MhaA+A5
xmwsLfeR+sWYTj59PjDKWBVqXyGYLHA4EJJDUa+niv/h5yBPMSxQr0iuBEVNPXZPTE3jAMGtbsZQ
yoA9oc2iWYPMl20vIvq3zhPpXcQfpNTWh7ZsgrwRIa/wHKzo+Ymp7LqwLR5RjZDAi6OabcAn3afg
uUv7ncHOZBoAenQWYif2kMSQPXVAbhGtCz2uTa0zL1QETdxFzW1bgmhUa5o1AYmxDqJAq+mIgF6w
emOXe6c32Ya4hT9WboIPWJ0ZtSmCsaYx8lAYQc0MgFaZZxCZ3WOYPk1MqICY5DfEHOGqOr1Hj1bD
/8Ul8ppXjuO4U8nE4wwCzpvRWSKV5jFo0eM54PgsJRSK2uyaNi5zg82hzEoXx4E1HLmgY59SSQ6u
rFk14F/bPhhlj7ju7sBepamciVV4L3fXAbUj4AJdD+u3TsyHCIkj/PazQRoFcy51/HjVKzc3fJgz
k+ZgpwX7AwvS6Xul/uLUdrFKCPV7kvt3/M3b8Us/yr/Ei56HGJsri5xxlvqHUxqhxZqsTGlS45Ic
Dujvo/x/PYP/JwAPp9CHkaB+7t1XPn5ERtkhuUifnYQW5HjaSx80dZjBSic3Iwh9sYA09XVidA31
6aRCEAVzYwlhdhq9wMtwBXfhCFNJa9ghWAUeKy3sTL6xXDNj4MSYv7BXJTpgLTxfkzm6N+CUASWy
U6ABtoHDlWpvEJHMRIk2HyFNx2MEFgd9KOfvcTFAt9JRbRr6jKHjdB4VozmuengM+O9Om89hlVQN
ELnOCrrA8DATxLVhzSUBtI+FKQfEyxvvcn6IHQTy7VtdrXa5nWVK0EIDmlxgy5R0e+58FGyNt5tQ
To8p2o61PLPgQpe16VRvf8N16gIMt8oa9VUedhqKsZqHWfwIOdga4R7IS15QI6Oi3p4k0d59Bx1P
YZ7fKikIzyTHRqK/hPVN5bzgsCsTU3NjiHcLGWN39bpoVerQaNX8P/mjVQDoHUE65N5PS4204qzX
7471Ur8uq4Fa1NK7WPF2lsczXAvd6SMjKSfGzK9ZqSJ+lvTU7IiBg5Hds8fgUKR/gdFssPfujLg6
HNAgwXHlxQ2bHnrSE3HO3zmOyWZ6OJ+Yi71tGTBdftyKxuqHabRA3723WLixxCLDlL7OFJ18MjBt
sK32BR3ftVqtm4erxOjvHjmPSHDKg7AmDKZPGfw+hCWGjGj81LMjRHjtApCfhsZtPF/vQ+/55fgz
rYdS4AguFD0C9Yzr348dBqR9g+rWhp6N+FYtWcptIfW4rXWHlcwRXwvz4J+xjowi0MW6eCyIOuLh
baLqQV1wRyAauDXuxVeznS/mPhjHy2WUWKe8CDFMFMrTsTFNx17yLy3M6EYsVK6U4EoCMpbFLd2h
QorDYJol4NnO1m88a6C1LoNf3komAHN30QobkGlzfHOnmP3nQFxfC3JUy7N8HYMbCbJDFqWPC0NL
BQ+a+iSCdUdBQ5ZP75lIchjz4Kdf6si+oUbEKA68bG/f7b50XZTY+ulvK32Mv+ORdv99sR0+xbNm
I1Fala0s17aFW0Xitmi9CPA042uf2UtXyHTZI08pGzA1GFIzuGrXyqw/j5hIR6M6CXIiQbDVGnj3
MYmGAODEjsmo7CGs1BFxsI88zuONeqz2z38AT4+3Ij+YrP/bPQEk6qwEPM2oIUw1VDyL5E0ZZEzR
SueUPPQ1qpZQibKPS7aY0ZqztF9E9EzXd8xUPQFSgrA6iqLJk501NWbJ50jlcxU4PuI/b2aUEn6V
1VPiOJmbkPNkUTE1UBsvpjaU9Y2tImozJpaVgoAIGMbDQRSOkO6UUHRy3R8o9LzITLULzQgt++tJ
exblaWoKPbe8GswgePmDpiEVqJ8NwTADOrCpjFFdrP2xdr1tpyR/I2NEkbNcLqR+1W2Yjjm0tuRe
iJbFAto2E8grkhaAr7eSHTv8HU/UjvpmMyEBdiVYj+B+UATgVMwbiCOMN2aDCuCTxZ2QH3AJV8tp
3KHELBLrMK1/w049LL8/GY96bhxvv07HSx2xpW/0uKeVrh7HayTuZu5hmq0bPmOWnVNWOUNc5Bbq
p1PadpCgkDiC9CAPGi2ln5YBOaKIrAWSdeGAL8YwbD88+7pPdIu9cLP+cAY+Qu9ETKqROFpSCgip
oVV0ujQR4HOW6Nv6MJphzA6Sfi3j2gOlSRAtoEjD5yzs/uqxo3LdTbzLLM6ToWzL8COBJ+tH9uAx
XcgqG9VdZL6q5kksX5zatbX1CSb32tO45uU3a8qb9EUd3aUEr5s53eq0zydiRVriUm43hgi0FH8f
QDXKpSRmzWYwqcCYNH/tKSqJbf7WyN5F/vwju6yGtzxneSzoxIVntuOfqpDXCqqLzALizQOB5F+Y
igV73YT+cIBjnSC8jgzi1bhdt0BXLWY0rftKiBn0DN6LBALkkvwIyoaqsOuEZxh8USMTomX2f8OH
qt9e5lj622owE/oYmsF8EmNgAzlQZTlJ1ctZvr9duv9D8vKEo5HXDIXbmHd+Wa3eg8uA1OcihrWE
uPerPWiwzBLJ9QuWrLXRVGl/w4/MkmDxU0QbeSN4Qo1YOjEgPdSnI2MW6ELPGEQ3QgwOK4C+RO4u
DEKjik+u4ok3FD07mVKbXtPgYip4/cGOuxMHKKqcb0fPTaOteOm6SQL49yD8FG39TEBvOdgcPqhc
ySkJv8CFEHiXTjPziUWHm2D2JmpZiJVEgrBtTkeboucMEs02ejK1QwdqTAN6igX6BuimsW4hCsax
YlitrIdiapmLEKnlnIq6wnbvjb3nXOPhdyynblQ969jrd7yk+bnBldfe3jx3poIoBbytwwgb0crL
nSWxokt7frhENyRT0DdD9nKZKjNIOAUHaqIXspM0UNfxBZtrF/LHQZpmlr6HtYwJeuTGavzjsKlq
+h7Bab9us80baibUk2sWm/RpbSs7HVsis+zRIdq8ocIjWLG8+1Q4EaaLg2rB92J78yc2T+SpqUGK
nhBRimJpAbqk0u6Hkh9J9QewPk795H1inH4EHiHBZrKA8CuZuAiZQeIDoxQ1IdTKH3to/dE7GDtP
bp2QY2jJ0sVXpak9rpOeJdH+HOAXP1AD9KcI4y2vtQsWLadWO2Qnor4iJu2USceIN9KoGySjuXlS
SjvqHNVdDhL64oqSJMu3vSkYjqgXpdn8zhSUyWuvjM24Tvx8n74tAVTbPnRXNYz59+n+WxqiHPSY
NjWTIa0mlGFcpkd3u/r4c9e9vIY5oiYKNQ3xnyPqrVisZUjGQhwRtLDMpxr4lJBZ5EkakwO1N494
cpriSv9TTm8HmiUbd3+lkE26QTufVzjxAA2d0Idit8DjGANCZp96Mgiyf9yprs5NwlT+d7xKTUjg
Drq1JTILfzAMUtVTQjSdT0FRh/0clbaCMFUKfGzngXX4w4k4PsdMa6qNtdDLenQuyMPWHrl9SDX6
+cjDcUebINuaNxpvi8QfuEZhmb8ecmyExfaiJdPdBxDATUFqgklVOWd0/wkT/32RoLl6/ALZBtA2
LNxRC42WYpUlrMoXWmcnQ8QVZAMo+kURGYpY0dpWCrLQQ4/Dem3u4KEPAluLgSf7zYR8m9gn5vuH
PL0coxhKSgNUpZcjBUFORJFc/wTdTiLFGhfTuQ4tGVuAlqIPaKjJqUnCEYiXSQhxeWquGAWRqD+e
2dXHjB975P2P8S6/OSaQ+mnARGsiW/txay4I4j+8PFAKL9XWW3AprErGF4dtPluc7IUU+/muy7K3
0iEFRGa6TaOVnB/+0iEc/FzmHP1tLJZ5VyKucL7+ZEKFp+e0WSccgIhL/D0SQzqaDl9PIm+fSi7i
nArY0IsU20iwvUALoHOCfQRoBjAUQnKmClNxzSsOY1q6Zy2kg8+HPFaaw+S1gy1bZBUyxd++jr6q
GM9NO7GZLEXZxdvEcNdM5Zu+ikKutJLj2tYHF9ePyE1qqf8yl+43RJcDAZ47NqluBP433uYS5j2j
IOF/9mNtE3GrqqzBnlDu99pxN2O2aTFlAd7qo+vKpGNzy6V4n8qRTF/NjV4gDGTAQKezHyIYxtEI
w7K5qwy17XRiySCe36LT0Su9twvwsdq6KgyJcpmx/dtT+3DzGGLi6619VILE5dqqMd2DXtJZtgfG
GGLTkSy4Yt9Ad9FVGO1cYYXNnEjJlQxFLEo64HlZEdfsY0TW/eD+73WWl5LA5+mwq4JdSvxmmyrP
Dje6bMEw3D0KKZZReohNXu5ak1nGYUZT5QJPGeHlXC+CPQtHWi6mpwTAqkh2kYMXKdMWtYKuRNkq
7Px5tzR4sCgqB+L4alEEIV2qghEN+0X6zIep9TbnkwWj1vXfBQjnJUo+SR1hF0V4q4vXvuwTYXQq
ic0cz8afKcxcpLFCtEzLgbT+sIeEGfqHQKY/rHrtUgzjoq66CUqq9goZvUR1Hg6h8TLl1Wy7vyZK
VuZXN62JfHW+91dgBgo3G2d1Hg9Xl5XwricBpOlXdqcuqeYG2VoZumoji2E4CnJnzjZQGCCB71XD
VslzA35g8g7IprHDcfLcDe+JZDHmxO3p2GeI/YQ6UHH1v8acTF/ritPvT4lMk1qLgMIVdwAONNXL
p0iX83hMJ18LaCwiPQYupAoql8OvML/qosNMM+a+USD7DSCMjYwC3NfeXLcEj+O2BJb8SE4UcX08
0zS2talun01Nam3Kpi7gIdh6EjzLXC8w54gS2u0fXQ3g+x+n7rAAyQyTY+Z4m7fkr6uAUVFy3pEq
jpj59Emm8igCzcJCp4w7bkTbB4+TKsIhXdBfds5/c+zCvJJZ+9YWdxAayd7bp0j606Kk91eaH7jO
znB9BgCFGtEeCtOFBsOxA8Rd+tFrWuKqLxrxUeqD/fkq+5sI7DZtQ1FFfk1m1/fRngNwRn6T3JoL
OSfW/OLy8+tZqyjLXp2vgXsYfdO3aZJxQmFJU6PtTcqXJht+npvTMI3nH9u5IcT6rbAuUmHVZdJ9
tVLZfOyFEqVbTHCb++b0PFHiA5on2Xjnt0H+TcC92biRh2X0o/avL56DdW8uw1IXVuXLftINthZm
71muiSXifP0BC+UuLVj7ScjtaU5JvVvwAPhf7RPkkFeH5SvVeMbAOZ9hxOovDk+pFBduL+lM0HF1
JMZr71qdC47Yksz4/stPszc4chEoEo5yW/3wVxR+hROwecAMqRVoAMloXWd8EriAvUYnFdljmJ8W
5+nOgiZ6asMONypb4Abs/jQ9HbmFW1IJGl0uxWU9E2zhrrDHUAci1y4OAkBmDpWLXZrpOfFVgiSi
PrXLXNbTeZg0eAjmKP9DTWbpAikc2BS02Q9Szn+UEINMVmyk777m3f9BUr/cEfWdPiIKy757Jnx3
TbeO/0OR4TUSOC5xR649vXMcU89ax2uGy5eaItbfciDB/Do46Gt7V1w33UEfRzE2BSbmikfxEl8E
Yos4mS6eXtaZqO5yGJPAuncb6zPzIwjZJs8dQr1DlQzhbsBt4bMlK/QWnaJ0OvIn8sMWS89HIZEE
jtRwNjtheSzbutZVAzQvbcHGRU/NYT34XbOf6D1eyEUL5Y65jmqnwog2kFMZet/uvcKa+6A8cbhR
avGbZ61XCchYeimdY147ks3Sxr1zhk0BFj3OYos+ubik8SF8pLER5akg52nrW71ML/NOWIiI5S7M
3T5TmS2mMITUROP/y6qZCA7i0Ga4wOpaXrIF6EC2QpI3jRMByIBdgxFqs/WhxSgO5QJaoRtKd22h
1VhvhvJ3MqUU5zMxjh0agIvibnU8oBMXDt6CCTxPqmWdTqxm2jbW3bwE/NEMV3lFyyOyEhpcTIQp
uV/t/oaIa9VVMuz43/mfr5lFx40VZhEfB3RAP7+GL7giwuEwtdegWdRpZsU2QWdxDZ4L9+5xXD6z
xnei3ofNMR2nkcfepWK04L5YzHObaM1i34uku/ejyQ1+2Q+05epgB0pOCGx2K+fbfSRCR5W3eD0i
9pfGkSWCbg+BaH0ibXtCbgl551/RIdgWeaGzAsRgGFaUB8mjwIWeIJli7aNkwKLHx68e0Ilyn48I
RztO7qM9vBg9bEE+X/vObppJsGPTwBILvLoR+QTzr1LG55rPeYNtv43WibqHf+ZQTpj4s+JXJS5+
jOfT1gAqVxZAalfdt4BXPbu05FKG1ZQW/fkhrZox/Z/kbX2BbtyqF3qPNHFp45NGkS5uLNz1oG6n
Ph30Se2nNbNOZkWuIH01i7qGX79Vwu1m9FqeB9UKMEBGWDsK0k7r9LRh0BMbjU6uxz28DPFO2KwI
iKDDZzgZuWymrH7sxRRf9raolwe1PozHoOvqyxN6IZ6ndbs39VDTDPgFwBgm+Ezi2gsedE4vR86U
gDOSJnnIeq3K8bRo8blOjbQknb8kGJqBWuLnYbYa+SCSXjrxVnYJGpnlFDUNKj5Pt423F/zXC/4F
O8ArWh64lER+oaAArz2U9916sER8+yoXndK2baTxjopxxkuWEet6jcSNNLb+QEB+dUvVeWpB8/aW
n3JRpueCbMR4mUv5EzNfPIFT8ciQxewUwYSRQoI2/0g7i//Lmwb07KYJhND0+H+Qr4c9GAAXtjS4
LKAy3xt/Sx5zfSLfjuc+ykIR3PYbIZexX4W+GihuuVt8F9DtYyYGi5sknN//NWDAZnuBEyxSQpDk
OWInXt7nEGF64zTkbJFxgfFeUzxzEJmYe547MtIN7bAAVa147LU08zYto6x/nRuvtq5VqfBO9Cwm
lXF2o1u+TuUTOwxJQAZDa7zSRh9PR06cjSB455YnKcT62AJpFyfKolOjcxUEmovUlYMRavzT+/N2
Zrhe6FJLK2lqaZ7gPHye7JFbhJBYcbJU1TlYB2G/4jzpAtLhCgXuY2pxXIIyXQ5vkgBUs54Fl3EF
yPrBNj+2Z08bkYxDJrSndca6Xwhez/qZUDDZ7rjkQDNol4GlPuMAa2usKQ2+V3d9shjrbKJKXcAV
EAnVDex0+vQRPlSisxfJjXqaA/3zd1d9sjksCDHWZMe+wDu8MaXdPLdzK7wv9XwVuxrsc+Ykj6jY
N+ITMenzCRox3YbL/qToaZxm1/EGbptPn3+aHRRzRzqvOiDwYBbTL1JM3pdKtof28aEVKYNttBsW
7w+zdOE5LE5yuLcw5Kacq102paSUBcTS9nJM97Iz66w6wpqcr8Hfh95oIc6U55/AHt3W9qY/U1x0
LeGz2uw91fpqloX0Xr4My+88Nfk0RuZ7ye5I7yvYiulru+idCOFvHqLyvpwFgGdnmL6ZNlE294oc
SLhhGoOT6m1UcpyYrkhPiLgVt7Tr3FRaswgPRdTV3i5H8OPFUbrlGp2sglTe9kIdasKWwzhyr6ln
/TbIHxnaM3kaP7u7P6Mzd3NvREFAT9vVVufexrHrZQkqPAM+j8ZIU5B3NZ2h6sdgUeAs4PeKAoQJ
d9fhjWslShB/0szMnPElWGS2LwMEP6W63GvUdJg8AqFkRR+8sAnMmNeM/50cY9LBlKnpZFKbfYnY
LiY3v2OeJPvC70zXpTfBS382TrcZjaro3GLXCkTULxHo1dUYKrAOWA8gnfWl625lbJr9yiNVtiBn
q4tA3L5V5xntRBSybf7LJtPsRrAZKciGU7utCBOGTAuMNWV1xLQ/6kI1oLq7tWVi+d/OgL3pCH+N
YJOF5AQmqnHdrVjTCRLkiOEQ9cS/xiM829mnd8NnKOef7EPaCb7nTVEwPC9t9SprViXdF0IGoAqn
Exj0+bVx7VYsz+c7wbPQS+O3cEmIpZiKw+MfIS4EwhSLUlZG/vXlXmq/2UjaoI+cuAvZ+CwNSsK0
ylOgMNWq3F3Fe4RfQ3MWa90L30WzpQA8pdlha1qTKqiWeAK/s9Zr8334OLSTY/YQ9S+Ves2SBpim
dTxVWZBcsLobtNRi8riYOc3DjDDadHm0GWJrBmASX5WQ9/ISXEKIcd1W/ftmm9uaBfr3izSrmgKz
32cZzAJPxnUTfIdfMHrbZIkEfXxHWC070R1qc8D+lbkEk2A7CbLeVPgEfCKXbKlSgt3wFQdw05B1
k7n7nD4OSm3mHEvQpPWNAtMNsH37tuqk7Wx4Xez/ENyy2Ye0h5s7MZqYsE+SJzuujw+dlsM3ARKg
mGLEQK5J0PLh/CNPN5rq/vkLtcx49IdcxlQB3M0xBY82B4h7VuU9tCu4iesJ3q5bYEhwVROydhwH
VViVCg1N0hJqvsbKFSKjAAHacUKPHZrhK/U2cMJwkf8lYphtTRxyCb5XFd9lSuH0njpEDYJOuCmr
s3FoFofLLNsqfc8/ar7EZbZTJnRLPgQoWfXZWHAtkgzwsBcB1dPMFPXOk/HeJmh0/6nRyfjCYcFd
9pXuf8s55EmNFAmD3L7+EIPWp/eZTzl1pdvMC5JhAmBf07+vYbuGFdvFZljVsLHP48stmGrD1z1S
3Qy76yt8XW3XYrSydIYOiWIcJkkt3LH7p+cRE9hFVoFzHl/u2SB4OzDHrwiSFsKqHDPZO4cbVJdE
nAA3l5Ps/U4edEEaHtK6PUW+ORQnoy2XNUzMFuyb5507j6oVSb+4NnEpmODsjmCn+OjWKDqMp/oi
ZLGsQswxn83ngi3nHvMIanClLShvp3DVALNBjTLZ5y9sMG6zuML8MN+OyfTzaAwkN1GkJON9YMem
yf1KOVPPLD5zTQWTqCmJdfsz6Da3a+XE/viwHc9SjvGJ50yAiQlwJB9bBn55jN8uq0uUMdK5On2q
8cCAqVnO5Ax927uk0fbPhOATpCYurlDEqfnhHUrtDFsWtVR/GTLXaOhxoxXGEsmsEdaM9vD7ZKKf
y2xDlqokLlK6PJlB70HHoxt+fmsVz3F2bmF+WGmzYYIWIFAIcRY1F+plIrOcxm3bJS5mY9q4Yvus
8jDFlaxBhwRWhGxd253pyIdaL7n3m6Mvxk9MZxJOQbp9LMS+agbIAJMf5ggD7aK1C1pV0Rkch+fF
NmgDQURpNh1F4hAzPgOj1RdFHSMVl9fJ1qj61elvFtI7E3eCzpwgR54CE7hcQ3ihLVikBxSx1SSS
ulovBdNrM51bI0LJ5XXu8/DdFwzKkQSVkxvM+cHWWF8jmMzFTXQrffJ8HaHii2G/TPv24qziqRyp
YLzwVqo4AseE7v6ncRdQSpb1Uf7CKUPPXnAir+qRW0Q/dOKyoW1rxTDrOeha5vwDa4DYcKov9NHx
li/iWj3S41brgAl1dsc3eULGiK4C7MRaXUC7vlb6+kp3efRFth6zv9nNXlyUf67vezuzCwlYaa1S
hs4TW6muSRBgVllRVLxIsuzB72krKvNUqjujTvhJ3RBGlykeGJUSAimq3JMJoS2HjF+ZqcWg/xHR
MhXFFUG5pOIPqVo7aFlfGwOun+2V0wZplfAwhd1EkGCooZGlhwousANtrF4YKWWsY7p7jN+Dw34r
+UTvm1eK6g9qrtdMhXndfb013aok1rFaIfe54EZwnV4t4AY9pygK3tc0xbswin7nOeYWIQCvEqgO
J8aO3rrS48dslvGEY70ARqbB2ANjuZYulG5RqsrOPXmUJvsCQbPWQeXFA8yZef0NwrUpPhgepgQL
vgvsD4H9ajWceDzQ1TYs1c8IlWaU8cN0qrm4bZFZTKdOsHm10fNII+N6uljBiHM0jbipZcwZkCzs
5bpZIiRFsYie0uKQXJrbsw6hOJzupZKZd97lFezcudumQKaIweJdcChpD+xVKTTYugiEzW8Zkfs7
0DOCC0fHhzZB3+KveVwftxgJgq2Z+VgdfOfpa2fbRK9moRA+kGN8dIJzlCE/HJfPCLHtBuYDFL7n
ZSmaYOhRIhy2QLAMozN5tvgw8U6uUL3fUEgrzKumynwM5BK9jX8AwAeeEIJ+ubOThwyPDF04yqCj
K/6hPK4rBjKlFmOxql4iKLIkqrd76qWMqaXlWyaHlkXgTr5pREUNGGRiwTLXovfopbubf7f6qIMY
sc+F5Ph8hJrkxjuDykNlqBq3k3mkJJ5z5vOt0pdvP/LKLpZIOwh9ERWukSca+iyrD7LxLNUqpUY9
GYmVL0O+ctI7NNoDpp8EEnPkcopqQns4vTaA8hSbxul7X6hpnR0a86Tnw5ySmVea6n/4f0+7kIpi
5CUgJHu8XnFamGi64zmWeBIJYauaxd4r72koteDh3nzF+VbQ3vcemf3Ek0O0l5JSbyPg0k4JFBXs
6q1H9+YiuFX3WdfE7HdB/C69OMZa7f43YUnNqupZmhvO4oBI4pGN5ng/Dx0fAIs4JcZkBcbfKy0D
EOyGuCiWcoZFZiWPzFItVNq4RSGw5WPGicOMN8bQ+GcpcvI8Njwb/Kr7p35P3iWbgQN+qFoSPgNP
Uf6kLjDTOdkgtvWk1beFobBcnF9NA76QouZwObRwKX9UO3XOpGov4+lWTHTx6zvZVa/LfR1MqgwY
XIruJ7AJIagpUZtEmOafcBMdvVfTqYSj3UvMwmCJoBeIhW4/T98awHNNmq9nSfb5ZuiTyKdk1vwb
plyzGSLfYbuc7F2uTB3lbL3iEpfa8yrUJ6v/xYy/ZgBzoo1/dnu8Ew9ly3WXy3+Ttx3sO7l9c4iY
hliXlpTHBqBGEOfcp9qYtf9MpsrN/OzAYsQ27l5OxtzIVfv1nmZlgjc2YN2KVVf1+x9EtzR3mH9k
AHHgq1AaTHShCMKUgehQwG4Uu97mG71qVzLIfsf4hqlYww/2YerCMRU1/rldrr4NLRWaaG8mmpX6
HGRJZLQ/zpXew1fiLqmiwqCJaVKRfNtpt/P2Jke7bwqAilwTAl2YgdoHQGFLDpjNA1RlzstGwTvC
+5UbVudE6ou9uE3fSDVRulyoPnOgTe++MtQiRrpO8ZfVr1XNRqW4JdAo7P0U9o3cPkqrYSjTmHGV
kX56DH5roQ/zts8tNWOuiV5KzhrhNlFxs4gWZRKQJXsLw80lgqbbGrGvtkCUWpOobexScThP3iOE
rze65YnuIuVE9u/tVE9/1k4EFM4fFcCqbe6ZfBXQakjbT4XERIC9He1UVNb4R8mzhFI014uYDS+R
D3slFuBLJtVc7YUSbxq/yS6bjvE5YjVPSWMqxNqnpoH5x++s0EHdqQFQZzF6hhJPCnqoOVMqLRLX
fR1Tcr0ZMvMtn4l2N0s6k+HXaDNnI1V8K3HaQ64rQBHhvJbB/grxiI5WzfgCeYnCrCJJsLJpEt4x
2N7iH0GrpxK5PylBNNFecf4q+oh5AfYmpK6CYO/TkJHD9zrjZmUvK+Nh+UJ34qwbJlEjRYf3u+fg
1UafN/Pfts0kfsLFn+4iXjm3saDb0bk57qc3+R+HK5tmZPusHgODmUa/PhzIgsGBxHwdsmq9/ACu
cANs5F7XT6OdI40wqAyvFcNEVuPgnEg6HC0rCUJW/MVPscDxfuz/oVkqR9nSfQ/y59qZRFc9JUCz
KDKo9JubVtHIwTJE8CIAbXyiRLQMqHpLVR+CX2B5yleb45t9maVfis5cPlOwJWeQzt4XnqwF8wDV
hmM+dXGhe7y6M8ISfUBs55c0N8CJWVS5W5vPhWUlziCpUTvcmaPSus+vf/9WfRWZMFH+AIepybfv
onQbga4035weFnew4O9R2bWWUnISNOqhQpQ83MXEhL1lsGEYOr1jxVk3Wed7LnLM2UIq53BpgfMi
v4UA+i/2AM2WULAtuDQp7/o62xvOtujbTeW31LFBkfX4Q9ROX2GCR2ZlL1vQDl2u9bb8WMM9Zx/H
2sWYerUKZ4iRLJmIdWJ4w28oLyCg4qpzFLCtfOIH9QLqY02sA5pKm+Q3U6F0nFJcLusPtHE+5K/s
/LWGUN1j69WkWfxJRNUsHrHbOba/CR5NqFnDWmGW6zLcUEDt220daELcl6Lk86K80CNcHPhH3u3i
2Tscsqa7wIyUsAtbvcf/H1WNtF9Bedhwr6bDQ7XVOKSZwHPqvvejnUNASERSync7qiEdrwT8VWMr
8/PhJncaASppok7C8pRpiSlr2Us6Pjt8/7kzxGu4hI98br+TI6R8tjTPjv9A3UgVIKCi2HzRAJ+g
4kJDctwBs/3d96oYJPWfXbWJEdyWd1XDVxykH+N/QSFs3obIw2ASVwnYtFaTV6IXfrEkRta5a3Ag
wK3V8+k5/Rgsmqprygvcenb8KKjXRhsdv2NHQfysqhr+ix4Y2LDihL4ONyC5lcl49EQBaXYEboAn
bF0tY5++b5PMdo47G+t3ucGpFtE3MmRU323DWR7sVxZAvNUFPDlCMBLXIJOQh3d0VjoTfB8H3c4V
Mq2JbMeRg2fJXx+SamDtoBQjtuo27F4L9/GSfFHRyg/u8oCO6HTdgjlNL5tCVl3aQbDOccTqk1Uk
CHWHRet/9G16/aRsQ4pwBl8Mfk0CWB9sY8um//8vEDhr0rPkOruOn/3LWjXkrQ6QOnwQgMx3Zi3T
yC+4XfYukFmN8xp8AguUeSu0jqCNwdXKQqjx6Zqq7AUmT99vbUWnqOQ83I+bNkQIua8MvuhnhgPf
RUkI8oNmTkLV6HpkAde5ip6Tq3vgvL74SkpD1C7FZ/cl7Qr/9VQYbjCNVq2CctTvTPYj9B8j4qtg
OksBT1QCBJKKwTx6wTqxN3+1N6akjWqvXNdZNS1n3vqbuuoX4JtMFzV/oKvwl/QigljuO1Dmz3l/
K0h+TaWuAtJOXKjDFJyQb+lJanyowGDSnqLFHW3Eay98s1NwrSB2yQZxDsMVo1wnDJZh/CqacxcU
kZOjXz8x7rRmvl+B8exymqfPRq2RcpU4oBulyzCoQ5qSJgeWyiHWry8JDhwUo386XTca+siEPkmZ
Gh4sROXfNdkVdqyEZzTMeR4UzgkSSyBjCu9ILF3Gd2dymo2Nn/L1+CZOb91Y9Ma3EYEMX68YkYom
4uKaef970qUI1zDA+2EVsERPU1OQ4bDTnoLwk+33S7gRe0O9R4kNEOLdq/0hwbbKbdbjRPRVr/6N
kdmNzS67DKI4UoYFcpIwvuYSpT47JgFhLPVQh3siLyKa9hQZTmYXcYrYIT69KcBTRVtlzybJgkdR
neF9Rge8q8U8QITPQdlin7itEQiYNhx/cC3oHpFXUTCQlLb5/Ug2tZgUocKYNIShY1do6lXzET3D
+Mp48ZOBeLxgDr0+TyLYJ/9a7BT9I8CRTqz4IYULRUglhhjviJfH+zpjIPTFep1u0BFTLrfDk/7n
WEgco9IFL22pBqaRU1G0wdMydW7fjY16A2ZGhShRKPGnVH1o6hp9Diw5SjieLj7Du4OsRIFqE5gh
i5/d9qCGb7P+EV+fD0/AvDKXHpa1gbWnDC0sZmQ8QfC8oVAqPdARo901IW2g29u5zy6Yp3BuF5hV
WYZyAzVDHpTYrjqsAQ0eW60f1JzqXap4eKvUMFRS357CdvpF8apxzdBoui0ol+EW1JC+ScHEk/WP
uM/1vpi3IwVYca+RG5KUNOeUkjzKEMlSFQC9XiXji0rQTZQ6Gjaj6znZQRGqbVYSzGpQwgDiUNTk
Er6nMdHpicEqtnOjHwobtKobCGCIQAOsDnA2j62cYCwcbc/Lv+d7s15Kw1aGntX+aINUj35R7JRs
nZAZvcsPEYj0douG43bvfb0wxwrQhGhErBhpBWMlXeWFvt3sWomgHYKEWW50coK7O+Jb80gO1OA3
uWAWXr+iJrasOILj9bMWaxFNID6vlhtVntrYhadErwWaG0HucYUmx65Tzl/GiaggPywkYxW62lg8
sD40+CPIjsRQEOq0HUGZCbKHMhS9ZxRoxUNWclSxTpNE8JShwJPZhwGlWrPxr7830ycjoj+Q8fIw
uDJ0BP6hNs6182sAZ0WzJ7bm+bYK9nJXF+T+tnm+yHmt13zrI9qSdy+cFE6/bY9bo04AtMj0lFHu
8I6C3xCAn3sIhT8d9F3Ur7w3B57OzafKWlRmGpvjRdo9GMbMLeFy4h7qZhUhClekzz4mjqKvB/5i
zTx5QfTb88R2hKeMsPjgnk4M/uOORSFWg/u8SSKecXmqt094wqN92RDkfY8xxAPB+9MA9gutAHBz
6Qf2IejIdprIqr67rFdVNHVEuhdO6CQhFnDnLvdIR06Uk6Fez5boVvF6AOeacpQRcFfDX1Hp0de5
ws8ZLet7EK3nKKZyVRI3n1iI1FWlUKTjrg4t7XI8TvoiBGrIIoNijqQCynXqGr/aHhWZy45Zxk00
Lh5vPPtjpiAywObjcXCAHnynbUlLEb5hNj1qAMcTYGczAlWVXESkQsMv66/Img/Wa+M0kopEoCBW
5OLB4s/YszQdn/xRH48OFj7CcitPIQxd3qpqJYwHE9TXF/+FU8wtxfg+y8mtRSjLW7GdXKO+r4ol
LyAardH4SF9E4w/1GiaA0odJf8T/6qLhkkwY7gs6IErvbm7+j9va6/px8grar6Xx1tk1/nzdsTdL
9sVbdljG4kV6GhK9DIRRoz/LZk0eiqPfU1dyjMjfOf49NhCavCTp0KdL+Hsue04B/aqr6zvNLvIY
U0Xs+0uwrrXKgauZ45D2bMcJfAIAtNXRSMjCx6F7OJRqnRfsz+YlBZEs7c7yyM3gkQME8m5RfSOr
1wUowjGm4xNgPAd6Tbbi44fO1Zpu9mZ/8Iywl/IDO0ZImqJqoj0EzZvSTOafn4D1eA/vyfUPnUgH
Tn4NxrY+wDZMtpULaXu6xlG1xbp9crUvVazy0Bgk/VIeebAuxHBBNRNKYwHtzd25mF82u5VCv6gE
pkFKTSiBvyUfY+jX+cONPjA0zHLmk/5yWUnFb0oitp7oTVXRURmxwsSGjCQB/Qkl8I89iv9W3wDv
v9VQWfuiU2gY8C5vmBZTlt15x3KNDVYzE3gWH7pSn040PDYCQTQn/dTT4BCO9HcTkFPR7I2QDv5i
4wQrHgAFikuo774sSlGK+8BC2ch8JUjeOhpa1D+Blc7WIUl1EEW/D/RW39kBJ559NJRQ/rpOVmPN
QAQcLeGWqvWjKFnRiGqabHYj2y+GmRRulVI28LLcp8PnaDPkp/oeqDh4Y238t6BDSc/WkmtWZQmP
D+QblI6Jwy8XXMaveVA56z9g6f7CDqzlBKULSutwfYJ/Nq9feQN2zcc8ES5XCJ1L1Kn2GJTBSVDX
PcvoxHgkh3ctPGI3jWnQEDaPlPv+oh+1sm66rfn0k3B7s5svDgK7ZlDup4JxLtAmla+BCu8+vCKm
etLpasI6FGNllOycCRDa7uhBJ5QOa0Smuf/VAuJfd/xKPY17vMWGgz3C9rGtVmPPoZjlH1bOcICN
1p5YTyHGnx+OzohcGYfKOMIjZa04uz093Kf2JWYTutMbh0J+n+lvhQoaLFeeKGVjEakbKFOBFOEs
pfrXmkBWw+oeNUamExwELVr+XyOqf82OI3ykNqI2LcWlTGHTQJfOkGpR5uz4NckVWB9PI86+QggB
7EBkaM1zqy+OVsGG/s4cLrtGz64JLjRTjFP7RooHlBSTbJwrd8Q9GH19NcvoMWmRsvH4YWE3Gmv2
Ay1TmYlG9Vq6rJCX8zEx7H8b6ITDVQmb9uzyjwxTN8iTnq9FyvrUdAsh1STzczj3Zu/pDJctAa56
hCT3gxqp1wjDcEDB7ySdnRDcSiNgY1ftvRHr0PcJ9T9u0v9UXyO1wVWDgLB2S2gbJ11fJnCAaAQ5
JJ0wY3y0BNRopDTrOsAMDn+x73tpYzx+ITW9QCk5jWjELJJLwf3Ze9+yCUSeGgP3wg8gbG3wCmvm
1pR2TgG9oh+QKfPMiMTDzTBmnvDAFyoVcTfA28MwW5QOm0CoIDpNKAgh7ThZ9Ry5gkpSdom9sHIK
9dHbqe2NWOOfZLa+hcDgrM78I9d2fw/x0/IyLZRXvHI1M4JNTVRUqmxwNiP2GoqhtBtc+uu38uAH
geIJLWyGGID2YyaV8kjL5DJyjyw/vvDl2xygF2Hh0hf2lFZPebrQqegbKMhuBWcV+IiuVjzl7GGv
lvjMoih2QXNQuM2oDoETXcQ3V0yQVW4XsFjNs1QVWpEbay/p6xXOiZyIsXZA6Dh/C9Ab+tx6pFDI
ci0l5A5b6UgDRRbuk7mxBhjBd2nc2HhHATmVx12qp73pupFO0+Xp35KluxjXnKcbPXTG6UzhPpzZ
uM4oE5nGd/PIW7b6suBmdMK8C0YR7IbmPOOBagXe2VHhETFsNS2vRMmFdTGESxyjHtrrbX/ogiou
3BJ6Zi8JtO/6T/G/OIrJybCSROjC5Gx2psSyZv6cO+P6xL0uGlx8PGOL/afuJpxPHnvbihB71+Wi
VT4+X0RmGVfpOJNlQ2fKax85sz0in4v/ZnfPJobJ/IVWE6C9bjcEyFIcEV4KktSarjBnYtPUHieI
tIC9N6Z1jdtPFYmO9SPvAksfFeb9w5PP6XYJwCd0HW5i0aKy7sx8h2furEjPh7PaaANl7O/FQF2e
orjuNrZIxrDbmimc4jqx+BOWxEZ+Ozn1ZTgPsROB18GPkVdGsIIHoVx3M1hhgZWAApc14n7/D/TY
tbrRr3JWi+vf4EpCtbf6OG88lx6NQ4CVugzhz1F8800D4dXq4kn2Ejj24vCbJWLndKPFHMxozlIH
R5xFnL9QOBVgM4OXDJmU0VcpOZWHm/rb+z56/ojwyra+/QjSQTwj1rzsLZTSMaH23GOq/jnxQzH6
90/BUDkF5jgo77w19+ptNG5NkTM0QfH3m2c8f0+psON7JE9C6B3ononTo87Jgi/v9IPlarJ75MZJ
hTulAzPUhMS5Nuhu8B36KFafxivezoaTQuB6/MzAXmXxd2Bqv4wjrEnCpf6NhZDdoo9fDiFMGDvt
Hf5tL/Rf6LMEvQfjIWAL0ZvBoJoDnxI/+YFo4dznvjPgRx59d7ojXXCbTHzL4Hw8e0ixX2qkyWJe
ls9dkyEVxixJ6yU7JPta5OD08aw2+bOjSLkiz+PtGvNw6Yxw+v99NgXidKdAQwNRCxFpHO/T7ISV
yoO/447DOh5VpEb6S2z/7Q0ZlzIULhZEmM7E2q3CTTlKFissSAxswydfMolyE2GRn1dC3dV97M1s
LFNG0Qc+guiEnK7jpeVcU5+11zqC5bZg+SS4O5N7bAf1Gi+6ARxt6Oi1ZO25DgOI32wWPy2ZtEHM
XgdrHCsIfVLPK/bKhitlK3y/zJrkNdKrz4TqhXhQkfnDvp5sXEOb1yWOZgLlW1+z+Fx+BXamuNHr
cUMVSfZ/zzfC/hKMuruJoR1nczXK1nWCaUhBlFPudV9sVMhcsHcqebu+sCb2VjZwDF2yvVoGyCvq
LCHsKKt4oGXmp8KRqZ9z4/XD4uCyAtxnMk1yAw7JujSuwnr0uI36wJ6goxdJSIYC3MkSpy81pC2I
7IJwsBohvilsQ4nurRIWJZ8d18SQuq1CFlluPBYbr8aZrZXRhf05mzL0KcSddijuWIPTyyY3eZeY
HKuISvCFkwEkE9zt2qCjQJy5Zq2WSoPLAjtt1BsIQy+2J09+HAWvqqvj12uQmD90HVpCN4ZyYBmK
EcdeCtVzhnrumr9jA8Nn+oNgxtYJhFUT+sx1YZcmsVR8rmzoh5luXrysVaKCZ0mLrawg51TLKK8x
PgDDoWPwzCp7Yl2xlVwZrzQY+45VBgG7zLoe6EHruqaYSnQ+AwN8jUnczlaJ2+LhvGszDeX0U31R
Og1mgPJkNHkxEQ0B/kDxMmjsRZkmNlh7rWLn00iuBztywyUOJvGSAuFY5O0hijMp50mFVc3sdJZN
la5APwnC2TGtEdaFfMDL6TIQCvR1yZEsAEVLGitgWCWUyDk7ilUy19EJsT3WI8XQI3/mK44SXskV
HilE6zy53Vu1nb09DHCr+VMFdTgddtx3A1d7bfuqujoHWaHj+rr3IszmU4SFFF3ePhsrm4t6K7lz
6lst6pxPaOzoGs4E3uvXDPA6Kt8iceIX5L4OxSTrdeVTAz0azI0afW08Die6aAaRZ0kj3r4gec5C
hGPQ0datsS6QgJmSw7D7rxo3p6lOEbvyLHWwYqGQn47NmrZ4bX/0I/JBr4X/dBpuHCQLtSsm4I3W
IHXmz1gBUex6m7DLLhhrTD/45iB1CGVLdBy1HktnIT5GqpdtjBIJg6gRFa6LRommPZB88sswIwNl
zQO27ndefMpzyF5juwSNGepEHkREc3RTEchqqQOB3KNCskarPfXvQOL1HACP1dP2WntwEZEkfUhJ
4tgFyt56tg4wtjaMT4JKvqRWnvPtcwPfqzEt1cJrtEJzWnBUYFfBhttv7iBFOtfYVvcq7y5VERQa
bzLC1MPqjv5OmFHmPnaTYvNXV0g+H/FrxugsJDSm1bAhY6NyypqBNC99so4F0IGsr4qmQF1HwwlJ
slEv5QGPMrnVvb163blL9tWRjaTPugpw4Bd/HjeM7J0HwdlW/DpdWbkDDrgf0xjGWxmfOmW31tmv
pYPfhkYYLSKKjuRV7BBGL5qTWMr3uHgxMSTu9dcScvJjZX8N+/ts5Zk3nAHRr9iRcvhLKq3O72I1
MD7JRwykjewN6SYWloJzscbN3icTsvPtP2fqKuFG0rARqbz5+2pnaD2YyW2nXX/ox2kEv4n7zFVl
WFaoElsqFVnHfG+U6cadfkQfTYTE0mORWlL0RtvXLc33kWlaV31UeNvsBnamSBUdNlkg+jb8mjCK
VqQVnikybtOEpiC1PFkg/s1KStpo1dG8FhXDSammzbwlalhYKo3h6b1Mwpdwkj+7s6veOQVpyIEY
QQpB4UPGbIGTdNZOfYvbSG2nrmMlK/8E2Tv77nZQCNin6KL//Tmspu7e4nfPf/AToMyzoit1BAPe
fOOqwDPtN87FjWdlqrleUa1CVvQ33YQD2v5bU0lR9RPxo7jexg5y7nXp/0ncLvK/qdtgxTGniMFa
3w84nZku/ZOiS3znIa9r5c+8/OyZB6vTsG6Kusi+WcT8msQsYdwDYTk17BgQQAEGgiS2BrPVu3Je
nSUvrvGY+1xk+2TSGlvA0/GrZZipmoOaVGsfaiULeFcAuvr7AILZnDZfQ2wpYBWQNf3bhy+LBlUp
9EekUsrdKf96zDpmICR6noMsq+GuONmYjsvK+GObfu/FseCl29RWgQFpxwssnpKvDIsUfH97152y
g+gxIE8PYhfIF43tj6P8IQ7yj8aU9Ch/EBQCC2d8tka7vXnS0XR+4zCLPWBlYL+oWzBk1zk6j9dp
y9LjgjomCbJtnB0+OUrOL6Yn07Gz3Jp5cvr9UbI9xx2mvlSbNOPv0i6l8hkKNfeDacSFVa4goEi1
ml+sn+X9eiWEjbibZtmjSyuIqN+t2URHz8vQN3kC0LM69lgjKlvlLqIZi/5DEmwXLxguiVGGmg2e
AFMA/cgs5upaI1t4bjiBvWg0XygbCgFTLlPQ6aksEPHGRGZww3O54skYoP8zL9f5eEasTFSGu+/1
OPLIjc3Ed01BjRhQ4I2gFgIceRVZCFYYZEbqI3KINGQCVzz26jB7jlY6Mrahv7lWWuQen8iY4eLq
k0vSPKEAE2nW2O+wcPtfcKuWVbICyEugTTwv1+/Wqskka6Lo4l0Z7LCk5ssW3H/PkQMpFNUVyTIo
Jvnw3jcZTaKNpCoslNGoDadHRR19TfYS4bua03FRXM6WMPc+bU+VWJrm6itWsNzs9jDs0Aby/N+8
w9/SBNSG59hbhMgTYOkBa7pVfMygPjKWgcckoPP1bfnTTaK9q6DVFXytVC00ILaBGE5tY12tHJ8c
SIfkExi/0x+vxfpPq9O+5iq3e70/F2lg/RmiaJh44zoD39bHxXnbUVqu9vNdw5pDIPCgeCgWvhsF
gWwdRKWfcwLcR57ANIe1XaCoHSsTtVXNLr7WxgbL7aOC4w+C1g3N92BEcSWVzxaZCFDdYnd8z9r2
TId1p1auUmj3X+YI3W/1HnPihLO9f+NTFqE+yFDL9bfKqIQ7t3YBNPGmmsqYxRsNVK+TtGMvcg/K
wlQFV+xgWQUETLA8H56i30mErJmFBt32io/AnkMNGVurCfc7JJEOLB46QWzARgxVZnaHBMKIIRrp
39ouTxHiQuq8FguoGM2tr/g3WA18RX197SKY54Dz4m5t0Uvl/vxSV8T5MwHCv95J/myRNQYNoRhO
rRhkvGKI01Z7otsmf3mpg2cF16sa/6/7MeNTTdeJTsEepZfPMJT0d4zCT6eOnwu4Wk+AlrfyO+KS
fMxQ9WFjGlrXN3GK0kmiXA9GdYrWDIMnCpxd7LRNcgN9HOgRRZwSNjN2M2sj5BKOBU7XTGEk2aLn
vY7slZV+aKY2ncq9N1B2sgQ26tRftKlnT9J+LxDLM6ayG9RLMG5ES7BjgNMmIqnCjA/hKnAjFsJE
OfXxxtQv+3qq3pTW58WIgd7VSAL1m1rPIIsUneTU/CH1prq0KvGNAMiozkSLDuyn3V1QqLHqpwIX
pE/OfD2PaHb7ehINQaYyKmdAzlAmKlj2/I5rpyeUmqd24lporj4Cm6Evj2tISOi+m7Azq4FUJT6x
aVbD1vki4imEHX9HmCr31JmiBre65J6KdUnoBjkzwsLQcv4PXM+qIbS21CSGj/SiIYBJ7jEUoEqW
KLDAKMc8hPbA9JaDQI4pPHXuQybnxKBJOL7BfBwokm9NYRzjAY+bkLmGl2l6B3ao6FaWAA3+Xz9m
Om3F37GcJc6oC7R09NJhPwToSOd0gO4c+Fn2lPCnEJ6dwENFyej8LHFz/7UAjurDyoJFQXwla7ZV
04S6onMJ66bGbEeeYthEVbsElE9JIUZBr8kw1mpfznYC5StRuRyckukgHAvEEGGeOBP/5gZl0KqA
e0XrXzduDX/+8idM6zidah5JZBqJqfW2A9QaUkVYyJV1iAhO8Naz+I1ILD/Nhsd2kal2vRq9p0lC
c2+Gs8yq6qWS0yoVcyaSbV934MUrz+04cfpxISKWSVVoSjKNUjbxKflArwQ0Mhaaj7R3swUZaLsm
amychpq0xCEiSTzl8vN0X4erKqpEbu2XNJLhAm4YZsCI50qMhluvwFh+BCR8+AXcxXJ7aLMdLAW2
4MRGjF7X0IUwdL34x4Z1MwTszSWX/vo/k4e/2c1yEaRmPWJWg7Jj/KdGahKp9qtpF94yUJCHkdHR
eIvIBkkcU0to4Ww3QmP+Yslf5zGxPENN2yve/jb95CunuD8DweW7wTd1NtpZlntMpDJDlf66JcQn
i+BOpw/1AzPrPYQPIvJ11ahDaqxnQF2GEgUhc38d4AarXds7+mm+lLLtacTKQWP1cwajqqGpH6PI
GS/2a1CtjrZWa/ozMjfX6VxtRojdLVxiTNVhJs/YQRVeDpA3DIfJnRVX4nAXG/kp2j5K6GJ0X89n
JI35RWyadNQh2ic2+O9HvOOE51dy5Ec4I6M8Ktwv/hcPcTaJABeoD9t3tYqJbFJDTUPuN4JmI7NY
317gl6UVom+soQmqeZnY1lW2azqcv4/c2XWfVFotx/brmE9/KU1JfRnxF23v9YR4OsqWO3A5S+5c
btxKxDRWj1AtoZwpYFA8TPiu5vt1N/edjt4VjZj46y6jXv/INfOA8fRL1yA+E56jtF2KktM95cW0
AJy8mcV1F8j/u2F3c9IP8NFg5lwDZB+JsUkryL1yxb2E13afCKjuDQOJNWTumS2f/3PZ6b5TjVUc
5SZTJLYZSe97bKWUygk6nFPpVjg3H7NC52tCh8/SjrWX/EbBl65ulOiRoxp3N+pfUHzrPGzkLPLn
sMr4Ywe6lLvrmlqfb4H3n6DGHalZu29nnxqu4Nw6XSvhNwy21XARAj+Cv/SW6k5M7vtbl2StDPYG
WjCufnJGQGGbsQGYuSRcna75z32zvefIRz/No+OUJikFwGaJl6Mx5Hx+BRaIBH0+OWREQweJWwVq
qV68kV8K6odSpyfDq/jvdickouP7my57Un3mzFL0h2UbC1Q1YPWm0KmtWBWl8Ho1Dx4jPhV4RG+M
ukgXYH2qxkpWI6EHAfNdFfQDEzSvj6R07ieDkmJ2MZlkBwKMNNQVPttSIZ5B+pdRsfZEUqoaGwuh
5+IfRqTw/snUAl3+ZhrFq6nFNGHqBXMmv4T8l8OiGfm7e50Ssu1KJVeyBeai6/w62WyrStoRtlsB
VIiqwSAXRTq6fpRScZQlVnvEepnj8P6mEN0qjv7woQ/KB8snsxZhCQ1XKqr8153qYHFliR3ZhBcf
yPCsVygGh/LTxXkWshYmue7bfMtuK+boLz9RUQ9ZoZvMTr9l9Kd0vcZSRiZj5fdkxG8jq/DeBZV7
EW6mymSeahRFa5Ca//CxTmQh3S4UYXIFdnFW+WN7IIu1kAo7cEfc8daUQ9imb+YV4Jjpe7MZ/nW2
23FtPmZfFSXivlMrza2YIU2ucyz50zmxhN0fg+e4AQ3IDhuvGS+9PdrhnVvyakCN0v/aIfGEeFSV
WZSnLl0uRABjeO278bFB1b8DdY/Ycd1XEL8AzlAIPxRCxL0J5ng9R4hGsCOPwCv+EEVGBNtCPtxd
U7h0a4pdO4xDNLIvSkIw7VxKSuxFMQ2RZVbuOzpKFL4+cQQmHsZy2t2A8ujJvIqfIwqHB/pamkFc
pLqiWhCxfZPmRyK3IICwjmC3gXmB01z+ihzuhYDeTGHuOtRm+CGGjO64OmXVR1qo29x6v6gzMn61
YYKe7N/MHCr3GOSHreu8gt+y8onkS5QiG0oNyFmwIXcvXYSD/S6md2YszOy1sdS+RHDNQyECUIi9
iBKU+fDvH235jtoV9nRe5y4AN2yPQakFbZ/TpM9lFaJnsKFY5HcdbpfyLbtlJ1ve8JEjZcDA6crI
o8V5UBSpERbPQLawl+rE/xb+oVHHwFPE/J0Kt1MUTLpggDzC1dh6uugYB4YEMR9hYrhY5g9Zlqsk
mJgVzboHIHGsYaaacGEJJtPsHciSYHXW0SEy1lJad2me/LZbAG961IQQNi3MTKCBiQ8XvfOVFNIC
8wdR+uejHHxOXQIozb4TLFwpG/i690ccWc8wLMuga81WcDO9aCiDQHpIfcvqU8poXEHfADU6yUrD
XHcfTzXEll87DvsnpnXMc2q3LQDCB/dYQuVI46nr7IkTIuYRm7Uodu3+k5RBmmj3KZ3H+2FzDfER
ZMPEWckTecgU2KTAf8XbIe+c96DfatNa5GnuTzFLNpWpsuoEwXRBeNfHgoJpQLw8A2tjUGnpUKNf
q0Y8WLFPGDvL70GTOHfcwNpOFovxLHuuPfQ/ScBRWFEsgAwwJUEh8R7vHrOPlj/ZkJ+KtuuSpdqf
LPKpxIRAwmhM9AZU6ZzjbDntBk7XcSKHi5Yn4+Rrzp7LZ89mlqwNTtzMP4XR2biRua8vGwmaWh+A
LyY9EKEZakPI6t6kQi1f4hzYVM0jaMJ3UOga8oleyT4FQea1dJTyTa8V6tjR8wbxbi9IHVL0kGhG
VyD3RV0td5qvZDkl0ZcxtXZTGWnjvRs3ZjXOIVtXLM9sYjLMsPAvti+QVXZiqTJVM6mglh6Nz3qm
68zqufJ6QunUaE082wtdDwiNiiCmOw+I5Qa3r3rsiR9bdmQtw+/mrT3u1jolzYBHxzAWz0k0PI86
o5q4qnqUoXtvAjEVmhg+eDm/a+/jBsBlbLjnI0AanhlYClCT9wzY8CH5QmZM3UqW3Pi+sc1YFPlQ
H5lB0LMtNHGRpJ1lL/LsFYK1u2SBiUhzL+3tPpVKPV/UvQRslyAf28idH7VS7aa0kmrdvSSEGgGy
gLkV8JEL4nn+iQxraPd36YyIgufWLpbhjsNa3XFcuElUTmsuXFcF7M1haThvt+rEZxKMLLdwhx3B
xI5/5xoYG7SQfjcBwDaUDT9tBVlRXuKgqMwyQNf4MUjz13EjG/CQn7p1lqaguFWISiT6yif/tXxb
p5wRLvWOL9Uze7uDLFQgp5T3099AyBiRcL7ERDGY1X4BzjLb/CsKAhG9a/B9kehZ6p9b8kDeXW7x
/n27nILEo4vMhb8v8dX2I2Au/tu2PjW2h5oNyyh6x8lXWV5OXBRJ9NC27/C1lSM9PQyUHFq1kwqZ
hWbv2tnshh+mg1o5yO8jSa28vMWnJhFCBLXRSFRl+9TfwstO0q6F6ewGVmvkvxoAXPP8BXS2Q3wl
oNpzFDAeRoMA3cqrGnXtRAuwi4G2qMtOIJ09dzscMYkQR/h2tKzgGHIweoG2dLem0x69+5PGd1Iy
ElxoNWBUYHUCjUbw50TArsRbz841VUD2JnIckrCKpIMMuWv8pHmIKEF0drnyt32tCHhCebpVyhsV
NzTiVpE4PJExapJ1Gh1/BWqWk1Ga1TnzmkT4Gg+rHliEhUOvYmW7MFaOqCYva2R6gtoeZya6zR4y
vvnPp6xlECc/goONiO5H2NJImSYo+5b69J0GKoCw4l/aBTL/86Xh0bcv+Uzf5JotMc7IkBm0FaCu
6Cnbe7tAMZ+jnh+q+AvOLV1/AdE+OtIuOBw1rVzSkwaa2g3+FbhJsGu6uBTPVMSTvaMrM2aOgD9d
UuN6wKunk8VOvbH+9agGg2BYE1typQOPFBJQFcBzaWbe5clkvKCk12BaH0FgCt9sb6GYyiP1N+19
smkr/0oLnZicj/N+ZUmGD/vs//lIt13zyQdyq0F+hNAS0eCXxXE+X/KbGkzHua1SaBKX+BZMRkxj
96SUhS0A+qAmltlIGD8ikaeePVb1h4NOzB/G1aN7c0e7lv3K6XgTu8N2FUri+7A6Sq+E07Vnyc7F
jh3mPdVgVN44qpjt7WIfyvkmvSdGsy/mCc+G1RCvNN5/GSSTS8LU2aC89uhJhBf5ywRLosi/dTX6
hztedjeTYUPdggcYbSRxnaeJYY4EmgXO9Xa4b4HRr0hO3IzlYL71OH/HAR1YTjEJyk07kCclY/zx
c2rgSgaT1TwZoXPwECbv13wqLKBP6rJQrkTrV5wJVpWPITtqoSXP53XgNtBKjHedtu59K3xnDkJW
S1I3FDeFVgnz56qY24AE6+c/42GirvFiVnrKEyowIoSnfDpvA8mPScfO9WwbWLq+ok+7I3adYZAq
bPYp57MR4uNaUrep5PWs+/eroSyVDY2zSK8CXuLs5uBDPD42YibO61zbB8qSNNpTy5By9EceWI/o
pXdbs7r2qRMn7jKUD+Bl80oTybai9X4n/h5oFW8Gu4sVIw1cRPUMZAXr1dZqOduxj6M8cBEUp8At
Z3vuOdZMTa8EAY0kgFwA/DqKDCjdKWm4RP6UdD9kM2HVwe9YQEfa2XtI6/mY9CRf5Aek095wV1et
dwSEEdu5bmkvOMGtM/hSgP4Fb74svl3NYUOzhSU/J/W3M300LfiE4ptSnwA1aJhka1/vgRUzQ4tU
3T4ecDTVm9HsQnh/m0wbpGevDxWVoxxDaLvDkFXn4wYSDwcb3SbeEUgX8OqRPIeTeMHiJm66qTU/
HinXivLQ7teyUcl1YuaqZqC050NyOLGUIID1o/RJ3LqiAFcZk6fg5EnoTv2sgM0/Yn1jn3qHfDrj
ACotkywKUUGcCKqIyMd7nLRqQhaGz51SWcLJt3428cYE+CMLOzwpAKTPrdD3dKWha741eFXOQW50
qyQHxIhOQb2Iv9SnKDOIqFV8MDSqOJ6sXR3aE//c4DJcTN2bbE3rql/yg5Ih/R1swOlS65vslxmD
zjTFiuWei4LVKBTfGYX3Izse6IRRBdVL/VbmVA/WshDbWRcQxOP9BNzbFozcWw/IBPOufFW+0l1f
9bQsCR3c7dyz/2TshqiiPxwqxK23tlAtgLOX460D+DpLrXfi+2hwXR/jpxQsGCBhQVAIxWaWFy8P
RrrkY+cl+eQBqWrlMphPqM7wR4JCo7Bzbw0P04n5T5dMSBnSg7MtTHA4CWHOuWF8dMI4ZI6QKN0Q
RcAX+NYnAW5Dz7pfqDuNKjV+AFzNh8rmvsyxFk86X+DKefPFJDGw0ZaBlZ29O0lBpy/JW/GW/JML
CNVl5pSyrEW+zHJFw9IPWPEG5zjmR7gAYrR0Z43qDinbNMylcRxr2HSyyfb+JlGlAFKuTOgMGFUv
SpUH+TKNv3xAogyvnKZenQYWUK+M6YKZKnIj6qdvy/PAuYbCq8Vh46cdo5RFyP+bwf5ytTRTgm2b
bA4Oi2EtSpv/5T7ds6WOctuAaruBrCESXWHpOlz9gSy+sB1kLlo4ddDy0GomqJmL7QoOKzHAZZYk
XdivMzyYjsORu+22yMevWaX6vMwBFHC+ICUIenYWbAqHDhg0xO8wvWS7ywDvXKEPfnAiCL0ZML0U
72YDBLe5tMvWgsu5fOUZdhZaRljMijvx9Jha8TFRs1mfbbbfUcI6+Vw24ZGT2rgrCT5F7zR7BEdk
aEMlL5Zc5Ad0rLV+gCdx7/kLwITTt1tkYS2pQGodIoKO+Sbnr+baygWAixbIgsN+TCKl6qn7gbuL
oaurnVIXz0WFQc6ux3zAOMslUNDNtfof1eMcPpQ47pmKKsYCT03zv0ERx0jmVaEsW3w6SsPZOToA
cUZTGerkFEB1hoh8C07sMkqArE7JwlNnP9Pk/0QKe+XbbRgzhJ9n8jnagWeDA6sSTXOHBkTTXP+c
Kr+jhffHrPpTPgNbajVoi/himlwmMZAZg5FVQh3FZuYbsJ1MPjYXROcBltUOKw+tQNYpD0X3uwlm
IcVSNM9x31VEgWdJH2ZfDxhHSBxFakRepxxlLHf8PK8kKdevWVnmP4zknLgaTpRJWgAFMLIdK6hc
uQgCmDSMXdhMG1ECE9vby13gh6PAo7Xluii6gRsNsPYnOKoXauY8TIR60W2Dx08SXORXe26e0eaQ
FHoJj4dnKSNQj5yAobO/YfE67gA5iT6sLuorFUx+ZvrLCdx5E4y4HL+YPzwhW3SGHPstsbdlEOHq
89Hu5j4q/J9ODudc6T0jDGVvFJFZYtl9jM7bOUGrjjk8tcZW3GY5oAkAcGU6qIW4qJawyb6abDJM
yaebFSKgfAB4Ul4hEWJgMzLHY6jw17MzWYKTxw3ZQ6yCQe3XNEDy3AAqU5FBP2K29tDoS2p4Y+Qx
iO+qUe2zTtWAnghjc6LF1rceBbc8Jb/xEekD+/2VYN/tE1i/2mhmPZBSDobrLXYQz4BmMbwxfgME
ut3nez3mIdtLHyn2BgxtpeiqdZPiMed5m2QC/GDoJ5ZlCATR49pIozFuFfc8UCcxExqbIuhT2bid
PeLixXJ+ZOA6CPQOdiMsw77CYYXVc66ySvlWsdxfsAwu4VWbcFoM5sN8HYDZgrmqc9vJeaXUbQjS
78UchWdQxKiXT+X6KHKJHEFdASwTpuyUt3Tom0FnmYMa1s3Wn3uqyW3clIokD0SXeIW1Zyh/OXOK
p8+DSGkfzbho/IUSAZQF8n8eLPguxMDMQa/PPDpIfPxaX07IvBnqe6dxzeOyC/SupopQNSO8WUpr
oaEtKXACTvYcJ/g99Jj6O2CRcELlAE732szUW0LGfzQKi/KTXc9EErqhTyGFjJ6MZ4p9VuweEsNv
+a7YC315k2+/SSly+lnwHC3TgcQmlvQ2bSap7rztDGmfMiHLbGLet3OU/WE7LKQNt0/KHIcBdY6M
iEn3jM00YpdHj4knrT1/e1bvhNxbRYsQdz5vP2afkW8cgIgMMaPWwHLdSpq0e90rzLsMaeRMljB5
QBLvpOJKO31dWfc8CwGzN3RBSCrxQK8RtXGYYXpEF5DkmQoqm37LXXCd+SNjS0e0QbnoIwLB5s9+
tVVietf7Y4/joGwwmE3Ytw5YjEdSRjDTdycK5uwl2v2/99b5TOefXIFdyOJujGA/e6Eyz83k5Inq
rpU3ruUdtQ2pqkV9pXPu42g8s9NLrjhJ0aI0lz0D1aiy2s+eC+1uTPAVU8TIJou+kvaY1fEAx6RD
UU0+gSyxxzcswY04FzEN4bu4rHq/d+3czp0rAj5dFX5IMfGlWAlWFmiVfiEKyhHxFJ82wNUWTAet
RpKa/1ag9e/V7pnjL3DhyPnQVSAYMkqpY1QETxvGQC42kwH4mZI8QjNjyg3yhxwl32s6DPf0UbgQ
4VGRBUbnxZmDH3J0y0xAJlM6DGcXgWxF0HcW7PWo1FIZK2C7G6gr/BKWdrPa2C3DXZMbhXYC1cdJ
ztfn6d8M7918WL35j+buc+Mgz4nHXQBqD/2lVtOqOasF9JVayMBPJZTrduHum8LWibt52gksHskX
dLRK2JqnU9WRRi49Pv0MiE+VYfaGdupfJtIsXn/wnJoZjXkvSjbFH+PXFeOc5HmpKqDM8Mhiudlo
Xgm0dmE17T+YVY/vna3dkS6VKsEpgUMged8Z4ZTuVwv/3KJzgsVLvwuJmZeR1fZ2rl9boq39ooeZ
miFy58pRyYLyKiBE6oefy1w/rxMzvzlr9UDN1vGWSfh5gnJTkeXkUKDfu6plRwoH/BN0FnBnptvS
SPIev3GUdqHSadpkqx0ykMxrAwXv8Ve4yKUacbidb5VCbvAxoZdYO6VPVI+QKekqKhiDn0EOCzWM
aejjjcgLar0QpclX89GZY9F9R4ohxFk6j8tzvsUi8i7E5Rom8tfv+1iLG1U3SruMYMgDUHljHSlU
JTfn6GPp7BTmbhB1jT1i4BLTpBPaougAXDa8XXizjHLt7PEYc8jSIIca7jM6qlwLwiUF6yLs/6Y0
LP3O75YYn2zfvE8ymuGbKsnqnJ2eXytUY69OWmB67/MhMgVj5bXIytLdgYHRc/mehy0bKHz6CFPk
AOPrWhYIkRmxm+RpmSso1Fp5vNKpTqhVGSw58/G4HDkYcJLmTKkasSAFifJnfdCjZr5gFyTmNcgx
7pnloCv47OP6IGHF7ATn4LCRVrq8PUIfGSMRy5PVc7FhfQLGYwYJKVSccZmnAgkiNhY8nupN8fNp
ZQBZaoA+Rj69PeFbrwrTbNdMFHYClclIEc5oOGmwh57rT43ThZKnhMy3GxUwKP9eH1B41KsQd5gW
+i3SDLWbGZZw8qWkNtXz942SJe9GgyuP1fka9aysLg36SYCLFfb3RLeWrPAw7WLjZNRZkOvgvgcW
kh0JHOx3wJ9EePswMYa6NmqLxVmC3yIobUYu4rrgUnhugCVPRg5vpNJY6C9sGEWxm9HZ8snAsKoG
jGzwmWHZ6U5cJJDNb4kWRszv6E2XxTGIDwzX3Oaz88c0pLW2qxNNGSGiuVZVLD+k0pNimWnEA7zn
tzceIp87zqTAClvGwRI24ToE5KUfGHQUfVdDz3Yc2Z2eed+9CVDUtEHaHstvpN6FyRXOG3QvQ7Nl
c0iFux536rHTmH5FWEU8Y05oI83mnNew+zt/EcRk/aEZRLd3TYfDQ2YRM5m5oCxc9QPTylqCXZM5
MvkngjGlAIMpeG4WyJYcqR6EpOHyXy8T3F1SJX28O/cjPun9GLtCIATdakBSMscQmq7fYLFQQ8Rn
MPzWSgxDLoYpk8Nd0V6Myx+0dkWbTtaj1uv0j04s7FmqHOu7DsZ1iX9YMWn2bgShswmuPWvECUZn
0K2FxXaGUYckEfR1+EkO+v/cmnPSMWBXNr2eFDpthkwVjwl/LIE9QUN8IkmXVTFkzimZWJ2TcuZw
UBWsMLiYaCJ2dSLtiWP88Ob+DCZzOgyKMNmXlxX6e4RNrkjM0C/hPC64VbydzOMZ4ZKcZsg5I9HL
jO9jYQ1qBQWmBRuxZLkALn3dxe7v9Tp31cLA/zsIHA6R9nmHJ0U4wdLtfPulB1cifd1pCsVfbo2g
nZeJdJW54O2BDwqYagUkqVGKDv2JGF8kDvKCTFoNtm58HYx6z2iCPFLw0RH4TEbwPMGTfA6+Uo0R
XqF0sdyN5orkVJGDpZS4E+Jpu7xSsMaGqAkZkHZUJOyp8tfBG6yqg+jHO8FLsi9W5Zxp9PH9ekD5
uG4HuYasOfbdLmMGzTdAFGoBgMxUoWb8iKgBamqYtpwPm+iq6YPSL5DXmquOoJ1cnhEFtN/oNYyi
ODvlQo0tVJhpi8Wxhagq8+o9ZAtNfBGJdNg68QLZaIqCG3wS98u0vxwgq6pcwbOoxLUn8pa/nTaB
0HfsNVq0evbBjyiAzBduyLTBvYOmxq0I2jk/1h/rnKi01HjD8bpBNyCJxwwInATmYIqvRCbyqHsX
4OTUwyDJFu3vKUdBJPZRHsUaP+ZOTaHJQ0HxF13YMBqsQfz+GNeStevcFT8ALFqrwaWNmfTyjgnM
yX/lHVUFwVXI8Q1ajBY2sAFRZbdQFOIycozJuTmp0KGiQ7ZlHTeUBTywXLtzogWBLBNC+5oOeKvG
BKcncPBotPGleEYS55XPpMrYlENAEVb6ZJno/l3BGCsbLkAUq4GCMYJqjqjnXv62gbJw+E6Uoi8G
jV8IWjbblW7eaXc6bHKIKkIiC/f7wIr2uLdVCCA4R0GOW1G9lHuGnjqkcsJMGL4kbiepZJp4idUp
JllP/x05oLS0+qSa2uANKILSk1S7dFMTExxWFGW2wqc+HTobSGKJM64GpMnxlvLWbVTdvbn9/tne
hnok0WMCxoSXQippnHwrpj64y8hKKvaPXt9H3i8SiJnxMm5PT/Xw66sapwyOylfYHpKmptznRFBQ
9XmiCPUXlEOS+BH9A50Ygtt80E3aFpeTLb+FZ/i4HOwnV+w/Wlr0wPLjpYqVT0lFC+C6iKVyiA+H
O0B35ijEIm6blGI5txH/4fHr2J8lwXBWoSca1kbnWSMF7lQjJ1UfZjmdbS4Kvu6wv6jNsLIod+13
6Fzm5AOYqYTntyvKRHeSjVTDHEFih3PCUV5qfVt9KvIfmq8luIvSfg9hrhv1afxY8zKbAeSWhl/y
hXuXWTtndUlCb81g/Mv9QSdXMWA+BsZCtjDy+g/2FfAXjjve3AUJRZ1rMlan4K5EslMrnENBhjid
LBbUOTbpoLsGrY+zgSVMNfemjbf7RqRfOVVm/dqH7nHwty0w69oM1Gkja+UKgk05CX1Zb3pY8k1e
iv9AyK62vbrE4YOhXSF3PalZxw9ZcnGgC3pKISP9q4HyVOOH1Wl/1MEYCyNIorJR/PNhbPp50gL9
/VjwDSt/H0y2pf+ROV/S96RV/qXzZA0GtS82gVO7XcqnkeSu/3NRu0GUnS/PfyY+jf4nASQcyYOf
jz2oYg2uxPdhlPpYxdKKU56KNcpeAt5CWypHjLrAxcV89OVE2SG628iYmkPMUQsYIOQ29a9okc0Z
D5aMQ0UPDVOCfZbaanYP9ahG60fL8rEBEf4AzFCKKcl4+PYDu9YHHZzQ/iYSchKAWC01rmbxl3wn
nftsGh35u7JBji/obmOFzB74RbawmVIFU/oONbvS0cEUJILDNP6CubEuXviojgDzqa3lyDWQ+A4J
2qR+UpAPsYEIlL0qtQEa45rL1M0wrufWQI4JteywGFweem5iBSYqwVRhqfzen5G8niBARrQd7wWl
yngQr1GdMD/TJ3cXwYGgz9DPUiBZ/tTI9u/2c5u1mSfZKRJnnPjOOKIGEy8IxdeVjU8csQEnCsF4
l8b4bI7L3Yy4JKELSK7VY9fXjuy2E2iUM0zSRVtQBqGWrIk1tm5bp6FT1fnEsMkVjA5WJWvKVJPS
Lrz+D0yB8d6UnM59Bh6XLbnfHbOa/6jzYocqPyo2rhPZtKA88mkQq7srV0J0kNh9n+Pp07sWqoES
71ZyVcLQDQs2K66fqliUZxAM01PNl7kmOttEc0Sq93NraTUvRkolCZgmJuAJETfpU9shP1dWos0R
Wepy8C9QritmEnjy2uptdo3gz4oXaSIX4h9pY9k+9sVpiP+S+4kAfhbwEIsvmwvtD2ms4he8WB5Q
p2auUaYDXjgxtfj7wAwlmNqH0eBufZHx8OCgiYLX3BofAh2aBxTRVGo/LYbypHvTsTJtL6JsFr+D
n5F14epCY3cfcFWeVcPFWP9Q6VhO2poAYmjv+3YBEOJq5vM/BVbjXoJ2XtHvuZfiyayBgqewIiF9
99umAMrHYTe6hBb8eJTnHlHUmoUqXXyCwfqK3e4hj+0GBVNlZeBfBuVRDuyt7uiE7pKUx/Ev6XBn
3c3M7exNOr0S9kPo9gYP0FrtZCSPEj6J+WXCrQO024/9zZbxqNOEJTFeMLZSrfTG5/ZFjmI/rAht
qeaQMnP3hsAs25YxyBBqPCf/cW3onp1lmOZ4jkaw9TkNfV1r5hiEsp4Augz9O6NEYNBsZcUU618y
StYXqFri8hXzhcDzT66fxCeeNZqiiSY1f00jEAKGljV6GiQsdx3eqMyHsBhM5lHMz462Vq7X3aXO
UekhRfFs+10aVlrIw1io9zMpJi5SdOrqMvR6Ws6h+ro9CzY74YQpa2GvOHxF0aGBmd5kDOWqArM8
G0OhvfaemXjSyoNCJtIGBwyGLsnQGCHVTMPm+XFh/+ZJSNeAhoeT+pgI2uF869FW7PxIx+JVQ+Up
RICrSVlIL0yF7vDeqcKJx3KU3ZEeK8rKtTpJjzFwZXbDvP9LH39U3clEwHnnMTwJ0dCLbLz2XN0Q
bHlEZHc8zaVsNxJGiXwpVcULbFTKvm4tEmFDYefZw1KYj+snA54UktzA6XKQrt/FGdLI8SoG086O
8UR2Al9oBFQYMdP2zFJFR+Pycwoq1SaQ0UCd4eGgZm62cpjyDwDiFyqD6y3YhxdyCZHJyElDsLP7
Vxb3a0d1wnAYK8P337Qz+moPB4sKaicTgp/johcd6CPc6rN6EGcpoEdVSwLG3Ubdw82yoK5pa3QH
qLP8eBZ/M739aSxyyb6C36jL5XuNUVHKl6uj55tgM0V/nAxTnQH5yfwiIKGz+xU9+pzqrdbRo6zZ
++snCgvglvYxW0VLA9BUY7Gd2j8zuldgNCaHXcLsGRJrf+deZV0LkzKgjjzJ9gNrF4VgGVkft/YT
T3ac6O8btenVFV4GVy6QXxRwKiOjP96zzVFlef5r+c1F1w+SMW4OFDceBlHxA38PPAu/rtX65q9P
rv1XTS00DakG9dDhbmCLCzBwOoC//riZBVVdd4TffODdQM8wR8ZfvFsBhssUzxJCsXK4z32zBKP/
vdbahvgz4Tg5G4QnZVU4j+b8DN8z7ObaFhaG61wnMAkXZ5kLPHTC7G5wzWpPUo8dGAs9RIeblT9u
UUphPNtAn4kuSwcZonDcUybDNArn5t2LsR1KrkfvLPpqOer83LFmYASfjHVnUBKg6kNNt/+dbnlO
K16fxEhWr14fsaJ0Tw9NjLFi2IZ5QT5Hc+lsflZ/Ea+1mQwdEcUVVIAp5cCXoU59CRagM1mJze6u
8wcirTvwFZj5y4/qEw5Le6mNgiRrF9EdiClPoTwOiOdlR5sYrF1oR95Mg5J1cOJsE16YVEhQXh4a
ewaRK66Pu5QEDa6CIGRiKAdlSBWAsALCzNBqaotaWMq9oqxnquGe9xtFz4PbIf+n/Z5SuMVCLe6l
TjYDRBWNc6HvyULh4YqCutQIMTUrSUawtGF+nbCJz0xMS3gwJUn3iXeNnYM185mNeLqof+9DQ4+F
kyoiOvSo9f5FAv7g48SEcm4zcsA3WZCvFHMVwPQROJokyB7KA14ux2unJp7SnpNJKN9FQH7UpvSp
Dh6oyIIlJ002rl4La0AsRwA9cCK6Fl5n7xOKz2RLAJ885AQnfrAGyPCPmK2/E8Jck/tn4lf57xxQ
6J00M5aU4JbfKy8Jq5Wy0ZFBWibOwimd+YYO5K5km3IoW6CGnC6BUkjis2XqDxUZ33Z1kfwhkZUM
6Y8OlLcDjn0Nlxrrh1P1pJTbpH1AO6rrmVDkATH9M/DFBxn6JL2wVb8ML+Xyr46QK0/xJioNfEij
TsUgmuoTV1l0E7BCnqe4rsIC1pq0E+mamB45CagXf9vTvSy8UIq6/JiuzrgVG07kRAzjT2r0YzXG
3xzPQ4awrQ/eywo+DZdTf6F7PtUH+K0SZ0uDPviA3gRUaKSwDfX5YzBltj0X+7P5jfjRfX1pRHro
pNWtapbYjMvpqty7ZCZ7nerd0zK3r2mXbvLulWvjxdgb6+l+p5kzwtL58WsJWabpkHna3a3OU4M6
sJNlY54B/uq4Le6XjzMUhk48mz4XLbP2ic/Npcu657VG72JWt0KGMU1qVjrvmxEh60M4GTM/c6NV
eCGqp7ZxH311wnbtGrHAb5NLZ0PVe97bNfPllQtdhNhuQkGpwDkV/NbKfkVY5ToPIjHieRiWe4Tj
2EVt7ooQYgRF+QRn+fHYSSlTz+zgh95MEZro4nXUpDpc1UyU5ROKhSx1vKnHGLQgzwHk6Q7Fialj
Jvr6ZaMqftHCd4HmR37TTs9Ekpqt3Tp4mhOUKhxJeZ4+5Opxv35iIUyky5hFtWG1Gw7G1oc3+yia
VnNnjCwnKsikHv+0Td7H0lSdbX7ilUnuOTrMw4uMCX26wL3NdI4wQg4OBmeM5uJqzT70wr3hj7p5
o9kUvTu2+3zko6CccYifY73blj4V8kF9HntPBDKTvAcxA5qpPRc2RjlHxaRxjn/A/fbXBWwWRXTD
WbqucpFxeNvWVKQswBzdVyXrPw3MEFYIqkgzoZGYI72sT8SoAAntJEI86UzApRy53jXGk0ESkUTV
KjPj7OFx7HYIfDbdm4EM45efpfGusVoA7briwmnkvjnSFpf7Tlpab9YzTFdzx9XGwxohMyZHZXQI
C8FY5Y6a5RXEphWJYWfuRNTuM7PX78dXJwoq+tbBFJNJ28+R315fAp1FzsjqN1wRUSYbQIXIVaP7
OtYVMdcDBL/DkX78+PQDBuxsEktGlJznVVzelXuW3tDNGNRPVCz3bBuex7Tajz+Ibw0mKi0HA3DI
F5Ixb80ZuJcamGW36mnMX2lCCQSNNmfNqDwybZP7ZFbpJrjjpwsxqt3wMxqmW3r4gqKCqLu26nZ/
KlhJYloQLFO0qwNvdzhyWxw52QR1yI+kadbZ3SCTah3WNUYJWehvfAvBLjuiK4YeIx4KGFBsfOQQ
0okSrW9mLeDkYaYxkMcyXak1PH5cldwbDD+MUtqi6eblmKDnrcNs2P5bm5zYWRcWecMUQXyaLNXC
aLeBw+itXBqrzw3ONt43myOZkKeVttELXxqgls0KlDgzB/3ySZwB4fZ4CCjZoEj0K2rxQFS+wTz+
bwq9UjLqSGC7E/Ae4/2sn3+s+LdP8Y2suT0YKEwdokHmCDBoFklQ0uxL3mW+e790jqDftEoGzWFr
gTK/bY9NOpsBGc3nasVray4ccMsiDRkCCyiB9Fv0v9cpkpmdqEzbA1pZGzU590uqUOURncjUn9Pw
2OcU+JomT1Xk6GwMtMFT4py+PrxpvIoaOH73DAUqIcy27rozhDeS74z1Wuqqh4eMIemxyMdywLmx
WPl7k8otyZRJA67ve97EC28ZHK5NT0nY35Oz3uAQuAIUMVSNe3GBYiT6n8yyJ/3aIGuZp7CG3325
RUxDbW39bcCYJpTZwG4UcIMk664szNxGXtjpGDRwESXhxVt+tr50iY2obGwKUFzF9SLlD0v3c4Oi
yC9ebk5r8Ve+l54DJsKXy4tqi9a+YfrhYGTV9edgqpH8AavJl/flsGv1JyDzM7iiEpBZVRXQku3v
yg9ZhKvNH/oWIaO33xUFsfBsMfYdzkA2PQHt3B82HGeoR+tASlVnV7CrNYzVwZW/lviAVTJa/EAz
agvUisNEneHs6DWKwExqzfPahAprNChNYIi1UQIW+p7La97uNYvwhQbrB1BstEaq57P8LCyHuJ+c
oajI15xTGk/ndalgXIs7B5E+ngT6j/ihS39cUebOIk3cJyXVdWjJ40o+SdVtmPYOzj8PyfPMQs7q
Y/wbgTGONtirAonsd8mriFyaaEq3Qugv/Anp4igFCIHTz4AG+8gcb6v9QrRnipZoYSgw8tvdCKrb
piR/cV3JlCExnBvuGYepNhgOY1OofZ9y/XmK2z9fy3d8eezohH1MuZEXpX35PoPqsIIzhuMtSBzm
gwMnIDmIC2y81Vz3qumh+ad5VXhKgds0IbeI+aSYoSMtkSe6FtQ8lgxUFkIXB5SbaE0iSTtTeiA0
DMOt5pgw/jq+C2Cu7SD5DBvy5rRCYNrSQS3xjEaqYwAP9UY2GuzIj0WWldkstau5qwpdJTOsv/nO
JgwRqbWD1Ae7WRbSEpfGSujbXiofrRujq1eGhx6QaMhl+h6N+U7LCEh2Hcue+Xc+btFUVpKVIh8q
W3HmcLQH04FDILPZTEpazP3wJYYAe9Xj9s4rn9qnYZ2PThvpJXmc5OTiVz0c0TczevzXxHXMkNYZ
rqwy7fyypzgCRjJJqj5Ookq8Zg9smfEgn6MRcUwFx4WvgHdTAhtfsplsGXjmQhztNkG9PEw3M5EC
kTg0B2Plj13V7DTbYsm+iolZHIXx1NQlFhLBqhm8FokUb7evBQv11tLsjev8wa7sv7KSSeVrZUEq
onGh06OeSrJjXWpfnNx8vlTxRg2f4uVE7d1zH+rCNpd/HSvfe9rRzP8j1G6rWWP+dZ1IVI56EpcP
uAMRu+/Z0CHIuh0AlWOS4CnqwoyoQbM6jc02SyVoIarR4mUOLiMx5RAzWzyWyn07N1SKhXDpd2Ua
SyERkvr/nLZLfcd+EqAASw7fs+rVtvT/OilnAfhjPm+O4aBfcHsIzUCdpvlVRkSTH7Y/7JgqIdkN
V4J1ucec+mwQ6QR5eOUCp5M9+EcHFr3NK6IkzUiEIX8i/dlrOshJnqLoUwBHaEBYXjLtP2gha9p5
miSzHhcJKrLCUVsgIia0U2/zHufeY86ASxhfh9YP+hcIEpPZnOYCKCGSeChkLOt9bXQZkMbEB1LK
N2os84C8Dc9lAfhPAuD07plQAwj3xC3qh/2nRGeX6APlMRtPl4wjrx5Dqt25jNMvGMwB+5Hqd79G
FuRkRtJPCUvwzI4EmqWMlmtpljeJEMbd1g5HuCHTDuv98hszVt68o1w75NOAoORSErJy3K47Fm06
m7ewwMeSvq7Rjh3qOcHucD33vBTeWFer6kph0gArJVnYoKglh+AhEq4eHb6+evpiQq1I7XMelmZq
Maer8TFI6B7bLP5C+pbnyfUk3U5Bp3U1BZpFusxZP+lidVzNtkQd9esqSsTnvUzlzqhV4Om9PZ3T
d0uSHZXL1Zko0coPwMMqa7/KGLCZIJDiRE8bw/Y03yOud7tskDejcTaIuTvX+/6ppIvlQvNjgLkL
35U3zgDiNJPGD4+RLaBzyoRLUngIpf9oF8Vsjj3SRTleR7wonY/7JL7cUNd/yIr3MPFynXEtHY59
q29E0eyeFog8YCkBUoZX8LzyuaBlOJ/ir612FiY0/QZrXrMSGDC5xj9zHN5jQk5/JOHDYgc0Zmf7
iUsyYN8bsYogsbNgRp6o6tE+aTBe0AGybAfFawjzWnCYQEnAkhSAaHixoSOFr+uitbVqgkmAQJHq
0rHfowhEtIVu/BFPJ+/v889mw6Qfp+TXsvDlAFkSiO5nbOMKuGUlW4MwoS1+p/n+H72Eno5QWakM
1cAYktdJHoPBO1F4rimyawtBaVVpjH4LO8ex0gw6x9hI4S/4uJaLIaZI6mSBKigO2t56WVNXj2QZ
+BobkupGZkKVnmbX5yniUO7AFVEX3w4NduDDPpiLEowkV9PHF3CaMac+J3rgWsDKLMi25kDBBc3n
8kSjejClLVxQifdAWhyA47YbJSXXKLS+UkUo/9VFrOcEyw2Gj4WwvTi4nK/cKLEPk06aouKD+J3r
EYbR+rUET1gE2ZvItEBZX6MIiDMziAYuZTuE7Az/Yn22bnKw707JjQHtH1z8bZ4KW8Afp+JSnxw5
IXYwwzQwVahFw906rN/i8MyBr+64yvo9XL7pCsrU/bbJQDAcuyonO0dxO4oLeKR8PDwaDngocceu
Q1dW2BZwkcm2PUHoCQJ/lvWdEa9mHjJyjm2H8JBussNwgtpQgtsOK96zJ4wQiX2CLbkTf0vg7P9P
hiIQEuZ4p43zm6Uc209n0i+8YoXKPsgSiYvdSuByybZMe12UfrHFhRUQB7nVPXuXVjzv6eMFMQN6
5y+DmGVyamgDBWbzNjnj/Cbn7fGQyeeyvgMlUNTYpyvcpN8dTnsA7zk2su1BjKjnCdoKeYsou1cV
e5DzzeqiuEmXVEsS+9Vuz7mqxvoU9uuANa7D5FchHOEPAbczm3sWi0z3HDJ/d4yGVHG0iBF9/b+q
DTUCAhuvSyGSSoC8molxNmoq2Ed208blUM1LGixiGGVEMQ/68laUGgCtX14yBGleqsYX+YIl2cSx
x7LAtul0Dv9HfgxT0MB2DQ5s4Zi1vvJ/R4gTXPj+ofJfJlJmNga6GODQeS60PnqpM/YGKqjKM0KJ
+DXpF9waGd8oicI9SNEwAttmHTEZP+CK/B0ONq7lfS8R7/rrQqDlrpaDqNVGoWk/zuaJt7hpupur
iKuKcN/nzaDgjkeDGrV2BRmmQ2aIJOaFMS6zWjr6R4KTbZ04OLHO2dnETowQ3USx5fE/2vfWJuXY
65TVHGAnv4PSpursQ6owqUBrUfCQzUXCWoh07aHhoUn+Ga5V6Pot8iojG1VH8kZ3LtQZon2bhRHW
PkRLR8cIAWAJSEw8uOsnrJzvy6wok5DPsRpih/YHQ+tWUP6YeSHjErNEJZMBMKOuU1tli8V18Vyh
A2ULFC1inlQG7N9s34Iizu7md+7Vt+J1StGsxdw8x+WzuCjB/RPCduzAl5hqf7hk1luOkFKYVRlt
6OcSG73a///9bcLemEJ8avRnN1ULgVQ9HMqBVvWvqohwErE8hn83u7rMaUW8H3w/93qFUCt6e6fc
REBzlWu5t2Ns5hI/X7DLct68mydBwy///29VBcxzSBCdLfTcXb9omQcPLWPhivUjMHI5dEZYHpjW
oxs0Xji2HjGDLG9mP3+aq1Z+IA/ko9ArnXG9/9g/YBoY7PI3ltK/Dac78rpkXI/CguMjlHeTjygK
mstlAsBsI8Nkm24jaGkoGOFD2ZpNFGgfmZPAEqlulh5rk62gM3KKECca7laB6tON5lZVNLmidlja
vt3glGRDC8q2dJjB36rnTwuor2MT7Ry6WZO+QodOG79mkrimIqySlxax2Aw0z2Wp961zJ1Nrvjcw
qqD/NEXoTwffBA0d2hFtxmR3nYwQfRsAWSxPUCaVb6ECFLTuRFmzgNuxPh2IhI0TvrsDodsbLuJW
HYx0TityBqahfw5pAaDfu0r4cLtuJor18UxAoTzfsWo0yjaSuC8i1pZol+AH4n0PnoJPDxEhwOYl
AIzSez5DntYxTveY8FK8n6DSRFDCWcr+DNXukP38xb6uHBKzwG0dVOLVqTJTZV3rJxSe2meRn2IE
NAm4gAw/9tRVGf8dwbfgS83AsGHkEoaobtLxCkObloIlnZmUkImBsxg3XjofVPip3n/vgZ1AOHlb
kraY9AeEo1phYlm7Hha8JpxYUHuaHxT/YRn4lSERI/GoEpT8NgqgNc3uZlYIXDvQymbgcVq0yKmm
jZcSIe5ZpjFSKPG3qRlouM13UiuenVTM2Iu7tA2b2eDRIU9VcIvoq0HjwPBsr3Pfdwq6m9jPGtx5
E8RaHPWcP8xJRQC6z9vJzblK86ZjZB17UjXqgmQJOH1ScJarCQvajUgDaSDv66783iYoOAdezbho
lm/gB0XM27LkxELAsJtoq8DBbVyUC7lZGwzswUww5oHeLb3uYKprcu2mbjBO366FOFTwbBpKbpHI
QZDTW0Fc0dUG89LLqz0SQnA/LBiaj1G+vo4kPb/5hJ8gH8k8JSi+m6bbhD1fBet3/5ehUgIIqZUi
BP5VUA8Ts/4uk70DLMONMnbmiovL9Z1N9jkrrmcauJveulJ9XLYHqz/HTzIOn0g52sLTV6wGaYix
8nGBAIcEgFGCLfyOmCmw/QL2Ev4bPuUjXWGDmLfhNAHKd16Rwb7L16zHC8yd8wmwvfgT7bwLmkzT
B7ArvgqQy/9mQIlSRLCbHr2mTjCYdoTmJR5c4I0WZT25im1LS5+LjdKzF0Y3tx1QNX6WwP1470pd
JwvSYWWBTpkN0qN9pUbRfjoGaaAC4RhBi5AjzkrzB2GECXxd4Dny0xFKpS5LjDGPZg7s4e8vLsW9
Lb/QIImFYCMUFxSXKVubtTlM+TU84hCCWGzjrXLpag1k8uTgkBKapei7Xt4/Um6/UciazB+hATjs
tupAZzYJ9sal7ydHbLJpHePitKVOkyo06uMyl7v/aDP7IlLpe26spI7V0yzJizIu3pBgC2cJWZkK
2/iXMITEtA4Dg1DPrv2bMOCTR2iEIlk8KL4Y0lF1OtB5hxDUlCCBsTwTBerW6G/r9kS2p24v+111
B+6QoqKDfbT1tIpKLBvwdDozTMRXjKldeGz8BnXo2LsQP28PI362d3WighQZsXuAh4r/JAl3bFb+
H46kgqgHA47FEr1S019LrcsC9heyVLqGxA0fXwIkdvYK4C8kSZ26m502wyhlQ8iumX21xhhmJ3ot
sOz08cc6yoO0OpeGEa9eUglsYHLwDJG1S054IpgmOql4xblNoqbix4hptDFnP+GZdIwgJazxoRXg
X2HS5P32GNbRXhIqKWjo8Ny8zWU/kkpPBXqOuxm9eZOUn6GtHirARcZkic9wO9ufQ19TfqT5UgQC
PGIx3+LQ1HYZGt8NkhgKcLMm5VI4gCcmLzcBFmdfU6LVps5Ba2YOizuiC/osiv8JzBfwH68qdjXS
zQ7+tBP8MsIUGRMhYq9h24oXkszQy1xkOIB29tvYImbBUj6Yyf2fxIfidRGAKZ0zdueUQYytOlu3
qNgMpfSYVa8JNZxQqvvGrjQlKYR1wS4mX6ohdmtGDU8GE/08Qxfb3o0Wf7+KfdFVDrwjH4OIPRyc
GjjOR/KAs6Bsdi9q3JKvTQRKpCtBwgbW3l3Ld8la2vhb03jdCDIqfK0UnOCv2MnxD7ExkmpncQYb
cjzKv4PSIAPv2V2J1vq6UECFEwXlduSb6/WhchpO4oujajkx6O+e4IzqoApf5pYcp9ArN3zXj0/s
7QogqCvm3jYkhlUgTXoECZW1VSzMMF+AKt4Mq20SAWdIpf1wPWXT3cB3RyjBkPi0wwzjFuCrygyY
obRoNHOyARJ5Hw6D9Xg6NuOqiBCj3ZVM8QdNBxVsfyuDAWsTyCMmGUnQgQYrEUhVMIliht69rQ+m
kxN9l/W/vTOgLf/7YbY1rLQclRthmA7vp/W3o6fXMLO57ZzfBGWOzdHO76yfSeN87LIAZNOS3htr
aJzm0hWMhPa3nBg5NLVY4pRcAczdh//92d44w1bsjsWcsha3bXnfGuWwiNmTpIcmB3n0NI08t2bX
gufK9AwdtPLN5JqkExjIbipgGVYpokJVZ+g0glVQnNJAS9ODmuQZGgFnKdCJkEc4E2aKdo54rstZ
bcY8k5UAYOXpcF0G6PPUxrh8z7ugM460/OT/zvbP/VwQ7sYkxMKqt08hgtq2RXXxUtPLfY0bOqzO
KqvHJFZtclrrMt5lHcGUvBLl1IHFN+sR/h9FDGAghuZgPBZyNyoMxcu0B73MlVGz9TDdVzz4DAh3
2NXc2ojhUCxxQ5CyQCAaB3eaFRl53BxrosWQUu42YwfqQkFBYY3L8fgCo5tEOkTmZk4SX3bQq97e
2eumCT6sFW/av2cd6KPRuWYnS23GD18s2FhkZ5vC/EBFUsgH+b2Wg1Vx/qa9moPUHdelBpSlKRHD
WGmxz2/ovAqch0iG72I9bfiJU3xQfhxXYCKDYH56T4/YEo2X84lniv6/wbL98v4muYKX6cJzKsyi
orvCQEWjy8GfayxOxQcvNfT7NK3N1TNsD1c6vdNDoBkIg2d15OFg1NW3oliy0YmvVCtU3kaItD3m
fb/5h5uhPL3+HYwp4a0jn8snQk9XnKqZAU05SMQXyD+KFRp7IVrEgOCTBXaDHm/OezuaY6Gf0lKF
klhl+B6D21nN5eY/Ls3m26rXGTrwO+6idE+Zt2TsOdaFTh7JjfgmgY0h2WwRfo7SHlbBpPIXgjFn
6ULP4uCUX4eiBQr23MB7xavfiiMa91QAnZSv0Qo9zdEns8GbVpISKoRqWYvL6RBhof3cuP1NDHAg
v/b4GCrJfbZRisBUx95Jg/wfhM1xfXy/mQgNUVuvbjYEku7hznizhnQRGAmHbjNIpl/Y9DlrW2Cq
bpiRirknErg2oFGPpBRlp2kS9Ig0VNNLl7Vurn4r5F2a9bbzMofDi0RggW8FxGdaekvt62WrBc9H
DATwMKQkmjnSypmcYizHCdWzy0Fjvl0YSEQtskYBECM/6nsox3OBdoV0K9F/U1fYKnQoqde1zGWl
oHV04ox3eHb2h7W63RYjknx04733+tfr3y/Nno492Z/hWymoNlPEBtM5paIF1QfdRLRMeyUt+T8z
88oHFYvvuqT0ZSdYK9o7RBep/JD0m0ry8+aXl60IsYOmeilGFa+x1xYicImcMjJgmfzsBySVPOZK
zRD9nwBKAimDiPEvisI9Oq+naRx4+CUKCblm9+RXmkbBZN/lUy3P7FFnlXQa5tStckl77qBpDUmH
Es1w+woPVI4n1UqzGlM8GgeyFhwqKVIBg8FaG1SjPKaVc3yjfDMZyGcjKCd3J6uXN0KoDt8g/7Rn
syn4AT+7o3eDQo0N2YINjBAR970yFAzcF977OcmXlJF7FOjI2d8TTQULoxvBe+Mf2weObMJRB2UK
sOCI0tKdDsQ982jAsSpS62ZOlL6kYJZaLL0+Q2TPkr2kU7HJT/9czKtP2VNMRyntS7v0urRKaCS5
9MXO3OjpZo6ddqF96Jk3YxFsyrWoKi1Ayz4fGvODUOYESY3Eiv8nrwo56UHfHWgSuzDJdCPMM67S
ga66qZ5t31FBhwSw8ZE7zCvIrrQFAe2suIQ3qpqbKzQv/ORErk9Mji7fE+P1f4GjFpCgIeyxJ8kw
K0LJZVb0J8IaZqPen5BJkO1qbaZVM33vZ027AiQcmnwcM7v2Xkst5H6iIthSOVH1umvX6hhhyWk5
EUiZDV6xPdFN50raGrS+EcjLg4n8nz51nn5c2tXTJkpmZ6AnAr4OVZqKB5EUSRMOsEZX3bZkA82A
5UmZGFMlwzLgDppaUOvI4lV2xmxDvkagO6GhF7GYRIHWiYURX0gv5UowULMHPwWgz2PDsrunCpSo
CDXM910R4sV2WhSHzPMWNvQZh8S/C71e+zfkYmOl0s5gjaDEzPzUvA/LGEqhdQ4N+Fn+pnZSSlKl
NYUySYLfLarjBUKhoiD5tzM+yblr6gvrG85wpGaY5RT3KSiQ1PvS311qGZlNGEx/SGuJsqjKgJN9
ZjQjOekVKbkJJUlwAtEGGgh8iYGOlLf8GbNNGl5Axa7qPyS1VHMGslfvMNS/LXjNacL/GTTT3cB9
epXtUlbqNVaEBEDs30yix/nx3Z8sel7oNr+D3eVrc3qWo0s9UVjjS/nsphbP+su7HpW2kC2PBWfa
arTxQhKs9JMkOn/7XMWhxJnR4aEwTTTVEd44aR2oLujG3Z8Z69XfhyEeBcMFwbrhEwRquy5c2/qo
fZ3RDkEgAYq8rwyspXPcul4Ttetpy0xlHjlwU2lUi2hhDs+UQXWFsGTZ6OatfH6x8zW/d6WXWL0P
z32g0n75vYJ2XSoLNOE5D/pqQbhECvLC+txOzjoHVVnkekfjvEac2SzUU3RmW87XoPmRJbawFbv5
mi1OzqUcowzJPbHCRowC56U4l7+zScVlFhRNGoupGH3oeosclkNYhDWUrxSj6ZSGix4r5ARSxrYi
RnVOWU+YBNtuXEYFipXJMJ76j7sgwurVsad35sMX3pISN0Ats7TGafNObC8Gf8Z0+TblSQyXldt4
SAGEItrn7KIx+zKDmSMF8zkX2G562mp9xBlOwTjNU8qAJ/S2WEkKl2fzS/Qdf9/LRTO9EqFtnww5
cBBPjuACtD7HwiG7pHsas14MfeBzqT+20zX0oW1cjNazw1ow9gsBeZRgyA+SYGO9XUpn26ogJW+x
TAg0/o8qQ9mF8oGs64HPngKyvCl/qbwC8byePAZ12BlSV6W+9PvRldAR2qtGNALbGu81Ix/d1i2E
TLfmJ91K//l8cjGn22SJ3S2qh0yv4OaHjYU1wQ4kSXaw4khf6mOWRUNzEnXJH17m6RF21KR3z5W9
FZ3YLZVGB3m4WeAIw7W5J8JS6CZUBap/bB6pbBuZngt49x08B6OQAgxSaEhQd3vDC0o3X+aY1+yW
PO5a50DW8fKEcpwbzAUuOB4vv3PUFYFFZhQeN0CpYSyyjt0yw0lvAu2V0hkr6xkukCx902EiU9Xh
XrVs57adypXJRqLDeQdeos6h2Fi3NVT1R32v+bWJ+n0IxFpiD4U1FfYnShW24jRqPISbKrf8MGQ/
tR5RkXc7bW7idKxzSr/hcb3RCONOKmUKxIPKEht8MHupGru0r+7xkpeX840CIeQQJJ/r7g64g+yD
OIKLjFczaN/qD2eejYvCC+wBU5X2uv6fxFck9tV2n+29Be3L/pIF0Ml/C7d3H3wfW+rptsqIxAYy
P0AMr5kyoTKWn7x9yMavsqIjBFEizLZqKgOCqWTotSGEQYTKK1mrOGsws9mY3WzpKkgH/qz6x32i
w8AMXellK75mybiTC81RmSIGqXVx12VFsOI9m6t05kHybLrGbMosHx0bpw0P385O73GfFJb+juG+
JmQJvXuHg4CgPgqfGh2/8G+hQljna3cZTRu8eJ6D7oNarSl0oawXu096kxN9Sw9szHO/ebnbNTIu
QgMLxfzUzLrLwiCt0z+ibNqPPVPtdD/dHlLNQcq3LCkJyit5nTra3A6iuG0wWfAawJngk6y01mN5
4svDaI7o3tEWU74fCoG8p5Ed3PdDgLEQ2yAHKYIVJvFn2hpALhUjX6muCp+nOLvifDwpGY4e515I
wvU0sUA13jY/cli2jGVikYtfoKks5a4APo1HXJCVsqHJTX7/DCbcJ0fvJFvW3j01lEevzITsr88v
3FIA0g72ggTCmJGZjitF4W1nLoLzs9onvwMRfkP5HyqwmS/enztg+fNRf0noy/al1nCx4cjl+Q/c
73dk2OMSbK4ksiPGVoYV8HZUfM3JirNFgqbqILX++Hf23IjJsnwIJidjZeTUTaVPkV7hXfo4Xon0
0wSwoZ58VoUEKyzhLEAE+vFYUyUIql0fv3tXMCD/kL7y0UKQyKq2pze0QKHt9GmekFca/i6YzU5+
pkkaotISFkd5tG0USwzsprrdmhV4HoggOESMjVLvWTH2ZBq3BeckxjD0/mcA2zAude/ezwNbDtRE
ktj+cU4MQohNOEhx3G3TNXL4Y2ynqpxm5LxQb2jFYj3K2yNmSg1X6NTO2TomBo+b5f07XjdwAhTV
rt9kGt3RIDEpgui4NQdGMn3heTXLtNU5xvJvbG6pp+/+pJGsb2r0dWj0hNzEscNKy6+KVL9NLsJQ
uVoKZNdqjjRU+TPwcNG5VT90DPh+FA9YJrLC0ok4UQZvx3kjZW3Tf4th5ZzSZgKWDI/1HWkQ8MHi
scWDdTlreRvSkTmbom+KC7GFx6C07g6q+bhsaqwnA5I1dGL47cnzMRNPi6x/Zvx3ESKH5a3/Q2aQ
iWlhCJ0elRZReWUrl4UZqDNZaKbjr0q0c+ao7Qwg44xpaz29dz3Wtx2t1kwOZbK5rGwOcgmgmnyp
rTBFEg8IOYNYsD3+clwFrPps90L7k/TDQxmDjYdcHzKD7As1qAWjHE33pZglwOuANrfS7b7ZLFQL
7qnLcSzx3wCMxvpevVdr3GHootg5R+4gNgQFXYmaxT1vhvfRDmI6vaWyDypjWyUmhlNbrG9ydZIo
171Wooz3lfYeybX1GSsuYA6kfW4hIwkx8FRDAcZAOpq68MwPyjSmoyqQCrk8QuYb+/be5rHju4B2
v11gQXHladK8+LZ4Vhz/fkgnQVs5p+ZMPrpjwN8/Cm3fWWZiTmH0xvU79ob2CWXxUiB5wxTdbb0o
r84+TvlXgvjNee8S2My/FGRBVnqc6/vzjetlroC0C3U1+qK4LwoK+GDdWyJSzz+YSj2X+MVy3tv5
10FmWPOYOEJqlGNCND8Q0Jeg4Itfd527AGUPQlqnBzr+EjQcjSZw9tQp2U1HPO0q74ky+oj3pKen
3iaAL7vRAvi45NAEalZWWdYAtYkUHcanbaJRrBtB3W+P2HCL+89h6ZIK4eRbb96e/37UgQzCng+F
op6vHeeNtjCLuvAWsTyBLQb5vAfmox55tOpDYDyBvp0MtsWZ8hYmcP6CKaUb3+Rk0kv6KRp4Kxrr
tsho/IksQdE74sfLYTlTPb0R/ZEs+G2K0xpX9yGO7ZGFoaJIzTcaqBsh30xmfj1geGZhKPv0Tsee
5xk2vjzXT7woglrEqOOboS+KPWfWaGPmQ1eqXjDtDg3PEYMnlIscvvoOm6E38SMHtfi0Tl8ku03y
fcb1wPN9d+1iurDIXeI+UTpY3cDibq0wtVA+67QnUO8CDGGk5mmjcaV8KnaadWCrbdIMVOQvFZDP
qrv805sO81c8Z0Bo1aVNBj4+lpdnJZSP+5vAKU+F/gl/9SixF9NjJ3MGS1oM2Oqf7m/kXOVkJ/ud
K6KXX+AmqyO6oyUANO7wSatHrCNTJdHL64u4gd7px1shNKVHaYhrzcMR4POltMLAH3fhrv7vOC5C
96JbOJ8/LQbH9Ykx/2KgmluCcIg4emTn7nYk7l8Vgj5OY8TnZEsx4sf2TMQsqtWBP/KTiiVBsr5Z
kUf7muciVCqgXSLbOCTSkJnYLA4JH40UPaOZgRzBppZqxgWmgnj0W5wVn4YW6b8YLppHftNIJZn6
T66tuRBBCphIgu1od6blcyEcnlggLlgZb4aX4xye0RzujJ4YiaMi9ZlmZni6XHMn2FVFCbu2yIbJ
nSA2WI6LpHHY8QM0HvxAghb8+W8/Qd2HFVHm6fmp434xHi2OUi7OPp+pYnevoJfTUNl1n9BUJn/p
vrPLWXhZsl1xKfAuxuBZ5xSS0L1eY7nVl8/w/XJDPAb8sd/PGpmiTQq5W465LvwjeuNKmAMN4z33
/vU+tShoqlPm4xysN0zoV9wv8OMb5WEHX69mmGy3+M023uB0XWzoNKxK2DMvj5bqR5k4WwteXz5Q
3AYGhCbG9JS5j1PUU+CdOuA3wirxwJMbAsFmy2dEvKtxfBx9qobRfam9Ete8geRKvAitpf7l+zxE
em0hpbwLYQGVRGKZU8g6+gHFbJIbZWBodUgHQdM/TKIRMxIopErNYwegPnqnxMAbgMHq/OQmbhtv
GVqLEOPaRnOvH+5rObJLJyCHTWmDMCy8QFFm0oldngAcemv1HtSVK1ow52kyccvgpNVB0MGS/LUD
lKy4lFUUCSo56hqv57TAsJcHEMOjcfIv07dJ8lVa3cHr4J8QVkOm36u7dwHia+Uy4M7aenbRBWZn
7zHAKEsrYIZrTH9nPdfYh2aV28R4/kJLXfb6VLoBcj4ZWtYC2t9TIZNM7YiCyTijcqhQUCb4PflW
RsEFqSuUxx3vD84xhJwH36RFHwu+ebnWKXdghwISrxgaKv06mvn0LVa3mUagkfxcmDpDY78tUg+z
7dsVvRYDp5uVe1jOhe1fEQSQNRqJ9wQxWTms+ksO4edMDLcYcaP6Dpz/PoOwco6btwO+cknJ0XSP
WJX7bZDo9MnPQIP3oIruCWFalSx4JLEucRCT+b9NCTusaziMOOKfntiKfzbD9YK2YKAcOmO9H3it
DQJUbuMcJNB+Yg1FzvmfSFIQdz/L20jC8C864AGjzPlKoqqp4Kv1B52xucTrdfAcYGD1TvHXNKYi
nUUmlT9omWeIapdvvNcTyWqZAoJ8QVrwR6Dps3aRM0jHMfeQrYHQjnnMO/giNLNJt5qU+oEhQtcM
ZtKEyj2uxjuu+zwBQcmBhD8eBfo1yS6N9pkazIN6BDWYR61UMzBjMvfy26zCXksnIoiFe/hghT7N
yNE3IAPup91TbN4L9C1uQc5oucigoPDVBY4sZI+igYB18MN8+YcetCmPda8gFsiE9ooRqm9aI4dZ
LrYbVsqtQSyT9C/0Ky+5G2Yp8E4TAh5roUuFyIuosQorOgIYWTQPm7/QqKxY02r00Zgn+XVetBBQ
gqVHmnYgQaRQDsMVqxuQs/OBQa7D12mjENg+n4BXq0As939hAbLzH16XsrTUEIBTV7UjrncEZfFe
4o3ctrYtOR+H8HWtLsddk4PUIUg+m/tOWVHC+IWBPAOYPq16rDwp6qjeUC3xk9wycjhDUBojXEoZ
adutXq+g/LzVMUcOMjvh88OZfH/G/Xb477gJ0wcqdamz3UBWd7ZD/dCUJljoVgrhdvdZEVy/HEQa
lHjGRVxlvqJRB9va8yN7a6bKym8KiphPR/7TWKrqztcf4hv2o5MoCVOigBGsir/xQ055fr/tXGlo
M0+JkBhMcMJD+OgJmfA4XYwMWe9qF1AKKK8IwIwDdNxVlmQnJMPAnRLlnBKwmA8EqAJkjH3b+hrM
iKT2aBmb4OS3elZPauOlzH3mZp+qXu7643+3tBr/ChOKAhbaenU9YLNRHFJDbGesAUcW7s68sx/e
/+t2S7PL38XNCqPHhFe5XHpQTCVMF64w5lNKrTUdJ0FIV5AoK1L8z5FxaQT4jWG6OPeWPTUZLq7g
y4kMiAs2uJOiGuXuHR9/mlZsexslo3A/v9r3OqevZgKr9jlotscDto+bx1mnsw41/Crtr83tVhKH
IPUHEOe/ScVNn6Kdgj+w+e64KDcDfQ698aF8l8W4vEamSQ4lm8N3J8+OBULh551XsVeXUWno6fV2
AvS9JjGI8Kbksd1cFY+HBOzw0ae9nAuUnkuQvq+d8fuI64L6iUvZ2mnx8tln1Ytd+UsDkMgPhlpK
Q/pqpIUQyN3E3MfKXzheMkL7YwZpkV7TFpUL2rMydCDtddrGTOFtm+33heKT5YFKoGrSQgKy8f4K
fhg0TnWP2NHC8G51hJ3vz8UtRzsC4qmXNpeXJcB80zsmz/UEQJMsCNJTE4H5X/0A0TogrCMrYJ28
bZtSX/rUBh3e8Lva/0k4G/1U3YxArfnQXYK2YGD4B/3BctfRJd7QeKWMYoDDboJ9ECahuV8L2jms
yNuQ5//bfPwygp44sJEqJ+we+xv6RHkmBvhfgUqsPde+yxnEu52Tugx1c7O19mcdHTMham8rpEzG
85ZQPGo5KmeS3Xobtnv/dNgWPJFW4UG6eucKxXWXvM5PmXVaPMW7QSQ3igiZouA2QnKkR5K8NBuW
YaENeSz7E5iVetl/0CvySb2NjvO7ZO5QJ+Vpq6ClvGRufvOlU7mJCpP4enlBt2UK5LlrXMWaHVU2
foPJ0bVcVg1CD/AApscQIJ3KSO1xj4Qt7V0feeYW95pL+fdPrr2ZVeYBbqU59FGGTf39F0XJooN5
kyC7XZ2ehwDvVB+GOHuWOtE6EThQ82NBRNoueCAcl+IqQY6kEq/W36n9UVj34KRgzt6D+6xpIsUJ
1KHl89M39vw9ZmsqC0V8604bOnJYwL0f7kHsOMNRHWyalp9F8KuIXUBB7CFG2nQ4AeRg7z2ojqqi
3yxajAzaQvlisvfp04Oylm53supIGlhddWn9krj/ozS6GswXc/lWwQvbwJrRoPdo+AQoAytiyhCl
oHHlrjMVeD+WKB0K7PnA3OrzXk7Y/eGHh9vE2fan/oHems93rRbjkzEC6iozJtbY8sBLnWLjBvEY
Q5GydRebIJfDGcfWjG/eYdU6AemsgrrtlPXqsMYLt/Q0Yt0nW4y9KDvEKLJqcdbFdZGNJ+XZZkFD
WngqJwtzECrY3MXz1GzvRJeYcm3/opsdRkAjwC1ICQ0ajGZy8oRll3Enfmy0Qoi5BGLJAWzK1It3
RutCW34FGW6hZdXDEOfSkZ4z6mrTQDdg2K5fQGoNMBydq3E4snExHeWLAAQBE4sYbY04s+sKiqua
rdtdcfwO5cVD8mU18W1Zt7W3yulYl/gko+wUU2gqbFw8+eacdNssw3s6gG5EneROtPy7jDGrOTGT
3zk9Ss6aJApzudvoA1ioM9tTa/9egB+uNyBI9xQtVXbuAXiqU4d94e3L3jZtpPG3/Ku9Erp3nskZ
CDkgayDMCHSDhytIR421FMhDLIYIr16vY5SbZRHuVbgPonkBMDGKk1c64meQiv79WFJ9OGuwY0vd
l81Dvx9CTx/i3yIDylgiNN+uBjkHxemLCpln+H8BN2rMV1cnYD8QyrrOWWRLMvlg92zy9fyTXOn4
HNxmco8Wm5mqzKV7FJOx5DCkIdLlqPnsJVqHrLdM6H/c6FusvtK5mLmTil6plYNkLN8IcRC7rWdK
VwoomQ+ZOviCQavpFoeu1SpZ2LwJ9aTFsEZek3Zb654V5rKpY95Y9v5Qcfmcw6f5AunftE/NcIZi
Lfeg2598lUSXzGguaUT7tHmWsZvzlB3uCAQRi7ugSISc6jWXIwSmP9FlYVfJdq3xj32Qulgy+P18
pnpphKvDMz/KtxEpElBkUdioZcj0/NsMc29ikSKxzrMzeY50QKUlCKKS9hmoRccNhwH0c/a7U4Nd
hmwEshkpzG2M07VZJGWOhAd4gZvo6vOtkulIc05q+WyYRHE64++qpjox8IJSTbf/aZMYbkuInP/T
sMqjmuKNpVs7KZ7EDjCeL5tQqi2EOXXkrVvVvTicQ7734jdfwxlIspIDoA762A5kIcGoEwlyb28N
SwlvCqkSGN9U1RhkyS/SQiy9B92GuHINe+dvGBVBwTYDSGM+4QJJAkypSQmFQmdr3fl7syPujGRs
dJFYM1Skq54grEyhWU37qT+1xczwklAQtoA6EIHG//+DyZV3mOLmhG3RVE9uSJayx+GAs5I+q/mV
Y5abg8NK341/t7sC089SgOS6QtJxpTfonKhsm2eT4uSn8ph/zWaqAuWoS6bDN2wnQ+ewPCo+6QJe
vFxYHgQFSffGHdpG90Z/xhYwNcJ7iP6yOdsQo2wACBv9sfb9bONNKkaEYVASdVqATIRIyDZP89EU
IAVTXwDC6NfRMLamPGc/bLymoxiR6+yr2u9u+J/7Jdarp77EEyu81lZp9+fWzGFc0RIfKWN3PxwY
V6/mrGZ5sO2bI+umncWLZSWyAoMBbVXak6oIDoFlm9xfJReIlkJ9Qha/Ve4zmiS/graZ8UJy0NN1
6o7aE7zdvuPKwtcb5RsR6omdh1/z/K2cgchtGCQuqA+EJtm/YA7ZQYNynZZjsHugBMU7gZa9aXOz
NunUuRdvv3c6zEbt2DP+kEnmKGlQ4+2mLFtrFT06KUiuGAvmU/MCg32hyObmgO/b2vy80QFyrY/I
7TefivPV5hmI1S5omJTQQww6Uy5zREuJ6vesumsnb5iR4Y7K5KpmGIoS4cI5pDDETuNY1p3yMicu
7q5UxfGi/6K4f277QXgpr5krrSVUMCAIselQiTlYeDhtSEraLV9Lhub+HP9igWUKCgmlvwhJbpsA
DbbBrNYu5Vytsa0qGCnkHJrTwlKs/w7OynnbyOSWHQe/mFpvRVaXxsCutYmABIu2Hm8R3VHitAtA
RSKSA/O/ihqIqd2xBPZ/hoCmix19Fx4h37+7CqUmsAZkqud0je9f3GoWhM9ezye6EuKS5ttMcy3M
7PT/JVkSqu0J6YlGs33GVabjRmau91DuPQroafSi6qGRQuHxMIeSyITk3re/ceACZr8JhRTwTH3F
+MdrrjpZOS3FWSqQoN8qI0u2t6/ayHxNNNtkHRCU8FMLtZFQ3R92Dtd0biPCAJjZe/r+vB0OjSDd
dBhGO4jlroK0/cVDZwXGGoP68rp9Q1PjEJlMtJ24STNEs4kZA4dcw+UDyRN6SnfBAB17hI7Fh9HR
5lbSYsZlm6dQXoSzbFCtKv4Pb1ojiGJt38I6wMO7HaevBymrEV+Gy0Mt9HQ9cRa+85KEe2F346Bl
+49fvXzf12+SKY//5Vm99Q7PPidJOoBz0Wa4WjVtXq7rUyfa0+lrSdPUrgaHlajJfRJatxyHmLau
6b2fOTdPCWelNtV2OFdj6NvRRd1lhruXU0sPGbp31G5ttGl+PK8v5Li9nmPb373T6X6cBb3m4Obj
BBqBuzwny4yjhJD8i/tpP32xC3pYnYCERfppb3clTAJsNrMi2jdVp6pId4PPbliWrxPoNN1Uj3Bn
aa8vPxr29elSA8xYWtEZmLMO1cuZIc2fq8RqN3KNbhmRV9GFSESd9oYHUoC1vkXfgKs9yqSaFckx
SZza3GDTHeNuFLbELdYUXE/RzxHr8mPDsad9g9fQ8fcFcq+02Sf4HUP1Ac8pVMMT08alIgxiqtvH
PrrzHEDQGScdk2/wIcDt5Esc4V3+3MnDCcJ9ikhT93Ii3vWTlGAbwsnOAxPzv9U1zsweWIKD0hOD
hGNmx+7xGE5LvcpgyZ2bjuc+J0j4GNXSZrltyF33JjsXAkA6hiYqEuUl9dTogMAzWqzMXO+pCgS4
FApT6BVwzNyXiiWQRWcZu2XqPRa1avs8gbo4gLL1EiVxLf7K5MdHm9jx16o/jnxg+sNN4JYL3ryF
YjgubySfTFqvVl1gpcPShg1a1sQHSTQdGqSYSoALyP4OEDF4/28CrisSW3ayrQe29UEVIrNlzN/d
zpyyKXwE8YK04p/5M0Y2hmw2bMTNGNaEpNRvIRYxu20y9yxtl2PNZAe+mjh8XdCEiIN/XCfGCfxk
YqJJEbtz9iDVU4DVCtC7irlhowC8Rm4Xx9jKr79uiG7Oc4j6oW/wtTbleymH00s/kQgFB5dQ/b2z
mHNXEwmEJ6I5zMV+qYBHlkjGtdauzHmjNFmxWRMrW8JULqx/JBmbOsLqvNIpH8BhIAkZgc2He/cO
edWavOj0mKHpJY9IjH0Dmc2mhDq6/aSi2iKT7rVYEPBwWOFhglsT7gt6wx5CVkdOT0ks12Qd4vO3
tGOiKsnfHxHVMyP91pRBGdEnTRtuwAT0XMkCsX02rh8AbJ5eEaHbYTYsDA8/BQBtnJ58wtefhyM4
zBLWMy4vBhqG4ar4UHhtpfOO9gU+zzI8s7WVlxL8zeOGP9BXpKyWrPVrAlour8Qq4BB3sa+wR3hQ
L5iE85gGS9AW6H5YMnTZhMiDEWrfzsSvIbuxNS+w7Sgic6uHo9CgZEZfuBh+rZWvMl+CsLuojnRP
Rt98GjsKn9uba9+hbTHh0CUHa8BOfFqxSUgSHWSsh4Y7aVYLu3JojVKd1l8OuMiuVLJ5w5b/Krxp
c06rXVsQBrFu9F2BlUYWY8WGF6hS3rVmxiPQOkeE7t2+UZYJ5/xBtyt0wP6tAqvppcJCB9Ar+gJX
BiceTYXb+8KG4XT8G8ZFbdmxZE6Rm8nACZS9aRC/A68Qy/izzjsUFDSPOP1fkl2FC2JOBBPziG3i
FEKDRTEdinYKcwSVvQB2U5810STBupq28dq+ZNZlhNZXBsPu4JP6Q8ggXifzdHl6CQglJrIVhqf3
/yTlmZRK2RYx7o/gvya6RGOFPYD79ItwqRoKHWJ/JWUgAx8K56zBfpvOyLb63wSmASe6eMjqFBO4
MSdj1DtGvx+t9iwGkqSpHN0vyUTZbcRgoaDg6EABStmTiXbmC5DKEKKMiu2bzDzUeKkOsFCvgYnZ
bticD33YdvcSm26fwSbsAV9iHFtH/KY7/LsuPtfGvU28pGSGmonxxS6aiw8o/qC6lILq8DWkARm3
SaXnW8cHCSHYBX4un0mROmD2L+7yzFQpHrrNeFetgGG2yqansEBqqZnCiRDeCN6RCFW0ZEOo/gou
AeEXVoRRemiE9lQQm2aAp8EUTz94UXDxfMsuWopaIcYgKu+Le1/Z0GUobPm4suyCwJ9p9rMuTQjU
V4PoBEC/dRAD94HktdfP07mXMBCYzNYyabaQXMO2LNJhdkdFt5pCKMfvZwcw0+lPdfWL11EZrdjZ
OuZATho+Ryf6mWifKm4rzfuL/EIV2mmPCpM7lsRjVf6Hj/5tGq2jn7/29uv64f5XL0hhAuDevzmQ
1ceCQGQBncXxlRc9oUwwMzstivMcaj7bYtddhaRRYHEx9HWQfmH/0k8vT/ulAfAPmnX690Sk4m3G
tzOsjPwS3eJUsWNiHYuijpgtBAzR9qw7MupCEtPlt0b1QauUMzCLio8TbK1oXE/6APSbsPHvPE/e
YHfLZEnzbKpKeHQn+FwpKjw0B/1W941dz8yGzXtvcx0gDD1aTnB/EUF/CVqcKu/ToDiioB4a2ApL
YLZUKp2q20ypnRvtwAdUk4+b9CNsb846rVVWOEn7fk2yHYHvxeHXpw6C3F8/o5RzJTFoIY7Ni3uZ
rvP4+AAsCcde1XA15grXmcIvb/dRnRFcppSyG/NJIM/s/mFf85AOqJgS4KOXYlp2KOYVU62Fczaf
7ql0dViftBRpTRguqaPI68hv2zZi1gLiVbxlpwm4Eh1FmYLcrEFSQKdDILB9W4mK5PBxm9m2fPY+
fUBFDMDeV0FL5bgydyeWgY6mNhWCtlJ3GSiRZxiqXFbb/w6J4Fkg9arjjtNZv4EF/5JZNi5lHzwS
Vedw+Xs+NeJW3/oWGisH4pqH3rht2P98PKi7uYDHiezCLj505txG6JGoqQtkWVeSSkEM6wT13tnK
gfQglMgx8XmYEEJG7qXlSP3jL7emxOx1T/RbxvxVNofnadi7oANnf3en26V1hAWTuIRuMkzLffgA
CLydkosebf3aW3yLEZjPXdNisBsJcfnqKVKnbFHf0YGjwzwgdmSCcBzTGTx/lDLElqd51PLU8I1u
of6DcOTom0OFAXZQ9PH7n4paeJmHszzWb140B2FQIbqmMYaZiyhG5BI1MeKEBp+3ZO5bc2BpvdRX
UTvAy4RIWZVnspfx+SrPRywpiBGcvcYHtoP8UkMXtbgceJRKFF+eWb+OSt5w37uqPi+KPzZAueU6
zbjcecVJcGEa7qIP1FtEJRcIo4Pg2X07k7oiyuFaSM2ZutYd32c+Q7jLfOU9IjV+n/+Euo5m1WcQ
mme8Dk9B1GfLLyDEKCYRiiptDBsej/uf2KxDLoM1X3//1yxBNHy92HUAtxSq8Ro7QyZVMsDgL4Rn
OcZk6dieIOrrkc3q8x5NprsU3o4oRBxuKhYlPnUs24ugTVbmhYGpPGf71CiXtCBsH9b3dvVvRAFn
cUmQQ+/1xcMoNhuGwORZRK+Ge+2aIiG5EEjAAf8KKdm9dW5nZnrbnWcjQyj+m5iRGOh8OoCu+thI
KKxTdYb3yRPCOBaAATKeWISf6I68u1YNpczw5FCCxYqWkFnM8frCOjP5y6UAR2dYkt9jCoYc6Vk9
9lSPHT6cst7jkqqKqNkrm5cAbPY/TllM8ixAb34LxTYsy3xi0qSYJiVKlJ/JhqDxiLjdewZDvjqO
1rh4TlSayw1L8vd80fIPiNx4yBzG8aXCK+CnGt6R1LLB7DjQhRf6fcQHmwjnVEW4SC6SNIBROyNv
La7agBS/p9OoUk1tsefDX51AZyvXIIFa3CKzPG4g7hRMlmEfOhrIjd5VIIn/ZlqWzzM6SbaSoaEC
ztHYfQzGa1Hb/ns6N7gdFJYCwNB7trGazRNlYtnY1n3z3HR0PIQeUKoNGtcu4AnbPc3r4Jy8Kmpj
BwDprW0Q7uocAz1tj9IyzlqzNbEdsqufs45Cq9/yHc5PhLrfmhAhNg6M4t1+NpaaZo+ngaUjR4aF
6zOGQv4LUINpktcDC3ivVf9zahFXEJklgQBxwSzG4Z+zR/qdQIHAQBWK0suZFmDItLV5HxNL9kcQ
X9n/P+GrTCsPGE8Lgg/cSH9PgyhlD0L7DsEEx7DByigIUPwJ0aqpQqqr61vhy210sPwzrZ1h+2PI
wCXxVrIFbcXptvkV1GmWticmb7Mr8UROR7tDnUPOVQcAhXbFMENvmNSinRcWzXGtezZRanOaUw+V
GR2irsihOuP30uPH+HPMLGuqTnrNeOuTW00j6jOt2P1E9HU2mV+ie3fRFzqxyxdx9zojK5Fsu/MJ
7OIiVC75jWwToAptnRCQm9mJMofIR4p4Lv4nGAW9xq7kBgy1zB14PrOnEVV0pqZRlHvgSV403rsR
nOsDG9A5qxtAft0Q08QmcVFPtBFzd8XhPBDOTEsIttmNo2yY0saocncjVpo3QizbZ8tx8xQeSFOh
VMOQGq7AAPFd+6DrpbNt0Q3D06MVNnEEQtsnszb/l3ekb+Yu2kF6OJ7FVgf67vx6ZJZwsJbGUWFK
8mhskgoebcrQak8SsvOAq5o9ye2eh7MBDiAbZnUGK21jOVe6JlyhRNxZ3dgRhVvCVVMeK3TbVkbd
c7VenhdZedylIKeR6CWfkFoumCIkF+BYlAzHqy/S2waPQWzydEafXnJss5CJBxFkfTCa5+HRAgSD
cUrARL6aicuUUF91qDmUn+LIt0qM2er7dHBNTZJ2oB/9mX8gj5lpqUrlp6CXbFmLrFWUbZa7LrfS
BFTok+UHkyPQCtp9weJ+3MfgKItaVaXaT06lcr4zssWrZtxuVi4XyxDrOZU7+Rs8uaXFN2IRws13
VhmnAm12fECEpcV3tXuilDcyeaUFxt+2BJWNVt7NUly8SHs63zIFBT0G02WxRbNBLXN4uELtrY66
bz/Y0akXY+DHh/IOnrJebtATBAuSJQ/xsW+9fKdhBVH5iVb5szGN+7E5Bfqp6SKxPIn0+pMFpeKc
wJOJXfQJyqPfJPZIZNmUPr3fvH69oreSWaLVe5S+O5yBal6IpiWt8w/fR3UALZI0freP2mSAQlKX
WqrSUscvzlzzE0xjlEDLxsMY8PKY0OVcZ7Llwu40owh3HgnBfD2/dY54Yv9jMBYNvtY1Vft3Wgmn
yzu0O85p/1X086cg5s3seZ0Z1fcGWaPIs8NFy3X1AFLcEMOcWBcjYf3nRkWBJ+wW8W5hkMmBr/Fa
fqH6dbwfKxwAVihYbgISBCtn+wMCZq3vv+OqT6Me9OfPrGR+JRCYE6XgYIOJaQQ2ljni4CLPwtDn
6RS3GTog21+bw07lkEfTwR62S2bEI0nBYn4Jw9KfC6bW5K5sSgclJpHEzStO+b5FAAICAOLl/ecn
VERK7ua52i/Sb3TmuSoobLSZtyGCP5hAd9DL0xpZbupSyMH1k8/Dz5YQFI4Y41ZLzA2K3qePKWrT
h2SWFRZudwHToSjwjbd7+ijbiuF1hlK7NyrZ4KnPmbcR75bIDhYl2qr2kvTpjpbcNfMDMdcbhtNN
mDv7mqOjb8sCT/gO/WXaJlo/mPW6OLhMVhSEUWleUITfeV79ekUSbyP6fwDdEHzzNxypWnOfJKdu
y3hUuVhou7fF/jCirv8N1rDrwYVWzyFi15ZW4oV3FStCV7XGYkxriNnnICku0QAX4YsAC9Geaw+m
HI7JeEYX9zmZYT4C+sS1NqO1l3540FezLKAukG3WsnvP26eDgBz6k7SSEX0qFeI7u8xjz0WJl7Yq
mltD7PgbvsE81d0EsW+DreOldRbt4lx471HUCtOPC+0COf+6Wm/rqEVy9IAHV+9/8Rjs01KTGNMK
3b7BHSkBh92h9KeYFMu26oJQZ/U6sGwC6iPukVMriabmgiMBTPhpLPJlcWg5NDdUB/uLKZfhNNZG
6Rjk1ZKxGaDRjUvfRtoDGSGYvRPyvnMqZaUkvXW2PsHzw+EjTuUo6hUCWI+uacmGttXcPKbdnykr
C2oftbh5kEJc4PsS/pzgbFgNBZI2DFFota9O2Fmn001h7GvfY8bpiDdR6iXZk7MrhmIA8fHnUZ3N
TeeE8g/1DMSBaC1YTtrGUSzAzQCEUhzaeR5aqOFwfmftRJrJdjQ2cE9qPBDQrG5PPRrTz57+TXCD
Tjuaug94rD2TatylwA1A2ubckvlnGQGO6548OXOKpld7TLA2aPcEBvTbFVhy1Gf/TibNqxGRG7N8
icb9pDNHIfBI556LUCkfGvsrIJhVSjQATijlASqgCXV4RsDRJFp3jXmbgw+EvjGzTtbapRJ8qgm5
htvTKBOGXh5jP5+S+kHXin6ZdhxmrOF16Um+cGJmsUbSsiYCFjYLPckUQJVac1JFJW9VAdnaKXst
iQz+PoXfkXBYmGj67i9997GxnIKHCU/yDZ90LTajFt0vtRGPKbUQx9ri0ENqTUZsJG+v/aeipMSa
CnuOhksxJ4y+reQDGeRhlKdfyKI5i5bN6JNxGgXNIjl87ONLJZgm5yHUADFMy0m1Tz26GEy8sxzi
esvAcSpaobZOskFWPhzsYQZcawHGq9KZn6o2vOq3OqXnCrNhsbj8LlkvQBK+tOOESk6CXIo/yQmt
rvR4c2zUZTLXY+VEmzGebY6s1WyGOSlvcBMRfN0nKCZiLeHtORj3v/VToumq/F1BH1W4/0qu9FaV
WqGXjBD95e5tU7Pj4t8gRt3KrHYi7gm8dpHwVk2dqwM/j+TLYiXd1XkqeqcmBZ/MUf9l82lw7Jrn
iVkWSVjSOj13eY5mw7gg77+BVRQ0vcIF0iUnezQlR4wCyjb+vRwMIRzrJVYnLxDcuSIb59lYaxf5
Ae2HscJyTHi1enbUVIdMa9huxLunxLXWZXlDEN5qkVvIBkXtIXp6wEHx5nhDv4LU0OeYf1R74fDf
dIAqvUXSIn+UZV/XPstbExq3vJk5dhvdCjfLKwbiQA2EiLRNrPTiWemHUzDlcl9Ixxq5SREt50fK
IC31yDQHR0LeLIbZ8A6vctWdLCNsRxioJtrQ0AsC3T9Mt8j72uKmTy7E1cuWz3GNMURL004a1+69
RIT2R20q2PUSdmZkMfgazrcQ756TnlFVjJTW16nC9qM96gNSGAVPXeqfM1D+gBQJcsub1QcXCTdU
rT/f3t5hDx6ALE9kEAOZdciTkaKUlePtR0LRSa2uPXQTNxPlUdkwAJ3ReRus4hrt4LhEtsPMYtcZ
RQkqjZrRoCloHOas2Ld3/nM99eTMnuo8s67uEaZlXMq9evGpM8d8+DbZxg+iPsuHGnTBVxSig/OH
lP4urz7knFPGSK8GyoRWo3icjqawgeE2KxYlN7f29Hxl2pzzvC94E81nfVC2U2RoXbXG4CVyYIU7
10fpNMUQqGrzpiwMasI88QYHb6k05+WJfkG+dtXwcJ9iWhuPM8VSExNd4RI6zy2JZsXsfdD1GpQn
ch5GYnMXkXhTlF5842aAtz0G8GfJ1xCaYrX0QsnrsZLBRu/Oszo47bt81PL2VyD0hZYgN0grjV/N
YWsvXnZFXsfdGE9HvF/cteBZ9Y4r+8VD1wtuljxOS208enGNM2c0IFOSF/9wDeS5X4Uxzup1kg+x
7yZ2lfLEZ+HMHGxkVIEEvCM0vznkyIrPgUHcb3Vlo7IOwl6qPy00c1rFGHLqngVtls/sBgZ3p1hP
2Bf7xth8SUDsYZipso0Dz8G3D5tWsA07pWpXJNgBfpzHi95c4S9LZfa0v2e40oIIyHMmOABo7TI1
qtMHuiblWwuooWpUhHsGlIPtQm1pX2UWCEeXwRwbqCZJIsXG7tVzHQr97vSqWL6ZTzEBtmHd3YCz
YmX3G8NzDl6bmvGYY05xY/mqzLtE3SzWYi2vV0CrjxLDvU1wDZj7yI+43mFXWvr1WiJKl4AxfKFA
tm1QLgPuWTdPAL2hGEiuMKw6/ANGzCkmnzzD5h4b87yPyZZKyE6cvoFrzi7GA6OxvY/KJ0E7hfPL
MJKpKH5VNHs2GB9u1CNRAo6HpbXAjhJ0E3Ht+C57ZptdSbN8xLotiLb64T6uzq2qD85obcxWdRAl
GH79oWwSNWHIGPFftnrhjZFi/je8syu/vcSL/CCifgJZkDUXYCWjqCP7GVR4/bQbn5aGDh+CcFpQ
x2tyQpLAa/5rScYwb1X11QEsPkRM0khF+LE4YkdYvRPW8qU4IQEcMckIjpVh7h69H/PX9GwbVluT
jfC7wcbDlOCL/yI4mgLdRZck/FCwCTb14/NyB3sFMo1zAvGf8/fGSMSS5G3BcDP7eRpWR5VZ7brU
Nbu2yqMydkg6w+tzrVaR2iLDRSTKfbaN2tHLLb8ScVtDVNgpzq6/u6d1wlBtDVmZwKYXdZ/Xeb4R
A5/AyvqVr4u/jWw9ydLAOJ3omO3buWaGv/0rrTbeoaegetRuZcb1k7Vx4tDB9PyRWCpxrR4Su62j
TL9I/WXutewLANZRKUM++n7MFAGKDux1vY03sRebqIkjsJVYKqF9CIg35VDswDhbnMpBFZIyV1TF
Ob92nFlwKqdcbVdUv4NhT06OD0XiMexp4eS7OaPyTgJ1tB8+5hzYYEU4jToo7A74cZSaKGmDeRWi
iAON1jOYDGBpvvm9xMu3JWuiRwJzZgwMMnwqRBL17saKuludlmayXX0t6sOUbP7oiNsCbPxjom5w
hTkTTgqExHNXoja/8fVDYuXOY9XV6RdpNfPdCWUoNnKtuNqbNGT7RoRl9N4jpn3fbb3SaTien5tE
d2fkdsnMT2YGrqFH4T+jQfWhGamY1AD3DV0Wn9dQMORVLi29GZHerk3LMG1OMtC+fDXPn+3UjXKF
eL5+X4LMomGYdotA2DRtrJIm0sj0spdF4qWBDkUSs2MWBC2jTRNf1OLZyA2sLopYBWhX6/RAwqlT
ENkS91U1QCBIcCR5IxYX4YFZIp52fwNry91t06JHGlW1shdOf8C90L6qW6B5yUouGaRO64YuQj6K
zGt4cMNNGdEXqi/W9m2posAkiS7DcSjjJjJfqT+7s2PeS5nTm1LliD7ecwwbwkETPB5xnFal2YiB
nXriyC5J6oZGa9d3iLBwQvfEg9c+8huvrSFkWhM6aUS4meZjHU5QXxW6Uyqjnyyim+jcS5rDcgSJ
jS7v/yVFsYP3Rqfcxu/xjsxgunEMz0V46Eirz//P3W1Rs+zUBLSNXF+4xJzzCVpXXAzVeFkHLUIh
/xNYM4Sn9Ol7AGO5out68Y/eWKTq1QQNESVLowkJkGpH4WwA/fLJROQtK7Z2Ak7Sd/uQSeEn82d7
X99sWty5tnfmy5vVvzTBMSEr3Scf4iJMdxbpkkXdWJX+4qfTY2R3wy7SZL2lNKljcZywguOlFPNp
W3ZkCiI3Jgz280r0KsNRTHQzlBVvEeAYjfsKQDDXtUdtHENHGMUkYVNIkJ/I23vM47J26gHIXpIr
ewK+FbYYQR3De2gZOmYhc5y0GojdOpGGQKPgksIY0AP1Y30ctZcolUVevqtEKAfFUx87P8h+x8AQ
rDw3MsTEkgr6tufhrbzMUYbORshFNDh8y7WTIE1QehfoKbNpW27bDbK2kltDNPTnv55ZNeDsCpdg
BaeBkMMyl6pF4sGQbcvhqvqOb+gu0RK6udpzx2YOesh5TNz1IT4gOiTzXVi3/5TuM2JLuYxTwiBR
GcYAWespt2zFojOxkG55IiObcuZJUmtKChjplXWjMV6nPH+dwcH+ZF/5m6qozN4L1HaYzN/RI1yt
Bdr6Yvsn0ej4Qt6EyV5dl4bRgn2ftHd588hodH3JvoMwzXDa85c5cw6KH5dzlHhvIn8ltqBJydeX
qV2qgpoNKhKeu7EMfpcuGtNRhLhs0EtvTH5CdRTm9Ets5R9v0yBhPOoqWck7wEpXKgcLSaYJjWlT
+EwoEILQjVLaGrgXDOCsQk4+1Pq1Dwssdnkcbzw/GnjQQtV33pv1JJv46Q+Ym7cTCgBxsK4XkWiS
BBFUyLQLtvBCLBF+1BfE5PquL2ALdJTTYaCX+HNKEYtmQ3j2HlBYah6M2cAuSTYlvCzdWLpXCe2b
MJdtBVFj+cq1yanyqxiX5pi+9g+TDpDy0r9tp1gm4ZlqpnaQZ5p/u1OytQM7IoKXvW2rS2aJcdXa
dDLe7qTPw0/b7hAaMgJvxgOyhUzYhBAqvsFnp2dHMFiuDWTHuCNHiCBKBUt1Pes0umaTTC4c8m8S
QW8VEWSSBmawXorNPkcAeli7BRwQBfUnSV02vvx1zlMzJChf/ys/GudhJ3EhsvdzgQk3xMpOFtS7
w459y8+5ajLTUEnrc0k8zt1WTvqO19YVJBmrFp8Lj9kpr4pY5XR5RAMBK+VN9yeMYaF2kDcoZ1jN
ofsZaTBYeWQ7OEH1H7SrSJtqvUQoCI5Z8PTiWcQevrnOZG7jcxtjVaSYIyfKrdLB6jp3N6Jj4ZEC
/14D3QAssRoyrbNyzgsbbaZ+YQsrc1TGhuZLUFnHPNu5BFtjomTCGuHyAZkFppaZnxkrUbswdVSD
C2mMggRUvb+eK6V1LfEO47uFrOEJ7240c51d5eGI+v5jBcxrsBe3hwXf3ER5OUVNcy4WbneS6m4c
3nJtPhGpJ3ehifKNT7oi7WEWm9wc6HxIZRQXv3BtRx/Wlz36TT1jDLINYp+YYC8QWNAd3uexOA0D
7tEtcS6BDL4J4CRDYn+tx3dsvVBi43Tb2i8A6voIy6HnpWU+XpOKU95aVUjJyXQbZNJ8o3SCy5W8
dnUJwRSb4VfS4N/z+UgJqh19nnOOjQhWdpfD5rWK3GYha0MdC39EPNvuNgu0tvC7+PO62w4nhNsp
TZFetoCEQzbHY+IA6Z23Vi8cPWTqZn87WSHgG7UJckn/5Dq7NpVT/sD9XNMXRTSEU9Tk3WuUAOIY
Uka4Kq0PPURg+sFce0TjfmFm7FDYgulUrJO6M9gQEp2T21spCuL5O7qwhbLieGPg9fb7PX7hAXjH
QlOf6GIxUoQv6HKcWEYJ0gyhTInwf1RbNTC27Cn64LH5AMrIrgX2/QUPhI8EyfMoJKLhlWHH2VC/
EgLo0A3RZJmM4bgsxc6H02bdkNVdD3S5afqLdHESww16CsMn3c+hbZKkK3lS6jCOJeQgk6v3JbHT
29FHfsOPFylJbbqc5itPO2pKL2CWM1hFzyTghd55CtSpZy6IJfgssvu5Fcxw9kHxHyK6ZrE5QcQo
gAZpk+jELKtpujAqecGjYKe5z/kP8lXsfoX42jxaYApeaDNCooSWphaPIfcWMxvlSSVx6KSzKOBz
Y5MfHziFNlobwPBJBjQEWagoUFT+6Or2chA+YWpxofCFzs3UW+u4v9l1Wt28U8oRlxQ0IB17tY2z
EgLIPsWed55KnpgMf6Meoqu66q3tyGFZZSGSXDLW0mICY/jKcF1JMzyEIvTFrlJsXRYS5cCvjjvR
4/YsJXduaE3emJ/+TS/zAdcUolTwffg7m8mf5afr+LZ8mR9zk9U2kIy68TizMDLEzdKd3DQXzENM
eKJGJXA5HcsnPolpjCpE6T3f7p3d/70XMPrKuzzgPhLAtc4WvqhqwzSfK1CgkUR/PDBmOB4DE1uN
lLhQpHituLyqa1DEzrr96SjRuACiyUWYKEu1xCSabKIRuU18QUDyVfShXq0jKSR50lUhzCovuGUB
MObssKXDBLvhmC874/ymQRc3YVJjlYJUnF47hhfvpI9eIOaHNii7pCcBt4/5e3oDYlJRf9BVUh8g
AR7W04ZyMQrPDaXDDnO9TPdk0HZhVXQRFZ14kzsPG6BFMy1BZTaZ/Wao7SCQXzsiLGlWwk7wJNrX
Fsoq0DjJK1MWZLRmcEdDz6zklEDLFkI7fI/22Cd6nMfDf7xL1YCIdUxaWz9TxPATTEtkHYm2ly7a
/2R3H2yJ/T3h95ap7dOzn1OuG/mk6/vYLMdYAONF/mJ6NqM493DmQQKSZGNqYTvt+U8xW328JKex
ui+Q7c9axaV/ov8Y5EtBm+SgFgHLpwRgpomY2OQi/COnZWtOgitMnBK3LaISKhIJ4/bTVBQeWPqr
P4+rtlxFxeN9xrX2+bswgC3gNAeXJYxj+VbYSbbaMrgsrntBfz+mB0wvW7d9YPQF6EtwxIHAlKrw
2TFBUpNePSYfjApi8vqQt0AbvJdzvnkyDYNboEcwh0kL6E9el4YqyfYeC4XSFHI1fR/L6anFgzKI
qd56nVXoEvEZaV5uq0jSdWrLZu8nl+XWZ9ys2ITBVCf3LvrBM+7UuROx8gkZB3d18qKir2JtUkDe
CCmJ72IF38KVNNbVNwpfwfjtDfttyNXYJzP6NHwog4N6EybhR+ew7c2HJ3mnsFOuklbkvcB3o1kN
bJEZO98Xw3QycF68TMFx7wsL7dQjIc2WE82xyzcBwURNJ/6OoQeku6lKZqhRXgpkW6ogQXIyLbPY
0mHLBMWfvNG8cISpaBOmSomHApoV8R6Yso23YkwoCKJnSvW0kpJ6Onk9uOZKVPWGFfDzR3dny4I4
qMZ4hqXMfPad8VnwCGy+ePXnSozhSIbK0USbM384hS5KRhtpL6UAadP4m+O3mq0c0wvTxKkb1m49
l80ZvFu3i9uBgTCX65aKZgI8ypopK7be04GRRFKQXE5cgNoPOUx9mrWUQsTxgfTrO7fAxPyv6Jdr
+mug1MdnYsGATuTgAJG8zqyj6NS/ButyDYvk4pqAirALBu67V2/pVbi91UwqesCXR42LwoCILlvV
3hVT1urE/M0uPTs296Xc/Ijxt3lrmYrnlqEBSP8Oy2HSquDRC5/kYDQ1FA5tzV9ZnAzuOlyW2OCD
ihUpjLTzuW/dZthjO2pPFVyFTA/FKNSRfSkmCIKnCMfqsU3FB6a5dG0yy24puZXrNIfnII7d7pNR
AGadNxtnHMWVRvHlb1dAhwK2ldfW93zBXF4DWdxpmDEjNznrHdVCMEHBeBNw/xG+zv4x3qOCcgyK
pcQA8mkBmUT18PZ+Y8TnxJW0kCgwtZ7u6gqPfXfo1sX+lA/5WBMco+scNZAUHWhYoze95r3hxhH4
My7FRN4zXfMocc0IRlAL9akST6tf5o340X04GUb6yiFmTIrJRkBuyppBjxEwg2ScEPxqY6Xyqs2e
gkw6yVs9VTq0auHppeJHyLOKO6FP9vsmXoJ4C9YT2d+7ci1AZAX5bY4tqIExrKWt9eUIHeYf8CUv
rIyV0vA6suSlF5186zOtrYg8oTQHOZhWbNkkOO6+Dd/YvEVv4vp6P7goHlsZurSZPivJTi2Yt5kc
F8rzPM7Yttr5d8Xebcq4ZQ7prppkxeEifr7OIrnug8GjkK8rkHc+YGTfAjJYTEMG5hX4ST7jC1/x
D1iNpyK7uCd6Y6nRy73seFo8L+2VJpujdekm4BW4+0x6fXxjtGk7EKH1kNVt9Y3k92/yUJTma6NW
XT5NXp1a/6IUXn6ZuN8Kd2l4tGae7k47M4KzfXY5fPO657onmp53ZYoBF4cYT2q4fKP7bEMgdjHx
Ip0AHV6CaCzTz41JmLww+AHGLGcgsDKvbCtAY6etvUNK0as31vT6S5b1yhtBKYgfsgAkgtA6DWgq
ce1Q5udciit4OAbXdtk12MYYuIF/1w3SCf5wmw8Qi2YhgzZ6OpEIogy/PFwpY976QQ8uXdHFTc4l
f0on/ZN7vnQquBtpQqsaPdFvwXWKxL6cVQdcECu8RWrmqhS1jEgB4avM2mih2mfk4JcG/G8Qj69X
9xhXQXDM0BBxkS7tMkvoikh6aF/hk0tOaWaZ5xQawjIhqEwoLeU+ePO1TP6Xw/INTxdEUwgBWoRh
HXjpHB+lGdP9b2CspaadMeAwZAMVaq3bZki0eIg2gqOBCHApFfL5WdtSrKYREVFkCTblyKbEsLGP
rWzGqVnJcnpmnpG/wDu7agF1WiZwi0kVZzne+CLAPHw8fHxtjmOUyQ/UFhFMU+KlSnIM8WXo+TXN
1T5FNrcpEUmicNNOy9IrP+Z36aL18WFX429lBEX6ZdQmG8s1tkBMOqc2B2Qtnr4gk7mQnr+LwOER
dGlPcAWj4IUHiGibtyJQoE/Y0vgSJizTtHDEaUFZe1fKx2XhmM3N6qDCNjJv5Qo4U4wCwGyfyAR1
k6bFWMpfgkd9hquTvGaG8VyUleosil7mJLOlCuY+IQIbBkUl1a57z0dr6C+S0xJXCZCmNe6yhgWZ
oD9noI9egv1gRkkG3XU00uNBUaRa7ESV8YVgiGZTTUKES4RUlh/f6nGwJO7aW24poBOwYu0TIMsj
Q5l/fLxmgkDjqJInWqgVAH85kJ2MESynTxMT35RdBqegSp2qoNsDSMP+eJZxG2ztD5ViTTTkeIJC
IqjUBzNjFW2Jqa/Rdoj0cD/ejo2lTJPRxk2kfFKw/WxwtH/g20SsYlPBydGAjVK9OpjSCeF37sDT
uBCmjxnDwIBecxHJG/t9e0nl+UW0wi7CLba+NVofVJMvVSSutNgeorfPzWuVxWBE0pw1lVmfmWjs
BIt1XoE8Kf8oW2ZuDModBMXbfncqf0bh3Py2ivsZSN1OV0y4r31hwmqmtflcobZlphJ3ZpVQnomC
rOxAMUu05tMTNVUzx7Pl2rJ/FXtFy5RtUDl7Duw5kjXjdPCX/7cHR3SeuD5I8JjJ/37K9E7OjJ1w
1zZgXXXyEgki9rHc2arsZoslm/7nCf3fv/12n1971JxyeCwPvrrN+jx6CiqgGVHiySWlLOAvPZU4
sMpBFh+tUH6zII8D52p1YOhTwF9m5yW4kFJ0nstlrnBKkunzX7dVsP2dhp82KWB0ma4/vHbOs11r
6s/nsNhPZlyfSEHoX18IWjJJBDXkQFqoKwoEDkwfcW2R1cDBUu270tMS5magMQlD60VyotyC44PD
kzJGVPNkfKXeexbqzbkKGJiHEhHfgDyt7OagAB82G2tMMlRQSQoK7ViKMZtQyl9Z41so6ylDQoIu
rbi3VoW8Gg5qGfOR/496fdTaamJivWdDxM2FJAeaSV6HfK1cBG7DdeeyvMTiKgVR2K7f3mOOVA+g
/DcCHaRCxGb1C/ya7SV1ULhPcWR22EYCadWKt7/QC1hNZyMPiOhd5ivILLBGF6tKpN6+i/D4APfg
532imio9l7luGtltGCx64UcOiwUxgPgAA7mVFK8G6nT5uj1yBBG9DRouxT8FSD7F79NwJZi34pVp
ZAfke2LURg+ZitRocypHvq9AHPmtopLaxeD0+GYKORSaqsWjtUKFomUZiv+3l87jrex4OaaAUyme
FG1/7I09oJ0523FqbAx0QWnH34UzGon6LudXNoxLPXY29/vwnGLtRbfBzKJ45/noblgtMNSDj1h/
RFLAsCyOwlZzgMrqSk48tpsOC0zyWShqdAhhxATdjhQwmWCMVeF3nhKrZsVNS2FCOw2qcPpCJsyo
ASfGbPXn1qmmKejYnGkPxsCp4D5E7c3OZJjJSWvkkDS8bj8dsw5ubpQwblcNYtU/6IbugXdGWHyy
N7TQ0XOS+vgziQHExTHsaiybRSlBFpZN/kX4OCYuKbOIQovnnTcPY3OLXH1YAWgD6BZySlNx9HVp
84KYDFrzSXQUefcINj7sw3ByfaE3Nob8DlMS+8G45DoECLIifaTP8mQoKD0eighBPqJyYygzee9+
KR1uS43LuDQgmZdXA4JRlZVKe5O+xGhW+sYpPx9xaxReQwh3JE21+lNEmRKZMJ7PQcioYdOkcPch
/AO4aJ0NYnqYjGb0iHKpxZVq4q+QNjBshzbB5Ax/klWKvktS19JP9GBo49K2iLmMlU9jfHVIGIl9
vPNPcfZmmzFeUeIu9OkL7Tksflny5Lho8YvVtAcpbpPW8jpKjMUfoTZDD6C0msQUANZki/OagIJ3
DSUAa636FPqPBxCJI6CwApRR4Rph6SE9vSOQ8AU8chGgBqRD9O3R9PB0/jZCdIJ4B8mLnK3OBL0c
5r4CAxNRVFWbhA2w0TDBxE2vBMj5fU6m3kpEWXapINCCAr7VVTvWqWH+LHcPHL3YPBJ/d0TejMxW
zUML6Id3C+Otd07bxMZtWxUyqj6+yTWkfGq9F5X0OQKljLiMoMSqPXwgoBqMCW/A67Rr5E6OrWg3
IIGi7FnTc8Sslc90iOWOvbPwG7L5jw/9ROCjK3e88TaolmdUQ+xm/DN94YLUwecoqS/fMrbE5NVm
TuYZvISD8EmNypCWuWF9c/vfOwV/twN5ahCje0knednC6hpgdmn7Wf3R+fRLLaeC17dyKxt0WeJi
VOyOpjPfa9D2lPfSUg9toxK/+lHE9e8TaOSrwuDYOwNcfCM53SS31XyvVS5me8xOThVgQ3chlbKh
DokiWJsZxglk9vyjFihT4b+Q7D7OdkZp2PXwZ92pwuIV/5quSlLGwB23AAg5jCMHbd8h79CFeoeL
pPEzqtU8/sUtFTwCh4pwrrhxigbXDx8YQT7egnN2mj97m5DCxbCo7oJmMiWTup77FO/6BZfZS6WS
B4Ys4qIYHTjHTt0ciWtvMuRmbwU5e/6+g/ihKyu7mN2KgJIPCm2k+/oZRNJDkiFHx8iTTKbY46T8
Bmn/QtKfP/9qhTyK/h/GhFQIYku3bOAJ+ZTpoZuCKjt2gl+oLq1P6ZEknasOBOwiaZ5Rwa4GE39v
fuW9OSnCwqR4noFnI0ZTPCXNt1QGpZ8t/r6k6F4mlv+1AuD/ER+vOOVZ0yNvRrYLSLcxT/vaPjE/
AGoCo6KP5SnrZB94iZphN2JEdNnX5sWLqfPTRM3QJ2b6D86DuqPxEscPbxb3e4GlttRZ1r/dybf2
QcrDblXvtldR9yV8M9C8qqj9xmTn32z/z2Dd23GKxACw/7SIuE5dyqjVHYsbCCoXQLDEN6iIWIGS
YarfeoGYnBSmgM46FDpic16pINXmcsQ17+bwco1SL0y8uIZ4LLwssFVe/GELIad3DBAmgNraTc0O
V/RBjfqgseiBw/Gl882VVxMLwtpW+VkUZEIecTZpso7jDIAaMPTnykHwtpcs8rnPNsqcKJUnqKHq
2lpWoRdxwnYX3YjI8Lhh0tPI/9IpCvYX7CpnwV1R3PY9PJgbrMo8IQ9JWM6zQ5aqsWRyYUjHOJ/6
boj/Bj91sHPcyA3PxGnJMSHc1rE6UGnynBVlbi3NoHiR0q+mYUxdmzKVOPNC0VBfMBccq5jSs9An
3E3M+t37JP6jb/s/QFH75XPXolaMdYWTINIXDSNj5goC8NbbGER5NoXSK7pWr6+jSCwt/ehs1jLN
cAF/OqlfWZ5CHDsCJmw/33uEFbMFIZmH6qqSOcz7+L15+DGfD0OyuHUDTeOG4OF2QWHlVRBMb/QG
1sURY91NoIMjaskpZbpZM7u5RzVl5TUtBMpcCxqmvKO8cTTE0378HfYXtVkuVmyTa/ypQHhR+2CQ
2ik6p2V1vVMxfdR9nq0miKMVIv/Q9A9GXOxaZ7fnO/Ta3vt7bJpYasIPeMp6p22jLRgM/CmMgK4g
ibBJH7WsPKzbsfwftp6g/Kd6tq7tpjzv231t+N9BLNao+LX+k4nZAZdGWrzZkU7pf2ICcBNpFZoA
mNNphSEt/Kq+PqfpGFuVtTPoeMhm/h2V5EJQMOC1rf5s2CM5wUY7HgswlIEMaD90vNMUbo12JjQx
5CVTw5ouo//SGwx5lWo20LKFxqo+VXO7w7mLzJLR/uWxAuv9g5AIQE/0TFykH9d+njr6+fQiEaQQ
vA88HeIJPuLaNMg/mFVQ06K71JbKZ0HBYgWGYa/jV3acpS9CsE8SPQTv47fMz3Tgg/yVlHJD2iy+
6bxjMhtkZrf1fKmvPoW0A4/IP0cz4bhcEFbdX068A/7rZN8qANK/OW3P0QluRaG8e3meLZcyHlRt
rOhhUtpPjp7kdnXPINg+zUQMCCcULTxNvyf9mv9HsifxHmlO+D+qzDqDdONI0nQcfIZ3Mt01xop5
riPUtN8Aol1Sw2nGveyMfiyZg7TqoPAvh9ndApQuRAvgb8NyVJO81ndgmA+2mNG3Gb7x18XgnzRE
eeN6JKUCvFeXRKpSwn0JnJ1tBF9lpVLz5AOBdww+GUaGZFVraTRDUlzkFf982O0CQok1bX2SZBN1
jD6x4H9IrxcI1p1jrDE8Xp+1RTVVeASGl2VsA+jjyoMdzW44d89meNxEC1KO4HzvBA/KAgvO4BSa
ABvblKKZPcr9CAQqkdozt3nr0jEiNzJQUXAmxkldc9FihG7xLO9M6QZLyDdaRgHmSymfD/w6daXh
ZDLNbrnlkJCUZKOzNx+ju0CYO0/JOchXgAOyPE6MR7un0YnnO6aBalCyEpq+OS8lv7vsrvzgmmtD
/xrmc2JIKGP+hn6uqY1mYSIi2OqCDKfM04ePfu9tIFbv04p7HveWqB2K3zig2Z6TYFIzPYb4yauN
o+d/FyuDhdaQWqOfK4QRJ0tQxqKS6T1iSy3GmU84dtlGP7CJjGe2yWxRy4IkHup/NILPJ8AId5nD
IYShYSHhSOJcyVlJhoqUs0UhV33EGDbU5AntqkxRqZd1tX8Hpw8MopdFye0/PzwtMhixppOMcy79
fnZWV3V/PPWvLkqsQwGeMr98+bO3WeSM5euNMRuHpf6Iy7auQk1WITVl/TybaM8b4bEF71FXMhy3
6fQW+OqcjmzPLHFhkhzmYmXqQ3TdrrOxlv5nzwRtCvvfXrUq7REeDtPZqhYGakaUQxpSFuTLklEa
CJ/a1guGEJirbT2yjwHe1dmL8mB3gewlEvOEWP9W5kjf/i8l+dhy3qK2ynn1hIhDkMUpxYU4UrVG
EVSgx5h7S7cXxsU8jmN9FfN5Rz0ql1LLcyFD8+D2TA2pMfbTkw5yscx3lt7S/RSUpgM3Djpi44I3
dfd00MFjEH0GZ9fZgK/AAjILtRmlXOEwxyERskmcy78dz0krt1ztt3zHJs8xYSnfGUgXU5uN2izV
XYTjHauzkYPV/8b/FTkcco1QtcOAYfWcWrvHfBma19DDsL9LRM/ufA+U92guHY1E+bvSeA0fDTPA
h8+3+WPLj4XR5l9m2niQI4E3iSv4uxVoN+5fN3LhA5uREaUTEOsKKz7kH40q+7UUY5F/ZOPFPMlG
hBPyIQjlsZaL1XnOkwmF8xRBEyNu0TVfZW0dq3v2/MXagYzPelgvzhTTYVriqpTyhfXX32r4yLAN
ATeVuDemcxMvr/hcrFOy82YBYUkrbafdU/WL9TVEMsVilM279i82lTT0skcqF8IQC3ZmZ/P5LxMX
HT8nwvisq8+RvYbwzY6Z3B3SJ2kbHNh08mcMXr4pV5o9n0dKoMm/jW+uFYIsKy8nKgz8uXDFcg5m
GCaJqMYJut4Bo1jgYpu5YueT5zLP5pBy1rDq1/BSKCoqAdccFk7HOYDtHDBMxXGUyOcU/pFR2edg
wQbRb+cldtttx9bINQGUzzwFTxg2KAdKBKNHB5X0NnMuKWc4GKVJNvpL1wliimWj2JoLc5VTW5l+
ZR4phfdRJZPOCe1bDlzwsXvtL+hGqSlwcI+cGugsOkLnkwo3r/SJIDv+dx0FT3fqPuPKlH4VVECO
9hqZMh0EKVwbjCvDLtKj/dyJ7OWN3gCKGPGNdqAGLqurnDS5KWmgfdkyw20FfRk9fQJeeXoLu2Da
bp3EOqqUufdLonxu0eYaOz7MDIC/LVLIgGQjw9YMdXKIoEsJCLwPOPSsb7mdfUXEHrXnAnUJaoni
hHRngL6fJBrMMQp57ny9oPngH1d3t90RtfHqvOVMwVSbcDexGl048YNUX/GwAtncwBH/jEFt8uUd
BDoftXgVel59GEkY6DEVwBNhrJJ2CoPzd/cKA3vNSQwVXGD2M+W2RaFb6Uk8W8rH0A7L8gVdRswc
KY78Fktei3IyCrt2zfeeIOKU06RJUJJwflzpwqb0wG985UnvGoEZtQPtOizXY8t3GCOuOYQeCyun
ORSEPcXGjVu8NkOPyoSqAVgZBJVuaTmU5qma7M1buf3KBgWV+VOaiY5pHt6jGHWXlsZJwirACDHb
XMHySlimjq+QHHF9nMVCGboH+TwfDDsz031RoNtCHQK4VaHduzh1pek64I+2dl7bwUeZB3vT19Pf
sTh4Dc5+YIyad883Ad5sj5hvzUPffPjAZv34VFDbhz0oT9kTJkUwDXcvNuo51zpWsR7BQxoxrzou
In43Fv/vvc95gHb9lLSjIQRQQ5jRIOXL1JYS+e3R0YuqXf6tDN03woOjsSVtXL1ZM8i1XpVHi/VK
zsAn6WKKAwNORsvAlbdKo3B0jn14DGdIMPYS95q9BZykxQY/vZM+0CvGCy9TPnWptsb6i/lwPJKZ
pYCwHBjFfXir/S1InGroAiUYypuJc0ec8GI5Lfv/P3nn6ed9VoJbex+sj857T5EoOFjYnBme+8Xq
AgDd215sM4s8mzxTH+PZdJ+K8ZZgBTraHJc48Y6Ld/DFymmibUTdYMy2V7BCGX23QF2I62LzJhkz
7o+zJJ0O3jvBytLZ9EOzCti9fYLDoP+YagOkhlE/mPXy/zDc6FZ22LRkk6qDQB6NoYw859cRc0PP
/HIyQVbWQ3d6E6jYxnwZ4nm//fa3o+pRiRNtRyHqq/ZtHHvgHn1wXU/0UJynjWx/9PFHmXIurG4a
J5DH5aUqWLkMGppYA7jsG7BYZETRcvw6ySQi1oTFCpaONFnF2o882vlwLD50a2aTgZj/ural+5vF
T9nuQzV9pzEBtcceCqxxclRzIvuzg7Kp41t7CBP+Gw9wY9/TEnwk/9fCq718SXYUysE+OVpYUo1z
slPBuFJtnZXIItdsMFWAJfwJ0I13L+8JcerAlZHEgw+4D6lWu7+IuzqWl+g/mHyQvhPKeHdyE19r
ufF6BB6GRAJRwsIuntPDFzmytMC1FoTCjbIxJmqL/mmBCZyn1WYekTju7k8Oi9S/gRju3hIYwbhI
TxdkCS+27ALiV01I6mlqKMYDzrWcbuaNatR9ImL2nvsAVVrSV+yTY/9no9jGqxlUuku5U2OqCIb5
vP2oce2ijQlvt1246ST/ObXrlPxE9eVAiUrmp3j3gIW07VukdgMeeGAosQSvt0//mRd8+tLmbGGp
xyIwfJFNTPMdbkhdrW+RkSiItnWJBWehCTljAz0upyGeSnOOWogRRU2/vbNVazH9gr8Se7O5494m
/BhwqrevIW6UP9HGCC4bGykCiEnf4NblTLshD3rbMalAYitLXz7aMa2A5IGT137vjNJc3E35vG8u
cU/QJk4DNqyfwCLfjdgTP1rWmwCktw2YQSDeS3nEl3PWcXly/krOSd62UDipQ7nWdDsCSakJuciT
O4mznjJIg/Xc95btZpwyIeWmUHQbQWjvWqHwjRkAwQ57SOxkDrEmX25+7kStkaIUZfHtgDZR0og/
f7nMZMMkAFKRoaSZwizq1hraMyMYZAXwELZvDT6uYjZX3lna8enSp2mKyvf+rtqcHw0kpjlUSDAZ
pI+J/iSww2fCbPFdY6RkiD7+35qwvrJj7kqtf86NCY24BXiuU1Ex/Z0hNHFIaC2jSIzXqvfvJzD6
2pgVtJUzzyxI7YRk0dryJuT6r/XUuqEC48/M2sZILl77zGl0YPFJM5tm+Z9l2yNjHolxwOzuWmpQ
RPj6BwQ410hPbKumsKH76DuJgYbK8H9ELI8zbNK2ZVHKor2n2k0V61RoyrvvYPRjPKVM73STx147
drIvJbf1qtIgncd80g4x0BraXk3rHuswfQdqKYvsH1j5nm5QKhbA5INwhYTOTobR8ELBilU+RKkl
Y6NiNOPg2nDwpEHhhQgm9OWp1n5SO4FNumIN4fK0i4+28QOfPiCm+SgL8rg8BFI/JnhDNV46Cqd4
gX80bSoyMBFMbO3J8ZNDivQzw5qWMEeyXNfRrPwuEHLG364KBs1KDtZTZ5yS6GfOdVav88OU3LzC
euZmY3Sd2yCNV4qaQIDERdCFur3WLiGZPHgOOkgAe0JFSG8SbfpoLlET0kXL5TYEVV3Gl/SW03oT
6N9UXVsuR7a+K/Pop5qYKaGyV462CDm6oWC5Kyq34oIYhfbE6thUg7v26ImkYhVjWboB3xkdXtVc
7COgg9vYZknyxgZZxW/Cxfawg8kDiUktkKBIj2G9Wi65e8JhgzwR73mAZgbZl9buKPlmVxk981ID
huVoZ/o42JmVq5lCy0DXyHEz3oFdQKNA16A2/LSS8hW7uu1GscyyPNVT209+RA5s4RYFr+0KmWuH
FEEh7XdSl7t3Eb/L07AXqvIoXe6tuiXOG5HbtdYWXniy2exGxuJnW4SK8T0n+p6ZzAiM3XXGM7JP
iRi4pZqgpDwwlZ1hpq9B4ELZa4tBBMGDcmZ3ua4S+RSijxJb90kfGQir5ySAOdYxCA7eoLmyTVVy
KNszHGblYHChe7NC+ovY82QgEzMLqcIDbuRlJI63Ilj9sBEIAwpaFIde6mJldafkjPKVjfM7YCOi
Rz8MynMYbyng5l84WYa64bsOdME9VMqw9B32cURHs/0e0Vxey9gHojxFqu9z8SZ2OMzp9FOxc5XH
0K1gRKrduWD+MRwA+3Na4PzCyIsED/OVzEklPsSYlL7tCanrSN/RFbkVUre3/2Oz4PgUIRZ2WyRO
B2JnARHWsSFgLW0WAqZCgE85k2Ub8scHPauP3MyPOdwvoWiuXtPsi165EU0f/TfiVekZbdpC6R+2
jiF/lulI4CW+pDsM6FK30yFwDA6mRXrWQasfWYHAhJwX2ESPqd5thF7zmm/YOrGCYO/nRfzr3TMv
5x/Q8xSMTwoilImBrvDD2d+2xd69RDqRvbQtAL8YLvpHbmDxqtBFPXoD1N2fELQO8v3MwKD8DpE1
5zR7tceOLu3Gn2FCEU96/5iVcaNmHbeMeklf7cuykXZwjQ46b5l3Q9aADjwRpcuQqsiuX7Kf5a5+
vPq5hbKj0X/YrldnOZAmwp3GgZDXjh4iRGsmdkB7KZBPgVsFzlLuqLkpyWt0I48XILY9kuCjXQ9l
6EA0RSWhAfZq50FPh11lr2ik4fBk6i2ooiPeFeHCnmxdGf8KZKoaMyKhmKabjTpr0jMAOa9w4MPW
ClAgheVYmkoDzoJ+iFBhdXq4IyohDDvPf+uY6vsDvFtKxLTD2tWDFPl2D8xo9Z0kn/glBrnur5Ru
K1XfFGYGQJQW+Sq/Uvd+kDrUdfeX7I8Hpwi1brPd7Vr9JM6pKsFZG/lz5Tw8zoLI+gcihDh+5ack
URTSNZg/ovaNsJ482G/wdc2eX4e4wOlvrDb9q3CcX6d3S2oBswKu8txlPS68Sj0SvL7+6BO8poU0
6RMuLF5ZwnKDBSE7sMvp5Cl2kzarAhRxwBRo0D5RAi5K01OMKMA+sr2ybSAYjVHhNMIKCZBYBBfp
RXKIiTjHfGi4ZwO4Tv5js5EwtmqCakmXe3lejFbjvhOXcpMMGL4PCcpJ3KeVw+go44WCzuRBHo2d
iGmR6UUYkFfIBau+HFj8l76Q5mdD3wNEzq7Ooits15h4VZArgDWNMCRoZWhg4EOAUlf0bcTkSR0T
BseQmsQ7XSS+7bpeXWPDiziUdVQnkS9EoaEGZluaiqu/OjhIp1L6blNf6vTRa9EBYskOrXOwCP6c
j8aueKQZ2Vf34EpT+qdFqnb6aH9Sjf7f7UtlMzZzQFN1scxuUORh1NkAhZQG12b0lkJ4Bt5p58GM
kWdGVKc+4hQVZCTVVsYd2soCE5zknw8Mxpxppkjn3C9aj3CPzfjRpEOjQaCkUGV2Vv2u4Ez3KXg/
CqiLLX+36nnOuCeSDVNUaD+AyywB5MRp5ucr78/eT/cMjfE03sSw8liQh9XRaGOgBuWFKrRov95y
hHilRQ3tsFqhwEH3VUMTo262ezxfvsv2CV4D2yc/G/vuRo2r0pr5gxvFMYWp3g6KT/XNkiTfwdbq
KCDcQu1dlKIRC4eo70dpEYJ9IfiviPiUczpebse7wC2FM6XJh7gzGE1LDe9NyuWtQch+nmHntyKn
YpofdvbRmxJRcin+XAsPS/Qn0ntAhm1dB5alwqO5MmQtxe/3pJSC0aODx1yZKUjXHzsfVIB4hRTG
w05Hz4/IRScb8fxyccJ3kV/JshPGVNgxMW+5rWK7bB+Ju42bNcfGhg6rJSX2ljnrpy3WxGXZW4os
LcrC108LixVfzKaPUpUaF3PlZdDuNqx4ji0hfXJgl8GLJutaCcWDyvC2tavpHMa9tTke8BZ1jLcg
jlhO/jUNhyn55Hchs9/MNbvl8T82G7K5e62YkzGgVbaDGbR+vSs0oNVWCV3wt71pty4C7FIgbDiG
aa598n3WfpHN1M/FtkoM9A8Ahp8ghjdzmmj/gYAGq69YUaKTTzLEWDx8Wg/IkHkfuVJZLy1hNPYR
PASnpZ9PE7OnqEgYf2KTa5xJUuP+2Sw8J0hQ+cLnLwDiGpAg08QSYCVSBhresEIKy+CCJ9JqZFtY
d4FAR4PUt5kqnv6I0/oCQ9MYsqLFDyhJ68zlRzEvaTogXSfNszQMUytf1tHoGlj0s+M7b1zMiGH2
iq0JkASEwy5ftcsS7vQSNdVtEgyQhrzKrd9KlZhXD2B632HVEZDjWI9ojnm4y/6d7F2C+Mw8eRQG
creadGUxX6xIDEmCZ6c/SnM+K9q2X+1/E8gxaGW4F9d5RO4tR7NTAAEB730LFNl8GSJJ2L3EWq4N
x1j8zn4UdOeCKraG0uNhQsr7+XzTYvMgb2IR7x5vZqT47hjEBz5SUcH/NQuZKmZg7VcGNpN4arYK
hP4Ov0/fQH1zsu7d1RDjSetGWFziNM8Z5E1VlnTFxaBCnyazhHtvN0dzP83RPWzjg9+gVbLexGBG
H890+JzZgTfoRngt5V1a4nUTKvGNo6guoz1uzzkc5KzGiQ0RGHg92UBjG+TqHDkW90zjTBvD6rwg
ThQGnEv7zV9qMygUakF6RZ7JiSvY1h8HjnTQvFQPum0ZNE1g34MVERd0csE/n8qrWTYz/X37XX3W
f4wrB0j3Bp03Pan9e/AjWNasLFHkJchx75IPfb6BT/Wd+J1DA/IAD0xvcYEWuxlUPWKW9zlUKR5u
YQDjTgq9+xulNZTFPpwwNiMUFW5PkoeLsCvuDbVGRDDPWpi8QcEYYZwVX+2rOwm6lzRmEcQxjaV7
mfcXO7S2aJIWFCS3J3jdhQkeGYvRpR2FFIv7EduygAHUGzB6qppcmEDt0pmXqInDSzOUbA5cB1UT
TeYzDyG65rwB3qs8NPvdEq+cNxyffFAYvkk07BYiQ4r3ioGuYDH/g9v1ZZYH5E3J7LZqlDBBOcBv
US0tqQuWCRg4AK8RBhuyBmszgk/RHeYddPa6GWOWmEcBeHKLnGB0RVK3tK9uRgMn/nWlwzpuAdvG
d6D030TqcbEgvI6typ+S40sUVe7VhAcRqMiyEz/75mQkDZN6AT0iWYZWz4IbJbJ8f9+rgexkJ7//
Z8fBPqFsFZqV/PIvvwEXAgOJzau//JU3TxIdn3/+osdkVURwnzBRrIiiVxC1l99E4VhjtvmNSUt+
qKjl4fXY6/zDae/lWatUwRz5BBxb+r5Z+gZuR7euwDX792b6IlY6pD1sIEhurpB5HjFIqwpJPYQw
cX9DnfbQkmZbK9ByZTPJFiuLwgmv5O2cz3lJGIZ2vrdNR9eELn5ch7fGO+1inUrNG+UR7usRZeOj
QDT64szrcIfMo+WK1uMGM7HvwglRJtfnmR34YY2NVXnQOLY831/x3hAElkgOE4P+ILbLjusb5F/s
oj2rMsh9Ffjjilahh0iNewyPXHnPT8cPpJQDbmWFXEsAgXepC8UsMjRjBrXBNehuviot+FDLZh7K
ZSmnasIv2l/xCzDDBMURmzn8Ih8a1BaTUvjN5TKWzcd+Q/2xDszew0/hzcuSgaDFwHR322vTqXly
lL3qZ2Eq+jLOEB1Rn5SdJIJxVAYeETXUc1iuLqtzvDNC10gaRxbf8KvDm4g3LcCyIh0NG/QhpS4/
2P3uD4CAHu6njU8KFogi8dkPd961KC2ewPrDuPxQw7I7cYNWAJkBhXWEsBjZgUdDSP/PbgMEa6PN
NEQS6riXSl1qfm4obVuN4ggNBZyfN/UW8VxzMlwLtfo8kbvV0Q/nnwauFQ4iwhp5upOhdAEwvozK
3Qxa8y/NBQgpZZMddicWengcE3RTlwdtAMY5uq9TB0CvQZolOG4xUhoz8s1zxtlotWop3chbBcb0
g3aqWAvOX7CNx9FtdDupO7+3wl7qY508yElmxOQgIgnUG9VFiafUmPm4KxSDKsMD4bQi8SJduwMe
7uR4xBWAwhnoEMPnTa1Gv3oE7oUY9KinIbvYXFIWDL2oKAPK5HMkXVxuAyK1R8wxKgc50b0BsZmJ
m8Hvp4fLd2fItFeS2faC+86hGlAIaXVfEg3qEkvq7DrIoLGxEoIooMT9Uf41lPFkUInadQda7YB+
C/g1koTzv5V1kMey8XG/ZgBg14eG01NsQQhnN4ydq29V44Ll14aR4pHGDhZkGvfnI4DdyKLiHUJP
ygDytO5F5V00Kevd+0ggOu/KeNYfgkuLeJUinwNACV9BZszPtcIINQ8MHcgjob8iGoV123LGIt5C
iPGqNE4mmSm+uu5rS+JYfZwiBnk+sReBJC8S63RjmqJrT7+G2qnFOqBVbylHlTLCatWo1ifIQlZl
zhpGNweWY0o86/dbpY/XUo75WkLi7sz5aMKAwe/Bxrc4MOUlRwpP8BxRQyd3yZxoPSzdYbsXolmf
whSokbyJq8en8huKlzzfwjZLcfCtctoYIB/a5Awi0uJyGpkUlex3nUueXoqM84n/ws4qonlilCiO
aR0qAjUzrwAJ+sua2sHjBR++u/6wps0HXz6bQvGpt79sW5v6Ho3p8p/ZSZdWZ2r1lw/uD60CejsP
5drUhIXaM1o86sJZ8ahtR5iqf0e5mHErsINPnbKISfgWViOZ79ZlRFWj7mx/Ke4A7x7WK7ltA4dn
o+lxIvn22+0o1APuQFqbuOYAj4Ew3QxWkmbz3MeyidOnjRwCumRRVSPLH45BCQT1ckvj4V2WHYsa
Sf9dJG1nTlql3owaf9yhzXKMLfcJHngGR97NhUj73OtpJZ1GSyN1w/0hnZi1uKtPLvTVjVc3u+E4
Rn8iKWU13Gc60hQep0VlL+qndM9TZdeBqxLxPpRv62rjEGIBJOcctrgnHxJgqb2z+a4Hn2VILo4F
SwA/c9t29o8V8W8rkuf+P2I6GhFC2KSaURwGuYuV9kXYflcMeCEFNVdIcUmEXDgo0/3HFs9Bkaem
jdCGLEE+UNgScgBZk5d0UH348hHcUlI7SvTiD9wQW+XJSbVAFF0zmRLDB5sD7bJg26Dh6Y5nZS5n
PWMiFmrtru0L1F8/RgDK2sLgX687roBurw2+TwtftK95Nj5TkUXxwWgHXr3oJP8hu5AZzeVMsyMv
P1UJnBubQyGhiv9xEuArYts5lHC0w+HDf/0qXJBAhkXpsgk3H6VKRDlq9cXF/SWwCb0kQyNRcS5q
2CPWpfJJZizL8NqPlX/SbxNdAPMSxXfd2Xqe+JnDWYiBr3utGNllDbNAA7mhO0zkLZr3byBeaTQU
2DwEHNfJGoTEe9+21JRmKRa85qzXGg0dkPjhybvFtFjaeHImu0M0Ry8kswLUoJg8Rz2nn1g8FIYC
YoTnRKaUR47uGNemckRwrcUa7QuOpZLGx4W40r7e7PVIiHpJ6ljVcP7fCeoPplhKSgcO2vNQVUcG
vhgKA4fJv+WrxwX7MYvUofpDq8cm2pTfmgVjc1pFc4vAOQDPRWhehqobwNQaE0MiWvTb7fCKMOTC
IU4v6DLjp8AOBSeC96VZZbAoLKJ9MhbV9f35Xvun8bNU/LZ1BUH5WqgXXuhGYp8Rx60JdbZAZ0J0
1GbQbWMPbEGaz4rdmWKh8P3Wt7FwIak+s8FKtnJD+MrmO9lb+JS9O7auiCi4uU+3yNvIMBkF8pPy
Nq4eIxNcfIfrHZDKXjlQCuRcjTFMNBMYI9huOjj13vMg1ouvKrUdfwAUCImip/P7K0NEbTlRdKNr
h66XZEeDFvVQXPsApL4N6JKjtkN/t9DhUzBYZkHt6CwHdkn7nJxDSmFRaPy+LNAUqTW3z+30i/cI
gtM2aSMsAg2E0puVqcepDZpP1S63VGV7t5nJpiEkMhA+SyHgHoO/JmVRsggP6mJB5cDVU0PFsM8D
qdrxeDOuU7yP9mdlak6hiNKzX7LFCb23zu2enJG7pjZXw5/gzGaqNkPvk4ECI7WM6ko3rEUujWez
swa+kgZDIEyApTDcvhsyRLzcEDizfAQ/jMcTURHjfGqVssR2o8U2edNfLAHiMVwUCSEepG8aSAKr
r/9Bebf4rmw9jcFqRbhoJR30d/LGBBwczdMLq6I3OycAuMJcpJ9Fw2o6tgi+rb6wI5tz2y8Kw6To
tffcfwMgAWNGTQkdAUYoZ5OKV5wXw4UW0+RmFvnBGVCEIriVtudVmz0bWb9LvagaOZE0yi0O7XHy
HppLvAVVY1e+12ANwXC5PtJX9gW855aQfW1VSduzYJrRfUyVEmCSOkmWHQTQ42aMtvlpIvOisDpm
epoDZO7TuZamym4mjnoj3Rq90EuBdCsLUa2HOHv+oOH+Xk3hLk51paDBkg5NUJ94Y6ukBkv46SbK
j5JBznn0CnvdvT/hKzfMBSGYa8ruHCouneVzLzH6cZrilgXv+tiBcr/ZvDh1rRT6PR8BBEj30ljd
tPL/VeXxQ9W4wBs+2FTz0L+T5SS/zCCbZtMfbma7fJu6kXxLQ6QTBReRzHSKEDuuwZOg7SfXG9fy
92EkJKBKAnFx9sYtT/SdYAHFQae3cKYub48OGt3rclXLV5RZbOnwT0eQLbihSfIUDQftegYXdK/z
kSwIIUFHGyUpMvv4X7VMqxa468QDZp3/zmJdwj1SuvbJK3uN31rvh+/6QnHzLx/F98IsmKJuAa6z
1SpjpTWejEgHwGRUxJI0UqZYeF/IKIPrELQvS0fdUEg+z+vOBI7tkqrv3rbhxCQmwHWM8/u+poZM
FYELN8CXWawYHgXR5oAOlgwNw5pYNx5dYmnflPXNqi5esUX7R0cUKBKwDWj0/gWsqE+sVdhfjopP
gRFOl9XkI75jYkfCr053r8AImXE3AuuLPLdku7FovsE4fgDT4rAkLjWYbXPGG777iAGz1aHFp3da
ZRlPhzT5XKBOoQuZOkZB/Q9Ux9fhxE4/gRrGp1QaIkg0tK34xC4MJXymn8+v6mC3SYwkH3iY6nTA
TLH6cmfjqqIF30RQBhaKFjxczvCC+TkyeMBj3Y4IUa3MbP7TPCiz1eJ3Xyyoi17dGi92zGM+hgLy
U1xfyDKeoa5NE+GXYY5NqRlH48x7yOm5Z7uGahFkn8j5PeOP5t6KGljaJKAGmPagBdCdRr3QDOtq
4uRDXkNcLuQtlEV1KXTm9cM9mNne7aCq46dhUxEDvUZDP3LIG9YIhLDovEh8eVAiIPBYav0v0LsH
ScwWSfnHH6fSLLndCgKgDoyhYbVL9Q5iWYrh39f2sSplKZ0DNFVMlnRGnGFtYhXhYmx/XcnAH7M1
9UV79EAgWB3wElfC2rUvuRdDmav3kEgLOHlwQYngmmRARYePssa3x4rPfEn126jqX7Vw/LJ2/Cj0
QjZk5wOpxbQwje4O+BRxQMzn9eTcWD0lRukPzT/AMibf2NKhysZEQEZl4QLa/UW4fO58JxW1ntvT
p+yJxaWetbld4jj1dhzMOmClXW+pYtwOzmZj8pXkcRmGmVKWlJj/KKeTqaoIeMcbKLx5MLsTpPMG
jJiuC396nY6t3Z4/Jn73F6/Tkqaq9264Z6oMrurxukO0MxeYe5F20yG++cFqpxU8Vj0cyTkosqOq
I60qqCNrY6aMD+76hNsAAtMTBj8ktNPOnp8K3jjHSZ9xeqGICfuvtclCPYkCiQmcSCk0k9PVXogX
Ra9cIBH6PiNZTcDdTqVgAAnJK1l+qut4fhPAjEFxMh26j5YU5gPTadGIzBcsi8L88U8E/TR8ar8x
JAYIaUpQjm4WWCt0mtMnV7gn9kEm7FBHS7X5Qi2jmDupAtNsxob6tEneu4AjsZwUrqu7nT61wmgT
qUH1W97JW4uEUiUOAOP0/Vaxfl3qGaBzB+CAqcy/smSUvYh6zvlDQubPAr8QJyBAksvoF0bElvRX
XXbEH5OLJeih6xpafg7+bWlH587dZvPIUEC1UV5mwH2vcPtPXJKOqaKraqpDFDfMuxxbuNhjRoAu
bDJLtab9B+mBx9HQe5S47UXBKsGf1q1p9esEbpwia2LSNN9OFz0weyFzoJw5bTq5SxijtGUQEFAu
vPb52fJLzVr2X07ikwHPnq0FsdFu3RTAjeyeoLfqQiU/mmSYGMeKwyQyRn7Th3Z2ckzmW1aCsaYv
OawVX8FTz+w45yIIAxdg6eRH4B2ndl8Pr1AeyilmuMbo8U5Qt7i+if15fSbAOLFi93Vsfk735Q5H
yquzyTgRdUB5vGKpuX5UCzry1SmX6334NJPa3SWMdaszx5DCthRZAX6WfeA0h1PHz7UN+5HIGdbi
XG/p7k2Xgcf2qzXjtLxOf53FDCRKWE+Xopk8dF1prxBEA39bdu3WQWv2CCYcR6dq8h5wjr56Zgup
q26UUaVSgWfAeYqmKDz6GGg9XKTLtCrYqewoF6sXlK6SbhyGWtUCn30hiFva8MKUcWnvvBBmYv1w
TRiLkbBdcqjS82IQSWLMqXa+QdQce5W5BXsEJsObkdP5dkUZABFqMdf73AfDsanE/zm/PPUFse0P
k5zre5M4XlQ6IItbHuh34UX4cVIwCsSntKSlhSr18zsOuID32S3+sd4D+umbIWZ3haeTqxjaWsgW
M42U/pt03XyqF3jZewRGn0Avep6d2JDSvjJgPgfZYtXav74JiSsAyN6GznblyDKPFS1YcMwK27NW
pXr4bO/3C7ZdLNRsOn6PaXAdxsYcDBlfmBpAR+uSAkuKei2GItGib1GbqLCMLPPds22fLXocRiKe
ODspDc4zp0Hdjf7Q2uKTOUsJgDxNzBu5T5UQ77f/UDA9h/80xXAekfNeRenbf+MIRcD9d7jCc0Ic
eu1JmCR+O2WSRTJ4hrZIJFGYfB46p/IEbjbxIjR8S0KGxsB4aXueGb3SeXpzRnzNWUuKQ/vbV/CN
t1Mb2midRocoZSNETpe1pACnKt0lTY/HObPzc3xta0ZmmiElicPhWmYcIITNEMb3Na5kv8mzvg+K
wByhjrPK02B6Q9/YT/lP3u3+ROwK0pZkrnGQXqNFUOnr4qk+NIj+9HuFoTuKPaCoZWPSA0O+DOu9
3l5bGwSioL2nRVYlNH1v676HQfEo6yxN2LSNe2l9YMc/Rr5CP9bMqeYxsji9ofBmasv3wpB/cq+I
9z9xIwnWzHd2V5IgdgILRhbxOPs4zX8WlljZQMkq0eOnUkrFVKb7fTshAU/UgU2TJ5uIo0lZe7TV
jNwy4/+0ObytHHWSA9MTg+NXPcoEUjskDoA7eaeVS33LWLYCPGpaeyMlUzMPIBgPXu3msGgwMmif
VEQ8GTyOUaVxNOS6hJDNKkTB3esNX/G5q4ML1GdzwDDulNGquSWtZWoOBrJQ0UisiemdAWXlX1kO
KEl2NPtA4DCwJUuiYphWuVFJaJLxxtkz8DBjdU4KsrATsULrK07Qk5ttBkPFIDWPU9jEukrlDjQx
HdykrZ0vfJC91K6KQYkFfAxOTp+QBqcZ4BiIXhVRPtHmF92ECtCLOQHbHg3TRL3GCiMu50wBfYS6
EhUbNan1zBr9D9oihr+5Japs1u0U5sKBIleSGfowN7iGeiebAVZEay1ksp6fo6Sxw1tLiIExKt/z
KziPR8iEETcGbZCm5IRWCOeS7bkyH9neAzPqU7ELrUpVsxoIa0U6ztMjEcgB80MzNwpWk1Q18ahN
FdZnqpUnKuDjCjBK9LOQrL7RQySffn+XHzWg/gkTcssj/nL6lvMFfRZiX3Sv7UJmjnhWaSUFDh70
+Sk5zodbVjLVDBX7iZLREjA0XOxiA7nkUlaryauO2Ak+zCHJKcLg9eIJyx3PWPdbvzD7x/yB1yyQ
R78nRdts+ZCFzWSg6q//0mHN8Q21iiR04kbiBxPMAON4kjtk6pCOoolUooQcVv65avNR313Xdq+y
LcZFMCiFZYR0GaRtMqCFvHy/bP++wh1/gqzHZdsNRxO9D9fGBflAh3S7XP8fuHsmnp5OSbf5KPcN
jbSUDLplFdV85YOWiPNYrFDIWjrEVEo09a7P5QVzutsflf/ZR6sQMEZMduN42ghGEs+IZm2/bHnB
+8VPMS+zZRrSMAagwYbL7E5xeMxdpH2q+JIf8Md2/h0pDNhpH9DToaoOI33D8i23MwUcA/9lglmO
pYYPkYwyeR6dDYCU0tCg59WbwNzoE7voYEDIR3rIvyc6C24j9ZLpdxOxEYXLzxc5oHjN3t4Cu08A
lfCW7YlqD24QWJ+UG4DTDPtP3AQM/Qy0eCmxNUrYy2kGI9/aIaERU8Oz0WKgxgTHSyMjaWK1wITq
99prxOYyXrh+aBDnYekgbp6YQPpzV6x5hs6+2WLv+J0+VnoVNUl9qkuXsuP5LmhiWHNqB8lLTB4F
GdkOc1wcu3QFgTD1JbLQKerk/dr/9t0x/4SMrO3lDjhoUH55OIwdktBjxfjONtR+wahTibYDFjgL
Fh3tJTYYvHLa8vks3cvA7qtXc1p8CIz/oh/xpf+mbltBolFneK1NGsIvSMx3S3B8Ec8SnKQVQZkV
OG82Q6fzuKpDwj7emNjbYyORuFTPNSPpdcXuz1ArGAn+5QnEGg2iE1PWRvA/YP3KUMSiZkep6rEH
OUwH4NIZOkc1qgV9twfMxf9fyCgJbSpIfvVpXkVZvc8YV58/R9EH7rIT+gNpTG/Fa0asYR6esaC1
HpAPeO60pj9YmPa49QOenPmjX7q3EikVLerYRrxxSxG44HX+cckxHwBXkPxcBQcetUQD1rG/+4Fh
zOs3heoJyNicNKfYfQuLr7unhbYDJ0oNDSLek/TDn7pHUlD83OISJkv2TjoUGwgowiAOpWpNbF1B
0h6tVIKd7RXqeVP5JE63X+e0BIPOmEHV/GQ0uM4IXJRAfTIejqllk6NOt6ykxCs05Dq89vQXsA18
DgJAsLKtD3QOPG/jTjviMPxpV8/ii0vBdVtHfO222muM5rFTBXXdF02G0qCBA+8RaDVNq2LihGH0
Qq5HeXaz+agOr/0sA9j6hgH7NbtGPks8OFBSJSsIjxzsw+W7+zqp3Hto+RCMW4Z+o9al2sT8nfjE
9odnGQXVQuHMAiAY/nQuHbLW4Wu37J3f20GMOrcZKBFKNylXsDmw63D5ag44pG7eA6Klv6J7dhWu
d63hYTSQyn9OArgEswPLdQe1f2Y8mwmkS8uziTwOg6hhJfdCV53D3hass+LkPvytQ8FUm9YfG3go
7vDHU2xa7s2fXSXiFX50zOyAR9wRbLXt4ktf+UU82fPTOB+Rdv0FkypNX9RYl7f+sa7ByhVVkv1U
H+KSIuMM8IGWE9GMEWj+ZyKHpr47jrnBuz8Z2f7U295+6ivX5dst1YHEJJXoqar2miEioWKIk2oV
Zoc5oT2z+k6U0rIaCQOZ0UQJfl7q8i1SDKFJ2NY0Lhf7i4QTsZrE3TMAN9ub5hjI/gre9kwHwgna
OadWJ9GgOxX4QyrBYBwJe4C/SKL8pzAJo6dbELYSV8GEKHJeqpPHfNOiBhIBrGIyhnycdrJl1wE9
oMedQEYb6nGq14gNDBaQh/0JVyUqWJ5YbrKzt1mOY5Y7TIc3VxPdPKfcsP+57RmmwLlKLHJjKxUE
aTgUq7yzdeHEjaRZ2TCzOTP4TS9zUD4dyWowmrMbl3n64Kc1HCr6ez/71svHaUpT1suGdqJRGjrP
fZy09NKtqsFrIuSKusJzfXnsxZE6qP8a0LYKOU+hpy//5IrDVNSNyFCb8vYa0SMOTl0aqMq3UV16
H5ObUEou5rKS+Bv8O1pWPNAT/DNwb5CcQE3mq37pIFCoSOwsjWcGbI0frHtXWq17ZZMb4WyBfxcN
2nbzlkc/S41u7l52M4rvyUSw4NEJ2Nd+VSPr/W5d47pzWgRlD/B7WaXIPhyfEOn6jGS9uCP4e+qz
toMRDWMkfa/Ehg+en8L0OdFqc+GfQ8zX3IRtScYvUbgi4hE2NhTJrjerwBcCrSp5qmJ02bH6sJOx
623wRP6Ax1u40zTFTNB72A/81RECw0Wv1wNy/ofU8E1Fw83iYppVeFAP2fYmJoLcRjOo0/5smps5
ASd4iohtJUcO46ETldqTcvLkusCnSj30W03H08Sjoba/jbt8AZ879n+EsTUIVOELISuUQPfmeb9S
zcpoGKJO/ouQF85cuPVmFao0hFr44OY/he/lhH8x7aaWKoKC1nVMYcIVQiy2akvhDXDrt/yagTTi
zYLpWZxQebUxeQrT4/HxnM25I5Qf0TVe2xbbQCc5dpOZS+Ts229vpW5N+o70xoIxr6ONp10NwP/0
3D1dxsUwc6xsM3nBiFbTk9NKgoXMCJfr2vwfxIGIs2fgLzSI4BkkRGHit6jeXGBS/XCPTv//mdUw
5ppYLafyWnNFqFPkeOpL933ZZep78YVF12fSSymGIQ8qTjIe7/LLydo17K6d/cr9sazkIFkFEhcL
U8Q5LYX9QQrkX/kBDJ19Jsp5izvrJNHoyOP9ZuOpkEYb7XsotD6RGQNt6vEaQ9UHACvDHQKtXK0M
A+zV4ZSD0R9lBIInRddPdq3kYEbhU2dJFEWqxYB5siVQtZwIQeJxXoddSowi576C9uThzJUHN+52
RGB1XhTppKfAkamyoLX8D1RQeZipSZcgf2VThHeiTo5ZNiOJBwNmfYotu21TUky5k7wD2r4HJiDr
JZoLfB6h356ILFmAGnHbVfXqbKPNllueT1dPfpHGts89J67MDm6NN3EXyPTq5VDwqawQXOi5cY4z
Bds/8/rgnVlP6q00c+xz4PkU2/4CD9f/BgpxV16bPtekHORXCOMm7pB+5zCP33P1MdaYmm7s/b14
XW8DzmSrUGmXXFpAxwKP/6mK/5LO2fK76RkYDWV5nIauTmqqy/2fuuOlxRPB3Sbe5ViEO7DPG94H
X5y2e8SSKbF2xN0ryhYP4apOYiUpf4wD/0VDgMxbfw9qnDTI30x7OnDhvAuZxeqfpx+v8dfC4bIG
u8JVghZb9TGHt9IsY90mfMYdtKBP364T73BesDohMgL/R1orxk+O6BMGZ5LNnlwkUGNO+501KShc
vjMlrurv2FJCU0ZvEwrlhXpbLr4XWrlfa5u0RBFa9FcEK18hwIP0z/EKq2oWxwkAPstXRWjL5E4i
SRJ09wiRIVirwFJP8L9aKdhE91doJN6q65fChfdFncESS7nn6iiGg8frRKrjXNv4Z5vDa3mPaSlu
HhDridr4PLlXhUhDcYOMYWiiewR7ILgcQA8qodowlE5fbXpJu195CoPOUl9nl6OFiR78+jmwC0Eh
a4tvXqvQ7Z4J/lOu4PP3UZEzE3ePaf4lHkdbUYZiCnC0dXP+ah5I/e9kv9j6lidQB77HYVanDBAS
UWgRIuHF1dicW0OutaQd/LFEsaacPkQ+ngXQsVSsZY+90nWubdDatuygNF2Ub0e7JwZNKEhp60t0
P1F4DzhipwLnFvf2622I/33nGiZFMJPKXZMHY8ircx+u1G/xJEvkFh91DDGnBPUSdI7nQhLWvfWs
DOTEXbQA33u9RJVKPWP9r4pwGJVQeCb7N18pleXtWR471bpZFIwvuxRfqyFQ6AIjJ3kCW1mTLHKI
Sc/WG5J5TXeXP+6DZ2aZOb4tHoEGB3fNNLcuIQBFDDrKAuJ11Ez4ZiUsizD1OAaDKrfDTaLOnL0S
ST+gF0VyvllAiqDKpWTR9pm3sQeSkcq3h24CZRvPkHzgIIp7Z15Lv9LMQJtpHFmx2WjLSWzPDesh
Jk0ZrqnIq+PdQs5jEwXoW2XS2aCHUeAj6IGXWhEGUPhdQiTu3xH5DYPBUo0GlEkwAuybrz4oV+CF
F3/oGhv4MT+9YtGpkci22IjRPP0zeWljDWA1Jc2kp+pOHh2sTVsJtWmK7bcCn6vqLVwkfxGrFBLQ
1xHKz1lYx9ithl2GTU0uacq8FcDH5itwePFIgPo6amDVEYRnFFQ9HY2xG4DqpxQquVmPM8lKyo60
D3l2obfqV+djdjAbh6T/aeHkUj8GfWHlCAEx18zMgSVYzgDAIBrvKUgYNOBkXM7FrSoWXgZYjxlt
XfxGT2qum0AvBQgIyW7daVIYr/KUYfF/8rRWwfK0U2+n9KOiQdArhai2QpNjmaYT/q14V5zfQQFU
GkVgof3p04ETMNj+K9DYPCb+RQb7+nOJ2swByUmd7BRBt8ohOTZt+A+yrtD5BHwwMizwwXoxDokg
48sXJP79rDs5aPQkPQPzaOAyy7qjoSgjIh4GiehMMsmFyKZLvVJ6vR4MTCNBe8pesrmlQW1LqP+N
P2kSlccbUaRe5iBhnkRFUO80+l+HbCp4cdX7vthQzXWTxdRDd3//hbpEVa6APUBJv9sks4yf/1Yw
f9z383GiNUBQGUFtuGFGP0M6kdsQBsdnN8yfeE4EOq9uV6j568GO//ToTXPpsBx7KkmACSUPHMmk
S268pBEwbJ3p7SQpAuLMUqB1oD4ZS5q2gjrG7blVjoCMVA/N+ign3abwL4t5ypdM8Ev39OUVE93J
nsSFT3smGCvijFHr78vmtfU40PkbZKc8Z74NDvxfhVpF6fM9Oxu8GwyYd7JQv7rqy7O15egZ07Zi
PyiGEaOGt8GIHy1yuAKO//qksqaHYcsSmelWsF0Ka8upTWp58tqtsV6ONLmPcc+Y6r2fc1Cvg4vt
tZN2mUxxgjcU1nv4Og69PAvt87oGPETHTZm+1hY+3Sm5UES0wD7YjcOSCp3/A4q6CSluH5wyYxaF
3QJnMN0yBqJ5gSJH9+tYtt2qTKyaLGo3qNxsMGhKcGgcwnxL1tiIXRHFj1Zz7Pm++XebQ+D38vBl
iS/b6RzOR/IifGjmmTJfXIHITnzjW8OjLxAk86uabIIYusKQW2RDdvma0tXL2Q0cby2DQJZ80MIC
QTtjotH9yBb3u45Dg4UoBd2gQCExOjNBmgShRAIMYNSfvXcGdyqAPrW5TJVgz7Vc8LYnhYPoJXUT
BgpnhPkOgFBMgvi81TDDiaVn0K7sQSYfgwhan51GNEdEKAUZt2y7DwWuRLNnhPr0iIjqerzPkspj
CZcHAPM4iKfUWWF/hfntU2IKe8iAk+P1oHcaomNJxj5sljxi2xRTjJ3ZajUzp0TMDrQ82YalXSq+
IaDX1GpBx0MvtT6MZsyBLaxL8LdA2lwVuq0ZHauBvxU7ltsKONfiIGNGS540cicZKx4qAuWVzb5Y
uFagIucsCveMs2L5Eh41p/etc8l0bNedbOayyvYibjujpHW0FyvTUQ2TBp4A3d3NidQ+Z4jBoYtY
ze05Ejo9qFncXHlnVhiPZb2bdnFoWg4qlvLn17Ea5IK2MHDf5ugNyS4572gehIHB9v15OCenJk+2
x1TGtYUMdKXfSvqfQo1jjNk3sscUASHFQJAPRAb0DDIoDsF9WjY6yW6b/+/mACMEFf4RTuREkDjP
mS8sIQtCEeBNmDOmwLxFnE8wvHt6IKXL9ra2+FzuSdJF7aRbup9st9IIWeO4hIgk/CeKZpoNeE7j
+N3e7latUoZkNZBn01AftE9YRNJbqC6/zzu6gXpXJW6OXNlxwMmmlMMWYId1km95lh0nfYd/2Y9/
jtcrTNog31JTmjLoFAI+KAAK+tkudkuzb6b1v3ZXzg0ihA7iE3yBtmJpIL13eQr1g5oT8nfsO4To
SM5+N1gpEuTs0RvJg7ywauiYBCpbpNDi5Q8Wn1CO1fSlbiwN9BDMp/QLzPi3Ypic6kzfD+VMxDTV
eSPSnnxPYCCldpZEy9VOSknxEv+FFrszU4A8E9s6K7lvkJ1YGqopgLMTX/c2ZskSLjDcA9UKLP1+
QB72gRmGdwGnS6hLCe3S2uee/zvDJix+L+ASxrCBGFX35CwJOV39DBJ1EFLN0iK9Lzyr5dCFoP+o
82kpfyZQExuPDGRzOWFaPsIEWVH8B3O2wroeYTF7JgGTQJ37tHPeD3jHvzmoKxxbXcHrJfKGJ2E5
/s6BtkxMj+BfWG4bJCBTMJQjgdd/6EPUs8/hBEKsq05G2CmEGxbU51Los1eY99msAhY4lp51udOY
BLS02yW1uiwWRGMLs1CtX39vLKO513Uo/zQWjV+xS4ET4ItfxDcFfFiHCVqbOG/XMYy5azjtTiSS
B/lzvtgxdgEatWXIgl+nBc/ZJvIzTCSEcy6Z13z+6kUfi8oXFYKQhOfS6shRh2NREOuC4Z5h3T0L
19A4X7ww4gluNFxn/wWZoyypvJeeVfY8pCknlIkeesrMz69ZQbLvAFEV/6f8uZmtQtCyRH6BZb0s
QQYfmOIzj2MibA0A3b6GHxng+XL7mF4GCOT+v7RArYt5QAdZ/KeDiHaaQ3gUW1d8Ehi0vp+1soo6
ofobPLsRTptfOmZVyaOUDq6IFFLLUpwyXtj7Dcx0tkABdWCRINmXeUKC63HXBGhCQAYHyKj962B/
dAEDmy0hNLk16KI2mRwgywi+/SJe63qTjLlYEwIxYgVo9tcuZOMxftXSMBXzmEVTlqdITCsTjvvy
qbpjO6sM2j5wgUphEQu1v1+VykDjQS5p8KTeHCj53/OcxDIruomIMVmqN0ip4oqbx1A+5k8nHz1j
vSIiLQbar0YPQcb+CtY07jeCl86j575OmK/QOEWNjL/DNbfutgvHHlRQv3m/rsS99BaBgWtR5j43
KvEtKJIdF44LCeZYG3VlGSbi3E4aRZbA4xp9PUr8pb9OARflm+temjpNVT4dNYr0h4m/zXjUAKfy
0+2S3df9xjFbfU1Y3Ng5WtRhNflDQ9D0ID/fQ3l0YM69XJfE5sPvmOs7xuZ67VmX3kelzBMVmSh4
9qOfc4JpUyBtHjiTqFmqUUCA7waeNUb9I4AGW4Yez7qaq8pM8RYl6RA4H1KyvbvNGQpuehLNn4NZ
G/EoyPExJlBgBAq5EMJkrZf+PXoRUUuRc1CZlemTJIo0/iaVVbTw//KT1ClCAVYp4iD9VDFVRCCD
py++o4VbGCEjQuRiAxhjeIl7RIRYE4NF5csm4wV7Mr38mmSyqp5IErNa9V882SQ50QC83hwP1Bmz
KgOYn8j5gbShoOIeGlOw6cmBkeqQLErkC9Hpc1K85Fsej2pKv1BpMsEjwXe4gnRAhFMGIiZuS33E
olWY0CiZ2oUOekGKE8pIb7kEuyXhIPkv6kzH83RsLVMNdR6BYc8hBsVsQ7P8q362D6xFlNv/+cyz
4b9kWDLAJseskITgaoSOjEHEYgmiSWIp2fT+vH7wJuvhrmJF5NuCOlXpZwcarV7DfAYpWm+0DHAO
6kHlIuukxq/2rSLT1jnisHpVwuvByGITZOldfMk8MLjquov8XBpwqxXfEjp4tSBugqC7de9GUj2n
0JpnMWIkA/3bwaZ615ME1HLuZUtFL8T6lvKWNkWnYnx5+CjSxCbasLPfbSpioeHM5LK3Jve41kvx
Zw5OEHjK1ZttM1CsDuDu7zD1Anf4trcYWc8ZFQdk0cVzOR/nI/cHarFYl77nAuw99WGRpigV1J7B
fYNpOwc2aIC/Ah+o8uekdlJVwCgTPT1u2/zJjByRX1EN5qqL7dIpK93tUgYC5dggMbeGV8clgAyf
STfsqaFvvA9j5juLU8pSSDpOvqIXgC9Zem+YrgXiLTmwZcb6MwHFgGafu+f1QmjOKNZDeZ8qa4kM
ZwqZTDptAep2/U8mIlTOXg78xUVx/IbYP/+DTQ/heXAXQMpoCo+wA4rlAPQcqAttAfnf5cGsv9gw
RkIJDZzKv0ZGYXVm+RgMbSBQoCGNvKjPGdAScsNuBm2cdsy4u+mx/JgxHqQAmhYn/WID6oR1moOr
oJ/P0lrIoBguavi5rcdnEQwM8TKwnadJIzzUfiut2AOZb/Ifij8AHobWvPrFhkQmFTfIIijl9vcy
A/UgfNBHUuox4YqhxPzZfE8T6LCn63xVQ3/u9h327bSq5dqLuYaw4S1ua7Gi3nwEvVnEFkjsjfr3
zwLpvVaDhwPalKHrP2T2EXRKromC/+k9oR1zEIjDHl4UGvhUoHjjN8yUatgHBBr+2R/yr+5QlY6Q
oBh5p1xzvVq3EiFwoKQGD2LhvCIvPVpTY4JCAKXLNKNGViuX3Jd7cePFQq7QKl5YXb+zcp3Gn8cl
ZDfBU/kl+AvNqlGBlg8Dg4fjWa+CaSCQ77CFnKWeAFGBs9QXAJoi9/8HHet5zDeH2h3t+Fr1PSwK
8KgYyuLphSlv1Z0qYb+Pblh9bozC1XUjwf6YsbU627R5Rra8BVKHEzp/iwEFPuT3ys/aeAao+geh
WcCmnDPWhfLdUK1zWvHwKh9H973mkUnkw4UM2CRB3mnatLUHLRhsxL2XLZ56KbFO3SwmrRdYlmfo
pZCdnDiadn/vEMWcAFhQkIQiTuhYsFQqej6tvsgRkeM7SE3KLZvxt5LUNScWc1v4Kaw9RBcytvto
W3UHXpBL8GmMqLxB+uxXGbmNP68n3I8aRQa4SqECIvzoD7XJBFUGu1L56mcNF3X5nqVt8K6jgaeb
DbnfPT0hDG0xDgT104YBcagKB1K0bd+0Bi1sJUSvabg3Ea4egpxBiUMWNZhj091SEOkjL273+Wfp
S7v2ySHglzERGsmJIxQw2F7QPRa02EikwQ7G9WGJbSgZIXQoYDuKBntVCBrw9Jk9A/cM5WxL8eMe
sDYn7eWeHyA35uj4NowT0H6yGu/OcXiPRnWdvQvp/D7Youv159FP0PRpziuy2aO0oRMhuASefLrv
4V6JID4NDUexnB9i4Z4Go62EQqZY4i72V0qCN1unt4mO1y84ounwObUiuLphOh5l8mEcmUHm4UgG
sNSCh/2RAtNCtzAHooyyKal573f4J3TsdR5zTKPYN4vwjZu70F95BOxY++spDXezDcMNs9q7x8HU
zuo9KwkvyEGrLuUjG369fewggFLXqjCPvTRrMzeU8RZbs9x/knyguvJzOA288tH7Cxo2ayRuRGN1
5oC6Y5uk8+vvpu4Ww2/IrxTM5WDwdc5XkEty5qAFDmDmilmossUBoyXC7j3EXw/NzHkVfoLvbAhz
9c1JM4Lnwjm59mJEAPXoQZZbcKQEytDfsUq9/BY7Qd01Jj94Zs4CU+3ORUtiiykqHNTSm8F0PZcj
s3yZb4d1y1jRTlld2YPyccklTskgDCyhQ2Nau2DXnMGw6MINXB+Ex6Y4lR4q1Iww4UNDF5/ZEi9n
FFKTCsae3kFsbECsAUXDncm6cLKL0mG7nclCjiM4Bt2hOJONcNVBWpX6TlvH+SPeMFP1vrLflFMw
yWEGHkzX46E5ZlJLLXX+Z3t3rDJtFpGcTT78+98pwYTOgQbLwF+OnVYsNyd0c+dndM38l6fnbaP0
ZvUXaPjdBqzoyDQs+PwKwwsYhRhot+CIn9vG6v2DnnRDqkTOACWnDjo3v/rq30whgOeRqltn4BpJ
zd+nTEhn8j/uPdRpWSj+lcrru1Usag9lRXa4xdL0s7F98nUXv8RiknNahEuAcW+n8owqCkNeHpTP
6385KV7VRUp82WhGvSayFtMzShToLptNRHpwoxfENBAQG/fTjCxv5V1yKlLVpon5h7wqETpVk+Sy
j4d4Mvkt9+XLUhkW/n4iZrEz5gA8+URS1GntXDALkcqUoS4OX12Csni215VN/FKnzEd8gojcTtap
TIy2Huf62JWQxXNisJcgTVTKnY66EhCOHj+lcnU6EStiVWQ+Z6EHP77lH1vnS9VRuuVv+FqFtf1S
+NGpHv7Cjfrx86iQb2LLPTSeP9hZra6kqjMjDEUiLdTOL21mE2XWVQZHc0u0iopzE+m0GaT2GnuH
LpoR2Ln4dNBUCLZzolTJPyUmgAK/IxxKUpKcT6m8S6Yxf9KaCMKXgOYcW8J7Gbe0I9JHyV3fcUAk
aaf5TNAmGe+ou1b7G0cj5A6nuYZkEDYmMs3l7v6BJcnbIsDiXqyYweBdiM6sEUhHNm5cH9rPqCRe
ofpP9md9kMA4A/876/kvzhnfyzf7vFNCSxzMdEqDsJrzYk9jfJpLkxtKcBJ31BAwZ8bCVyttSZ8F
ScR0tQOEjY0NwcP47QjC+WmksnNqfoyySP/kCep7iH1fCvbQTxn6PkkYGsedqfJtFwgpyQgcxUaU
aaoxwgB/ULaG87y/3bSWGJ/yOvoWpQ02otuTTu/M7mhk268HkC/k2G9PFWdgqquUXle4fANYlyjp
ZmDU0mdygqEAYZ4M9+bLfYCz1UKrR2YT+1jZFUJ8WVI8vo5YLifU86TtuZsVStqhHxKVII+6sLMw
0dSrUgYmwEqlG8XHCBO1rB5WzGos/XLNOnQ9NGRKCo+BTnw6ml/ncKhrldv0t7/NeMnprRRFlmOh
QgBKrkXkz6sLY5sOnERSR6VEtQwmU1LebGgICWYOVxgVUKcwq4C+GlJ0G36RJbTriAE8Ek5Uk1/f
1kww6i471k8Om5QA5lIDBmkzNq7hNATqD/eNI5k/wphSCs9765De0XqiOLwg3Ax4L13u2hILyqGI
0SwFyz/RtnZmqk+gpCztEUld5pKLZ/J83l/MhYKrTkzsfRXe4bdBp/cQ83zPMeeqY3c8qWIJuc//
9X0YEPH8bTsl1Z2FhWbBznP5mTu/h4K/snLy4hKOQodI643asj0jXCS4anenRr1lXbFwKtj2kRwJ
GW+D3YwZ4vq73MDII5fRbwK6Ay6bsiEUrM5BStB1R7VhPPA2pgbuNATeL3QG7VHkj373TV3ok7MA
3UkdsOLqeM09pAHwFqhcJ3gDKgqxCjMpd9I8/dtP/QV/9fvhDT4IdOX0wp05Y7DP7QV7Q7HAXtr2
CS40DupPnCYLe4zbGHIdZ+aP+FdWcF1reSJUkPRxoTsFP5VTj9HZ1JQQODKHooJHSIcisRvsAhHh
y+Rgm6ADNoAnrQkNWLpFDiatonKH72N5GG08XTFJHDtBQw5GXa5o/cN4sP5UApbHDTqWbNY5m0dQ
8SAo6Z/dGHPAa3gnfHDrm1KtNefuuMR/dAUn5w4X1ZMUaBtbXzhC28it7h8gYmiT9mosoa2vueuX
3t39xt1u/KngGtPUdAucisAJw4glxu/XTh3WKB8662MZq3tULCHGj41RfZBzTBE9SsUWyjvOSMwD
UlEvF5BW2y/YTV8DiSRJP2Bi7s63FLqw4BH33TMRksPdyVxvsLUZJSj79XX1snRRTXFbR8uFQOdJ
iKYvuyWLApwfVimfomcdPFF+Qa+xOnB0Op6Ukpw5DWAStMfvH2lSdYl1NOZ7lDE5/+U3eO/EYgWG
xUvo+N59tlddf7toQAlrk2TWJUXlAfigB+IlWR0p55slUZHMQ12fLIuwLGC9bW8btKG1cljZK2hb
6rcwiyOhys8JbJ8mvbip7RGfJUeMYFANCdIjkk46CeR+pm2AQnwb4d4isEleD5iEhxHPLdVODxWC
Akshky0W3PsMVsFyP/gOte1QD6SdkbvcwDhX/k4JAq7T4JJmPY30r9Fe0fsJdHVgHfLofiSeZSj1
kONMjNliglh/OgiV4hLTN+PeJP5c4pOR1eKUKZ6Bv+Jbultbix494Kh7arVCFh5ruQ127KmVocvq
VcB8uyLzloHm6Tok8OlbEDaB9Dhvss8QPcb2uYdIBwa5bra5Ggf0Z8sEoRKGHn4eMGZW8VLStkSk
5afI9G4D4KXbY5PPDGZu3KZh6lL2hxGIa4RTapbRyDup6zVYWs3PLVsFAT47fxv/CvJDw44iqNSU
NBhYhSc6kiCLUJ1yQJm44o/I2PeGzo7KaY2kEw/TyWVNUXWEcwJp5lAjHl5TKauIM93sGqnJsAAJ
w/KGeRACJwSiMkAH9IktV6TI9aQpGMoAKashSZxQY4xMcmXeVO/BXz61q/KFXFsPKx9X2ro0iKK3
5mUjt0TyRMjWGVji2qstGaD2TQFw6J1WA3+LxviVwsX9PHdON0lhuUrRGFjuhw2UWiQjHJTqK+mN
E+e4pPJpbNSdd6ewSSN8N8C8iO1zLp5y27fymelTgtx14sMUmBT1UDtKWqMKvSQvmt+ga6lDnJEJ
AI1eqOP6F7fAMvA4Tupy1OS0xtiMMKWKWmU6Ac493xvur8zuyllTqMN/0Bld42ebIzRiU9sJeMG9
l2NAbgmsxhAJKQKBY18SOio5pnBNeJoH/GVGaX10h5MHD3PcZEIhZrk8HvvjPmEL8cXIBiUjWGwF
XWqX9IYTmYxz8Rmnwbif8tqaUbR4yVDfysYWJCvAiZk2WJtODebdLZueELqGaoMvB0pTsdmcQc6r
eBn3jhTlvfQkGvLStJ7M1d1UP5ULDCKLhcJU9Bvw8fBLV7GERBBWONhIl5X+EA0aEV8O2D//RAhM
31j/vUzDJQ6HsmL6ApBDIoWIKKdqiDBvezwqHm1xFHVjpYnKFyjf5UDgJMv06FRlyThFR884A1Wa
Qp7Y22GektJt75YaMm28R7CB7k06UH0y4hcWNGzSNmCJrGuHFy2KO1UwdZJKorfh5t3JvV/13D9F
lJkfAdADS8q/LmY29qjJ5Gd5Q1HJl0xqiwv+QOy+b932Wr+gzU65r843aLi3W+aWWU3WvGq1Nbhv
Gp5GMJ3R9i29EN8nMTyABmSGU/Dmw9FekxaItISJDSP3PmCtJ5BEXFswQxgoCk22CTM3/35C82kX
PlZNwCrcHPrkZN+2AaXjdNuMGU+f9h+A/6bPNbLBVQ5R0DFHqGhMvqKo0fG2v9jvzAZS5zs1DuHV
AU25EWatilalQrRyzQGdkfzsTtQmB4cUGsQOA5B3rumppGqro13aoG72VhIyA6gXaAg5aNagqpnj
06OOAdyH3W3CgIpix0Hq4kod9CqaXK4EMXXmsEo3x8BrIcgVf3yZRdwHRwZOyOc9U4mXrWtMT2zb
FpxBmqIpKQrjSPDvwYDf1+7Iu5Gu3SukEI7wSUPbABD0IJ4EP557ca6D7n8Y7nKQly6vX06YTc9H
h4KI8owZXlkTmpuNoYZnMiUJ1lRty7N0wrpjOFIkiCLEe6tTdHkjciblzN4MW0XCSG5wCXA9R5ll
ezev7XPDLYqpGxBRf6tFdbVN3nqozzBSC3UUV8AMFEKL2uIkaYih/K5osuL+mO0f4XRKRk7dcc+W
dYetEd86OlwPI4qOc21w0F4MtKPg0GngHLtNeXl/IeWSdHRXaDHWsW7NvEuiQ8YQ7+cWKiBFbz7+
rmnRsJCS2OnMpgmT32esxsS6fzLCqg6DykiUYuuCsSd88plFxkGM95a/bsHUZaZsviFCjYGlfnLn
6zTVOFU6n7h/Izz0S7QV9bmUhwjb9hc5up8o0yx9qlwuLwpoNdV5GnFhyo+29dCrU0L9sdwx8gCG
g5hWDfLgGIpk5htjAYHvR30cytDIoth2mSLaTX4deo5G5o486gLbB8ykehV3V8BaL13xfaXjah5x
Nv3k5ffDwCFLPDMuiL72uWvk5XZyGHjXQlNHJuGFT/NrQMRYNeKJmm586BGKV7PTO3KLJVQ49UcW
lED+YCu0KaIHvmZLtCVo9Hca5qVUFgjFYUwjS7yJWS1cpAYyAkKM3uBh/keCKDBK28NlCM1l9bQE
/+doZ/jF4DUtMlF9/lZJLjKeAy9EDf3nWnWyDY9rckFJ3Tkr+YGczllA5ymf+7fmAXWTQjr9VTus
w83dhInioFqKK/9k3bz6zpCsqzUl55lI4m2pLUJDIL4sJIGq58sL2WnxPrtmFuh0QWD1HCAB24Qc
cZ3RL78MduyCBOCS/7wx6qEwaI/ynwc5s1Uo2t1azxxW/m8xV7naZENNcNDf1cYdmhxcmtjSjC0I
/F5fm6wu8rBdvLqd801Lx50hAT0ln4GlnRZ8CfXjfl6qXpXHPWqn07xxfLdDJ9e8/cbV4qFP8vYn
nUocDRxtmjPT/h7dA51S3AYl8Q0gfjy56BXy+nugRYxzBJoY6+j4Wrgl2R9IQGWCvvLYhJ6vzXBj
pxk8kixuEAwNNYZhj92S9vO0FXYFcX/OYvrTfNyuHulbk0JqyE9g9mhQxyAfan9H2MQeR6SLqCtI
QmAgRUVIRlgk8vXtAZ2huRaD0nKMZwapw91iBFBC/2OwjL6sA4szFeveRkUZEHJ/5sy9/xQZjYv5
nj3+55fTQJiOXQko+2mmIHWvw3y/7QzTAz1XQg8tv4sKLVllrLITTU+8yOdWM1sj80wjRrvAZLoj
fLoQNKQ1YbqHVSbQEPa6YB7FscVFBysA9WPZ5DfjKHWW/3XuP7yngVrpZi5IZRgGW2Ess63xxSv9
3pw8uUKKZl96n1ABFUsx9kdju5xQMh1qdeRdEeqhZ8GD3a4ohiN0TocO15Nn4OkmvSawPV5tBHI5
QqaZ87mpROCqCzfQdnJj4WjYUqZ7NS7+Z/wIamLiGAwb3c7ndkCgx91mQb0m8rZEvveFUB8TSGg0
fWfM4vLFhpNbJ62QDSlIcsXpNLWPVXet1tVx6+ydRTS9xtyd9dsoKQoJlJKHGP01d94hXpTCZwaY
TuOzFcZd1cRD8zGVAo3rKQVhOhfe/R4p1hL9JG9xEovmSiB+5GM3sD5xEI5/dt6L2xRmrkuWHjjn
mjem6zE6NcQovGZKS6FS8sMNqGONsbk0koPpCmnk+QgQ6DOJo2lQTaOSnww0Dmje6FikTBKuOq6Z
x6wfm+Ex1Yr15lWZdPYYbypMo3P+gyXejYGkm7IA6DzmsYiASEL+YqTAFg2QEXOGSAw8Qa6objl9
BSweWdFPRaEqTouOS0JT4Or+Xd/UOqaN3pw7joAZ6xw6zbkWD42kRypZx3rDEkB/GGUbBQWzoDcv
S7aoIUjFGqrq3dcdPmjXEf07RuXJMkg3D1a1Ra/gNZVZPjHs9M1CS58xPkOlQVUwBsML5/DgWsku
fpdrChI17M4hGmL+rn+q9sl+7QbndoXgs0RemSaJ9RBMaQDlyL+XAbzEcy1x2PCB+SLOMpbAeB+d
KJmsu/y/o5rEHHZdKV2fzi8zliY/QDNeyZebL78msxPgndqn5exJpFbJ7E1/0OLAxXo3spqrufDS
EqrWlr9SI7T/mayk5n+4WBFcaXX/NAG6zkyx05NgMZPjevoifAlJq9/Ee+TFPUZHwDJv6tK3ziYh
3+qZ68kLx/NdcSQsJD2O2RvG8z4TvUN4zECXYWXMoiNIJw8dz/xMQkSIFZZRHD2z6bYnf/FEHhdQ
HTS0uUSKhpOcak4yAzoadrgJ1+EvuXyU1HAxdA9gpRB/VkeBYzTuqCeWxpbdNsBG49g61rx9eR6j
3c01jv+w2bciXTltUUppTDCCel4QUlHB033gq0gcw9uhyEjljWp5weE3trYTCk5YBE41gAmsTcFg
/n3n19FfYL8LnTt1LO3YXvAb/fSsA8JXdxjFxVLY4jhJJHYdfsHRq7c624ehRgiYF/03UIoa33qK
vdEfAzk4FV7p1GqsvLKtIGsWJ076I7DqR1bxAAROiCMRURv1Nh2mR0jHFt3lfCG2rDIj+cWX9Xec
Qu6R5mmGEbMiqcxuUILuzXYMwv0VDvx2zNAIO/Pekz8CWPUIy0dOXvqh40/EaubW1HmujmV9UxqN
l82KT0PSOODqV1qa0lL42INtSDRynYxuZYFwR9waSPqt/NiYxSQBfPm72ckj6dClECenS0tkm5Mv
TX5i/yKuIKHoW5cR/OMei9sjcXqvtR7hs+O09UK95JvDwd8qtfLSVcogvHYNBYvFP1iqBgUVCyxa
52kJpf07dvLVQGIpNnUgeoPW4gyjz+qOFFYWZ4N5tiTLXM+LyQw1rN1/rco+xfA+tK4k9i4pPrUh
rPhrL5nyti7cT3Ex2Emhfa2D6+1qPHf+UBR0ZWwWX5c1PUEZ7xKg7sH0ZXLvirVS62vNrJ4AtNfg
eqDGLpTq/LmSapXK4QQPVH4xR1AxVObME9i+KGp2Cdv0jAEj5jUdujENWVkjfKz8l0H/sKAfLc7s
O2VqGCWAhnXcOz+DUXTe9COLFJeYsRT7clwA/pUCbXqrBG/KGUTFd/RuwsevtlM/A5L8Xegtnk5E
phVhScqnl8clOoLc0AH4qU1Ge/ebdgPsFSns18oiJOgDQkwougHNqJLEfm99BvnYx7D3Vh7TEJzw
33VVMEBvrtjZzHAta2vRWu+Wr1o5MHLrt+ED9yPx2JYLQeMqy8qtqmHXsDP+HAzMqEVzN98vCTZZ
2/hGPv2uUaAHK/UGJluuGa20gg/9N+5n6Pb6Qal1Lgk4UmzKDOQyinj+wR5RuKVEdRb2mnkSZesH
eGEUcF2z0XjHG7FGriZUZ15DHWkRzQ2ApKL3YroEP3qy3eCUHam2J1gNHT4X1iqKyWc0CK8gPxCt
jy98Q+sTa2yC2GMVhvhur3sE0jbxucnQKIZJbctY1E31/U4yipVS+PPAh+eicAF0r85KBG9ZrGir
cMZuvYWnG0OHP8+UIKgs4qg6dVe0jsbbZb8PjOMzPhosWwpbk0KNNh9ZwWlrhap52f5Cz3ZvRzTI
pBlC4O5WiECzGd3GSR+xnld6PYv//gPlecSgeZ/eTYI6LYMUZdO+56aTMqrLVPZpNKSmLZ1xJibR
3SfqYCuFhe75VkqvNFw9rLDPNl9K/P3/hLF4+y9wXrwFRCTaFTuJcfvfPXE4/TeLHHMjt1Gevf5B
5BPL63zIHAjDpi5I9NSWMYPmjsI4bqen789bitNZ2L+Ydp/LZhR3DW7IOVfnef2VNIkEoE4vCg+i
drfqIcTYUrl6d+EpBC9kdmrfgWUehlDBi/tmy3PYquwb+mPbAkB0cIQ+D1fp1lvx3o7K+Q6VlD2d
WiB4knx6LhfAqH/waaNSAZyzHaAOy4N/njuoyfr5An3TygoN9BZq10IN39hD6dTo5cl/6m/qSGb+
2F2UNahwmcR1ndRUFeYruDpNezQ90fy1BztFl3DPrrCtMxbzb3x6O5j3QfbYOl4Ear55GofRn56Y
kVyBVlE7EvYnJ99y055B1YHp4elkofc04k7d4D86ij9VmXxTFtr14MrHtLxxYdH+EM9RMjnOksra
GpGH4Jk9JCFuKJoClHmApqOBAyFK1+dytFR0ejramx2t/q7TkkOwBIp6LvSN+9jwAKIwiAZxKMNK
NfD0hrVmC04OJOLdJ3Unyhiq7VWTHo7coo7vh9T8zl4TPOAQ8mitJLmwbnQaw0NaulMXmKhRIHiu
kXItyLfEguMp0gTvJ05yb+9JkZm1UD76l2ekdu7LjmiSvtTf8urV/nH/b5r6p+vE0dXgfESSDscb
u1kkDZeU2VGr5yX4Hj3erE8j3SD8Y/7XxArpVZV+LHAFcSYBLJoBUss8elMade5W8tRhC8AsXhLi
uwFqQjoAjGod/yBshDzn5+lz3xgNiuqNSDtwGSaHuPkttC3cyriKZO0VcD73hYT9w4LHKxXEQ4eS
z32L4E6KmdOmSDvTtW5ZJY285nQiddOGiYXn0r7Ycx9jymCqBh/paglx8YQWVyKdA2+kU9pv/3NN
dZdUgY/7AQMR+3pXCo/c2KaGw113Ho8GUUAkylV+nKWVVJGSYqB6gFm5QHwiRYtN3hRZCM5dTUWi
A4ZLa6LuLT1btrGl1uqoBhKMOGzak49y5sP+FPdineUNdQVg8akbxO6qE9XGmVqfoPF9PbxMc9cH
dfb0MuB2eKEgyDjE+VgeV8Aq/9R/rBqYjS2JX+ecZOmwYsGzAF5uYGfyy59daESXdH/dAYgGl0EF
C7ZWpLvt6fp2S38ysjwypyJ6/Fdshjz3YmyKkZ/apA5tbxngYpe7jV5q85NUh3v5oHIqObnBSXNL
J+6BVugo5hZ8yjr2QvebPg+3oB0nh/EMPF2ueGysZ+XB3fVOuKLpozlWnGkbzfVFxdYRYMz7o04R
JPTnr+Hg7ANGH+QrGJC5f1lX1+S1luN64GRMZ/+m4Nu90p8xDfth2hlqHx1m4ZYYwDDqaXm4nZ5k
UxUop2aOoTQFr52Y7VihfQPqO0tpSmNrPL1fB0QnaVpnk5mvLTnoY+cxTyDLgx4AnRjI4b+1veWE
TEhmSY7T9EgzLCS0Z3SwDP2c87mdQE60c8mCLsAU1y1cIDaQt9Y2EKH5mkQ39i3LfA4JuRaDuk1w
vb/Vo6ITayZ1WrX2MWjMUt4cp963M/t30crHI0gW7pOAzZGkGdxNjRW9a4qd/lbqkFnxYvar6oBa
kq3fkPhU7cNDOyOCFXqGkxIr8Okl6a0aSagAKMx1yfhlwfk45yA4EWldv9GBI5kJQckDyExMbxEd
CRQud5VW/+y0CWA7r672pwFuee/Y9z5Szi2vphSYPUkxbCWy60805VYoRME2Kx4zhMVYAT+TGcAn
B0rPRWmHvOnr2LdSX0BhEfyuiwcFKCpUvlVI7H2XfrNDT1zAzc6+A4OvQle2M1Xt1TaxzLBcfO2s
6r80xLByMtUTMJ79+vtHUbgAQXKb4GUj3DghX/J9eTI5ov4YYwrfB78cCiXauoXDmCLhhKUFbqXZ
V/4IeDgKniAHbMk0OmD9wwyF0QDFSxq9/rLPoOtL0iIro2auW/COnsNvsMbzzcFj3KZCoHuDinMD
UBXQs4gV/ioWMk7p55piOevfqMbWPLOz1UeLUBZqsMVZYXpCz3NbcaDwXxSlGYTJnifDQrXoAS3p
8s28lDNrrhBURN4dX6OlLVTCdmpmjcq3jhbZ6xuyFBo7LViHm4uSxVKCR4WfmwdmzIIAeUrli4vU
CaLuuijxzMcJ0hzRYVZjEc9o+Y5i3zL2oSFOSQZM2rJcqiEiDb3nP99sgPQV+JXumUVUubMZKmA9
oWUrQN+Hud32xRRapHp2Tm6MWFFeJPOKzqbS3oKPyPBRhyRc1XcTp5BGKkS+dLvvVd0/y4T1dPKL
oS73kGyKzUsct8u0dXkLC8rq8w5M8901LFfS23QZWbAXrt0+loai8mbMtTsSl7KhhbyewIFQeZHa
1n+bmQqszdClCkDBR6KhUUQmIkJlMDNacpt2yS6+pAjZ1j+LE7xAbMDit47Vn/0pK6IJuVn5d5tb
6815r2wGPW5ULLoNGyy6SWuZFp2mmvtqSXDgRiU9E4c3C9WbtrPjSoyXb/f0YK7Yj1kJGEibtGB3
SZh1OJXLvwZv3kVeyLYrvPlyT5Y/cdBMRRexIt62kBq9+P7gn4LYu2UHDAkeG5LM/qkyB6MU5a/E
KIcd+yn0WBJCECifWNqjr8G3eYpWdlNvnmxnA+8ccOF8sSqWnkqtogntUeRUexyfyAo6vuijswwf
yH93o16mOKKVeYA55dPkEd4ftm//4/pK2WbiVbgnv2lmN3xtYB5FtR20WxN9kqYqlrHptOc/BMn5
wR65XYN4wGz1peqvwTU4iMnkjgZMaskagIrEXGdNpXS0bC4aDpMXt63VZWLGx3/IvJ7hYiwASiWv
qKaCEPWSfudlOcbKwb+k3wCgBPN8Ws/Fh6ju4+7PHwzCjwCb9WgZKuI3yy/hXTheBgH68+YmUmkm
t3Nxjx8Mr0cNp9AT7k+27JtA13uLLzejZMv06AVU3LuoNJVewyk3r0bDTrA3xIM/zhof++D430nU
jLLumsPPJWM9jkergl6gPe+TNWoIAij4LOyFxqdPtZ6WCaGWjqKH4deOtPfsE58RzWJ2+Y7lx0Xi
uRjhnI1dKnFVxX3d9AOtrQ1qOfI6puYHG+70luvX7pTlAtXhUds3o875AQH46eH9+nw2rS86MD0q
Dqg0mr2xTg9bS9MlGaxZYsvLBwkxBTRSvjVftH+6vOGjxfdUj2t89vEfX7tlx2InPFQhoLYHzX4D
sdKXeWXEUQLSmPsms7bbkTe+xSi7khk/ATF0LQ6Bqo2B6+O1NqMNBJFM4VQ0aq3z3s7zNtOlSjQT
zWRzWjmK4kJ244b1sAe4WZhnRyIVPboP3JXrKVnWd0GRVwJ+NFcETjmp1KMFkaO95R93YNf8sGxo
WQYm+zH9SMn6vxCgdsTB58GBPatvkt1dNe94jco8dLPpYbCkFMnzEJJkq/TFNOQoY286qtp2FXTC
AU5/rU/w7WjldVmJ2nNmUX7uTq/ebls2wtNBB+NZnLjqrY1pQaWtYGEZvqFifkVaoeaxvfNEkdtG
9Mj0xwShfJd54cpSlM77fqHDx9L98UC8NZSXbymMG25cuRvFmCas2e14xWy/0ousdkig28Js9KJV
EsLJyktjdOr9UGssQVG6IQQVlZFQHAi8/TEpM3pMPMT5KBYldr87nrc9CwHDBM99BpawnFqQIcnX
Bc2LliozYP4kSzyZKsCmSmv6C3JmggpfV7JOcFcChfoO23jKjhwh63r2497wSLmqbBjGjQclLd2g
TaT8cwHkTBoSbD2moxEKdyGxtzG/fPqpUgrKKDXGd9yBs1+HsIvO+/q+i/7NTe/4oYZ6PE5HC8An
jLPhjKiCXixTug195MzOsJAI/Btup3S0z0ViIaXyP/22pwMWPOZUxbh1VKJ7SHsPA0H8QlYIT/W1
WCoXjFZEbzhR8ZvAvF9jaA4A4ySE3wusT4ZG+gSRJC5nPPWa0rQLgV3dHOZ12naV6APDVVHvdr6w
nT7B7OwdrnGl6yFm9jmCOqp2oi7Oc2O+DnYyTxPCV9Dy+o5OWWnHvo6BD44ipzU44YhYZ5/RAwK+
n/E3gBpYeL6FZBXfFNocF18k3JuvPN0BoTjbomxn6foSVYsA37owzYp09W2F2I/ExnfhkgUy2L+4
N+MbxMchfNnuMKabnWouwp9TM81nT7pFFwu3DUtOuj+EYaVOPMfNMor/uRF1oRzb3Cf2asTPvdCl
PPF/e3VDbw8YBTrBOv0hJFVkhKRos8QOia/ongEZ/pkjjfCn+TgKD8C6cC/JdshOIudGk8yaobpM
LM4DfNJnLTHcN4pMzeRpfAfYgtYmo6rr3Ov7EYmXm6CYkyIhzwI3mTEP9gqfWP/KIXu0aDjjD0VQ
6Cvy+Ihn0O6LjlJQivOCvkezvR0/wlp6oCh7y2UEZ4O18IZi5O97/INLN8Ybhqs6/pzHoebqtiF0
Y95LAYsHeAWzaRnpjNyavkQ1UWZbr1HSRATCZiDd+Am3Fg0IFU/mR12iLLBEv05Vd36Cuw1ZhKEp
TCbtNZqvQ0r7/iwbLcZW1hNRAKQ2Tmcc0ywaHd8QRhtc9ykhCnmfjZI34lVcVHORcS44U4c5rfiO
tCRoZMhTj6dx0fwtCKk/Qte9udo9R8aNqU+xkBouKCE/CkMjLamzwgqFoPa3Ie5OaWJIvog3uBck
YElEhW4fVmn1JqU0b9OIT5chk8wQUcu/OtJhcosRSggiwpQpLkRJTQZzv6bbAAh7yOWKyfrvM92x
8hjWlup6emau9SMIW9CKd+xN19ZxSjxHMGe/h+72UKJyrxbwj7XXwOGCo9P5vF9BDzBzyOkEv+FA
97nsLBFxWQDg7bhGmxABKzHYDthVbhKJUtQQ39NGR4W4cUBOGb8mH23DfnM9k/X2lPJJUhV6rzYP
2Idq6HX9d+1gXmG1+mjivxUubFYuAXrlPepXsVbh2OoZW7BDb0yhPCpl+KMFVcAnl+oyAiFvXeTt
fV9OdLJXUNe8vJ3yE5r7J03HNZIVUCovL40aNpSLtpJA5QP8VSRRJflk+A3z+n+XcAzjD+0uOOzz
SQN814FFvEcQVZEVOtW+gOstNSKVwMyflzAZH7k4Sy0LMAQ3bou869eIVLWh7Uy+tD9x4+z59kfQ
mLyxLMcLiTpDt7mVT1bEnYYcHAzDCcOZOsFuVskx0byVYsaN2uETcqEVXt9HduZTjMTrHO358/zw
xT3kRhfVwqV+xWhLEojsXPln0L2zxbyvONL0BFol0J4snNGU51z8wMUUA8Og8q38WA5QEoUD6LFl
1JFEZJe7ltGkc4tfR4ZgI5q+LfhN/4KQwqDMNgfETgLj6IXTMA1HjQaRDHMxpTBLeZbsC9+Mpd3S
FPSr0wlFD0Yq4FMOjH5QDMCYdBqMDdoVLC5vJgUp/vK3wdLKeq9Zn0tnjupeLWVjfHagiVH0ijvp
j/Twzc6YcI5ROp9hBVHzQ+t/2feEpOJyb30pDUFAnp0Fyg7GZ337BKSi2AuAQP79dNkEYa0bWAV7
S1kk/MiOUd7EPPXwtmDgJodBdTLZ66MLu04/xDzDvxRJJsyYqbzaPg2Ny5G+29npBtVCzKVTgUfr
OV0I++Vh4mOqAzulvWGAApTRSq6gVXvvxpG/aGOJSqefBoY59GU/S+/W76lmZuBl3KXDHuLX35To
+AFQWLznaJHxGnsw/tOnz+ZvoPoyh6sEwgcdMuUhXbhofPHz9Lqmg2FS2GBQ7fWdjbwSLBOCP5rt
PmvRhQlUVw4GWNfweQxNZFjjr+S+K3WEv5dznlaNtakYDGV8I6yvjLWC3K68GD9RUiEik90kOhFN
5BO90xFc5TfUKFAiw5BuPsYyQG1X2kkGnndSFZuf8KrwKNk1e6U3ogv4UP/4av2OS83VqeDpJHvj
6puB2Mew9bZ1ZK9XL4TFwM+F9zbfiv+UPFFGIVNYoXrHbWnHGf5ZLI6tFdLc+fhzzDo/iXSRmMa8
LTAFfKtjRU+qU9D6xtzx6H973ZycUYxfey9sZifBMMmMw4x6ywJ2ZDv3B15uKUJ8M9e+T5dXL9lh
eKM3hUPht1XdzNu9+JZCV7DXbul4Z6hUOtQmlTo7eq/9iB0JaZw9UikQ6cp1Jv2iY2Y+fOKfK1Y3
C9hQfDRVYJxDYApuqaMli/Z6LLn+qIzkVmEYxSx9CLxU8JhI4EuU5jrNNRO6zf0Idg0ZuzS8PjJt
PouvTwfOxoeWiPOFGb9OVeDg5Jo0x2OdqgHp1wXPBIwNnWmCpwWZS4l3zvPbukRztLz33C3iQ17g
CMItXlMvsgxFA9iiIivlfNpwooxqfogJxWRTUAwu7odRDdM6N07Of6z/152M7boCW8kcJbqyRDRj
n60hDsJ1cU82vwByPfoCdihL8Z1q8CftnMrJk4gkf03jlQNzLxMqNwvcDMgDSfIp2EnkGJPY04jW
KRPd2mo2j7+z2XPRf5cjz4bkH68Wi4YEE5r05cd4PeX6CUU93/P439SYmgpzugaQ2XjA4Age3hVM
8KZOOMs2jK6QesqRtpDPLQjYLR1jYiX+9R4pGe5cDjiWi9MdY+46o+dMQY21hFFHnWoAKBkvtxh/
4Cme/ONRoWp7yV7uT+B/RjAuiIqmrJXst9Hg1Q8PSBdpCbJq/sSinj57UXJcqEjMaYDXtyClz4g2
UhLJ7a92qYdoVdwK28V1TrbAbr5Ztash/SAvBlbnhRo+i5XN4CjG/ejR/7iE0G/BGGBk/6fWPOKd
AJfuGgF6Z54LVnifyn5rpyTTlcFrmcHryagxai58lUals290skdBCqeM5fpxUoF+vmh/NUmFsEAR
dFgw1idSdq10qG243IfPT/bNu2AKoIL6FfTUjD73KdLpqgP1P7s0aKrpvBehoUzce1KhvRe/bZX2
s/ZpcbynWz0czkBW+45OOKwgQwCSHj2Edd4FxSXBXIQSggLWWM1wB9B5dAX4rEMX7gh42XM060Gi
V2f9sTLXD/fBk6ydQ1pdeNfwMPanZe490EFpsxqiTNXoMHj39nem+bQ7xI6MFm9owvf8CuZ32OkV
lN9VftmdzlgJnehzgLPcllkXBWAQnPJ04AQaBF21zwiHUiiRy3p0r4VFg8N7njdPyFKfsJyovBG6
0db7BT2PPInyhFgnHYq8ul9zKw55PoXyU20WpEiuAB7Nx5CFPQEyKV/zKiQ/7qbV+1pfk9Ev5GXF
T4Al9k0sqwPKWxuRQtw4BcyF/W8kEPTlEWyqqOpHcH6tSz9VUg7mjtsJMJ6DXx/fjIH5JzNQ5zyZ
KdpIquDkauKWh7fp5iEXf305cSnWRRwCj7Kmk6VS1kVmog1B878bh2EcnI6SWWqYMil1nA7OWivt
e1lLpMoxJezFJNTEGUvMTQ128f50hKM1+VEQop7ZVKV07OXaniDbLWzuXsOGmE7WtnC+38rTC17/
VEzq1mvi2QGEhslk+AkYDR9ZLghSx2XUQZmkx9Ff/42a6xMlvEtMJ9yV+UgOGKuIblHgEASs0h1+
0luSRfIZ2yID4NiWUiBNZPNIOwUY63kSBTdi2zbtzs069N8JXiRXjVuCs+2Cnrgdlimncpq6P0gI
uABW33W0gj3/wxh/icrVwhwTgFNG7X6jO0yTl+/7QWBDy5+Q5/GWNIP/lsdOIsvxEv+FKPGdoYCx
W2OEOWgIWM+Sxsm0belVmAQQP2lxdD+gm4VDPdRJsuZDBE6WfAMOWB/HDMTPeRyqQ/kEdgK6M0jB
e4R3fB3TnVgLNDiDAGFWFPcSUiQ6RbdBtS1Vp2vC37gsYIcqsb96sKfp/48wI4Y/hIwG9DfqxDEP
PWZeJQOpmwQ6yJrVesfLtjA9v7qlbDoPB775T/unLUlswyzUwht1Kc7AfvS641svZfWqexVp5cR+
IIkfKi1zYsAu8u/5uwlqLxfsg2r5C3go2rmewyJdwLcJ7C5wwpuXJmDwPgaxsn3772It+IP/8dQb
rbGgvpuG5p9Bh5NA7nJp11+BKBscNsfzqbtqaoUWJ5aKqH6JItB1is+q7VRrz64KXClTvZqcOObj
IK1VkjzJ+8hdC3Ki7Zqfg6gAFkDcAdGFSW6kvYtavgb10gh5f/rosvqEVBshvAJ3BUnhCWTSEO+M
7p7PIdi3OPa1OKQHd+uw93osibaQAynKQRA2sBNVSe1HWwldYIEdhYkqgIE8k03nWwlk3b31tnQH
c00IETMP6mRT0iORqpfmjx621zooD8bTSmdEB/nldKOScS+VUHseQTazepkNT5FDatCwdKiI1AO9
bBTij43vLZ0glSGG7RTIIrKBvuV8q+kzTH/CvoD27eerwCMLsUtyqMuOwAeQSZu7mOsmZVTdOElv
LQK38QIYTHyYO4az7H/AbQOdELs7XQ8FnrCsEdjXLb5Y1lW8ncH1YegBtfkmKk8+QQ0Og60b21mR
wz+opOZU2LwHKQ5/OjjC/wVRT8WjuixKztvLbSpFJFT7wpv3a1doiuvN48UKE5VdYK8aEpRtfFZd
D3S4RCL+JzyHQ1fEHqu0yZNwAEmijMayOh/qGYAUXIdf9WuNdT/03bPehgpxdJ7j23x+ieM0MyD8
+JQ+hatNp+FFWv4cuDehTpO3mOMAP7OyQXFqWO5rlgOYaLsnQAeKxzp1dnvekMY5DEp2tLb9hqta
bQiLDvPKOnaODQSGwpIdO/LD7l+WGeptHHX6DJN6mefCdQggyMsHjOJURjPezqJlrMTh/KCF70lI
ZB++Lf+PV7AbMD6WGYG8C5c/m5z+zQ9a9VpIoMgYfyaGdp9v4qUE5QIY9IOU4rSDQVAiRO8jIS41
jYgIV25bO3xmKOzPDKCG33SfKljwyz5YyHC05LitXOAe3V7Z63zCkJj4UFYEj+kmkEq+55Zjy3wE
tHAclGKOow1NpD1y2+WHVNSU02FoqIFejdGQCMG6vimsCQ+IGM3ud9BBdlWjO3tHYP+bMsNjPf8c
o+HoCE06m9foU4jswD/SbYS2KPtYVLp88+tCkQ4//n37uIswGSMdS0k2+n22wzZifZKcGTBeEfg1
9RLvKGI2mxfanBa+kkp7A11MYewlqS6ES5KBvmyuh5HRLcfPvmtH0T12r4EZ8nsh8vFAe5b5QLrH
E8AhffAGirIE/3GGI/AoJ+6iqLQFi1IsC1nwUg6HUjBHDruuFwsQzRQhch0moNVbN8VgtNzSLjyp
bWfuEgWA6gIaNkaMZZ3K/LadYgbDEC+EwuN+tjjorrsRO6NJR55/E8P+llvFFZ1KX1VWjpSRQAFC
yLdBSmJ8O6cCiPgVLrqnsr7LVBSZwia2CZHpqvr34993oIUiO2s43HlV6AFlrdZbVDcEN7rMGdLg
l3sL3VBKFGEqlM4HGM9hbnnR9WacsNws1fGxi/DOA7u72gszcaudhfIFNUYLXPnysfAt4WTQbag6
FVjiCf/f2KC6j4jfXW/zptNLOlaPH0DzgY9xzx6n0ajOyDHGq6hvlRe0N+VrIFm3sZMuo1zv2U4O
jCQUgsY3eShdNw3TidQhYAOnU01bEHmLpVtDu9VgACZH0lvuRsdTtMIbqmtnZtiPARZ4lMQUJa+c
f9RT06XE00TuoaVMVhQmPdDFo5Jgh3APHlPyx63PcQRFEtpRN98vQGe6Q80RnQT1+OUZAfX3hf01
1632/CInsa2WJR4Gd1JPgdWSnBj8afSwy7El7Ahjhn0SsZvF39oQWVAQD0cWz4OfKz0DKOHJYmbq
sM8JDkUXuNHpvnYH+ZszhzK0aGB4RRErQuRl0gDYhKs7KNq+7YII6JpgkSyjnO/OjTcHURimfly2
Zuk6TbLp43gz/ndgMaDxEWbWYcKz+z/IlSKPYweM6IvK1T1oCHx1xvzg0YBQDOKNL0zyVwjWvLRd
psqv8jq+ADU07uLLT4U3dQT/Ppw4sNy0hQvJ3+WU4pfi5WupRRbS9k+RrJ6TvnuiUqTs8iRWKNg0
eKManVx1EuBC3sI6TVPa7V5NjHnsFqWx3AOglCFJmvXPLCtPvVk06AzC8ggsweW43qw0bwq+SVj1
J/3tTQt8jHRK1pGawc3rF3CqcGHDcMKhi4UAJnLR//bmIL0FfXFAx2xA9gSk3qzPIJ94jiEUGJJe
DIMIA6ajW8VkqBtuLg7bvSR3MtZV86Ga7LZnfXzhTvAx13TMo/u5Xo2fOAj6QyqGuyNSYoGzAjTV
drwyOApX5hE32FhVwVcxiO1UGnxbU7mXJW8yJQhpeXnvfSTHuodmfdBq9xJb3bsTrgaP+yNfansX
SM1zxduMk2b8z88FEMXbd6qhLB+9N5wReHQctaGVIQoF9KyCOP68GbTDHrFeacAZCwwCjADx14Nc
aDnWN9jGRA37bgeWtHi2uU0Olw4qMflnKm45fMudEo2aVn8QyJaVD+cxl6f5eLDBzUZnjKnmw8Mv
WR0jdPkgfNhueZk+ktoDv4xyyBwSfHoKTP9qCaS4UEM/WA4bCVMy+vRbcefuvc3gfQ2Dk2IdxRVn
E3D/FbgZq0AobM0TnWZ2Mu/E+eqlfPgcRR8Y93RDLn1sr55nP+3k9C06a6dYEg1AviYj+fyJs3Uf
GksdM8iQ0ptE1O+GDm21KVfmDbETJtGYdPchdxyu9WsNK+l9f3yWmI7GT4lfCX+QeT73RujEbRfN
WmQXfCxQDAokXLB1jFl7MLo9Zpe4UKzPBHiuQsBVhAcG34p+fGXIrpO0sfb4/RwDcsQOhGo9kxQ5
T4civas1MMZFWNH1KZU0n789wxsXSfMkLDIFik50ybE3EI6oZnZQBVAZNkPl36SX2vn9hdL6H5fL
6OFHhmerheA2O2L4gbucae6Idmezgv2NA9XkE47AsKsTPEHJ/e2bxO3VSsDeHzNhmf2wLBH3zm1a
Bx69op1RDhELcBsjVDyPekggxKn7AXQ9GLLPXu1d8rlGt+ocMuWNX9uD4XRGN8Q4nMgKtlXCRvKA
3l/XWYlNWFxqlbu1uL7MiXIIsZfhf6M/xqDlb6oODkbRp4eY9pAAe0zs3vKu7/JY/7v/D6uB0wur
AVwoA4QdvcK6RyikLtkg3px44wmm2LM87I72d6KAO4Wh3xlvMTqaHJGIE/n1nxPxSFHasbqrfqa0
KzzG3tpBhF+XMPaEzu0mD2iP07/cQMcW9yedIcnIuVzXBOBGDKYXd//gVBj2b0OzUdKjmVcnNu7c
WQK4y5fyQA0IIT2LCgXxVyvpkQx8EETZ6ITqD8O4QKVG3hAnTN3vS8HE0H2I8RPKSsjpAx8hDbzz
zYslIkgvwmU1gtmXUbOMZipKRUrNah5VqhCKCHOvx9MSjdrR91kGexkxGxt4mckaSJoEfUkQ1R66
BUCHouKc5GFQ/PtK8sujMUeukOx7/WJTBDqvjGjmmNS1QaK1pf8QIiI0sETealOijbVrmFKyAB0D
jyWq8+dFGGfKZ451ZWgplXQZDr8bDemNt7uXY5JBBxUsj69WxxDMuLM9SiBduOdhLu2TRVsufIBS
q5D2N0axcJHTtX7IOYK24e0Ws6Xf8IYuKxqtE5+VAJuFzwhqXlpCNHuXweZ7Pnn+ZmpH58qNyjiC
D3Qj6h6uPOJh/fzOAZgxmlasEI7QOEokRuRXdR6Q4HeTeONXW/kO+QC/C/iXMS+bVMGyKiDJVl5y
p2ysJsZLs5upcv/+mf+vhZCsxS0/jyR/JKKu9l+h+2AvxDIWw+0sZ/xDj3cc5Al5fIw8z/7VZyOk
gVFR3U0fN2p0GGgFh5oz9ihjGXgncqV4cVlQxH/VgKxYxJhCr1KaJYw1I0FwsIlmIyV/COHlr3Nv
q5pP20m1S2I+Sg1kJ01bhKMsZReZy+rAtZwBAc/FdlVZfGgO+lQVzXo2w1wLgUdXLlKwkCVuRRYt
GUbHPWxJOcHRElJOAStgEVHI7snq6oE7ib9nQlk1XaeOBxymDBtBGjYHI05saueGYyDOSxdZpSVG
QRSAxXzV1A0y6+o3g0zO4XXkgwj/DtIbZNgGMjq2GZSXu1hhHaxzsIq50woL+cwqZFGxqXrrOEsa
05kmCuD/3c+4h2xjGHrMFcIoKazy8VRWeOPe9ZQzJCanY6NBrVyoH48fO77JxnsajkVCYTHJG92u
4DE5Yq+8KQH//pkUSASAp7pFznuZTmL0RSoY4tlHyjg3u8rePOwY5Hv3kjZ1+xtkbWGdPkIkC3r5
0VNEFOkAugAhusiXrzlDFQaLwc4gCpfsJrFJ71LOXpzlE1U0+lMyRuRhw58LHRl7zRaz3Qktctms
Xi+Zu5j1zN770j9TmGDN6B+y+fIuH2MNasGtobEygttLuNi7V7mTN8622aLbYHP5fQcrzjm30jMA
L8RN7aB68bg024S5mO47E6BM50haNg/+9B9aUc6XykVJcoYNBKmA8xEPBp5DuLtDcFFcIjzLGF3H
8gJT/31njJMj0kw/5jsRUOVFKa6/ltrTu37+lVK15yG0+DkQrBM8ZpKRGJGgOx5yCW31NFem15Vr
P3xw8cFFR9td/RukUp+PXOLzaGcv7TeFVShcYbYDFSHj1Mq+QhWDs1ggKUox3HDMOeDIuej7wTHC
Z6AbWFXEzH+ZN6z3tX+EXQSRBshkCddRGvASwvGb2fr+g89WXE28lxinGJ6pkRBg7jTvt7VXcZgD
zwK/Eiwi4E5y9dSfvRm32Q66EpL2Xy/ibXlFTgE/lYUzZVEekhdVx5P4E2mF82Wdry3OhU4Gyoox
/4S10nKTnu3Pbn2NX3zeOh1L7PLJnToGf6vT/C23fuUHWOmgX93Cz4s7raGgt6QrIlke7gNuuP3T
Fwu1dZASyp4lupOT8uvv6iezn0Az/9O5ipMzwUXh+KnZq5xPm12VIXl7AEYElOgQ0EO7Djou0oYk
rZkR0bwzPr5/CcYyDew627ZUMs4rKK07VDPqinJD2CP3oZvZeDcdxWP7J15yiBNcQsJUh0he+RcW
8uQiaLaT+9Af/UfPQHDqHP7Aacnk+xLlt54gS+aHMaJ8+0kepb2h1ufxAuxSbApjHHapLP+YCg8t
4BBjgsxw0H8pczKirzfe0oTfndSVZLO+dczbSFH5vVUMBDxD91U+lCiMRWrL2lX/9EAeHX9BOSZd
q8T3UXwYefbpgy+E8Q0sN6pX23npGBM2VJgQ3iBtTjnidt0ItgwGYl7gsF1husjxFa2pSZBKKeII
Op2caqilbAo2JA2WYWIPsqsNmHSVAxTH2d0XrU/ThbPXCcGYvfFyeM3QoXIilYEsQCBWZbcaLrkZ
oHYc87haCNawkeaO8kNcHPqdinuf1jI9WRXU6/A1BPbeCwWIw1j/WDhzkw8DqNm0Cv+CHnstcwiK
zIWGjMjGcsau8glOfJ+0d5l2F7je3goh3MEFr/rXGBN5jHmYwDjoU4W51B8P5If0A+jOdkqiD5PR
T04PMUoN2uPP6eEra+dp/u6LYz7aPRETngxvohDRbaP0s4JkgZSSZiuuj+kzAYbMdRYyvVbaRGDt
44RVmxK3jnR2JMxfBQC2j0DXzA0Q3b8TQUkOKL+PFs2/DRGq5k0eJkzU7KN0enh/MeMrHt9t5JHx
O+NUymREI0/O0fKCWtm/G0e/kvOEXUCrUcnkSZfE8vqHXtcJlKh0OXMWZWGGvPHUV+fjjFMuI81k
MOFw7IWnCOrI1JXK8hENLpOTLVIbqx4HK7OTTnv5nMMWvQ3UeUWFLknycg==
`protect end_protected
