`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oYYUZ0MeKqJUJoI7DJiuvSB+q5Ix+Iwj9N3EwG3d9aznfrZuw1+Fc2PVy4cVNiksbh9EhD023m7N
/1rZI7UBsA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BmgMGlUziZwp4Aeom40PM0gFb+Lk4HIg7NJ8Ke6/iR/nzJgqwxvBOYZHlsOO/Hp8XOgAeNb9Zd4o
mPFcvStSgKrLqxBJrTC4jOtTOOUVOGECik9X7RElVDiKeZuCTuuYfKks1rnTANMNKsXOPeJj6Svr
YyXA9D2NRP6YkUNuPRY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1jtnTjcMZBAylJ3gewlkrSdkM4rrC/SF7w+2Gpl8C9SK/D8Tzq+D0qrZVMnmX2MWMKbqqYu6bkIj
sy7Xox+kttnLUyhBRsrBNs6gr3T0xsxsJ7Gnyco/P3Bde80gstdJ+PNfjg9uJOXa0R4ym9WtfNGf
swawtPDRNO3XB4oPqX/YBORxc12Z2+Xzlc5kJQDf1WM1UoKUm0j7+JBzjmig2WrmokL853BM29jT
4Ht91JL1B2bOy9A+fEpZnVLxL5NzuQ9svrSJluHfL94vaMxePXlPq6InH4B+XQp0TAFlIitjElNz
4mBAF7U6zb9GPz8ite7f9+Ofg2sCbTc7qhRaHA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gQeqr96ZiBT2MmGHCpbhB9Ma/ONapmaS0FJH16GFlg7E/VRDUjqbqiiC9oovpVsOBnNDQZNmXNgv
dI/YoLxA/mPd3NXizDTj33SvvwJdHC+sPFJrC6pT5rNUHqY3WkLW4EktYj3xtwACazlM0R3H+N1W
ZL2jtTv4hCIZZw83DISHIwGMevxP0unAXWFpAlJTyOmzC5wsjnlwvjA6I18++KC1ECVIFCC+grSL
XEAA1xdZCU131f12m2UaGi1yGaQH3scoEe37TXsoGUkWCMAn3jD7PddNt1X5zhoSRxPsOfUDmtSO
kCNVtrnPznMY8kVS/SdMToJlnwH2sKbHJZ6YoQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aYbz66wynlNa4RYsWnE11uoqAUkMOGD1rK3oC0qHnHAmOdMhPdz4cV/CAQENwbN3ryQY7/k4qEBR
2l3bOqYxA0+CBRl+jt8CXXxWU8WE2qwf32lPVes4/pVAbKANmE02/Ysj4IR7MGLvUvtr934XOsBK
cCc/KqvEbWgnnzkEdl16nzyz9Je6iY7Ni836+/z9BA/OYPszoNI5lKgO/06ni9esrcL9aCuvKXjM
Vplsu70i86fjOGURYjM2YFmCk8Xng1M6ROF+0KD+TufNMvK1W5if6MPJr/BsB83OF/hzcDKyULpB
p2+Eliq8StuhC0n7jUXEo6ZGATEY2a8DWEYVhQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B8e2xR5DNyjb6SEEOPCOnfB9/yUC8O8izWpzVz5s4/hfcHkvr1SHS13gqMQDj1DN3uSpaoGxcSIv
a3uLHDL4nIDztAAEPOvl5rp/eCLKhGUauWJKGzgIaInIPCBXw0hsptiyzlIicQEO3rsxoS+LR4e9
ltN4asLfvR5i5+Aru5E=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o08P3wLx4KXr1Q02DiaLH2vPxf0H1jXIwF3rbwsiMxYgYGWIJGF4/mxUFC7J/WeIjcsQFoTUns3o
ZlNZWWRR36HJ1r2GmZoMunV8HAWjNjCUrk6RBWvB/4dYllizQVzRhb+3YUjmiSEMr4rkGsWsR9/t
W+i6luLQskwMDbMnn7puINFUehSDaOzDytgvFigNs9cj7haJi7XjPeMPUBa/JbbTJGFnxz8xzl03
55+BSHF5m9JHUn2eN7uDkExSgYolpcYI1EQnoCH8U6Zfcweg7A+n5SfklkTKUeWInYHoz9tHbIHA
y9aJwNoT7f6uxEt4GVf7oKjEfFlxUe/yajXHuw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
Vz8zyaOyF+PVAq6J1AOcHrVAt1M1YJbx95XHSKFiCMdQXX7pmw7z7zZFhgFzILMu0vZYFHxSGbO/
0tsnpt/XvOaUYOlqq9OeVNgUYwow2PnoEWn7N4Xq8OMq11dVK0uEE2B1Fa3LbYoCjuvrLyBK79rW
1rwrg2tpQ2PTnjF6OXXpWRowLVU+bZ/egH0AP4tTimjEEIe76UO/RUzH3d5oxwwdxbN/ubWfx6DA
Lk2yp3auZ+Y9kKFpWKBFHIIROq0gt/M6+78n5aswEHoXVr0sJ7w28z/rcIrZrk1Bpywtm9XfbTD+
3NbRkv+cUSumvTLan5vXDBGKsrICgw4FQwOFqoTvwok1W8YgIFH6wWHqFvwlNhssnN4+hHj04F2X
2iRpkO7YZ/2r6zbfPj3WiQDqnmYM8/+n0rgVpYR3Q9/TECQbPS9RmlYTYgOAnljDXdEmZEtX2ZXo
C1WQmvnLmxGX00UcAhP18pzhh/uTy5MV7yCZkfsyKqBMleKFW5ht7eSaPhQ5qInXMnpNKe/nEhV+
VLlc5uiz/kxcYWo0/8elkSoMICNzlorcMLIAJC+ncLmKNU+w3Ti1ByZEBAlpV7z5lP/DScQFpJpm
vhwsm+o4ZSiotwXlYdqf0OOz2p8eWSGBb8ZHy/+dp9XVH1+dYxAT6ernZzooNge09Wr+vgkq/3ai
yNyD5l75mcxiUjHmbxpBy4DaJotokZhoDh/v9ICNLfUsz5sZd/UDMs7qXgN8aJodlOPG3xNJrLmf
iX7EnnCa5RBeOac1gxxhmyOMnzuBC6GhGAjE2Wxa9MdEckTze0ScExQeRrckQgANhDlFNh4ceVqG
4X9XqrnDEdIfHy9vF8daIaFB+mgygMLAL7S3fTaI10DK8piNMGfN3QQHgKOOmBzxUq2I16fSacPq
AvX3zLWOWAxNixBzZK/5xxk4uRoI6tnsBhRtmCp8VefM6GKCI6Cg6PpIuW2h7bjMSSYjYisUop32
HbD0pLXddxL+r5Vz9j41bXa/ExzLWOwJQFnLbfl54QHlJGOW62zuMDBgd1AN3ntPmZa4RkbNvLy8
m8MYKEBHxgEKTe59Bk3S7J9smZQhaCsYHiHUxgoO3uucgnns4ouMzxBZO2b5LoVYQUXR2FBOu3EZ
RDlEd0qe4e1LnNWWsOtUIjbNPFjPRLJe7bKvDke1c42ncNMzTBYT9z6LXDchuflS46GzuOq0wRYH
VH7d1LbZHxT6rT5oMQr8wNCsT+XlYBCDqesDiJkD7xMfnjOrvvQqspMISXeheS2mYCtXtm/bPaiV
71WiqqaKsCNhGy29z6fvHLFDRwEI8VaCJjbiNu257eFxG59ilfvTNQ3Ethbbt6kuWfEBRExovfGG
HpXzXsVTRjx/Ub0exX8dP5kDaIrk40RnKwjVpIaP/neJulJZYkwL1mki6M9pIcLqQj1CdbQz1zii
AeCSTqbf28rzLgh5ANcA291jdy4nlPW/WRjy4sLeieibQkBQTcOOYOUoxN9qMXpVOeu8VAEPLqKZ
tAlDAt5DoBbnNA0RK08pzRDYNDoYTfFM4kdCwLQ5jv3XGLRYB+TzbvMFMU+f0Idfs/JdIq+jBHkn
p2YEbsSfiY/rYU4IMeoysAeGb88wCRlm2kRLzn+KMGeoBju1V8owASMTey962igrWQk3DEKV3enr
JDVOgjS7j2oXIh86nnioJzZuR7P9VcmMldXCHLwya4fs1HPWpM5bJhl8n7xHJkKwLabBJb9BogH4
6Nw3lkYE6KL4qzlD3L+zWRto/VwpykMNmdtLe/awPXx2p8GfaTviXistNj6qGE4PSMvRYNB0Yb6Z
5hiE0oETVVFEHMT4b3vPVwL1bM3Rij/ClRWGJ/f2ILMfPd6YHPcTGvxycHU9yRARaF45SKb11ixT
uIqBFV7LZURsH388H8WjDsGqLX3MhDTRHsCZF/WLEJm6NZCisjCHBXIiYJliWvW5675rpnbwKbkB
PuaZ467Bhrj9peKfbznePKDEF5yceDv9i47FwPO46Nt3SwEmHwNiWHK7AHS21uE+GoGg6JLBY+1V
n7L0OzrLmoZ8Wj9RLwzk2YBqj6repl0rcWvnwoXHha/MH8xdY9IPUGk49Rph8igY2ei1OD+EPDWG
d9JsuGjYPbQ6argE8XlNfVCdLijbNCMK6K34JGPJNDykZcrBUTmyznzvG9t3Log8wVycHfGz84ek
tjELOXDW4effmJdX0j48xLEHd0VbF9UDTlTeBC8Kj/jBykLrkRxAUOomZmDP5VpO71gD+bA4njzV
zFROTvXFCxO7lO+h+j58zNaVtJfDNkKJQcpzfSktVBtroFKPEM22PBeKytmq/z/1N/5ptwIo7o2G
Hn4rlD/BUZu+OmD0tRVsgXSDl5LNa1BeRNEXYpHTFFUe32E10gkKt3pXLLAzYPRGvMhMc2Bb81NU
UaiwXDdtQOcRHaq+gUjamYBwWJO0s6ATAQi2o188VbkBo8C8mAGSmrSMnDt4luEcQtOJl1Qtwd7E
NlKpMFZaRiRjAMzNpB2tIDH5PJm9oansJZp4dZFICGQ0LGeWtVAO3L0ObOGWfahfO7xaNMPw8S8B
JEbLlKQ394ZHHi9Uqu2lIG4ZtxQ/ZF8SdpdMii4Q0g7tKF+hjB0VtgzxUop0jSQI5xqOCj4GIgv/
Ugmwl2ThgCGME+eWEsZQWmGp8bv/1tWAKwbKP+23kuyYhPTG34p4HSA5sHb3+ModSyUtTzOee8QX
9bsKUD8aH2wJtycGkF8CFIJJbOu7hfyrs6AgLgJb7Lbw0eXd5IbbeDHUmkbxrKvWi9qJTMoTrp+S
lvqVgFhPtjeb6DFmS1vYQGr0oWjEw6Ldv++AiKCnZNa/ZaPMav3VNGybIDWcuPDA2iZBq/zbfizU
uqNcwEkI4t2H4HqZ4vbdJL4JNtlt6GczbU1UFIYSegRxPzNH8SK/cvbyRxBLLwuXDejEGxZpI7nA
i4jbLZOaqT2c2B1naRsBG88UWFf4uG75l1chrwBQthA9ls3Y5GXqv+9JDAI78enAb41SaOtEcOfZ
Q9AgH214hckoAKVNH53vlcSUWInVn7VO5ZO6K5ZPB10jZyKoDUuiB89O6oNn3dFM2/uoz2pimWgc
2tMs96tU3qlyx8P5zUzaobulheMuOT2RPi7myWIXu+veutieXmAYbLKagHHoKgL9jPNSNmaEnVpr
da+ELmMyOLHq0n5ZpE298G5MTU1L9lprxC8m/sQsebyVxnmIuSHw3O/aV3Nlv49EYuT+X3w5tO2W
Bh6/D3ulzYR9zb1XJej4FQsEZZCzxLOXV1I6akgauf15koc7miyjO4fl29WbPSS5xlQCnRDLi2PF
FnzConjLr7eFUTLd4sTAI2shBiABiFsBqat8rYLtjmdRJXPDoR9dQn66pEKpZt1HywjSx6b4oe+f
+Rg6nYkMjfNd8D3+BSu3nawQjfJGKnGmOJci846kY/64uXocJvz0tsPRNPCcxvUWh7N17Xf0wz6Y
f57LMiTygpiOpvrBa4EisiVcpqeDrj6rH33D9391qAuGEXcP314eSgZFF0Z8qymCPel4lmYpO2Oj
CeBs+xKLw9sMjfkjDdAm3BqOLbN9GvNItPPCjPjSMMPZWIXYwFO1lAjw6XyehfxDVILBi6SuaTNh
0xpEu8d6y47MUKj78uSVitLJ9YRQkriMwaQbhVfJv3Cq3eDewcqh/E/mMfd6Ad2rP3T7a3c64Pvu
OzFOss0hDXsQxCHg7eDd98wBz0MKpQRCtU1JU5vBRRcMiC1k/+4i7W95k+r5Nf6+iukHBkBaDLMG
WmHNzEKqfFMdtZNYAxflxP4dBz+U/00ZyYHk3WUmBRR+Eah/oCDNKQ5UfUs39y4nHYkkLoAV/al9
J4+n4QuKDhpJ07uvmLWsv0GD4Vag77zShnzLdt3CeOzL+NOYutgYv4ci17CJ38Ijc20N2zll9QO8
gSGcmWzSrgAjIR2cVtou11th7oqk7/l06tZOFpep8myRTk1Fku4QMHbB1z78v5wc7fOx6MyeyDPW
MQReysqkCXRIDYqpij8GzZjqCPP4HM4mzDV0ZpN5YDwg07drSW/CzXYpf3lPbivsqW+gAi+NztWe
L+tns9F088PDEhqFCMuZK2QbdBNm++XddP83F4PSFkXghwNwP9NWrHkpxao5Krbfihqx+LjGZNoT
UMJCR0nsYyKBnkmYdAxYQ9UJGXPmAzofPSWxZCUGNJaWS583OmeWgv+T6iW1jLOlsAQNhujJy/gB
4tgdy5R/ZawvtV7l9oyf9JUzbkNcjj1hi2y3SV3J7UTvUhO44j0JHbM9OyVA40d8/IkpuyAbrZ43
EeTt804xDB+Q9AIOrFTL7tET9hEqkDdFE1hh9s9f1EzYt9j563H481oxlTt5mvnqruqkJ5MZ5fTh
JrPmMkXboHgdYN3poK238IJ0DsWMFymtMvvYOudM7jr3OaTo5Saef1IF7o2VKZiVNXIQ3o8JCL7H
vSNNOAY9Ac4o1BN6FqRCQK6nxC4iznyw0SjQTmG6lsf1ilwSIJpMCCWh9AMi/I/wdYfHYYPMwm1f
TMR6p4c+SeczXfDY3bcHiGdMVmrP1r1sl12mSzqBcqWJcQC5ELsmPFBqFPHv2+4C9j3ZGeahdDAK
37KtxFCrkrVZeqT4/9jnWOLgAqMOrrehT3gSUrFWRxeZo2XkdqFixlKx28nkxEL5pmULe3RSENhd
j3uv77/QPhKoR8m8E2PZoQ63bJ8slLijOoFSxMy4VXwT4FbZEuhNiXGAlV4Nlwy9N1MGXAhxt3O0
R0USzHi8SupEG/kpbMLQNssGOcE/lCgIiS7feexu5qUGnaBR7b+AN21SGT/AndEOxuNaCAOj/zyN
nWzquicUha0HzEMx0JvISqMPEAXVuJ0amGFdknGVd0mCRO/akPpL9iLiOyRrJv3C7Hatnu+FfXcL
pxNcdUFbp0krH1t3rdmlXQe+AsZlgmaBvloD+dO8qzM+JbRedLKNMvDKYs00+i4mo9CCDBN6qTI7
fKbQPfYPZB9lLSSnXghqdieNQFc0AE4bPD5kiQhjrwS39gRcMYUmi9DALsji+r51xu6ZS7tkushg
yHynWwWVNQNe6bjLIZFwmrH8+KCxwZ7+w2NeySyiRkprSGnLJJjc+WCSUvRnNzgrr15sgQKc5f3d
WSG9BJd+BvMcZGyH1/j0N66JbVtnVweNLsqUN3JyxhjJS+X+SsktMUmSb0gsYwZqn4itSH/TljY3
qHm/dnn18p1W4daZM3pL1bsAzfWrWoYWM1Vjf3UQD1twuQSwcR1qTwARGVo52jzL32Me3jZoY4Q6
Mi9HhguX4vPBWukvMgiTItEkU6AWEirzffSQxPCwv7UTfWDORk8I8CqI80QnggHzhPhC0y0CIQri
A9jixZmG5lRmYSZBZkBHt3QDNZnaFAJel2jz8jW4n2IpQd9y9uWDHX6csxSJ23tTlewpPNMYAM50
QMQVIW16tn/QPU9EfdTj1RdY9XjVq/oUNaNlCccNItJCGC3qs1ncWt301Adnyb301HeEWdeFQLF8
b4iggfrIkBJjq+3jACIYcz290NqckumFx4BQM7u7mZsvTXt2YqU4+u04WWCov0Vu+bq9hcXhQUQV
Fg8rd0myWqOnm88quecbh/vNquOcuu+8PLC7/hWUR3AHBpr9WM9ltgzA20MqK8HVSuBM/h55pPFA
+9TUsYQdfZfP7V6QUqYc+AWYKNmmCD3lVNjnylc66s1X+pOLlkV9r0xgxNZRMEYvJ8CxHnTdBcSB
aywJ9mbBt0pgcHIMe/ElVr0fL2yNhRT+7R1TZy/LVaNA5U+mqX0NI1ZDVqGm1ZYrk/Ox/F0hVC7y
PlXU5LLVkORG9tLIFhydu5vBa+yx0TRg5MGPi74IMiezL3PpJAAFInjZBv8vnXKC6nN8zONxwAIj
67inGPZuadQW3voB45p6MjnUH3CpGJfSJdmP9u7godpoVQJTAXGyCU6tiI+E58KjH+kE+a0vQwj1
Vumd4g2tF4hEDx9ujqtrbMjLtqlVZ6phjIhrmQ+whVxhUDuEr78PVM2rXnk8BJRdgxGk0DCtuywL
9PU7dL8IGRb5GZNFAzNQn6mzktuKMdkjVA+/053ZepoW6AkOoMS0wbcFZqNaGEiDeFLubPp/3euB
nJx89RZPMs7kogT3exCMQb0EoTTrGLdW2apqUIUvjWyrIl2vIq9jzFiII27QyBlsyynHSe3/5jyR
jar7TmtukccivvQAqCVboof+6amW7uvQoVMawTXXkeHcC6dPj2K4sTdbvSE3OHBxsn6gzdRtpRAx
iFuPcFXRRxRjixJk93YIxrhSE6UeiwVJ24I534HgTDjNI3S5lFtd78Ad4MMVP7vxxVMK7kPvZrDc
I9+RvLdxnjLR1wEjshZCwZ6ugj1CNaKrgZPP1Xit81a7tSCSlydxz03+U9III9qQ5jw1L6Hiiagl
SR1oqMbYA+AsGSa1UkJLZ7RFJGEqkzBV45LJj349NcO6Sjt7arCBNkvw7qkU6v/C50lx7waHq2qn
yN54Zk1ERr9cQywbTWLI3eFmyacflzkbpzpONkWGcPibOPYNWgNJn5slr7g3dsrrB1tO0dKidMtM
221vq8pqwxX4OsJ6qP2agqNl3xZ48bX64TPxlg55gsBdodiA08bRxQw4pycuOFbBHInL2N85Nk7m
gfDTY3LHaF7/bc9NsdWQJGHXnBMrpzZLqO+bqic75dXBnPDymsUilulqaN2tl0dLO5uF4Qo00X9N
ADVQBKmbr8XFfuazhkpyP/caSPj1AiQZ1ETugtGgfsUA1CpicAyeQTnLZKhRNCdmsI2ase5pFva+
pFvK1tkekhzrfjAqXHp61F41VYmPjBSeQzJ0M2u3o6k1NODhh2Fxxi5GAsBnXrwKwY3Wjomgsegp
RyhhoNGS5J+4ixHdOUW0xBv9RsR52zi15iQ1wCPjP0GfflWoOvlXGQP7+8mkotrjpeNifFa7GOy8
7hY9lYVvmuX0LqHyZkCTStJpJlGVfS6jpA7O4LgQniee2tsUxEASGzYvn8ZUFOqD84Vp4jfwGP/4
M1iuc8FMijjWNM479kg+MUmBMvSQVGPZkRWXKirU41h2DoBgBdR1Pss373Ga5r/+OXLgshe6hZqt
12IEQKwCaRqHoRU2p/ri/KJNcYoD4/JxLFxQAyxtCWVhiRSe95CYcBsjdXR0nBpwpl112sCJkVHj
IhjZGWsphpdWu5SQ0fCh+iX7EQCQAopaxeF40CWopYyA4uMKJshuTdZQlMFvvVdC7CBRlvbmg24Q
EEFh+JjlmsCjnbqzZcPdILgKuGNv45WBh3S5WMkGieGkOCp6MKZwyk8MIjMbcM7lWYPmSpKtNOTN
L6fPGftAuy4V8h2FvcuKVaHdmUKiYaH2TSs8vaOJ+0dhDaVAnQiqrxX0QgucTgfiyG9bqAJUize/
XqxiqLt8+tiEK8JmqoFYelcrHuCKHLVJPKGygmuMERDF9To99TaUVvXVOPU4xshhOEwewyhgumCh
z776xjgkLnHbUTenSrPekoQEOMP740LOnfGxN9ZSxeqCRRhz1ujkVlS9Dv1Ch/9rklVooTTuT6j1
d6DOCtwC+xy+PpsHJh5R32NlujtWdblmFDom6XZ9riYIQGO9ybpayAVRCYk6OUr6D40KKt4xGOzy
5A1A8n1T1lz4JEUKcnwRS/ghQLBJULAehb8OckMjSl1igr1bdRLo2Hrlrvg5bPjik1EJCGgesYuL
Z+61XL1bDfHRvHbqzxDkJFhXgGch2WuCunM+Mur6+KfPOHEUhW8Tspz12Pcs9MWkG+gvoHadLv1y
WPoPBNmWsbw8u9ljKQ9sdT2gczca4gqCQJ1i9zqKIjTmLBcZ5ubH5XhsGUAgSb9o9EgNYs1I1n7B
JZZek4H/t/EFGvJX/caDw6peVm6fclWPB6rU+hv2owMWcMvtkTZz3ZwcMthYPgDE21BWu6SJhW3x
Lxu2YRlHPJkp2sY+6pu830thXiXbdHAHS/cuesQd/E70fZQ+c3lbBjPDdBo0gsiV1ITMiQ/wOiGV
DjV4ejAwJI0gtsCLT0BxqtpW9R6zXG8673hrbcIwJNCTv1+jYwC2z3wBUKKjEpvpz97CrDWB6jhp
iIOdI2nTM5hBu4dikSu7WpCMf2xDsKltjePs5ppaO11zZ4j/oEw7ltptvLw2t6CLgNln3C/xZb3d
vEdt7WJi2wGQLI0/UQaFndA8oJ7nKJ97Z30O8rZqgYCKw9Cm/1aAUf62jyRSnLt5kW9KfEPa+zkd
kjxLkAyU53fPG051x3cAxc8GVPd0zJ3/tUeo3psY3tgq7guN4KIz0WqB6de3W2QK5+Em9FY6g5AJ
/+hr5QP1pVsKlRqxe+ldiccHG7h9lKTdngEbTUxi6swdeyqcADsTYUl7HcSe4dhhyBMQjDzHig4v
8UAPZ+Kb5Ofd6CFCYxQhhtcnAJU6schDuxpiaG5aTKlue2g87dudzJmLp2OFwhz7NdHMbcLMdtJV
9KZjmZmRXqrsyzqQEj5x0thru07KyHFQuwj13LjMADkabvEFGq8dREDjBGEm5J48jNaLs8K2savu
oT3PlsNSgcLrmvD6VfNCKoRzOflBvTfwm7Z+V9yZXGetSuf8hd3dtQTnIzk+1jCz+9c2Z/5AIpuq
JKXrNfRIRlK8zuNl25eyqFictt4Gi3DNWWFoWvrVsm5aPeVmyYyXROCLchn03+gzLSdbctjG49K/
qqVaJkdo1ivT41EXmUr6PQQszKwkmGEl7kGKz/5fuUGEd0hLmRoo5/e9XM4Znw2bKj4QjCFkRWId
F+kkVWTtLScuWQCtR1gRkIW2DEiM2ZsuMhvOuoZ4OJ50KHjR0k7IFHvxqxXcQggvhwSRZ16iuhc4
CuKBtps7L6eOIK2tnysNYLLL+gZnP1ekrwuy7oUYqGXK2VRxXqaV3mGif0VOG+SPgqozCd47ru6f
EKaUcgKwrIbPPZnaWdeXeMlgtxZAkt2YxekT9GvIMmAzlB4HSvHZB7vbVVYyQ4OyEXvGT03OOMPx
9m3yQ+l83dTCeTeijRKTmt4GCNnS8S9SAlpPUFQ7OWH8R1JpnYieQOdnJr7Y2tMRpCZ1PDWF4ned
4oGDMRpY8AYnGjomi16slJVZoWTe/Xb3r9d0VcobxG7kQiv7zOCud7K9IusULCbgmYRTGyOX2kLb
KTNiseEpMXVtvw2DemjIf7+PY5NfJhEjptFnK6lVfsEu65yPUoBSaHHXuJ+FUixHdrVDTOOuwKvf
2ZmX8u6WvMy4E0edSTsZcUP2xHs4t2L7by18dlD1/5/jQ5LoHrdsIQ7W1yHc9RgbYUhVA/lrQmv3
2V4TM+89Ww/VA8e6iKmwpPGdnHkdlRSuN90CvV0lgD3oZ2or0RuUcyYtPMTc0NDRIWYqZ2BZwXp9
9hiBnLa0Gcz9/cOd1QDUjvyNgXH+yI6WiOKQ6uPZ7et7at4x5T6fDI6HXGT2zsvW+5A3jJe2em7a
/pWd93/r7lLLbVpBBVPMDSa3/nSkYqFZYDgxBD+A5UHyODwBK+panysOK8NXvVaiq9q0ZDc+y9v+
oEjQaBwC9GqienyrQNZNd9nTmP2Drc86H3Gp0dSTsARbmRPeUxGFqh3VOz1akUiwKhzAQ4TGsHrU
bPWAJaAPuaIYWQ7H++tBpmhiBTRYpRp4CQKsYTXdBsRVIyk0QfkmOUcvZZqfNoHSkR0At6y5AR7a
ij1k7xUIcvw1OCUTlmeqqUhzrnHUFO+vDk870OgcLxiWYlmFr2cDvwBbBE5zZHgrbJ8LMEQDOyGG
S+YRU2si9rBgGuu63GFD6DL7YEwc1qgmHAtGeU4H4AcglPSYmHfcsVJbFDOaVPjahpKT7CO4fbNd
Le/REyB25ve7uJGDKphGPgt9H3VXKPENGilVs3ihWH79CjOd9tmJqCgZYOjvwRMvkrVNrIegbkSt
frO1RPdM8jWwPUEHJ2HCqq1LP3Li5QcQx0dctbqN3bs+fQNlmToo1OwaZgVYGtx3a7WesnAN78C8
JpthgaPCvvo3Pddg21XSZZN0+qljmaaw+D916yeVeXGye754gi2+9JRotWYDDF/2/kA2/r4DMV9M
5zhwpBRSi4IR3QvvG2vOhW8Ham6cRjzSQ/cAMVoqopc+mvx3sMakzTNDgulNuxmKpDIKZDFAGJpC
N+rUFe8++Yn39v7xJb+S9K5j0xOYf4o7nm2J9YDLmpY6wL01QwCplZWI9rzsj9bOkO3gWvMArb/a
zCpaynK5hfte//8QFEIfLIk+6PKObZlU74Bfa//0l2nvAmmGB3MsukGrjZmaqwJXNh8dZPo25xnX
ON0h3gHylZRYVghFCRoKWLhGULx1kToex7xdZ2wMS0amSDXI4PHz4qdEzr4dufMnlY1PeMmrNEha
Qks6qCl4nE5lt6u6W0RPyHTFwVBYbe6s+Fu7ApFsBS3/y0Ag4vXkOjCGoM0DWd6vKZFRmO4Q1ZJ0
nmHqZ6QUufa9vsjsp4cUdJi8Df76DugONluAfvVenzpa1cIpSmsWG0WOrS95gd7VlbeJidQGYiqf
drHvKGupcgSoLgExcRPejsJ5ywtQ3Q4SjgwCM0cckBsN12PaA5WqMHKsi19A+j1/8tWl3fCzF6yZ
Ou92X9dxHIyqDty5IxgG1hMY8ocADUwhRfjacbp9CCaiPP+Zp8Wlzk1vKVLyKJtzaTOmx6CS8d1W
7+JfVQSFZmVYtIg1WQWK7VCnQyZfVdGKejJChuwTiYVXlGKvXFaEXTXUS0ZbxNvlc7otGL/lyYZY
Icj+UJtMEUj12kA+O1SZdsxTRByieqMqCnDdh+W57RAwOZzWbp4HOkWjhV05AYBE0tS7grhvpB7G
p52RPX4YazwkClCWFbPdpkkEZPcCpTQOzsKliZSXLNY5JePhw6nrbukJasQDf7c4zof4nYeCMB/4
nBfFyAwy52Uzvo/0glp6vQC7JL/QHZeAghENea2pBjBHHKgO4knlvuDw+VHDvIwRDL+t1aVoi2Ae
qZk+cEbosCOgM9KincA/68LMJRl3EXprsFUX9C/K0VfFGJnmyy35nvS0VtbVmBUK43aYJg+XJ4g1
YRY+JeeTea4mMGnrAsw2RoKMJaztHfhJDuLHUkhzDtLUx7opHNBNJ3hu85EKN6YmB3K58q6nSZkL
3Vj4Y73w7rHphUdqkRhS9ffdeoVK2o3sZSewxTjCw2PkjbkxuJsCmrHHpGwUmnAbkNLrfB5iiLCs
N3uWiXPh0lWb1YnDz6q5EOYzxpM0cRDhASiJl7f9Q+3wN8keLmYFSRUQHJ6qFrI3Ki6UF4JisIg7
qyhLF/2H09iY0pRwRg1YTQr3qjb55HoXfFYR64OPreA92tUxBS0zqI0kbNM1eW2XfJDXs03yO6YU
msp/aXYzy37X6rlPkGIsuofy2uKdde6ZyrguaK/65rDhkjAmZNgG0zJYfSUOCwZWLlsvnLTInSSw
vyT/zjSEhgLoIy6JobT5eESZmkmenzB0kB8xEfV15w7if7LeVVpSNJRtSw+SoXiu5kZ2jXi68O9P
rGL9gWV3HBbi9jkFWR80Vz6hnnVRkIJn566Zs5n84bwUeIVbK7XX6R/dB7ZC3fE0wTqkNPjHHf1Z
69A8LbjGhYEeRJDYaBE38Sy46FoBNAxk2E9Dwi7ODDP0QzMSD63GsjgeuKvc11recc+GFiE2A/ei
qK1ZxyXujhfUq9vP9Bo3UOZZVDrNQtgSoaeygB9Fu9o3AHPPGJONk/27qmvJJt2znOUmr5Unlpml
s5i2vkoeo2DNSWZIZ0OX8KC59m4/RBrJRMSolBg31v1AFlxIr8w3aPIAT8WPH/4ZaO5dbdZBK6WS
v3XuJ7g3G7PlAW1tzwIL/VXt4/p2yAX8KTtQ9ZPujtW7glMZTno0j7Z2zMlNB68zBd3x6VeFL4Hn
FCp1gGxW6KBD71XXNwKh3q4me8LPFCJypb7/UZAfo0yUjwyVNntly0Pj1uAgv54UHY+mEtTBj63Y
P92DWzB2dXaYOjbC06Q0n66Q5vs3SN+bovuXgprYfbl5VwO5mRenbKPC+me4c52bjMPtlDtwwDHG
4A9HPFCr68/CWX2oFzDmqX9AqBcSllgClqXDq6UWxeHKMo8AwOSkxNqred13lvtVCDE3TuOgPvrN
PYunHU/0sg2DfxxTV1Um2AQ7STp0y4hgFhXlec8zM5fKbQVnV5jF4KRp7ieKifk9umk1NVBm0DHB
kEiwXwZ3Vim7+jERh8L2ulJmFoRb5YFYPQt9BC1hwUIv9qYVT4k2K5g9kAe9ZUSqhHa2VQpbhhbW
BIMUgrwkFfloKzojlBzV8i9zqNIp9BxD9VuqoMCrif90Mff5aSHD55e60KP9YiRhMwWykOZJwsKc
R4+LtgmGzlg+7cYsU5S1UggHv4jF33SHHZWGv22+yfN522tk3qWpYuOplH1etcXs8gkX8Egy0Hiq
4gjBa5CTZdrl8ksdFJKXofeZ0k4fS1tA1GHvu2Zq+5FaVWBtz5mi5c3dDmS9XgKFJlsaytzXQnTm
w4Kb0Oif4JXLpxHeDAuN68EJqG45kINr3I+P+rcCjSKp0ulro40igta1V+50yOLWxKNBdRNWDH4m
Uvb4e3+X+QWhLhtTtDg0RDCjJvr+bJhBu9GbVyL4C1O3SNrekH/C90EMnPpWp/e/FwigZYQ4JB9T
XBGcnq1Uw+f4XfuUFuoM7jItJny5gMTniqEKQPBaxd36AyDBUD0GSKn5d6CDUY8rpK0zj373u9uE
f/9Td+zFekZMwD+uMdFjYBNrCaCccu77pBsZzvEL4h/iyyf5h+HUcKYHvByl72Ez2HHcyZpYiH2J
B3mIkj6VuryHksmE3p2GcyS1LY2eCdfXI2UXLL1U/nBHbvCfiKRPCrLVV7p50qaOjXMTBmReaxh0
iHQ1aGiRXNd8Ut6vJW2+9KGh9jJbVNKNryFTKRD0iZUpLeLj97Vn0nWVi2AYiNp9ynJ5yuAaPFll
mN4hp5QsTTncrTSu38xc7eOPTNHVfRy7eAFyjbH/ba7Mz1GjKk/xjDTVgmnQ5je1DxE+9GjAjqOV
E9FJ9n0wAYoPVqgtMP8v9w0pkrDLYTpl99qM+ITA4hOAczio3EiUBZlvNLiQ4IpOG0YqGo9cE5vp
aE80/3KksX84oRC+JhVZXn+dg9sQA2hXUWZM/5azgXiT7K6YUUuZ9k5wFNO5u4VN+rjIAIYCpIjl
pGd7CnCJzOlUiVG/taY1xWy3ZPIaeDJLJ8w4W9O2tyzBBmAzxBuxsfMfMXsow4IbGNsb/nNizqL3
gQob4dzChbJAsJTauI9ei0elvLXGSjEO0f2uQJiBHeetwoCwZ5kcnfXn0fsjk3C5V9h2g9HvesO+
DF7ZxHha4G3BRiIiuybICA0O4K/1swHWWMZVhaxTnfmf2ss4NSoFn+D6zMZ6hqZqPGkUQkOlQudW
0TUpktg/NP8X7euggFzw5Y//k4/aa2q15isaOLGYT6l0oqzn3Af4fFhuaZGgrpGmETXF6+TabTJn
v31j9CtWC+HQwbwT17AggmAcuh3IcmD5BLrzfjMAOpJsYsL62E21/a/wsqBUKh6rAEsHUBAnOKlB
wA7p8xbICy5a/GWKGGNgt9gt/Ri1tePTxbHLO1nY1LVazQEuVxf5xY2cKGrdGzUNWmD4Z2dj4vhW
mLjhJLflzw2+yTsqUy4cW6rUr5THSd6/i9JOXPladw3YJIk5vXPFXYihlJGgfa1egEMp8SwgjKfr
wNf4DXjCo9rtqFbs2a65mQ1uiN/Q48V6kFRaZw5qSanPg+XpLM86xSn1Mkbb+tviRjuW22coZfpo
995gh+3eByO4MhlK2sSJQ4VxzC7/50gDIyQ28uFxoTmgNTB5QX7SfW2jOSrWofCnpRUqtcVm166H
WaWC8BxmFxw5td2qThIN+Mrb4ti43iL6FYsUXXt6D4tRtVtnsCLWKWBl7wuk9GXum36ezMI1mo2K
qo3QC8qGx5+iSTq7KdHCRurOCU+2sQ/facT3mwBFT1E6pney5EaymUoyPgz4acOpui0CfE7us94/
tKYQkbchXX0HI1D7B/xGW/1zpBJ3CfjE1/bxoXCGzsQklS6a+rCBagJJzi2WBC9Qyb1/bC1LThhV
LrLq45kA7mnNtj5dBrGP/aqZNwk/8/e2y4WFwFb39UfuI6XALRvJEMJEEb/ejRMfxOwESdX60eV5
gHstZfs3aOaOmcROTUXq995snZWmpE1WKsGuDbyaP4evU/MBnBJFTdfHzx/BNGUn0vA5FP+pi4Br
zPJeE56KIW+tURAfU4Ll6MLSX/wqzOKe4zMtmPypZl3u5uhBCekEVW0rqtPwfhjcdsl+wCnrn6rR
2jjm5Ufq2qduTbT2RqummGfDQ2l1pYDkVUNS1HWbMjvT+0CbS0gvc9rLWZo60+Hz3PoguBdE+TbV
VtQohNGe6jJm0nHqhuLO7pEiVAkUDSyO5zTYL1Gw31rNwC5jkqGDm3aWfNU9T1Q9Zowns4vV6Q0o
9T4K8/2MlKWKDGSCAmRRKDpt8DJr7Vc0KZJlabwdGlLUEXqNJPrMv5NzY6kZZp2ebr7g6JnAziDG
Ervp1MuqsLIPBar8Ms+vGYGrkaRtkqoDfWJizXit95eDmGG9jerHzxqjjwtKCMlyvu5Gjk7QGnVd
gOCXwWQsFPorcrUD+rp12DmVTkzoahfWvdAdx2dph3vkKrkNRtwc6K3E8NSbjSLCd803IDIPt+w2
RAyOLfH4DgsL1fJEdZ/O332J8T+aCWiKC0MQX6u5jWS+8kM5UGtdXrEtLjm1nqKrNI4lupuP1vdz
au1qD9xoL0zfypQEytVVr9wBrd6Tx5WuJvUr74T2H6xFyfMUH5+VrCCP8M0J/bUp3FOpeynUy1Wt
oiIK7hEXVsV/hEOlXMvtUXC7Xmmf0Eov3KXhR0ylO2+/LuKj69YOaE5lStvjO4h610kGy1qd95tp
FXlYp5eq21vrAvW04Ft1MZXaagwPuhEdLctPF3885Ij9NDxLhCjyGU33UBdhqCGYusmB1B/fddKT
2WQta6JyJoQpvbFGDEN/MnNXQS84yrSdbA9YiUYBb8At/uYx1MRmvi1y4Gb+n9gfSQo96WJcweqo
CM04vzsKNCaFYCGXL+lz8eA78W9kpVs+IqUnvigw9DPoi1CAzIunvpe27shL+ME+Vx1c23rmcagq
hI9gAGahbaGmaYYaDduqciBXW17JT3VKnO+koGqsLbVBwlZ6Wnh+UZCsX3Mr7Z3uQuT5UrhC3x3b
IFoQ2mT0CiYLrosJ2qaKxyLu3rs0rWlM8FX1wXuMHOj7R9JpfBz0sI4NFuWUVAE0OApwVjwFzBtO
iDYTc9g9W2a2yF33MFzmmyiG2qPxXuRrYgSjHXajH432uGolm3IAqgDltMd87kUs4EsHP2LUcZyU
tFIguCDhflBraGNX1dYXQWwPveZ/95e1LfAppRi+bRAZmCPAqNrvSqTCwfZp7FA5vDcbWrqJo7X+
bqc9EKtmPGvHxMU58ifDKcQJh7sj5HtXtaiVuJCp/4gaT0y+hGUYE6vJVE9wmyF1D5hO1Aj0+VHa
1YjP9kxnLkUzABFBwBiErn5yLoOyldKzFG4e4r8PeTGJMSowDZDmIcZGpvMqGGqY+5UescmRXRZx
9KbnLvmFyHRIqoHxr4rxXwHDkB5U4gL82PykZRHt83Mns/jJ4/3GPwVjRwUkXeB2ekbdRrPa1l5O
4L4Fxu90NEWc+DM6Og4pi7WeoFZRDCjjhjI4002BTqt60PMIuvsXW2whCyMSXZrczvKyNU91/7j0
GEkTJQHBc4F4hd6l+J09kFQNZ3ne24GWPpdl0BFBln6UR+BKi97N0Qhnwawp3Lq1koVykAKqnxoW
2tTRyJ6FmVAO88S5zVJILauH2gXbwOc5g00JiUTZYdgxq9Et6p702lmNdu0guStC1JtonvRTcm/X
QZA8gh33OJBQscmsFCvRAwVdjgJTclmvjbTloex9STmXqK53DRRkdRywfCFHkn050dsuZfPtcfnZ
f9maqlsovi68yue6keM6EIx3jCRcCiyH4KytBfDFgTwiWyIOQM4oZyHb/cuNPJ7zwZ6uu+YH1xLD
WomH/ai/4+F87gO/s8gUyxQCqj3Ozvy+MffU70zrOI2b/FZSzvVE9vM0jTkkriKN7VuLJCgBS8uR
Temk770ZBzRu+NQK/PlC71w7vpai7fPzBi6B356DQJxal4LoQ3dWDyqsX424gFpiycQMviGeOLwr
9Kf6nMNF+T9kx/y68nEOWO/BnKkxahfN/8W3P2ug8P8TPAqZWhIlna0cOg36gSvhmgDVBRTdY5gI
kS2t5dxsb0JMGv3KdDmXYYHTvnBz7QHD6XpCHsfS6hoxeF6xZnvmkM+RtA7Gjzvyn8dzeps20Sio
UkDEzJj9xVI5/uGgHHVKlVt/v0ngz38iIo4qMmBi0Ma5pvMcKqJjvM0OQFnfrxQgMhRrBzkor/78
tWhHqGIMiMhoE2XHZrYeSz+KDMEI0b92/2xGlNJb3L3HY2Hoq6Cxo5akTLaX9s27O00bUMdnJ4+p
lLF9AEDemY2w7ebj1vTEms0qta6EtRe1yFRpPUfN+j/iFs/QCHgCqvnGptbOtWNmTrg1rX9Vls1V
9FUr6CmIHERzsfn8hnkSPP/JtnDZdpZa2qWGnmzLeL4HwbtxRGjKPKMY5EyoiKyA0JkDE+h5fzWS
hrSGVKzr9vsPi1w/3wXzCNuD1wXc02cOmETDxTWa4+WUmu5B9hq41i7N4birH7EpzPVqJFMaMF/h
x6LL/i+Oofd1cvz84rFN74gd8+VPPWiitLe/fWAVW+UQ9uMzjzqSpfn45XLNJg29rh0bcg0okBro
85hPajX2OjhUuPLTb4c3T0j7giy1gRA4bh03hUHJXG4UUEa+geWP7eMZ2aule19mNb/Zzef59p2j
GeijOiifBqi6H8GdFOTo9RlRAf2Dl03YMkKs5qcRC+FesjaObi0W+SSAJg2quLlX6Qt2krHolB98
IVJJSmPwd3/ExscT+1ouziJITyDKczNtD1G9JDdrp/jZoSDVvhymHv0bxec3NWMhr2xj9li6MGQW
Dryza2bu9vrOVIz5oWc3osQbIiyFR4PCimfAGST5GsAu9mGyz2tYBeH507sf34xcgY8PajOSq7AS
2kH467HASvoWyDadmJWsn7/wS8i4N8kG0mrFANgyLy5CRzy/I0abpJ8CFMDQlnPVwyETIhhDC4ZA
EElSbHPcwCUeKbxnfvQh1pS6gN0QBV37VolYCV8zOvRjj63cHoL7l/g8l83+UXKuXS5C3SqwTFzu
JDQh19iiDyHGm5y732Apl76P1JIoeVZUX/D4cURJADURF+tgkh4yLs+vZ8Hqg5hKrUkPAym/P4zF
+2ORwkdSi0Hwlii4ESbNXpVcRL1NuyBZ8QdXwWcdjIfccHnGC539R967n4AS9ufPmhwzSSY3+pVr
CuJSRmoaOgdlUGQ5A6DJRop8e75KDrulM08TS6RjVDN3PW1iQ177g9fPjtJ+a+U1nQNPAzjHhiYT
urcQJ4gWgjraT2U6ZiPhXuzgnq9EN1EKUJDa7x4/P7ln0pzd/IHfVXUf/tDvD1ROZ0RK5Y6QECFN
tWrpVZxLiffNb8l42DRS5ZosLw/dYErooo7PH+omGFU2J+HhuNqw5k0P8KsikySDcCBtdpwqX/qC
gtAYfcJ0TtgXnSA6XcnndXxcYlgKkrJxiUYNJfveSjeOOTZMszScuzqM+BDMv4JP7Z/BEmN6ae9h
9HTttBWOIHa06PLeIEdCY4Aplg5/+uejNuFy/R0hvlaUyNDnPDswBJ5GBb2hbiz+WycfY4pl0ZfF
IjC94xvrkVRvVwOlE8Ov1ZQuXb/7RqwJT0kDPT1xOxq7OXurwGeF3WNe1JDc6rwxRQ68ryJKt6a4
qg0l7iYvqRe1ORFjpLxDudLEQwlOjKk8XleujDxIn4jFg6YsQlleZTnukeZm7OSgRX25vtPYa/Zo
6aBBB4/nsM6XYGh6GdvNiTu7YDU+F4yaeejTLAoO46tF3XPfF0dUoTl3WDa4HtQTARLwmhWCkZ9L
jUc1MqCXvs7e1frObl0ErYytcPkGjXoLHog5Cg7Ek/MD0wyOTQB3BtjyfzpSPnAPUpkZ9EuSRjbO
m6X1SUErE2o8W/6WqgGgpGu1TMsu6udyu7hmq+4lwDtBY0psLseDOp/7BpgaoI31qAQbXbL7YVWi
+bzMQspTgiDjNO3Opk0woDsdYej/1VmB+xwCK4c4UwCIS9fabEB34msZWpw7Odh6gJSfh+HNcxvb
GdfJcucYrGvrL1P3Pw6vUPqP9bWeyS7pR/j9uipQChZdswzcgm4G7+2zEpcvAVMprJZhaUHtzVU6
Wj5z4BbUT8tFVkaF89hSmwf4uHpI+XH6PbONtcClWqOzn558ooJlpM036qR0ir72Uuuj3ptpkMS9
5U9scFtKnIcVGSdAcLdM8qItphhjkZ68Ri7y6LEpBnbA2Toq+pG3X/Mcnq6MgyEOseUI1GTX61v4
+QvQMdIxTjl0cmJ0egg660qy6wciaiU/aV2uGXByMcaWEb0heBbiBgI38AQkmDT0/QwgGSH1Az63
aRq3gyHO3jDYlJek4OIUERxLUZloMkQi7mpONbsXc78gx6P8+6fwDb7l7l2SFzjbP2PuaovTlwWp
ZoLa7uc6bWHg0sYF3P/cpLYe8pyHCB8Gg7eHV1Q1V2NfuUsa4RT+L9YptbzfNAIucpPsw5GQGXH/
hpHT1dDQPRKaR3qsH3O+ySZVz1W9923T6Fu7Zn88Bvms9QqcGnQYyRsyCLK7uShjCJpH166mxHpN
ZoW1DXb8M/v6PKZZTQj/+7LVG7cp0k8xVMkUz6mir4DWe0JnQbAX+L2NrqtfvXqnRmson2tORrf1
c+0FJhU6+cXQNlKTiGP9dnYBTDGil0NdTQueEYN2DgTWS1/iw3r03wBRzf02dn992bJteqYNnEW+
ZPTdWtA1nqXkqwZgoJm3UYyitojrwmrZNmLPioRY9F9vGnIYRBueVwbyldz/Ybg7/PAXhatwzWHg
wM58WsymZ1BD61LoCFf8Z7l5bpIinHtIxlCXFgypw2BF3Gv0E5z/dwOJhV3BxLVtZtvDr+fCSZM9
G0WDTUqvqTDRTbq6I6n3i10DOcVrFUfhPopjweVHejGvs7NuwGEDo07mMqEMDfrgwmE/uCQsCytZ
49DXx///jsErqweXAOnfB/3ZOpLMIBRXp5+k2k6ob5vLRjeU5+91PfHogyb1CCJCRKHqvoSswv3B
vdt7eGAMgfjN5OLE+YRtO9n8qelKeFrO6/P4k4wnDubyY/XsIT8tOccuK8iSKvXWrphotEXA8Kj/
MyH0Cbhd8Mg3EBgRTjWMfvhIBmMAbuKIjsDH3Wh9Oo2t3CHYj+vuKxiv5DB/YRcv4fEsx0mxcWMW
2BKNsJ5N49zJzOngUHxhovvRuk5D4SAzhvfJr2+w58SKekcRcXg/8UY1VDQrFEkqV84/xa46O4J4
Omu6YXE3Qw2ZyC/JOSn5b363wqIWKRKBdzBhOqFP+G3S+btkkReAnW9vAoZ/PiabcFkrOif+A3i1
C9hzU7WivTZd4tZie3GR4I2mePu+NU+jx6GsqWmdBajRflacMuStGPBI7kw9jHHMiu97EakA0W7j
8OWE+HlcQOP2QdUJhvPUbpGDoJWLfiz63ynefE5KV19/5bXRzUiysPwY8lsghwKkyMHO4CBUEAma
8KTcUJnyPxSYs4FK86PpzIPISXmzipoXqmLMrMymXNO8Qkm9cSR7bn1Gnk7asVGz5IsdNF0Qisu2
NO575LCXClCujPAveOUxKoClYz54wa73i282O3XFk2iYD8mLcjtA8jZrs6KitFVK4u42gTs65pry
q8t3G90vkKyVfjtje2XKeZgO0b83PqPQyt3E9FelaDHEaHktHA9NOIzPE8E5wafrKudjMAfvIvmG
M1xdtIC7hxaGe9tOMJF8M4SXco9Uve4O/VcTUS1Vcy7Hi8vb7d5k1i+Dzzkgrvo0MssmWhDpVvcm
Zl/EThV6SNde7PczNcF+3lzv/puYWR4cFJMf7UvNM4BR4WL/R03jBr1Y7AchRtfQ+GmM0Nxqzp/j
H7uRS/bIbUvkZjMcNKt5jH2+yhkCGLEWAn1NUQ4qC9BUAJTmW9ki4iXqbAmcmFLY+v5yJTNQntys
xsBrqErLxx+2Z4rNg6RqMBGc+jSRrtAqthOFmOUzfQpQF3SKD1qXBbtjoZ86zYDjm0H5on+E8jQZ
lcJ9PN2xnf5A3q4ZlH3cZOEnG9p7/Fwfid3XHuJaInHXYFizzqA2km8+JyyHPkJfWOtQLIhYwwBS
PJrm3MeaVsosv0rdln8gsHRc97b+2I8YJrKI0L64K5QVJXJ5ApjegY3HVqjeUKbz0Kk6xpnedjmT
TgmqCQ2aVKfvsVc8t2YUyu//ybxmFsxxUANwdX89LOf6zSP5U88RaAg+OhmCyZw/LflKXBo8hCQ3
y1Z9VmifuccHxKANuB8077C6hI8mCO3ch+XOdS1KLxwertVphpsHIYHnPC/0FTsL8SFcbPCMkGxi
Rf0moqmDT1tNxq7N9fcO5yxyKA5Fsxl/D03y/ctgT59AwH/6DwaIBZoEbmLG844Yl+qJ7Qg7+5KV
VQ9UKjfMJZQ81s9G7Z4DLQBJ25bkuHFpK9RmAhevSPwyk3IzxX0wQUnnABRjSdAKuV25wM2Ewq/B
fuELbUi7Das3CnuXsgEKktcGxf+GSJDdhtNQRcRj+Ge8GxVg9jo/MnasmIb3hw8LXbPoeCz4WGwb
8hwmCbcU+Dd4VmOv+ypr2gy2rgXHmiZ3kfb8Pcc7KVJxKaEnH8FWImagwRbM2awwyuYpejs5F4eP
OFUJ/3Rk5SqzZasjX64uq7ZlnP/qw+iueylZbE9vyLCV60SRY8nQlHOvF5uN10yR45SEVVtfcmwP
ziBGnIewjqFa9yV50dmfmOOgUbsGQK5OOh/I5TmK05UcqmkAGaN2t2zIxWftnDHA8rmytFdoJ7+n
C3/kN7YyL4v8HfLVYW8jsopbiqPTvJuZ8wdu7FyMlwrv11l8P9A2keUJ5EbS7RXDqV+4kQVKLxPm
v6wtjL8ziNGdGF8SLKeFD1V0BZG9Se1QvkGiLZKFSssqcbHlaSyXqnS/oYeXCRMBcuSsUJ4rotHc
1OdpGSNk4c2qe1/VdKgYvUrKkxVKuYNs2UPIeq+IZJtB4UO/uEyOa6m74weqFqYJQflSxYAvwlfl
6aVKbE/tS/NGuhACvKwcTi0j1vu525lO4UXwC47dSZtj30sghmh472MOgN22PiogO8V++AciEIJ9
FcLCDhSpz/2/6Oy/iHKs9h8NBAivfK75mX6oE6Ca5K+WQMm/rVsXFI64gpb4FF7VqfzCPzBd6Vmk
vIn3UscE7pelC1+b0S5k8xxQnewQ0VjErLHkueFbHUqW4TXBfxAcTxe+yUkBwvrW38Ebc7zE/eAe
4MvFBDOXdKlwqZCDkNow3EslprPLnvp3Z4LFa7WS0RZ/HbDtcdWhFch7xAo3WlYQlfx2+ZfhQDYt
Wnziq46R2tHtTWhv1BUWKH5mbhdxWNfQC29EYBlsP89cJSaM0WqC24HOhwrmZ1Nq87X5XsYnIGx5
Xbm3+kJYVkL+6aunJ6OvqOERNmyY3V3qy26COZyxCMoWOBliVupMjpcpsWy8nmCizglDMXyDAQvw
xEu4kJidwAat3HXtjYOKDvpH7Vznq7i/KNmSf1VIJ4dfVpixwnHJ+ay06Oe/zmBokALl/SLQ71kx
64mUQCfpqNkTLN9yBkQdq7My+KkRA9z6bydmb7M2HCQVI2BtCO77B0Uqgscnu/DP54lVAsAfRcJQ
WmngydeNNGnyiZOU7id9SO1wu1PzmIZz9zMnZsc2meWI0n74c69kRk+gTfCW6UTMTBM4kvRTde7q
R1AVQUXyg++mW8MME3Kqw8AgEiL2QeYMLQv94BhuS/ER9xVcNBhcFokkz5sYMpZSdOHbAZTRpd2s
E7B0TtI+3b5QDtjZxFJz7oavLoiuHHLuAmnQZwiBkteomA1ZMI/ZmG56g9AGVOoLzNFzc205IHdx
9OyuGNxIaWjVT8aA6tDDgs5P4hHc9eSg7EvLL7KermwXd6jj05hANAkJBGooz9239VsKNMMRF0sE
JRkpbRON5Bi1EFqZouqmarCrNy4w3q0LbZektRclAg4/+9HfEpgDYi7frS06ix1L44KYtd/wGIHT
5Hd9om49wCKkdLRNypeQqCEZCuJd0v15o0rYcxZc+nZbhKjKPNBc9Kh7sP3SZGNp0jE3LIqcqnkc
1If/2nWYCAp8DAR/BZYma3A++yJQqydUYhq+tGnNfZO1anHntE/fkchfTVANMq33zieDuEtVNA9k
BopfiZEfia4QwM4V6t9GVzb1h15LonJnRrzr9YPLFoP2niAxxbmoTy2JkYZUyNwh1d4v7zbzQIpM
NKP/WpBjHzTohP6sXj5MBynb23MUjU1Dlq6A1mnLz5e8IvObuXss/Kb8wveLN2y6MQ9aXLPbHt6d
e11Ag9TG69B1+AazRYPPUNGV+0/FnD1phXcyqBSc1mAXZZpjAC4mPuQKo2gRVvHBhUjlhVEtc3EW
A/gH8IAT1iLfbLj7XUfL08NcDO6u+q1A91QKnd+i2OiqyFOj5Ku5Y3WMkJvhUj8sIZpO0XHXhL4r
iUzbLZ31HsuKuueuVeuUDq/SI0plO2lstWXi1cPHsWh/P4ljVAqDuxY0d5vDKxtnDeyzzyzOgPbZ
FslDTI1bMbM2Xgk5IQ6o12xSVfU+KbUAWPokB5k2f4kU9/ObWCx4wi088WDk6YqodsAspRMjxA5D
Wc9CEovKez8+ZJsFq+QZ5TLvXpowGuTM4JrFT2XUdneH8C740mF5fujyyi2OCwjjEy5ljEspemwW
LQbiZhf1tCDM2e8DNQ/pwOW+6o9VdsEverhHtCUXUImolnozBw4iQsHaEiy3gLZQ6Vj+4+OmC7I5
PYR32Hhh9mEGf8e3Pxm/fpNh8wH3BEOBAIh1XqBXgFJHcTbsdIzCzrHW3OLyBVKNzjWNwaZq3d+v
Ysbdw+3ROSIEqqvMJRmNE4kmuYy9NGJlLFkFpfXrLucjKsVq7m6xHAqq+NkMULtGdk9MPHdQiu6P
hpFzOs/rP2rU/WnUK0PZbKlI+KX5ft16yKVEpoJ2FD3ciCQxIpdvTc4LpIdoYhCF+eozyKK5huwS
uAXS9qmdB/Gq8IWgfOCbIEPMaOKPopbVHsccxOn5pr5/BtrRzEK6m8q91AiRy9mId9mBbIFUtEr0
KUdPOPkpvO734whAioFIElKBVdrZrCpAlpEUZadeoKZvP6PEcKXY/eftVBN5fNtR5azyg4pzKusp
JC4InWDu6rm8ny3ZY7nMBj3oBIWizqqTqDmgBIaSaGSxQgGXO+XjNrD2ZAJaCoELgXxbq3W5VUgG
tk/HmuWWfGhUy8EL9O5c3TdB58Zo7jmaQZV/V5hHDWyWBvhbm3JahlcCtFHR2bsMh/KHmXjBtqar
dJmSimLDrEzjP/4JqKZTme4MbGLsygwAZCo04LBplHx4p5KYHkD7xsk4d9KVRqlR67YODehIognq
9/8G7DjGbtJN+Q+QybyeZJamUxMwaxYVGPtC9D9rd/NxZHGZju6NjHLXv4Bv7EwvWmvATCEPCEvG
JAEF0HT0W7EdW3xrHYI+b0f/BREQJ8MNi4BplGQET87ikgTnwjBuAPEg6MUsADxzyGGgEWPYhkgE
Me7jsXBFziz48gaE+uNGENuddZbxhesaQDsv+/dADyop21eZvciFU/1SLYhV9z/9gA0iJxoGAHBJ
ds+TgmITTUmuPpsJ52RoMlueo7VDY7DBVyH0Th1jcSNwq9nCNBwOPZrZqu50z5RyQ2XG75mNMwC/
XRvD+pVxMiQxjMNkMFxeYsI0FiNfIogXk0xbfQDMdx8fjhAQZdhnfO2fUyZ3cRv98nmAQ8cv1vZK
VVkjFcxCXTPb0hD960ITwj+lhUVkZyaVhLtMEEdCtv74Hv5qHUYj0fOiBm/Q97Df8HFovEdDnGis
CBKvjxeGJZ3AZVdtyNL0AINx0ZHxmJVXDcpZi3ChFYOIaiaJ3sbD8EBgkfvNgsW5L5HVYRAY3mZ5
MBVNlKljF/ynIn1R0LgoHvEsXLKaTaXwg2hO9d0KiRJJxIGtIkzHxtXN3iUWuUkzd+ODfB7So2Xn
GAyQi7IcuVT8JYCAAH4tbuhbTx1Z6ZS8ThQ5R24gEGGMkZdtJ/ecWjT0ehciJLxnorWv4GHoLEqb
wcu35XBJ4BfqFqys2+y20pqjvjBTIdJH9RY8s9upKjcjJPipaq3YLYQUoVqxcfydJCBRFegU4Zaz
GBDPEX+/QIgMt+a9jCyIFfP4PxaDWdqeT2bcHapLHJuNaWl7nCKvQsNRnTEOgdLlTpSd62/ZBxOs
jbhd/JxRWJfTHpGlc0jirC+uL4PbeVCjl0zfegzov2MvRXFEuMQPzJkHnwBhHeGvb/nmtE2nxWi1
1IIUgmnve2RZZBSnUGUv7JCEx/Qb1FwgOjbtpmLkGCCpx//PIKZvX/9h5HmsdP4exRRBvcWwY1v4
It9lx8SPB6Il8uu76ReVYBDHTYtPNzLvWUF1kDPbi44Lv+raojiBgvYhZd1extuxYaV7ZD8D/0o+
KmRZ1EOgqTdDj6Xdt2KhEQFhmnVAe+zX02ZXbcoLXX9MmOU1x0cSuA86VNppU5psO4IlZtJxPWJD
suqYf1syEUAj6vgI5drk9DAGG0aCbV6tcqdXKhGzJgnklCEh70dm0KMeOmCL6xaLrUEMhavu84rM
qgedK1YgL3JCSHCVkYLRFb3Fmr7Eo+KOD/swaqZ6tpI2djBi6gshFogNJcagWN6ZrW5BIo88IeU4
rv7sv/aauGIjFvl5kOK4jPAm8c42rn80UcTBNtRT3+hcSvvJijJFPvgY9MXzy0mxEf7yW4RV8ls5
sPs/dQ4hcS60chrQkz7pm5hNYRqJ7uTgfy8WZvmAgeW/EgUnBYlzNeFXlV0yuxgDX2h6BnbEWB2W
6hOR2KDH9omcdnemSfbZtLfunYm18TImgAVUiBCoLh5i8CsxA1vIfcAKVEiG7EvDnMTYSZRJXdMI
+EQkRdbWlyjt8SPmpPNvsyV5d9ZsIePsD9F4Fc96p3DKKcjNdD6X9pErGpLEVyeFtwd4y6JnFrIv
81qi9xkis4QrxQIXJMpcvCpEwZ+70oz1X2YKNZqVa6wJDrmCc8jYElwE2o+6nQDNhHy/bluyVzrm
fX/hwAVGWZNH4zpc9lJSKk6hm89k/uIGJxTdGvvHzasKnacaxP0+HLVGHqwt4AB5gLK4wYvvXTfI
tt/MvfIkQPEor7IJvgVzjVOP1nr67mcXouWnbCw2BnuDSdWuq/cimhOXY1aQESnc7HWBqrEbo4Hm
M88uYrC0jLeQm/0dATW5OIvIi/fxzmhtXrAxuSjZV6JEEC0pubmh5yp5Top6DN5VutsWlMVO6/Pm
k/RK34XkW18N3NdOF/wNNb8Age81zv+3mK3qg17ssJ31quXeOesYgQldOUgipgRAuBnvqXQTSMZ0
ss7aGpXEWu1I7V1eJdMthXwq3i2flIqjfiWyFLuz17xutrAZKGRgZ83UtTzDGMqY++nCycLvktOF
E4Jyf6Na+2eMUzgr4Mvxzvt1TRFZnkDsF+GqZQy3Up3A00A5f12vyW+QrZaFaZ68MZAJKl1i+VOV
NOFKMgE+3XqKTIChIMuHnLediyh8Q7XkIQ7Pdo9cAvVb9uTG1ESvGAFMEkPp7GUylU7IwHE/65HM
TU1IJDELvcpPnD8u8kKVjupWjWHZ2oRJOYd4/DgtjiCCpQ2lfn2biLVItP3aOfNZBH54kWyLWhra
o2+HuF61twE0rKp1C/oXNK/FE9udF/LkNB+xzjf6WtSAiYaTMwcs8a69mplMLToyrOZTxsK3ADib
rOFFqnlEEuMeJG4FFDtF6v5pE9H0cfWnoZz7AThmIsqkb2ZWOj/fm2jmjFpvpcFX2w63EHeFmpK5
hLHKNYtd1rUboaN0BJUOoUtQriGV2LfzX0RU1WKn4bNvIKO5CPUMlSErcQBWVsqa37r92vu7KPS5
tcfjkmPa84kW1Hw1LZSYWU/ClUdiC30rXKHK7u/JzErdD6ECBJGixiDKE2pvR5IEgGKOLzODqFgp
g0juLDZzQ8cpC2E4E35iTTgmkY1+k1flg9EKZ3XKhl9V+4p/aQdfR9mip20RrLYAkJQgHb9R82c1
T7tJJsL0jO9OHK4YD0ybvp8M0n2Jp70bJCTX4ZQ2zHhoKXWpCObYiqh5UOd7E7vK7mueMhoRqAd0
qXGlUijrRJzg5vofYPIrtMM7V6wsPyi2CFVQKe2uhxfCg15N7vq0tLYYVFKq9S1bB6cyTo+YIi5M
V9dSnaoQwSup1mTQKU9npKKzffa0PUruBTsHngH1RGTgmq9u93+QD7clabgF7qGZe3p/xjf7kEXb
Ez3EANO1gCkKO46IANom9LnBlzievQRTKJAShBjPg3cR+aG3TAdKN4/2CtnYwE350UcqHQ9nE7Qg
VqaPdTjO4J7qOnszrI8JMWYFrItSXkS+2teuM7Oho+J0Cypep9teXrwed/QkZFNWJl4LDpZY43ZA
Wo9BhC40uU06jqLA2WSa/1A8eNGuVczGkPDmCJQD3jGk1ejDAN6EYV992a2E1csmAShDmNr4jlnO
XWseDsDIz3wcaxMkFRM5Jf+0vAi7tpL7m6t7QodaTo901m1rWdQSuzeROGZQf5jqFlb34+ghGtYb
OoDwRVhTJ28Osx44skdqmfe1G0W0iRtNL3tJVjr4HIsFZFp0arnTXSTuongL1oJJRRaqBljaD/sV
mKCeE9gDSN+Kl4XpZ2evJxvOabcCRkczR4nXaNVWIQUp9bWTAH5Ht5M5x8GsExh4pLrkhSylt2gD
DP14HFwatIoPHUs0hT6ADLAVQvhphqz+Z1zKY22TRo8XVXAIpyc27PHi4zqX5d7K4/OE8GprX8aD
pYAq6q7kB4RXPoCrm0Xez5VrfC4O+ymqoQi1cDR8rFaJYJ/WhxBQ2ChJYvcOTQmRMNTUjZd/l605
DMJcuGXnjhKQtA5g0tRo8ntUzthDa0V5Nc3c8EwirsiJGmZYCtHMkflbSbxOln2rA3Eb8A4zh3WQ
l/lubtWULjnBjmUJq9hbsJw8zdMSgLH0j/0mh/K/xp4gy9qd62qXc7Mbrre4pu+8Dd8G1XHFrfn5
ymoHAgnUpLgNSzhzKcFI0kIgnGbWgfKFZR3ODzgHlqKZ+pISQYpaAA5+tanvx1h9yg5Alux5k8+U
Arb30VMmHXtbz335K4p9UJCODKXduaChCKQ/Bqvu7+aNMPxe0+dB5n6JQLRDqD3Nu2/+Q5XsYlNQ
MdrfmiuLCKvtBj8JcnhKjZhMMMX0Mq3aXrBDTGKD8AHmj3Kg/A/8ticFAJD7oJEKK56rXBMzubCK
TfaFc23dxFrMG9uWOOcpjsv3ao7nbBXPxdd+lp8tFK4TE2HgN1Lrjwcetn0hNb9a2TA7KHcKkIa+
liKdWBYUkdk52AEXh2KDX6uwHPgW4M8rypMJ3nkOza72GxIJHgi3rOZMO/0MHh8w4b8xulPsh7Nx
ssfJbYFHswKjERvvT3frATGQZq+HM086Qw3RbDBAq9gMCfGWn+V0aatG6haSwCbzXZ9UpaeYWgFa
2jtgqPOx2xnzvoE9LZTXT+xVFlYFkK/sNheXM9Qh7JdN8Arxzz5/KEEwAwf7DdCxwoH5pBTPKWaS
+/hZvtDM6RkqW6lxnQtULsxBQUxAczMX7qNPKBLinAS1LbaLWLf/M29m9QqHyzgG3FPoSYjK7SNv
7G8io0KO84KW3rE0x5Hf/dyKckIt/h3x22Gj3c0+OpYju+flwEDr8L2OdOLvnmTqa7z1DW0U0QMb
rHlo8A0ck3F0nbZYYV1IKQ/kLt85y9CAbSs/o1EAGFBs+v2AlqLdDZ/NWK73KmFSy8otIhEFAfE8
+8ag5fZob+7rU1fn+KTRvVcLa781y+UglfoCzHu8wWRvqCnrORN5Ra2u9W+Mvn8Qrhx966QOzJxd
ZQ+h8B/2ERsCcn/W6NpVsSO5+6aeKe4h7S0lFgtyxvZcEwQWTe9Bt8w12HivEy/Vm/JRkcserQNr
bkGezs6Vq5258npi3hkjCx0ibJFMpWXUOTpARNeLRLsJuAAUJF1JrKflgRw/kslEbWSibnAj8si4
slKrjDt0x76x3qnIMCEzUv2vxaz7mfRCncABERzieQf8K0phVaDP7iIR1E4nD1Cra9Rqflwr8MEe
cgr0q3PQIcdRzCbziXsCMTmxIuZpQI9f2h0+XeoEhRWVFqMSgY1s0J32c6sjHbYvKC2AZE1PEGZs
EWnyT9IbTnG6x5KeWgsEIZUssGO4VYr6RdoNudeEKPVNONEK2CLQ94wlQdkY9F+Wp1IPkEMPABD+
HSxWhO6TFaSXFe8eo0DzGKWb820HjaicSFniXPRAHRSAOwHrEgqvVHPZ8emOniRluGyCx+i+CWtq
SzE//rEtR6GBx7jljdOYgziFdhhyYpmpacmksMyOwEKf9eNxQ3cLvGA6xMW1zt92GwcLxETZkV6H
J7VHwpkWV6mwU3aFNMjHsZNzG6TKuAuGVhoh9rxjI6a/VzNAlH8ew8II7xLQLq6DYS8ojmqGK7Io
a9gLCnyzSX7KaaYNjBv/4RgFYImFeIEqE/R30oEW02nHaPcE2aeORaiS/8WKfIq7DeNKHs/OiL4K
khQGPO6sXAQCuIuFRSnGNyZqlnoGXR5bBNQzq5E9WOhph08zL1jkcdLujp6/NAk7tmZlZzq7hlHc
E3BaaQvLifhjz6mXFEkwzLZTw3kVjJiRiCH0uYP4Ul5K5IaYREdysDrU/peMeh+YQL5/1HwkDpMG
CvfHqHHMEXA8VDmsmOc+bPL26Wun8ACk0XaSKuAYIYzuXESjy7qkXHMFUIcQe+i2W16WnD4fGvU5
jqrnWqSyO+mH5k2/b4+Z/8SWYv/RaaEw4XycJmu0YsWIT3qkxUeeDWZ4mzFiIsEEPp72pxWfel/q
u7db1IVY/udVqSlQE4TQp58+gsBTKTDI6EhP2RGPYaXS6WiKJIRx/lPC+bxvNHY6C3gke9Gtuxzs
trasyjHkAOXxp8nWgU3GWA3kNxYPVuzrxpcZi0TBuRq9Zm/tBoXHU62urVDvKG7YYYRweY4EQUII
wUT4uQXt1omawaWGju+YQsaz/wImiNIK2exEXf2ErpP3PDkhLq0UJg8j4pRQWGomBC0neWYfHlLE
skBvZ1gHh+fFUy72FupTeyjIfIVU1J8CLFQ4h4I778m/xVrhEQyvH5X563yWuS74eJzgRS2MwEgY
3+Y9R9dYn+WFF7aNhdOL1eKc1A9o0eAVEPUlopRBjHB/qCEcyQOOWgycdm3ZYrsuyl1rh08UgpYi
cX2azwfk63z15cJHm+f14v4is/F6ItqcFWnzUpGNYDYIofRwtDesqjbRjFebULWWvQa1QUD3POs3
mqtt7SNMRCD+cdrE5YCeE5HuVm6bYBA0pe4eQlu4+IHQaxK75Ma2WQWVq4uxNrI7hTNjwritQ6/a
Eav81x7wXcvratcbhF3v44Ep8z4of8v/EHyfu+P2vBU+N7X/+R4wODLeDLZS9CZX6pzgdEd55hKB
kqkOrRWDKu4BQWjVeZHD9UAog4bd8jsccwzzoUfl9ibPUQ/eNIwaM+shTNsPg2M86HscBPiLgpe7
RQrTsY3cZq+MZYQNexSSzstrJUEBeLiTxk/6YIh4ULIAEB2zxdtHEHOX1+SfpwjH/wJgkCdE5KDr
zSR5mY+aeG7RlqCKIsWa3O3+6REG7hav1ej7Typx1AQjGbC/x8Bp58FdgqTj/XWPuUJJYAoYUihl
d/4D6Wcpa60RAALxNYL6kLxvXFKgy1YYjITrqFaGonOZ8P/c+0B+dF/Yq6r5qtWty6nl8LQzFKdn
XKmrb2ZNNbLchtLvfI/2lK44RZeLB+Jx+vlyAVbra2kaA5/EN0XdmB9ouSbpJ/LOz7CzyRsjRkIo
KQD4DvlXM6eh6PiYTzFPG3fScY7R3v8BJxIkqp87cwB0qbp8cqGulf4M8e8QmfdqbwQQbQJRKhIN
MVvHa2jNFG0TPSezNerGrkeKZrv2aYJlPE0c9Wzg4+tL+WrKTl3jr1X9a1c+igVXZ5ZSTJVNvLfB
vnGqiQNAy5kk5Gmzv+65PUdYsWJAdsmW4ZGW8o8JP11h2q7xsyC4yAUPWncpVh+MLLhCj7LytNpx
3T2+fIzEIr+6VsMeAB980J688TcoA/flg+LXQHEyGaGHkPg7Mu1v45/VPPWyK0p+lZF3SMCCOaaT
pCNUiqpU862uHzopaTCl+VEh4AtAkDowfUno4wGOtAtznhlPBVphN10LZFiA53yCdWzRPgQIf4+V
gFDcl1ASTo/uExROCeznGM+EmZWq9qpjNFnRaxD270LUHFLbZvDMXguHHbavmcu/qJhoj9onM74s
7ghUkl93V9FfesSBGmkjZVgrB969axuZKzVBOxPGZ3u3gawFCjQp0g3LQmIwQH5JrM+WNjPoGF/7
KfWJ2gpMvLw8MWHLXzxqyv491/tRUJuFPK5bOLnXNppX9NWi57kXhFUufsSYbI1hdCO2VwIu8PV7
2WzKwRt/v06wnOKC5QXc079IGAFgXLcjIUTRF66E0x91RxKWzPlqsT7aUIik+C8gzFTiJACYRQty
Zu6GI6iw/Rgz2EQ/4lN6aBYnF2+dnYYrsAZEfRtSzTZU4K6YCU1/2vCnLQdI0oiQtBrXsxyV/n6k
eVJV48DnF0FVYOCaHPkDNeSiuNbAlswc2RpqtELuhAYsgSFK8e8xOyXx5xFnKt0w5sTWjk7GmoOD
mdczexLhiV4NAuQdEJIRPjBdjlEcclLc+N2xbmMJCjiX7Q2KGx2X7OuGWo6+bRMiKx/YtqdKK1Hl
cMYEyDewOPVsZT6D+Ktg+4u/Eb11kLGk/X+zuNqaTFwUxcuou414S6TQaw/DaieHn60Bqj4TRgRm
HeGRPiVAnw6EBmOfluU8vIPcA2gdCNtGwrVPMWv9xsehtJvb7YpUdWh4bjO+9KT4xoFW6VOiiOvi
TuadA4tpaQKo0TtebfJ04btqeODc5PCyw4hUe1GCzBRQ5sacGOCuIb9b67dsAHb9wDw4f8C+W4Vl
kXmZYA0mh3fmEfQSp7ftSIg1AhouCffiNdm9CYDAHD5y1/Myo3ZvabQmVZfaT6dcXvjrCkW2ZhVU
CAT3gkKp2ZJXaa6XnNh1k3WdZWmzMDIgyB8Hf5rlMn3ZpY06QRKhMfUyOCuTIXZXOczI2cIpRPQc
PCnoBRk1UweX2IoWOrkmlmeWBFmFA8AD1s2I0xqil/150Dhz9LQPeAaNPJu2hvDQnrEUB2i5RHKp
QN9ixNu08/2Hez6YrDhx1re5Z/Ab0YyHmAiM3iBAGigQQKUXq299akSvPvO15ZZkCI7Om7tF5wQ7
gCh4ZDVfFge6wMxYO+jh/MQdvbd3FIvl+595v3cJpzY7RRAG7dEtW64JYzoXKM8oqkTCLLzrA0u8
b+cZgSLva3oV7GQ7jUWmkmLaeWGtbIXm/LaJRKu72ZofGHyMUVFTQ1ROBKBXgSVlLHQVTTcMdtSz
WGl1jIl+1tQCzvYIZC+Eim4eVs2rVAETSsJ8qOFqlUPWiJu82JJYZUVjsJznDS6VoDBaWkGS+t5B
mU/VKdNw/I+Dg3UJFvU0Usuv7jutlvC1D4YuLJUAiXCxFq3kNBmPlVrHgAGrmiriV6nGo0d3RJ0+
XY0/xconzI7qLFVRmEMbcmRqRbXjmhYgSSTiPdbFtoDwqC4OcLtNTHsVPdfQyfjvWw/QZ0sii2ON
mpgpu1yoZCvXkqFgQwHNl1fwP8VOPIU0z6N/9oQN6G/8GT1SX8rSker1ujyF6AIb13dqf+Ene3z+
TehBABW4ffHZUbYb00luumrIQPH0BitlM01lrh+tIwwHDdOf8aRWiZ7hzdIV1VhyF0Nq1bi4Rxjh
JjwnSPTWgUPuL97NhUI9jIKB6PMuuNrgt2S5MlU5wgVPklwYzMP5UvGqaobctUX0UqrNriuSz6r4
0Jtkh0Zsbw7yKgdKzYrXNJiJwlRcbjiJJRCEA9tye2fSF3DkfMtSb9dF1kyCRSKmAN3SKT1EGSz3
pM1MVc4fXT1nCEy82+0fgcYhlHIsNHq6rnDJZdXvNU6MsiwAKqr49/4CcoX076GOhenx6on5rSBl
ZhoNnYZlrbtTpHtVsERF79BSwdpTQgOhofj8icc6BAvWDfELx2HX7Pe1jMLuklXlASVpzNbqEgI9
WbD9QZLIULjoh4uWUu3JQrVWuu+FYGKAX1R7CDKbOrIjHgXPoEGzxTnaGN/PMeuCvlqtDAfNQMyu
7kjeNMMRAnw1N6TDPOW0//D6adRJ41hCJ+tHJFEZdrz+7pB8bI9QtyQt8Ge/Mdkp7Rp8el95DPdK
JU+lEDh1MOIqSQrvpi2KKFj8+/Qn2fwLbnBaMG0GJQi2bDWJzs1FxTYeRRqZbmVQ5DHef0tEBmoH
dZjFPMY8uK/wpHG31WNv6wcBJ2V5fJlFqpnLkkTGv9iF+pFz/kpwSezNkKOV4LGo0JFOv6G9UVep
zl2zHv9bQHfXUbfSiT1CCxmndkvPYGY4hejEhXK8jS8PZ4s2r8JgZ7v+2hIagghS1zYtAeOVQHT/
xCN7nskWiNWWuMDnHjMdRy+DXyutugc15SGAnT3m1cEQrwuS8/T0XQZ4fRmutGFx49v8ZWbu4k/S
pYWfakHCkKYtk+uI4QvRxQdS992tBnRluuRpOAU+4iJ95BeKzNcKLGopA8BMOxiTmyzkcFNpBcpW
zfcWTYNmXcJLYNlLnh7OcbFaAQnTjPjyOaQ2fFH5ECSpfuaWwIAPP6Ijfg4T/qx4A4OYgDe4Vi9Q
xDTMBgSARyx2yacorBVxfpU4dN+5FG5D2jzylDuwcelFeLWygGZpo2vhmA8W6Evy29NKSEBzwOEz
RpGESaosv6vS68EZofM1Gfgf9440hHtiusTUukaptkqwntpDixrYhBXwpxZDO5QbsrvV4mwfjJJ8
Pk84ecPdE+Eggok3C2pYhE773Imv1fqXjEZ9DAmdjiCNa+5MmdU+CNwgNlIKD0EmNrDmeZtUFDW9
md7OAkGc/IQS3kKa94qQzRigy+3rxe6nEAgBNzvDCJJQEPEk9SSS+lJMI17nmgDSA1nJ7JIIR78r
6/SCzU6Oa5Mn/8UiPFpOnU66INq0nsQAeiUIJU8wE68hg3J+M0ZmxbIDQXE7UZpRMP1hLx+NB2yS
lVNpHjAjaGPjsB13yjOc+hzGEuM1gRm4KbKZkPjwWjzZmdizMJ3cWiw+ZaqjrJnSUbHE8LvqUTUF
Bt0QdHReFx+gtRDVC9ZFtZGBEUVdTiV2EIe3kc9LA7MdO6gc4eyvWlqR9BW6CTMgvIwOb9fE4OeP
rlnfQjLIycsNdoYO/zlxAvhtctneeIXCgBnOfnXckkgePzr1mJ/a+chcJRZ+3B5PqdZTC+NV5+XK
v8tPq+SzWuDOdMbpJezxf+Mt/2axs10k7bok1tAdkZnGAANIuHMCmDxhqtKc9MpEwrL3kPgsjYZV
vKBrvu0CrqlnEYke3dJlmGefq8aop89X3ANII+dcdJS11Auq4guFXtxyxKQrk+4pgnfDFI6XbNwl
DNAjVjRWZYRU8k1WaqBk7KnSGncDoEOfJlFtSYGMeSA85UQbGru2UH1IoduxwOPUsbit+3x5rfOv
VPWGJQqv8kIiy/9lUxx+hqd8zAx0kyWHTJ2rFlyh+pLTRBf9Pa01rQLQJZ7hWNbqtpXBefiK1QRf
384crLOfbGMwUJgv03uu4ogcax2GaVT3+E675hR3r/BpTtKUiRHCoWJiL+V5fUF+1kB3oTSTz3qe
okaXJJA/Bjl77X20c+AQK7OW43+oHLb+3jJHJikZ2Xg/62jGgLARaZm9RiW2RHjUlra39jcemLFY
7AsSyod0mO0Fq28N5rTHjWHmmcy1OuT1StIgENAQTqHS7vjvWAVxBzXIwa2WF/4aevpYadPTc3cA
S7jhSsuTAo7QVFXznnRFFUsBW5mjQMOwwn1H/3s4vx/0lsE3AsI05IB1+PDvkJWHgsolWcfJpejQ
0FED5xBXqZtJJDwtrwbIunMdIf6v4/3iOf0QZzILnZKXAgtV35I6jncW0u4ghZdfKVxWPzKMnHAE
sftjtGF6FcYdDkncBqfuJFJ2y4woAE97KiDlKYNFnKJ1m1uYsnCc3XmGm3dYtM7vfwEVHqFE+J88
tUpm+kb2l+d/BWHtOBjXagd0xPV9mSFl28qh8Vf5msczw6gAVHs2YDltX+Deh+P+7g9KJcLVM1oD
qSevttWeYrqzlJbiyX6JpcsdpQRVaJLi/But9kWEWJCfpy4TDdkjhcJtYDEfNrbvKGUyXcL6VTAh
5eC+96CsMKnwAgWef3Eem6EUWg9bEBP3PPxetyKCxlU/qtiW6dlf3tP63KT6ciX4Uzc37GEmuCIS
H6sgOJljlKuXiLxISXk1U4LtfHCPqWhwfhWDv4zR58w8Nb7B1spzTsaFkjkqYLHVZgcO6ZU1Z3KB
X+vcPz0BwgAEWTtkq6/sd307HMbkdFtcei6jAS954KLWI7U6qn2qvA5NLUIZIia5C9Jz+jpp1Fil
AxHLgYHf4l/IpFngAHu2cWmVNhXWqb340m73f788kmyrjvqxd9+UXLoF0zjBtjLn0VmqZ8LMhxMZ
2KVWKWV6bt1MSx6K73lJdpeE7fxFjlfmRJq7RGUb3D9VYh2FoYY/SyE/jgNM7Hefb+bNAx0MSHmt
/jLVcz1DU4cFgn9N+I/VG3i5sIe0ieVKGmDv9XwZ+7nuSn5hFbj0nnmfd5YyJkYav7EMBgPeXdMB
28pE6TqZCbEwcU+nnqMdL0atYaXJCuYbRnpvjl9Rio0ZS7poSuzggdFmnFIppv5gMUGg58OZ5JdY
bKcfkfzIOkOk3YCzRQezHFqnei+OOj1L+p8ximCguI+O5sZFpouGVnhqM3Kpw89hZCQNJKYwZeR+
Ipd3brNB9zt4s0SCLzzF4oziemnvz9ZcFVRwzc1HXAuTifZcnVeKfP1CbQL2h4cXr9Y3hb0y8VSO
q8YjCcx28YpsUnaHAJ/LHMbcIPPeuiLyb1rZfuGf60KbY9eVCMQUwbW2UR9aNJKtrxmzaaw0DnsQ
GJ2BQd/UraAEvxRugoOe7+3qetc3Sf2wfeymnKUdPcqPYKQSgI9eZxvshHSaENhHaZesMEJrtKFf
InSn0UwXXuEw1coYanaBNKWo5CshLBfppR0lZVuc2lRJEJYosfWdCvJ3WGiq3WXjPfGhJ497xnuu
6K0RgRE+VlgAXjwnfJKqbahwIMkwKGHvbeZg+z+KrK1euZ9b5YA9Tq4KXeBjIe+3NaL3txaJSrYt
i2I3OeK+1/ppteMztuQvUnMt+9P9DEmjn9xrwTTr6WU7x66VYW+f/y9L2F8HpD3H4Yuq0TAXqnZG
cyPcELMIgErxXmtLXg/w7R5epBy4aCCOLlWgizKHnrzMLtpwMI+YAaqBSUyV1yvxqxSEF2Nqg/jW
8PSVyL2BSZuJXASQ5JiRZ+iAvRHza8T+FlNuqwvOIEjAmKcTPSSd8W//c2LSw1W/5UMt4yDyFaGh
Bz1P0dxjsFXIwi5HoU38+nM6dhtKdI4HLjinb0lYxsmSDvWzlSrtW8+FWmk+ZqKO0B01d1crh8zT
vmf0uAzuE1WsLmquO3lpbbERsyTOUvILNhObd8/RAmjbpLwuDDHEoqpLmPXVBFlf9hYSRtZ/oUd7
XAtRT9rSgAOLuP8n0dBNW6XE7jxcjj/Ig/ThAbdWBtCO/vl8DMosynAx29LACc+K9iZ/6UB+qnFi
nRZdMQ9lNYhFG/JP4FLeYeNoQxmS95wYaS0HrLqJga5UaGDVrTIsnyb7B60UfcmBN+rlOrTJBwfy
etNmfmlDoVm6k8kbfjC9m7fMBRsYipJZow4OoW8YBT5LHbC1JUQw2KfM/kPMtdzB+EQPC9aydpz/
7U60aBO1thwCNP7pjDBXzzUr84Kpx5fa/Qs80zlE/6MXXXXBz3awWZR957gJBILvn+CPR3MlEWvN
w515f5L0huCsLo4Mp5ogGwdL60HtdfPcB6cCIWRmbyRYk56eEk/pPbkJ9YuXbNV7hG8/j8nCs6S0
Gfooyq9qx+iJudyRQhYFQCKhSF4ksVcbhSw79fMSOJuB7CAgTJBXczP994Qj2o+UREEaI/KVb8X6
Fjoe+jfrU+Sc1sT9qNnHgtQGCGsM+2qdGYlu1zp2JK6IY0GFbdDhvea8kIdp0erI/eQboTS66ZUj
r2iH8UVhXttW6kgEfWbqUZv4JmwCazo9i1NRHnxt+LtibGGT5nQhS8fz4hFy114/Tbp3Gqtkdk9M
+JCanQiRrLYhyygTJ1zd32mCfK905Hx6I5R1ghUkm3DTIsGHr1qmVdbdsztUQKkd6AVkSujXONzQ
TgaoUJDEjxBfYXE4HCVrqkjKZsSormRKpIqgpyspojkZ2lHZIY2h39iMxx8DFuQv2Zy8B8xkE/OZ
j4ID4RnhC+el/POD46SsbteT/2mDSzUdM0IoME4uWO7gpDQJSlH+qP2tyhR0YASDfD4aNc9ZyqBj
ukgmPH0QV47wj5d2HjYZv007idSooE7ML6drLSYFiVlsS4gF7RuAyOUGraadZfCqX4p5vg4l40Oh
BwoZibjQLf/vROUc65fC3cYOcRR4dFFDzDcVgAaLlQ+yEiMdWVoZ1OWjPIYAQEzLvGwMq4CNB2KM
+MQff77WEhTqmG+JQuPG8b4sk/DydtnIbTH/VoOzfubB3AgW0zAPlphHP/1RPQLX6/LP6IIlcB4E
kK6Aps9a6+XYrd1ydzVVG0JAnLBG59bryWeJ9FgmM6jCzr9ATyHVVJDABuK/RJ1BQ4SJ+Milmsoq
NjQfjD31Z3qxdRKdtSex08mFGQXKLO70W57P71GzISuf3Oka38jWkrDLjbr0UErJxuYXJ0Q40RIf
wogPaKndNsfchI9SaqH2xpS0/gzgmCENpixML72BQTCnGNZsehTbTvNloPjsiPw/MJw42KOsLAP1
txahtrMAtalm3LpJ7m4Eu8hunvfKhgGG+KcQv437clAiGvad+w0c41BiSWuhNONuAr1F4kPCBJYu
Seki8TVZXrSy825xlxd6rJygpqF/7TtLxnYopeqje3iKLJqVywn4xCtyU17VOtJr3ZJfgTS1eoJ2
FueBlMj+g4RRZOiMGhYaFPfRdjT4/z/2hywhvztLV4VtwP7GOgPUMPPX+ZlTKJo7wY7VCttz3P7I
8r1XUS3gp8pAsTBclWF6qCllJLN1yU2x6HqpvtkgzCtWWpPIMWucc/POZAHCBn8FreTxg4iwllqo
FA20SHzHk+VrHBIa5+wAVVKJmg469N3fw+peTBv32Kk0oLWCZL6JuKOIp3+WETA4nwqeZRykDVbF
77a63wryCOjrMz4Q8oaoOGk4WZbfabaeYfnY0+yr6Mnfo9EqskgzdUrpaX4KfXVSzD3TcDZtcfE+
b6PyL8gWUzXoIr92vnyWMSn4v6clxmaRwQhMocbKjWo1ZKBp5NyBk0s95EluC6ZQpbLto4CS5pS5
Mw3oFN6h8obl+8cltqX0o+JE5wOP51S1K6/yvdHRh19hfBy0Vv9nLafDgIC1o/HP18XEg2brvQKq
9zFQ9Vww4gNyOef1cWg6uS9WyknMx2//uaDoexih9IzEUusPGS+tqXXYGrPThJR4guW0ZwhnQ+dp
sBhOhpzULm73a2o+wrRVZmb6rJtlKlnH9N/cW9orDIkwDEcVEBQQ1Rg2LrK77cybqJvP+waLOM8O
ABYBKEdisvsQxV2U5IjSGiINApKRcNMJTsBan/0oMQV/Jp+sSPuLPlWSrBCCpQ6VnGIONEhNTQdt
3IXqwj57TqgT5ICsG8PL9TvqFWd4mFFsFqRDl78OIpzPjxNEzUFwttZvQyUfjP88wN4uQAWBTD5G
Y+md/dE6lLbrRAd6k0FVHg+b+S4ZNnH93y8b1ssoW8tAtPCe4qte+9qHE9bjGhl0e6sCHr/8KbKW
vHp/v3SuvrKo0kHimhPMCBbYsYUF1rCTteYBHF4bBVQEPWqKloDGh+qS2lSX3JKFDphfrv42dUC8
Rh5Imj0hmIjjJbRu6MQjPsv0ak1zYZU9DnizeSMc/u7XFJ3YAvV7nfHmqOOeWR9Ds7zYWKvhGt2s
7hxNLr/Rl0viXkFeIoIYDfAhw5JMTzOwywTfHivDr5pfQhiHaEQ/NnmmsnucHNrXTsJBxG+pGVgo
VdQYPHWFs5D5NPhgbYgmgsH1tCyncDodRtG5pLnTnEvppZpDhsvuTcMVtuzZb6yuqC0DWmiv44bn
z9d3uvfntfYZ0s6LY5l64z+HAknNixHWAl3Rf/QW80UGFUSn0vz3oRFPdQI4xktO0QT84b2y6AXQ
xcZzYdo4QLmt8nAIYGfG0zQRlx8D2ArsCjtDLDdGDdt/tKKEPcuby5qks3pgKfZfNnksRRUZL3k4
7lTUHeRuJj+taVtk8PGiIzM9Xk2XET2FpMiCWPtXbWWldPjsqWOIWOLi+CtDroL/MnhDD+M/2uqH
EzcwxMPelIe98lxAf7yWa4FrHBzAArkMG+UiW+VBOQ9sfgJEYL9aQekziB/VdEavGti7VLBn1LZh
CET7VZcOzfXY/dXsO5TCfF5ox85U0D/WNfne2BvBVH67y9MkrIQcKFDnfPJODv2gHwXu1jHcHALV
mTWfw5fEGQw/LLvyAnZOaFVpXmegnZ8kGe4zsOtYes6A1VxnCX1urkgXogjtG6E8vNZgAtpeWH1i
qfq4yE4UVFSYVIuPkUBGrzD+Oy1XoLSkul8Qf/RgtcScnUMdkGUu1sBh6tzgqK+zIofPXkq/HryF
F/gdMzZRong6gSV0gsspSEQNvRnWwCKOYN4K/PdWlayhFYq44YrFCX/1ydOelRfGl0jPlvXGjiHY
9IlugrABAPLMWudgoYLah9kHd4UTTQvx6YxAdVSho040/SHE+zk1h3nB6QEBMu2pwQu20SGYSe65
rsckSfE0Tda6acxcL8z2miR95m6tjXhdspfQoLtELH46xT9fKnx7PrdoDC9p19fcoE98pV9Oj0qy
opsHdftPldGOFqatr1cLEVMlooMQTlLHxTLgbmY89erqde8Vom2v6L9XH2IjskXa3ASjaXJPrmqB
rbnIV2HcNxYtGnKzTazDe+gDgVeXph1i9xIKq629aFCM9+gfRF8PWFm95NMjyNOb0j79L0tHqs9y
Y3vVEvaOdWe5XcEdUIJDupHkS7uqDEnHvjoktlCSk5WWbxDXSOJ2/wwdUCRHDkLOJ/pBpQL9gHJ7
07fGUA4o20U/LHcOYR/mxnGc+aQRiPiaY35zmE6F4RKx2TCGrd27TZp7dVeUfD9I2BxrHNPrspXI
ykUG69kqiv0AXvQtOHAeIgHlNPM/IFQRZwqlvxwmKn3mtRmRat6aJmW5Zno8PIBURgVMO9EuZrsX
IQ1N5MwCpPoLCz4VEIjEshtdqWkJaRpXNHXaZ5htaIK+W0cpbXXKvRUMkrm8DdqhbYh7QbsWlSON
Maf26vly6ZVuFub/B6Z3mBwaomw24XvkzuAj1yMJuO7zqMwW+62YWaBoC39KNant6aPRGMjU+e4Y
l6y0sJ4yGDbq7f88HWeF5KUgSALY65SlsFqwzc61AplWGXnzeO8gdxOrDFGUCU98C0AN1bXie6Jo
nEkP44ybaztO0SkJZ1kNMvqB+zyUCUO/5hBRGV4zDdK7iK9IWLEhUBXW0hpR30/xLmC4c2XtKekb
JQZzUwfKqtAqbc7kwujdj6Mb1Yptv8EGcs5q96Vh3Z4edaKY89VxznaeVXNBsiCi6WTPE7s3MD3c
fzY/QmnpI+QFPTUctDQ4hS2skYevgErtqolLwJsKfg98LJHxJXjhGmMVe5nxKHM/tpFoQlsRIA2j
JuUrs5gym742nAZhTShQX5X1SCYyAwB4xWFfhLWBCYRxz2QGHhazMoxHsJNoV+1tB/YupHTG355W
eFbuJIrCJflxt5Huhs1FowdwnOrurEpp2qC5UvjAMIW1WUyIlUFCI/ydhsDLKK6M7pvvgqdPDSrz
bHrbUi1lcmRcxuwA2j/z+bGCnFteIHL3zRhJLHabWOOGcyBn2fVpu62bf3N4Bln8etFpTjRmpkZu
yd0FwRB+TS1ufPJy0WzBT3/Lc/B7/TqZnYQP8aWAn4yawtRW/gae8ly1VhWAt44kZWGV6lGP9VZj
toEdfBJoEZRRCR6Jk2Pn0ccir9Mud45wPmRLe5kmT1xM9ZeAf3T4n0u6qZ5bQjRNf6nhpgtrFVyw
qg3tEWD146mrwn8WA9fjhYfh9zZiqspG+B8ACFT+IW8gMEkbxtvnLW6OM/TS1QPGIcfPuPaMntG8
8DDnlx6ZXCiQMZxAYrFyfZTEBUXEgcer697wqr42Ck9g0DOIpEaGZEs/Y9noDqPIv9cqIuToU10K
8913HKYqRF4ZfoMStBHqH0eE/cmkunbosaYmBxYbb+thhL86c/MFlDIzGt8EMKyFyR6uuaP5XyYk
0dVHe7LioZzPyPoKQ8x1OaLBHVWozU3/e4SZgWoJXzF+O3Wn+Dv9C7c0uQHrvWQskYqsvFuG8MDX
n8MKmTiKHxV5azEGMDS9duJU3Va+BhBowIbXdsUbli5WtzaAzbMdysvmEplpzGhP+hXULdK4OwNJ
tkCuhMebI42IkKYM5ntCx/wj5+xHHmMGMkhJ5GRyIZYuFDNM3uLzT7yV3lqYcGNC3Kq/HKaErQKh
nSq7c7m0P+sbwsTBrTiXsIfjkbUpFOSBmx7J/kjhxexfZyx83D1ulSnfLsPpDwrlpCmMMN6mJ/x4
OynudHHug+vy2qQ81cGituND+8WpVDyRa0Wnr4mMK0ckXrvaCg0iUgRceVExOq7Nure25HE9LqPE
IoYovDCW7DC5w2104OfzAVj12X8JRA6YZ6/LJunArlJ3pZs9RDowT+y/f4/qbMdCQ/rB0QpOMKEP
mPFL7loJtXHoWf/6K71x3A6jDoBvaYT1TBGAiz57I+HJmPVetE6CplYxSGfdaITf5c6NG1wr1MN4
iDfGMkA8coBNadRKT7w4+ZFbG+UfZ8vgyYj/fwuXVbTNt22rXRhFC3FhDZd30vi1rwRUKzuV0+s7
XiRoRAdDOd4sC05a4V7cRtW35hlJNhj/hHFcrbmBs6iPQLO58txWfraxL2x6wxTh5I18EikZcl6L
I865z/o8KYP2lVf5LvSSLEo6ecNOAb2ctFHZiwo2+JUzsujSMLMlNIr4lO5IxGaf6Uf4ig09LObR
xxnTczSqtELFlbDlkwlauzD3Gv/NxO3QnNT6FufBpijOzEiZ0nIWT6xC7q9P6NzTrS7WoVeNJyHY
+M/IzHQs/LsxTGhO7CM/DVvrkWyYBHyZF6tYTARP0XaNN/z6TD8dneh+/BT4py/xkmCLzLTkk02Q
lwus5XrMN3SH0CajT9U3zpaTs7cVUrlLdKYOgLhDv+KlWHr4cEvwC/cJu8SevcJrz2DQayUuxbvt
vAvJXhiFUN0mB04FnmHkitj/4XVUST1NYXIP50owlK7AsbnoDEbVWcGTVy9f8m11fyOghcaiWERj
FSam30LzRNNNCWBqmRpNGngqt1anmdWCS9Q34RSCexpZtgS7Y68QIOOMBUt1vtsZewhImIIk0/R2
GI0FN7gAHXmsT9JfqmVqvL3I/sck/O0doZYuo2Vjozrq4gtUrouVMhOVP6rkwonqPX8tCkgR/jsD
aUJ9wbmWW4EyQ7rTsQhyX/WdttW5tT446fe5GrZggTQ58tZmkHICrH3XNd1lYtqjFGN/ZEW7dzhL
OmIUqigtQX5mEV53aYoeyu3La6BK90oCniav6AzgM6/DlJc6kfYKBbXHvqYRKEoAVtUW8hcylxnN
AlUq2rn9t2KqBA3SQZgjRrnxT5vWmAVvM+M+92+2veX80lDag/4r234BxGxlP0wmpXUP4i7DyUff
JpJ3ApoqWN2qRr/Asuzq27UZY+paY1UTShLFGMP1MvAeMrMD+P/JMdEV3a60N4resArXxkNe0VAZ
XUAaWPKBco4v4ebQ49vwftpVz8Mie5FWV9Th0jaKwmzxnU5349kUS3Vp/mc87oSI+tNCVj67NQ/s
N9hROomMryma2cJBbhDlKVJLSDrFijnRolLbL5JiN3V2IkkSzdwlc8Og+wQSWW4VDztLyUHFZ6N0
UB5s4HmoX9KKP3gKNnWWJOpJ8kf80iLR6Sz7qpVefmqTvXDOI7vvk4Jqi9lw2d1LKqCWOXU8MONO
LYlKEnBmZ4CF5AXjQ3rg971U5fY4DiCGogM/zkKpO4dRqZ+zTWB0RBgUN6rogvufyEeZwmfdiCZ3
M+qX9GV7lHbtR+aNh/vDCv1TwPMM8nCqPd+kxL0dktpVTitmLsMwBmVmlmJVmVIcMsqHJt/J/JP8
DfShc6d4aEf9o/xnurZ9ufyJfMXBuvK4kXl7sPzsay+yOFe+4p+70w8dL9+Zdx9DNNCFgD8f3os/
kWIUOs0veAgqIteqcA03BizG0AWAc20qpDDlFDT3kwTz+dZONcpLhidMtyYaW7uKPHu3orjwPO/H
8er7yBV6F4aytnF51imgXE/I8PlZN6YE/nFnbBqTKItH4/GJbAWP/w6SI2LEF3Wkxzu2IICkW4sj
tZSAUwCk7UpjgvpV5pn6n/PTITZ01BClVkxK3bZrGe2KEHzRADyUnEAKFxp7NErrWsM4wS7heulN
HvoiXPfSVeEp2WrspHPf0QUe970BlJj70S7Kpg5Qk+WdDDCt5jyBX4lhBNrVVlofwhaSsUIoTAmI
9yBm/Rx/nmotYc8MNogSB9FHq99CRdtvdbEiozhfeu1eFT0b+5al8ubM5KHiW4MHiomSi0/vVVg2
KZKsyUpwxrJNo1ZGf1eURTvA1na11Yhl62j73gqOwzOmIE3+NX9TEwGJAh8OcFxT69ESm4spZwfb
yNmK0KNT4u5cFJYRdMnR8tBVPB6iJz0wJXmN/LX2B/Cgknc+n86l7fAYmwkZ/n+d2Ve/OqAtvTnN
jwjU02UASCoZqfaoESxp0saM7tY9tCAvBz6xJi8/H1zyl4ZUSkAFOBIoFjJ2GREFXYqAVQAyi9/L
z4Dx8Asl1R4LzorLyX0ZAT2PF9estLPBzuHeWvA+081wdq40mhukIP3ki0mKwt5XdA6z7bHwPtjh
mKeRH0oB5xqxguMnAM3HPl6R6h/Dq8fu0/3xXkYuX6YucvBA7lQetH7mwyfbZjvdrjsc2l8lSCxL
5ej3lzFdLgGKH2VGMwasI04FG8YxBIZ11Xt4j/Dw6ztPTgQPetQE+5A7aUCiLtPTBlvj8Rqjy4ji
7itACC1YPgHcXrhPt+Tr6JgtQPVrhwOMmXvOyS7nF12rVSunZ/l0VyE+QX029u+hayfDwSngDQJZ
Z8ZbleU8AqTK6H6fwJRfMxx4FnV7rNnFtfY+hMKn6YgREOH85FcVCF9wR9ktw9aaJ94sxI4JDKs2
fGw+gixymsAkiBGYdoA70HW9yRWGF86M6EXEDpHrFfCOb73wbU5ZnIlhIkyV0AcacVK8nf+G3y5L
HyqMPEeWAR9xp2ONUxgvKsJ+5AEPTPxcBB9+kb6v4tsbRAliEBF0nPQGcMQLWHCfTuXErTBjMLEP
ykEi8/c9WgD720XM0l9T1DPPiDxqyYfLoNGgmPVvZS1RjtGqa3ByPhVM3wILYfy1jXjIk+uBBnGm
hmi/N1fITLpU8UJLE2V97BGptXzCOFSqp86VC+g+GKDji7IGTzVKtUP8zSF2mSAj3Z/YxYt8I3Ss
M9wfT20IzAY71tRn7kAlMHo2b6lTBBBx2x+R3R5tPi6BguP4V/XcSaPVTWfFiTbK+xLbSMyaGQsP
FqouLogcGOMUfJ4vJ+FldzkPoafH/qOLfGjIhVM4PCrtw5KUpgWCzvMtkcHhlG22hvXpEUThGgmh
Xe85I9wjyl87/Z6zgMwqphPY8kmmai6EDbx2goK80szRcKzA4j3h+wJe/wDLPK1wkPN/Ax2wFLS/
KlsyK0WH0I23PVBJuswh49TDhdLLGREyLRNroweK7Cqm9o11VMGK7uk+THBXuqe9sWg/gckLyK7E
mG3sufUEGHMhlOtc/shj/2FNduWzgdjH3ZMt4Sk4ZDPPfs/N0zGCE0lDTGFwZvBSZcED1ZVRUm7z
rO/SD/QN86JFIhq0huO981TvkddG6zFMCIebK/jBgHnnLNR0EZO03zb9cP4uPRTeO6ebheZVvBvv
ljg3EX5iNqmq64qtdBfF9bDtrpcVJ5ExWUIAZbx9pIxR5+Ha8gHiQiM+8OOER6AkrYnMwJGkqbr9
LebiJ+CWbdt04edx4bCTHCQDLJKigkcYxRPV4ci/VrcV7Ppm/bud5I5YYZUaQpBHyW47CwZN3hwc
yUPtuyP21hsb6rjsWIcMN5E0yoPYXa93gB/N7wKH4UYPrABmoFPwsxXTMf1Oc3LWpOLecmenavFm
B5DCJK8FlrZBVUENNezFdam3d7WCY2zfUfEX9tMMx5Ylidb2bqRiFlKtE8oHKEgSc1Q3H2GBgGI2
ZG0xEgLg2ObPWiRU0YYqgeBNpmzuSPX0YeRcLQ/aboX48L/jHFopdwgq2EivcbQiy+gzMryD8stF
vjHkkq1uVao1UXfgcCQYZbNSS2XUWRQ8Qk6iwlz61PKhupQCW6kb8xbPD5gzTx1ahQ91P8H++j44
nllHLCnxPSdldc7xd+3EqRhCKii+IsT2cCBfKPZiEEeDsBBzmwFs0bvTzynUqHPbiBBaLISAlguy
LprfcWd+q70Pm78k2gQGJC4DphxIh8p6FG/0V1mNehWrgUvY+WdhzFC/1h/b8qkLCakQXUaWNKdO
cAqLtQlN6Ls80HDebIKlR+4qzVrDiO7p1XTBE6dtAkSj4Sc6fqjseiC/WXgD9S7v5m4KC7s4AsVj
YlXPDJfNX02s8sUn9YH7CW9ESRdFUPNkPMagnkwHBxR6rl5cvxF++3P+meLTBMoWEJXQlRluoDY+
diIS8HA2frQRfGac3saWqdWWMdvu5XmxXlamoZw0yb6N0z/Xy98iF+cTz3HGj+nXvmZa1VY5akml
+khuOLG/SLllko/KO75edZ1BfGdpw5HgFM7eoC4qiZ5zSEg1MF1lDulN2xgzUCikiSGxbQxLotGT
Kxjqn11+DjfBPdIDkq9YOQTRbQDX/RuH7UfrlXYrMwSkyAoEIAWYG3tU7ytsU/Nlvlj/02cWs8hH
Qy3jNGfebdnQosSrFi4jimfHRR4jtVfutfJzy91CrslUTlfabEWvL3x1CpF9mkgcDSMb09837ZII
3mTrKRrU0Zioc2XTpBSLc8Tjqz/ucxelGOWq6u/dojJtmcDYzd9Yne/m2C0klp3jE0cSn6bRwjUt
knL1IsbIuzJK0bmj7doinxoxVluLfPJ2csbb1ghDgF8Uy401WG+T0f1egLey+CadSTnyUZu3EtFS
Muxwd6nbl43q2rNC/puuPeVst6O0kSvdTKUpJXI5dtLCkilJ7sYd/yQy31yjmDEsMSkF8bqCX6UP
kw6duBe99ybJfpJ6hNtARl5sg86zPAiiIfGrE89RmNRSwb5tyXfMHUyP6NCfH8Uwa3pTgW9uuWf1
efh1XkUN7/OECZVoJ+ADjNmnKMOD4wRXnXEuyLWwycpKtodFI9haIF3dzVYzvdNNwbikQrbcRBHn
18hm9b32TCuWNPgNs/viBJbp7ZndmRLzSkxCWfYi0nCNQiOPypVrWp0G4/azyjdVhkIIKp1leiUq
clSm0FccOJlI513rXcVOEKj2H6PlkGAg9IlZ8FRg814FsBHosh8/NrA5qzBPsV+zYgya1ks0soMH
TeSTXgcBLzXTibTQ01ejwaaqaDpMaaqxc2oHc1BsehH5VJ4FcxAQ5AalQ+/+NMEVq0espiHRFiyB
z3Pa4siUAt5HFZ+Pm39cUwykbHaQ7zuY6IaUDByVZGV0ZuP1AxAVzYMNs4Am+8LnST438VGF6JtP
Dt2mvjqX88GZUuxxUNGDSkYK6Y4N3E2v2I+Qt0hyCB3UM02BVcNUBuhFHSwDqeOjkYuTvVOKkNcj
EjRhEHsU4NksbJMqhkoANUyokp3YXcxsxVyT/zZ2z8UklLv8g5lqvBXvi4xvd/Nhd3mP2JgOgRIY
7BvwLgjOu1QORaJSk2wjiuYnkFNaaDxhVzDtgYzrtbyXlombvHEB7IDhoTjoeTi6ooVygeaVlIoB
tcwtDFrc6qR0+YuzljY05nkFXOHHClcrqZ+i/EbYtaqw9IdwfTaA8OjjL/wtVEvX6AgrGlUp/RGt
NAhGS9AOLgYwDgRl0xsyJg+U7eoiG+ABtgmwUORUQsKd+a5u37PPodYmZ+5h60eaM81U3MK79JzM
16SRYuKgdNLIhUW2b1n0agIgeFTpAfgGsvgLc2NWUnzcQlIgjT2+FkG59wwXzjBEI8BTiNWYV24N
GQ3gprDIngfLQV1FNiQlkSmi3fAR/K5fIBb5G+4NFaLBUlioU/7UkcQ3VF1U2nBklBSe3JQMzFC2
xyhLYz8xVOUsz2/Xfv8hP3UZMUk0Cj46PkNU5Q8yEHfJgK3Z/6wV54rwB7alNTeVNjSWmp8wDph+
Rs0GW8uhp0+TGDy7o3WubYKRwzKh2P/Bx/rWPvtMPl0tgEtJy+TMCgfbxqjNl44lTYu6/0a96vHn
eXUDnVCB2qr77V6mFoWxKwGmAbcqVl2klEsA9CUxE1hTVPfysfz1bCnKD49Nd1x7MoPEjpP52bJo
+0LLMs73WHljkKsZTcOheIa1uNyIOQnfD8WFsffNjg+pUX5YRlzR1ksO8rTLsD8dHPggp48Asz4C
ZO/quHxCS9ygM/EWUg+LyH1EixJlXFTk1gOs8OlSvMQE7lERPf0aNULqqb9V1bnboA8MsV5Vu5m1
+GM0jk6ujR79kt7ql0ZK09J4yLlcOl+UsZYxvM9kSe2dVGdspavZU1/SlmGDAHqUmvbI+dC08ubG
tCag81RJD2yJfI2n3cwoLsFn6JLbnqp1hpcr/DK+lap+7AI0+3AWb8tOrrhB2XjzyiZbVHbDw53i
fb+Ie6lBlOMCx/aghU5Wnu7ezXRCCSKHI/HE3zE7U0gMwge2m768qJ3jW4vLTmLXr14EC0NV7MKI
SaVhGszLt3siB5e1qBNnFZJStC0hJYuNIOAabi+e3wpA0C6OWvvIKLBQx7WApRznOUP3B2WKHlAb
MCEMlAD7CDHAS35yjxUnTBadyg1c3QHMKiqVpFMlsziXi32JBW6bSSiU8peU62Y7Fu7VK+wVF2DP
Teyw4iRuCD+cUDxIiwWQ3pFcLJJmwxexGlRGLou9oSf7QMykYMKKsQslmU8K4AhoXdcRTJvR25ub
gJ2B18xJXLyWntc134lJTU4xH+EOcDqIzy3LueJ1nvLFS8a7uc/UnTWTh9hGia8a7JIJ6Ruf+vmL
5skVDvTc86i7gYPBIJQv078TkFO7ktcnJQgQFSqRvPOuKbWOItKLoGUzjiqs1KCyhMGl3IKT7Z1/
1Im18M0bai06j+ApHf9FoOWEXbSUw/TB76Yw9/1WDkw2ChE0Wi0UP8TuXcR6VwZX7YaiALnj0GCH
RqAkeDLuJe3tyDoTW3tfYM97L+nnZJcZH2P0ZxyxbvXiDZoXdXlzXA5l64M1Qn4iWQPWGUnV9tXA
43L5gXGv2dayMZngX9nIQN2nevUNLSS9+6TGQPEsTyuEIBu8KAI03Y6RowUmowVUANO5ewAR50s5
PPK8ZNnX2PlUGmUcNo4ShCVkudWEUVpTOw1CCZRONzlxD1JtgR/s/sDzWmMZOH+3l3m/D8eWrE95
obyOEYegneSw/kbcl2IUAEQ+LjnLMmN24Z9TzlrqL+rMPtZWMd2nusj76tlbz1aO1r1FSyJs/722
9zzr9betCHxuYMalejeV2HZ8C4Ss59JDPRg7q8GX0gDOkhqR1O/tGM0usIpaFyB9Rjdnj5l9yBqp
IV1strUxf8SmYdaaVl1U0Y0QiXCkd5Hesem6Pip6q7lDHCzdSk4bfP2zc6MLldiqpm1Ge/LIFyf2
tVggbxnJx1EaAumWEufpnC9NCzN3uWyV7TBJ0tV8HOqy15Ofl2E9ETpC27VghbuQ8y4j8xbUWw/p
A9WCxd+HfFVEFFfDHeaRHvAIRPr5q2w6m562bnwTapWTPzx3iAV3AoIl7InvH3DWdnyeemr+60+B
BY4e6xD8AEhyiW6pMNh2DiUXU2E+rda8OZuoTiCllinUDk96jKZjQS50wXRpfR5f1oc1l2QySY9o
qGYKjUWuxYd0sXFyBJ66J1MQkvbkbuEtyRJ0tHLajLPf+yGqARIuf/JmKdRGHPmKacUwX+COA08B
cGI/g4GHgMhHutP2X5kfBgpMFrrtSaZC0qj3yMXhKVQSlBgOUQc4yQ7LHLVhQuWCXDOd0O1na2Yy
L6M7XTOkep6C617hulDGYZHspENYpjXuzRi4lcFadkOAYUVpXv2QIJGsHa+lIeE0kBGb3E9xisSZ
Fc9IJ1D2JujW/Lu+9G+Z82Iqxw1M/nzgj25eIU/IjIK+1g8mXN78sVacBzLvj0Gsqbd5WT9A7zG+
bjTZkiskjiV/YsyPv8WVzQdBcCNQ9AuJpAgUY+Po07NNn3caH0IuS5nFzzJ7y5FABjpG/YFhzzwS
i0N1K/oNJChoGof4lzYx1sMJHpbzOFK7ZrBvQrUc6Wtk0B6kWEgDXJSY984k6A2iFu5offU0IMvx
9J2HseMZLFfaCUknkFWFg7nsPmEP0EafLBJWEB87WeR631+5rth0Kwkt8wwNj3WRlpYslCTmuekA
AeZqbb242hwW5aphHPhwWjXDf5/dQmDOnT7vpaRiMF2lFLY//catH5hzCnHRygNzcRgsKDbjLUE6
UTuOzGFghtfSmRfBg+EWvFTaV+Xg/EgC2EEnlOEbmi64A74I915dvpxg5xqZ+VXbzVZ7thDJe0AA
Y936Lti6r+5aotLm1lLDXifvHYbXPehCyfM4aV+KnYJprvJzG2Ak+RX7X0QvKj0L/Wmq4+v8sGVl
xpf3F9KF1h0I4HIUiryLbGgXnJmJ7jF92DBilA5TLgwAWnm8V+KSkdIM4Y4TmVkwXU8Q3U+y73N2
+gW3UM2C9wG2WsGslCTcIK6etg5vxWZhEK709IeZ5KjaaxBwEmRxfivQ0AHE3kcaE/X0XaHdy8gC
Cg7QU9j3YeySoP0aM2PHG5BjbVA7BMqKZei3tmyNGZb017LyjShp27USaWjH9q9mfNPwGS5CHXdG
SN6qsuJDBynKecEnGuyAcGK0lxixUzAapdTPw+5iDd4FzlwvOcPm6GpnYZeqP73lArQFchxw+sMU
X32RCmuuusmaO9I3wV8vgQzs8Ji//aVVqMg17f18+L2MnQk2BIop+cNaJAttjExA3AbDxyhX/IkR
IqLev3tz3fF/rWN0A+8G7wqlzayIB8sNUoHS95gve7cEtp+ccsQrKrGtqsEruJecpChsySaSvnzq
jk5EY8qMUG6Cr/X+9GnfLWRTVqXsLa1FyI8QeuG1w3eac2v1DwJxxlMvI3XukiBmgJpbwBSFRZQg
wbfcvxiRRvzkRfCfbdIy/vdlOrPbxPRjNjudNCytquNOm7FUsYod8S1EmmW9gmjATWDFNRruFvdS
EANSJrA6BkwXh4RS4VamLHmKF34mKi1GKeqzJC92DF22Drl2xWI6a1xT5mzbr2tPb5lLixDZC2x9
QF2lVwPublip/n9QPnODDXrjwExX/YlQBcURg+0RpRoTVx2s3zj0Har0Zhmj+DhwszIhe1hKcp6b
R/5ZP5kt7mhqrLKSgrC9Sa3+TydFHo85dgTuvFEMB1H7MmVuUmm5p1nXkooG2qSBMkrLrLWAYrlS
R0EonkW67VPRylv5iu8UykkVR9CG/AadiU0jPgcez7n4XtxwKoHCx1JgBk2ghaBMcOEmhKhvJCBy
Bw/dpC16rEWkha3a+ulNKX4h1KaZq+zAtpml42ff/0jBwa9vxA/hbyhyaZ3Esk3I8QgKcp+mX98f
chPYw1MIedd3zszo0sc2rgbNMHyjr88EjVoABIBjUvwZWbb5p/xx+QbJwcpCtSkczt/GaHPSGivq
yaGkNnmy2sxGpUEoOMBAtcWi6TgteC2w0v9y+q/euLK9EiZ8iJIgf5UuNvwuBTCRQ2Pjc7kLltF5
IWgkjWqf4SrHnVjccwL0hd7fx6RZRhwiZAvNJMEbVTo+RqG4LAqwRrVboxbC2eLWF9nVukIH5zE2
naGG40AJB44TLeHAauY0plduHKLrA2DYQ/SXTGKHqD9xZboMnKXcvSlOkeOLOoKWXpVKp8caAPHw
LujgwqHyVuUSEccWrZLWWailvE+v9gNRwv1CPMoGqWSVhsOHrtlTkdn9UZ+3J4OT2EGcqI6+dFr0
9uxtcpH/0yz0zg7evwK+L7edeQ5Ow1f8q847rQQINwMhUhxDX8T619fehNxwNTwsbQDRKfXHzeyy
P1a1mz6xtuj7Lqr5or/7ALFELJmE5TZe3TiJe28B6oVI0z+h4H5BMd+51ieYxQEmXhO1vbzDCgt9
RP0zrX+jJGkOlUQzVolOzKCqMlpvltSo30FgxB78RxSqQmn7gZ+GGLf1TkFGhIvGx/u7vbK9gDy8
gSg4oQqDLOZeYnq7ifdqsVAFPyYMO9wraUy7KBQSs/h3nV9p7q6dUl0773DhKVPG/xVff+e/lDFG
gEpxntMA6iglAUanWgqJe6cA+JclgYramV6P+AXl2eN3oWUr6vpKVogQPFCpJbQqZHjvTkyanE7J
BoCv/yQz+9/ZWl1r5HNhFJrgE5yjM9i1erFaTo27lVYpJ2bqVgwVYq7lJnOOjvN1c2nltc0Er10i
gSAjapWnwqgr36+cdF0j5cohOfcqU6c5o8tdfA3aQkvvo/XllZZE62XTVTd8J+r6Ofc6rNKP7axQ
B8rknEuVscT0REYZhs+Mr7/o7MMWWapDEBCbeNxuSXc/sinGBmYQaQNNXtY0ix3ccHTPeDSyKbAg
+vmeMrFYgSEgF85K00+8YFPOYeCeS66qOv088xEqiuWKvST5ASmjE/r53bPKlHs0UeBt9TqwIxli
FclL8lvxoIOdmZi3xNZivw2c8Pu4c77QGAAnLwLZ2UNjZte7a9XzblIUEUkL9RFv6eNpGzqo/t39
yaNWPHnE3KOgc1klpu335rB7Yg5KJgAzTt894CGcS9imVZgcuEJws8Fa4vYNtoLNW9vHmJVkJI+W
OOxiWy6LK/mKuKOBbp1EJ+EKm7r1LpVO9UpXT4kd4SNAzJlPuqVRyiF0cB/VLw9hZbNFEGkfPOku
0O/feSmfKJz37VhGgWRQJj525JcGwuROT99vzi4kYhk7j1oXM4V4qmdGwIZnxTt8y+uXegGfiet7
oBRA1E8dW99C8wcxevwpVa5TipVs244MnUHeeADuq8PHgVAa306sxHzGC8w7QATzLCq263kfF/ww
BvuXRkWhiSqBHmMuca8m+VoU2orrsfhOMCHzriWzfxwCj8/08fbAueNbL5rJ0pdxy6J1aAKNVnSu
YTmH5BnbTUXZ1CEPE8CoIQi9dlYwqIt6CGrAbnPFgPJhkCzwovYTM20K7MiwXXxCKhDEKE65ZwGX
+OeWEpUA6ugssZyZbVuOQS0gdqXP8s5wh2/h43KrK+6r1RoSIhIwxADvZG+FtezohFMoN76UFEZ4
dHWpeoyQsQwxTnhtd/eUE4U7gBNK4djL12SSAfSKrQVIaG8OCQqtVpdV/kjNt18PDpxasSoAdYvD
cU4WLYMSEs4m8D2gwZzgz+5dFP62h5ujMOd3lVVFQkxFg+QahE1Mfg82TirrOj5chrmNA20qS015
SvI4Rzv7qCtczYCI+xfaTcBX55q8BKmOI1A1iZhQP2MauvBd9oulrPLdF2IzUHBhAb7wGzsfG84s
KcnPdt/mQ8nWOYc71/nrR8HB9gOOjvHm8wiT/Sy1Ml/GfltqNK0QNWdl0+czMJxKEtYIIrJgWATL
+/ZNKtclFIm9hFlaom83ktDL8Bdnrj3li76YSMLB/jX8LhqiR4V4rlq4IDGw4HHLTkPMQaL0z+DL
kUqu8OznxP01RaQPpv8fh5meRr/sv/dbfHPn5mTaBEoH81cuTxL8rHr3olHCAtdmAYqAsHfWmiAh
RmT0jyuWA96Di7jdzh7G4j5RFbDZrekDVZIZXUeYP7kmCzJR96b3TErdYwpOB4hdJj1VZGMEY5a8
jRXgR1Ltdn7Rdb/oWwvJUG9rPKgO72DrK25PCXRp+AOc7GKdArcm68U1bw0weD5p4WjdxkDLq5ve
3VG4sZwYUEPOn4hOHiY+BcwSLUbETvTKspwjHC49khmVGI8jBmA1A6PFI9DHghx4bgrm3CEKmO51
7qcDgQsjBQGyxf6OtVDolZfpve68h6Hne/e6yqzx+ZGPja7HPDcB6MJRVeA9uc+PsfYtkYBrSKE5
5Sqft5ggdQ7izaQoo/TzT/pBS5JmZjLvsgY0mZdzPDA0EtPTnUVR7ZSUg3bg7bYWyVev2NdHmkuo
D5c0ZkEgO4DClEl3S5f+fDpeXdr4odZCs+H7DtYXhfZiToiQGWzUE5BSo2B4u4r5JYKHTtBc7Uox
/Ea0s8jiA3T0Iu9m5eiVuZdz/AEMRRrHL6INLTNOvzkj4wTwNdIZuGgzpj5RorZZJ2JvKoxmyiqt
eOme7XkR6yzk++bvO2oQMc0tgV140NSVGOk5wvAFybgrqQXNM5nAcxb8XxiR/BxTkAFg+Bi53iZL
2XPB8IaFV/PPjtU9jC4N7siFfW1hveKKQbMxDt1WJ8Wjty6oLk4xI+qRgaGnADAkukwidRl8Nz2/
8Y3nfREq+vL69LVwrCRpFj9Gs0mB9Vtg6lqlohhVnJ17SAeZgIn5F98kbkzal4b+Xn793Da2z2ws
IGG6cYKLuXWKsQFoP/cVve95aI0WxTqomvDKxtfLR0oF1YHhP6oGCHDiM+d+cCbtaVDmajlz86Ig
oDTbaY8jRwVZwmJ76lpGfADWHbVgty3Mc3uWh1SyGzzCUzxXiqPOACez7QB9DmytOYb8xuDnmgk3
1oU9Mb3zR9KcDapZXs91ksgnaOmqljKPp+bIpYYt5vXAvhca1ggMItqBEKUghDLLIjZAafHP5rVF
X5vhcOkHu56LXmqpDktV1lZmLui9ApyqIMkApHAcBpe26JrEqJ8eC/B4umbO9refrEnHV+FJ3DTG
6I4IWPZ9NYCavTEQ7/zrGk4hQDP/VPbeXtwJqvxwevlKGWOQrdI0moXJqvCrN5w24K/p5NjQp1yY
1oypJylAobwm2pE+DW2Ng9wnb9gbf5hDpsfPNOBHt7pA+rFOPPk69y23n3PpXKZYXr8Zmh1AK9PJ
/8GK8kd87eRya1fK+/PbMhuxi6J0QvRPPJ23bq35A9sv6rFVVi5KrJ7jYXkBoI2W3AFXs/8J4Qd2
cH8nMLEtEalVr4E4VMRxGY0X6pILgZ7YaS7yHm7h/jgumCz+0+HW6cco19ONGyGIXG80D1DmJJgV
ZPO68zOIg1wWAOLGPX7zDPiy/0S459F3eSBsE5JteORfhKVx+4QdAfi44jvxmQMCa+zpZ8u2C0/H
lzirzFXgXM0qqgC25EMU2Q4l+h/0lNOZeOP7/6ajU7Q86Vo1BBySB+wPXK9QkW1VGAq+Y/9atNOc
sJspLdolf+t8jrQyAAbNOw+F1IgfHhCfE91tf6fZe02qPThkjuNvkdGzAWQbCTKG+HcXNBike3D9
OGuVqlU7cxeLdHNuDCgjKbjboh2tFKztI3mlhUTcOLo2OGFx3uX0idOg6UGc551qx3tcQ83Chfa8
yK6J7dnTFhnObxs/tz8Qw1dgsbUh2O6GgWaJFpG2IyDlIdRT2WCl+FVlYVENConC9HF7lmz2pCmZ
Ul4jl8XcPBOLkuiJJuhNnsN+WcvZJp6U8N6ayr8mmhk7KW7vVbUBSgr+nsuijdHJEMEhk0BzpMlo
1/hCa7z7O0Ule74PixpP6afVoeC7jjBEBeyi6nNsiZu4mn/rERXPERHgKo1j8vHb/cn8nKP8KJS1
d2Pl1r+igQzlyXWXnAUPcsLyfqP3HCvLc+1/LK+joElb3DlOTqgM9T7Gs1KFiOX4KMDmde/SAtr7
x5vFInuztGIf3f0Mlg5ld7LNSKacPX0rnwQjmvN0T96Xm+xnBQ1zG8HGC5pRQQMaAC7yQxYoi6Vv
dVNgGJj+qRTDC0d1dXXGq880UMdFfFr8EcNR0/9wcNKF1DnEhhNadGxERtnAAaA3ohOc7nuwktH3
PgCaIf1vJ4bF6ZlMdRSlYqSjTnBZOogceP+Hl2LTCMpDpEb08t2il37fCgbM7wIQYtWkZTThe7it
ZA8QDJkkQHIkYgohBmG56PCaBiAcqLXKYovd/ArHVv+lgGOaGRNZS+DzFDSL65cjktDoG7fRxzEl
dFUcp8BYkwG+wQ+SuaveV6x2r/Mr+C/K6cz88nCxXrGS0e9ZfqEXr6dEQ4Mz+RyjPPqMlZJMo8jp
n+ccPb4P7JsJYvCzbuTz35g6i9XzoHeDSjEtDNrt49HLPBIsHbjQZmqcjoWUYBp7k+6/JmSDvMwG
MQ8jHtUsLHfUEYbDr4b8l5+VnMSdFSt3ogREsRhy7cGgkxPToCh1U4BoWa251ULgebuYouUUd/j6
rldq1O7OHbNltvWz/2Q5xOgNo2v+POLAJ0clWiEjgimFauJ9ndL94ZEdCQs4NDxZ7SzkTmz5xk88
LKO+f4AR4adtVYh6AU1qJV2uFqnOTkgT4AWoQZBnnIrfIC3auxBJiODq2EnVmMmZX6WI+NUQIj6u
3ok0V7jU71oTHq6vA+WWrmBORT1J/DS07DaSgxtAmCFQQ5dDYsWrMy2Z2EU9T7F+V0BTpu5PbBxp
qlCP9t4WkA4GMB7bJ2WHse750oK41dduPea5uHRHFvnMrRUnXlOt52D3e3AMcnn0j5JhpTZEBPS+
Jj80MB/D4AEDnA/MarrONYKEkqxvJGDM708V/iureYJcIEHVLNCnLSNuU/or7I2y4GVbij4N23Gq
TBdLt1LUQaDMngR8WYdGkLaIvHoY0GK+cD/WnWPN1kTV3gJfxf/gXrA152jDlddHr7gcOuD0rAv5
gdRRICuW0rLVinOo8QyTcKuePVagxUKzS8KUN7MEJQS23bk9MxQfp6W9GOdPg+pm5LSlXS68oKzJ
85O5b3Wo1cO03s9IABO07JSemrH8IT8IbAWAdGeW3tqCi8vwOAKkf/fqEwZnjdK2W2q0uRtE/U7B
WsDbvUYC43DOcBIgycmhNkQo0iNaBdO+2BlnBtCT2UveCrhTVWA2VEI1/JfkBATyOf/pHpru0uQ/
uCwl90Qxl8lTcj4RarVjElHs5iEV3kUEE75vaCX5EqWgBVemMMdItq1yMzt3gl6cqkeFNrEF4XcX
rB5p/eoBg5WvJhiH3/TrnH7FIIH4YMuG9AvEBwwZoydgsDmesKgMHdoL3BGT4OyNTL4MJkPAYAlg
rjrpWDq+kFPxJu8f0ngwTUiuRr3hrCScpPDjUMmQ9+g8WoXQ3Wn1T78H3chjaN44GOa+6SYk55dg
h+hSmV5m+5ad/z/gyS1qZeCqRrewygWlv7cuWYDJ4KoChAkRZGJ+MVDh21pBmSxYdriJI//9WPmm
yMvcS6mJiNSm+S+BsPCn9SCrO1PnV02p4bWqChKk3a15nI62YuwPL41rVYuKYIaCIXP+DRODk2fA
13tL+ET/ke/MK1biW9xg8s/R/YmNPwQ86uONLI96NyKe9KihuLFPqB3F8EQNiSfdA03uXU9rDOFW
lMXFa3TR5OUKeAH3MzcNYtCdJXpqWpINwSoNxAMSAASntyYRTMD5ta+lXGjpT4rCI5HI9kmXj8HE
dbaGD91NwE0YOe3fk9o+EnZ2mKe+/pDQrZqJjyAq+Lv2pngOAKpbBqL7C5+1CX4Uxjrxs0bZx5jN
X2GWnlLGzPWKITVezovUyR8PiX6xFjO7+fXxYw7nLWAUsyZbJZC+IV+ZXhHuaswK1gALCUv44qi1
Ocn9bXdPaq7JwV/3kEk8Irw5qHlclNPIb2qnIBLTUpDylsf7Jvoyleag5mY3TVP9Se0bOICH3uUN
NCOaXzzdJlKMhrbZeWGUK9KZwFz3qnABLsxkH7EeGYiJaYk6G/QpeA4VFKB1oRnZTCdw/gSdPxho
aX+WshzAtrE4zraYca+H1VfOZAfb9r2DQbfLEr4cpd0ilqGKTxODUtxyS4Rp1+hF0r+m1C0xEDLH
H1nI2KEXb3jTIn/eflBaeRa5mIFlK9uFugaU65wDzSYVGKgSsl2THPOXw77ybQ3w9jvDvqhZjKCr
aC86ikqUNYl12XzS5dF0EfjvL2MB1RTcddsfYjwWhFJKHaU1xF0Uz2122gnk3xTBuToi5weamhWh
FIiwuhP/Wa5QUp2a2Y8YosrhvSg70YSX+xn7AYlynr/FTsMki2rpcLre/KrbPFTad/r7BzfeLosh
F5C4Zt6/NgR4+E8wazn2mf+VLfYK/888Xb+OmAXwayZney5LsZS4hsCQ2r8XTIENTuhv7iC1WM3D
CO98FXzhO3N+CT7TjXBW+myiKmGCWItvSeDm6PF8lgY4Rnbv3V7lhBNOvFnNXUSwpnFSXC1pFsdN
xl5iDy74GidHLzNBH1vMrOwEfOf6mUmUFJVGiT+HJcFIMk8cKZSErh5ZX9YXroo0FEfKPN2e7Abu
ggzLr8KqbNMZFXWsI1DGBF9A0rigdfJFZbMaXCE60+ryHtchpJxG1S63qOUe6Xgf2N7jC8XKJ9eO
jltYfyUuI6XoTlxsM8OrUkFu7u4BaYzJfO9WZB/vpq6LYuEo17UDIVc7EVtYQEGz575zRdQ6h2Fy
01S7qeE4sdYIqQOz5NNS3kOFiKwfmxjg4soHmp2gG+DWvuBRWqxAuPXeUh912h56kMOpzCSP4EgM
zNfZ6OFsD9npMbVaA/Vm5qfLKqWFcDooMwvXHhsVAYtByBVE+b2rCuDkNQg7kKykyDDe9NusolIn
Iql5/Zf38ziphZPYgkh/anrtwtBAuueMFOOI96L09dVZRmjR8fenvUHiyBOUHtqUIF0kkIbmIkKN
RqFY/yVYXTtXHBeaYbQfb/gID89yEnTmLhc2BL4pc+OpDBtRcycPUFQS2zHqconjIduvLCdnqu7T
8aD2Mbth8ON8bWyw6nxQyHHc6kwuxjChyOAhiK5l0DfT6qVFd8AMFsOnEtGBzAynxhYeGyrpZjHX
UR/bGGjE21IFJeP7wqFb96uhEGaDKjDRx4VykXFAL/jumyhsLh4e10y0ECXgtNCCpjxxjrNKoaXT
OfcHu+Oi1s4Wm7tOCtvjYFoGSvsAkG19Kk+ig68o106/v/hq1kHl7T1zNpSSYoudQOJSRmuU8Kfx
CB87Ny0FhLLsqi6axmDSlzB6DQDrOosdTuKwyyWxL5hL61OP6Yya1OCTfSVn/OHTQ2eR3PzJTlJm
EkUhFLHxRSQu/oMEQgeuqiVSYhtGnB8e/qR+kbDYCRbjQCMUZ+x0Z5P/1tsPY95XYqQZG1kmBL4c
gkp2THKV7ubKM4/Fkov+1r+l15/pQ1sm7VEy3ANHFmOwbhbCzNpkGAKFywkoIgPb7t0X89TYlQ2b
fipuzhUeDA9sYEAdhZnqnisYOz09JxFXZFRbBOC09JX7sSb5OdPiKr3XmJ6WSbm6ASFY5mwBW4dX
doCDbEsNBckHBFhjKkToVGYSNnBi2rnfhgBaiP4osPgVqbzsNbLNuM3iLuO+b6rmrB8RhPZoX+HZ
BkMWMwQln8gl5VrzccmTp5S5iWUviL7k90YNz5bweMGy6AZ+BYDfIbjIN/CbgjaVbKrkCyELXQCF
MIyX2z/V5EnfLZWamL6hBCftJdSPugSwFiNV/8KnUo1Lp2XMhkcju9jgF7wkMdnmkz05Bp/KGEwK
v19ARe+h8xNWxz05G1nRQBU+uLah2dTCjd8uqSZF8LzqqtEsDj9XVWmNHfILTKZYoN2wEeYlGYKX
xbKTgdvohq9g51uMFob+IfYAf17h0uFSK02Z7jEGro6Kg3zhyyRpycOnP3cl4PacM3Nfto7V/uZ0
gSbspbqN6r4Oj7Y2e3Z/JDFLaaBkOFOlNZxznJR++0kzXOgf+nZwiMwqOW4fd0A4rEocN7o9GTsr
H4sDCJIEjNcLoKUcfZ6CEcfZ+2W55D6KjirvxY/TjLEvvrxs6hSURK4xaQYEZVs7WahNcdiZ+GZV
DcqNcH79jnJ0i418T/Z0cIEUbOjZp0RId7HHE/3xPADkFTKfCFZXaICg9ZsqStIQ71Beg3FJIGrC
Y3fcFjE6sBP+bkW6tXi5OgkUQZbZsLYuSN6eYWz4K9gU9PVcQVvqGl72ULnjYSCKGzS1wC4nQ9MF
4GHefpLByUWVM1sKeldlkX3INDQNis7KqIwJ9Rqdm4ohPqmrRbVI8aILPco7kpRVFrldxd6+tEb+
KOIyoHm9ZHaGW1k2cMbSjMmZKb4qu7ajrhWqUK96mLy20lLwG9AXraiaZlHsGS1e58QjJ/W5zQfy
+wium/4nLrt7VN5lAlXAOzbkJev299ykFSBHAjXDNNRIBSzPtalx4H2gEbMmNgcFTuJc/uZYGNS2
WEyDAzFnjvaKqFYTdcYmxP1JJxMjMPzdTG4ECE/MT3XM3ip6c5ZeYOSh5BZUkslbcOtlTkbx1UmY
nQ1ygToIfgbely73ZmF1xAX3szvmkHi5XctlLfg+UyxLTs3S1ZZHkuAF/neGTIifVaCReNyMuNPo
13usM+GSl9CAEG/Wcgihf0NjRSeNz8ORFHqK1fko/tIzCX/BSBaqJAYUmJBiMk6c266w5RQ5mlmc
ua/rWYWDevsURsHiho6JS41L/t7xh0iJuc2JE9dx0QDp7rrH/9zTrfXvfDJrtybsdjQHfl2iRD8I
EMDBrwD4gZxtfFThLNPdZQxxmOGFP2r5M9SUe393NVQIMRgnWStRstfKnWmCptFgmAKlGgIi6s+W
/QPoOdOlUT8NW3hXU/OFxV3MoFqSXEaSDajNe8ge/Pr19Y637oiFBT4g0fd/pt0uAinsknKutN2f
YaU8wVKGFRv81uEbYPdIu+JuiBaiYHYrHpeB/t8YMeE89wDHL4C6c8aU/C0dHQpOf03CIyRhni98
1arZZPoZxvRXO4sEFFBUUqoJeb2biMAoDFLfXC7w6gdUwWq8+LTkwfuLELImxy7SJ7X4LKfeIUJF
xMyueEIkStmOTgjH6Tu9iYnjylC0oHXql3xmVcrhFuy0w414GbXmzXI49l+caC4MOQ/MT9kC5pOw
nGjkSxixADaei/tpodkhFC/kgw3D5nquakZPT9G+VY+tZqfQvFNkcfsfrSkPPSwfwhewY5HRj5eg
Zta8BtnvUUnfxWoB5YL7KjZGtasNARvZd+ivu28+LJBscW5aJf0ZvKFkr6/VxZkN2gH6RIHsA37j
CyBPyOBesWpHKnj98QYRG3Iu6IXavKW6bZJqlhbZTeYxeMPVkRPxEhWsEaZ4q9WfNJPf2SD4YxDY
LkOobfaYSVlZQpRe3Adm2+yVIDed36qWtnvx3bcCT3c4p9aZ9zbE7rDJM5MmEDzQNGIzk79f68gu
M5e55lhhkFGJjWMJL6BA/SSYR3dnJ18OAwFceHEg96kFs1FM1+onKAtvdnvL9r3PGi864ryUimRX
uWChiiFWi2dER0aS/4wbb1Rhn7Sha9tgyggQHdU+AW6oX5VTXLcAGkA0pSXncO5QxtBderSGsWJE
iC7fisWralqzEWJd2RGKH8QqcrUVu4ZSoZI1s7puLReTRkV/pEyaiCbgjbtNwxnK9xbuda1I4/Cs
SEtUJMCRC3MGoXqFa7mlxm5Fze+BsIL3+38jGsIrDkMx1dCQhqx9nzPSS30A9T0sxT6UtCmLGC8B
QxD0ow4paDPxcEpSM0hKdGOdvLeo+rjsZ+h8pwtSGuWXjhZwY9Qf+zBZkAtokk5KVl13JCm2VdpK
zHK9QsCOlsN0iBQOpozlmjbSskQR1VoWepiHrl99pPB3ZKDjDWwjyshz+1rPW5g9GI9MF4GTcOuP
sLvYLeBsMlDfuPlzjJ45mZH8mrpInSF6QmahR3lxRcHvK59R9gVR1jwaJOr3kCZX5TclLjocoomM
UBAFvHXCCedEK7mNe9cgVYottAJ4qJMmkfW1TAO6Sy8Mgs5iF2XB8q+mV+sG6cOMWaPDtw5sHth5
16NKu63FsQiM4n2L4ra28Gn4L4SQGT/e0JLWsY7aNjKRtLXVizYM6WDXF6geD6ODABOMC/xijU2f
IX9dNB9lbmFo+FUTYXHpcc7U37AcQf0PprtOYseCpaEmtNyeVTegsh97oS9fajfcMxDfsYnLi3wz
/1U5lwLtJ/JfWdB/KEVGsl7/9nhtEEwUXf7/3lt+0RzTpCrlnY5iVMRgFxZ+YxbHdMDIRai8Ivj1
XTncZ7ZNMFff4kxb6kLspdPP5OCj8GZvUBfGKFyjVYqWZ5+mo5WZPoyb3ybzhuoiqX85/SX4LZno
l/bH/y/N1vrRZY+yJnhG0vTPeN6LvE1lmTI5j7BosyWehXKhUkrachhV66qFef8ZTfqGdodEvISZ
ATta7ZkZDOaneawXN6IO9Br2ExYbqF2YRc776WtyygL4jKsK/w39ZEkHlfQ/QBHp4/bpqI2Ruyhq
voyHVc+gCkLtETxozy5MFKAPixUsKJdsA4uxoYPXGfNEC4aU22XjGDI2NJ5gpWNi9h/xi9DWiJfO
gjPAjA1MGVqwuZOKMvv3EOtUHlq/OczZXwEDq+yFi8LGST/T532TWuU9oUki9yM6fgWGwgfQtGit
CLOZ2n8McTMVWlP/3lLameJBtVTzrFJ+8Y/f9HHHZ+/Ph3ZvcWA1GGl3FItVsCaPUjJNbcWCV8Dv
Gb2K7vkhG7LnVrf2e3NnSCYE52Fo2ys9qCTkCCHrlYwUliYQruFbiDXLujWSFPBnsBgtxARAWqc6
MTFJ99aK8YWLT9nrSoV1bJrL7zg/STbpcYzRBh+RIcr8hGWPDZMlRudp9CTm4XvW2GhKav+TOrLt
iGnEQUgvqiWP4trUmAFS4kaZo3WuJxKcE2vUAOEXAjkd9iGjqlUryv4nvqhVNV+CpGVXyekgwaxe
moNON+0NjtfnFD9mNvTpAdaXW1BVyqQXOY3neOwq9TaILB0GMu9JqhVlnYbLIyaZTuU/9xVflpHM
EFK0piKkCERVOfdxlkVnrKJrT+V1IKzfg/g0boQs2sek7QiFzFoxx5Ud0ubAvQV0Fo4rgvKmerQ/
rqMEfV5nf504cGGzktG1Xmm3YwOm3Suw2MIK/JIXt+aH1WJbRZLLiqETEiH7wH3wbfsOJzP+h9gT
Yfkf+DRD6do/WTfpFp/MbQPkRh0w7Dgem9ZauPEgglBA4fPdKxK5Hn7BhiWWqNP3ao3ITYk2Y0M1
keDD6Z5qAQM5G8UeqWwMZBMah8ITrqPiTOJXscM0LQJ3MmZCTmAWMEwhRGFeq5OxmvQXI8///H3L
aovt1D7lQmAL9YrbVjX7QNB/ptm4fsL517KNKYXDgQiv43rh5iWiPOYu5PoMA8WbMiZzM43d27QN
aAZk5+8rUtrNcWnFQoQUmzrdRJ1JCBaroIyTOiwXfNQWPCbfE9y7131O6HGVPYfHc78q5Sfi6R8+
y7diXqKG3aIVqXwfKh+fp/tmtO/PY3fLpVLDgni6xKRNUjRAqh7sj5NrNVp33woAP3QDzEY1vEpB
93Vmc2qcH+GaqlQAmwU+7ESrtqiKP0dgQgQAcI7vEEC6ON6ALZHVGhJqd/3NAn9zkkKRrUOvrYEw
O+4oMy0nnbtW0i4g9FJheqymLyeIXararvwc5Anx7A1gh6cjHp/Idd5W7hUHsN/1kDgfPZeJT/Xf
XAbPyI6gcK0ZE9QXZWoTxlKxDvgqcO8/UUDS4hckfmi+PceXO11CUlU4fgKc1ly7sHkdVFkJyKMA
6yPNrYpKVptts2bBm0CpKzF/gEuKadGuRK5Vczay7OCYuaugY4UeOcp3Zx0wT4tBth7vNu8iD61n
hXpAIWq5mwGP4u8rQCDiiIMSa0oLH836SbXaIkfRc9FyStl0k/TSmIPyH/UlpfjwU0G6MCjV7wXl
TH74wUA2G/1djFltj1akc3OYrR+km5Fe1fu8T0pFW5pI+e+gOg0+blrQykij579OPx2IBbv4H2fh
BzuGf1K77KrNFFV/qoclsaAFgvpRd39zxN8OVVZB52J7oQ2n4B93PET95wWxhQBfUMKa9qob9Mz2
0Jvam2vw81PibngKqveAfewO1UAVGUWXBpFtarasKCH+sGqApimiEfUDNlRxk/UYjkhfnL3rrDcu
OKDkHHiTIZcUgopuSr6dRGYoVxX/c0mdIivDcATwQ529yPokkagEPeMPIu38GzpYLZDsNVxXAaK2
8Lc+ZWaAdMZTmvFPJAKOM5jSry0vZOCiTriyeICVjt4qXi48KxGeqn1qgnivhTZk1U4DW/HlCzax
pwodJr1+Ylxw3hZmuhpyIJuytbJ9ZvjorBoF0Zm39ZhGB1uqlzBzKerfEYQO9FqCI5BI8qZUQp9M
zdK8cZZMojEDuFxOxPjjkqRVroML8REKyfHVu94OWOcT668S1dcHQUiV2G1QtQBHxFu3yCBBHkeU
zYdH4b7EedrA0MCPDFVSgu0OMS31XpIzcJFPXFL7tUxtNQgZ7/4PoikU6DWAChJe5o7rIuimOLoQ
mRvwkSxqPMNR2fb06tYpXIjravBpSwqluy5xxM3L3rWagVrcybO7GCVYtQUJpqiS0zkKozFvkMX7
l5CzmWGNtFOqakQi2wUlRsvWd6TeebvS1cOAzwJ9NSbt1MVINqqANELkxkK9fSgQY+QCFp3XkTWz
4pinAb7yZxolMD1Xu75lNIEzqNy016+iGrW6m7hahbfqi3L8Y35Ug5zBaxZoWyKi2diB+JOoaV5+
B67EcJ/imNTXxZfpEujSz2NzUn/+Gbisrxu5sEZFrf62XTVRaMX9it4FPW8hAfGFgz/1XvvqrkkN
kJnYmHHi5r1vw9m2dPmneYF01cnsFvetEUVS7LAPn9XXYY68VxOPia7ArF2hjTeewEvNbK+gyLAx
buG7RhXc1Q1oa+vtnliqvooEgozYRSeoNs/wC+BgFrXWS4burvR23vJ5KaA134Rvgzck2gyYwHQn
vF0km1BNA9Y8mTD+e7A2SPtkbKI2Zff41jxbLHpCY/w968ps352abuL33t9qkq9Fppl/AKaymDXk
fwsH+04IDda4mw4IC8hQA5y0oInuS1PvNQNDRozNcbBMW1oKIrdMWSS2CmK2/HS9LWUca6QOQLC4
sYwdEQXYmMOOwed8j77AnzSS4gpMlmAH/Rdpbdz0GzyMFXOPdzboewjhXPa8kcxO6pznIsVeE8Q5
5DCEanEkri/a/B/G1Gw3dWrQQtCz0TLqhkVfC2B9plMpJa4/+ToPsyzeofRvSIv+SCmLHXZpj7Nn
SmLSri9w9PUE5LFjWoB2Nz8X6O32YW7htntGWXYuuuFmqEDm9tgTrIV7RmkfSmem/kbV/G8ORWCi
LGdzezPdRvEaenbKVypdpzOjORkx5tCq8ueZ1oJHjf72eZkph2pCj6dRE3+S2axfniv8xF1+rZ8f
LjLcDGyHIiIYxGSd1Agn7T/2ME5nPRxX4vQ1L6+OiKrRDpWWJYn62qoSO0NFJvXA6nlTYJqo8LWN
M7Ec+lHWEP3y0GFmfx9r20U8w/ZEqfjC6vKqPabpQJqOVFB5lU9W4U/EDRzk7xsflzHLBcuAmbMc
n3bIVN/YDHM2MA/HfSc4jtFL/NAni0WEBHjECB3ffUO/kCQXyyKWOQ1Xr1Dw9loMvesNGoXPKEu3
IcNb/k6Mu7MHplz9nzxsEK6CVz9cYzcMWh4eXPy2HUXWt4BhFofryk/YYDF+4ShiGb2KPYAxN25d
L8a5yJh5dOVR3CnPVaYAE9VT3dAa3KwBTCcPMjXX4FeaDyONyF4/xSZPWqxYXmd+UehYg7Wcbify
8aBp3uiJdwI+0072KZhsEvDSIDpMtVIw0aBmcdiIORY2HsTn3fmqLGkNgvHWIrnLo01e/3bzfasp
o8OCStguBGD1NqX2+7eSwOIfXYQCGq1tw1B4efCWZSv6GN4YFBTw3C3uen0vOOLBaAMZZIV5nX0k
7I4x5+UY6LvexOvNtt1GQLjEv8aSrnmgDL4PdvS09c4wy/29Ka7Dhcul8UrQlwOelWiV9F0m6ciY
+ZwE3arEJVwwa4U/A2ZAcec/zAHAThrZFapaXwBonRvS+5tBGoABApv/odKyH8LyAMcnS/NcPJeQ
UdGbW6xXQArG/VWzTiSLDLjcL0nYBWquMvAlaEcZUZ32/hssC9Jy5ED8xBv5Ox055Tg0CuB2k6m4
qqKrZ9vRUQEA8ta0De0sUvIySbiruW9NS1OfMwkMUN8c73OFsc0rmDgl0rO2J70lj9N3WP9KTGhe
Q+7My3YlZiIXAWIcB643/+UcG72YfBywPPnEq/Oedn9jjrQUck3URgYrYRwZvZxtW+J2exE9q1//
xY31Hb/1p5xj/rsBzDkdyjN7yd5XYiiq5Z2DQ6cjSbXfX+S8jp+KBeKu5UQEhyuo7MPVDwI5+2Kw
Ahj000EL+BKPAHo1ydOaRNKe2F2C0gmW6he1ggqpwoOuqQvJDSOwcoXjWYDeQQvlXIdlEsOeWlx5
O3vonHohC3Ct9PYtYx919YlU/LUv7hjDG5MtjN4xMlBNZ96DSTUAUQkF5MM5DuYGug3h4AzMCDI6
Rzz4e/26ANES+42Mh2lDiD2aiXiw1++7xoX4DpYOrKOcWpeMJYCuzdTFJIIX80JDqxZYImTcn5le
8ZlDsX8mtUKcA/6aHHCYF39uTMzswERp9egCNhJIHBoJFCbB8g7KrwOR9Hm7EcIs70n4YMP+G4+c
h0r66Kxn+IHkl4lWLC/TMovX8R/JRoM3JMjPLbv+ZBvggTane+Z7rTF0bqG/jh/GkHaGVcKktiBZ
0dwUkzBNUvROQ/o11uLVC/aiStzmdpPcR5vv1dfrYtmvhRxRdBkcNIRZtEKZgf8WjqWfzre/fn45
mQy7JstTVtPUWIVpXEbSXiKJo4+hrEVoO0EiB27DeUF3FzyV9Jb0O59z055PRFmS4gJ942db7UGk
RvU8RPjD2O7wnG+lIt2I4pqwOnU1G6uczMvb+WBQoyvtY8LMWNtkIfHtwOw6btPhe2AZ583WEiQK
HDWBjEqWqTDN6FaoTC+VP5XbUiPDepIWtK9Ns+LjBPvCDxSHQ+3SG8Rk5w2F4fR2wsGyTGXoPdpq
Pi6Q2TFH0eV3UWDqIln3lAZtLId6yKH3N68oLP40yHmiHx3cJq7BgiSKnQV+/2pQn2C6vXmUOcEj
dP8JfCgv4FG2L1zWWPDeVcMLrzcA5wD/qgQNWf5XrrqSud3HCNRDLfptk+rgQQQ2f56Tz48crE3J
l1fyJvDC2RCEyFF/pB293QidAbSlDJlGMGndtf+DRzw5uLh8UCNvZTjR4uz90OkTxxZvgZ38Vsdh
IhvhfHXUrzNoCdvM3wDRWJIBc+yu8Ey9BzhuQSrwod8t4BhGN4a4ceRk18LiIP2N0/eWTcvPDSGj
FJCC0h6CowDfZxULqjGjtQD0t4MDC14mFNw4d6P53+4ZBmQkauf+kIJp3j61KtFXE8YdZ73Hlj4F
e8LtWpm+XfYkrdqiaQwrXv6ecODk/xcuJfoUECHrq23JCXYopIPCIwn8Maoc6qP8oCfAdV/iL9qa
pUBGbT95zZYFaLCDUbbr+jFdp75UeKZDDjJWYSIFMtoAgGZwyF55r8e/o5qOq0+Wt+uAN8RgAgBj
MK9NvB0waLDhkJmIk1b4M1LxPRNovu87zTijbxKAlz1kz3NmnG5OKmF84MtDEg2xyDSQtwnsjeAE
nB7JabfOH942zAzstuf0y3pKLm4IFxvRpYLWaVxb1PTl0V9vITcI/JBLkvDr6hFctpAm3RzlQL/i
iHij2K+Z4bCGY4djjn6EGphzfGMWmM0Nx4kAJlD69rj67yMLyfCeR0bpPWwvotp+a0wC9xLfL1XP
v37HZNX9Lmies92MCPGlsWs9IBBzpnpvwK06pR0eNeRSvtT7fpIVqgM/BH4b0ghtjV+EgKmnb+3m
0oGyuTkPLrFmz6WyxO06xmqE/E8JShPtnvVCV6EQpe3cVwrL4hix7GVncRcLj9IocuNpqIVn1ygI
um3jpo4HIm4rSTJ/mywmsYr0t4JHqaZAxz/e1BsbFx/jcO1Pk529AsUsgml3PtA+MVTdg1WSj5HF
wmqnFemvpPB6Tv7zlhufN54/GZw9JFpAg3gmwmDIN1fC6C+/q5bRUSVJsw3dUIt2rvvlizHF3znH
PATV6KRocmG1jdFE7O+0/Pg4YphiyStMzNBkFDSeduM1s4cAurXiUePaMKc8rvVnK2414VpWI/9G
t073zfFTSEwLrxgWlokxbS/h8yjhm1z97LTRcjjRHrplK4FpD/LMuK7yuVFpaoEXawrripLZIriq
RctNi1hGhyC+m3KuLtcsh+fV7uezs5UOAfckluJoYXJeCo+CNW9i8gvn0AZj+Y3CA+hKZnZ/8Xw7
GchJhb2d3pqAGUQaPofP+VNB61aI1ml+dsCCNgKdYKYLsUOfPuEIBen58FBR2dXL07khVv5Sixbf
6vZd7bV5Dp+w6a69ZBe4jCJeO8R4Xe5mHPpoFXJCQpYYP30lleH9ryWJf8D6xYmsSQs6pW/o7SjN
9Ge+CzmksG6q8jw6MwtBekzeMkFtuaObPbnUCQoCv+ghbRLg+fiIG0NSZSDmQ7CEp9gXkgaoaOwC
tHgYalOmGEBghUMqL8qFNvzH3S6Wrwh4huCFGJStqHZpsl3bhx2YVJDZKOmLrxjcopWj5feiiVPM
Bq3JthXm9c5JaOZFmI9phfD3lZvN2Go7/iQXIiypGs+m0K+j64fRmlHfF3PX59LDmtlDTkFgSjs4
Mn8n/iiOQ0t14vcws6i1NLkt8a88GDNevgwqGtjtRDJlfLD1Fi7+ynOpFNdKdu4BXe9T7uynmAJo
yWmtj+ygZM7ksBjXdyzu8ZrInw+JJDQxM0RgNBtUH3RnkPTBzjidhJF2UP7+T4TWWN9P5FDdFY+K
QWUsCM8CBORiB9fCTOKfsKAuQl9QL5v892tvBl9p9tclfFNPdkvMgRiL6DvItuKn04KK40aoF+Ie
AmjH9yXLDcuh6e7IgyfhtmXb7i70D5AHlrSrOQmpKlfRbmi/bXJjgaqc2g+ja/z7s2hfr3pdFxDk
I6A17Pj6y4aHn6DqlhOk7JaEfFyUCdEogeEcEpevb0HpkZk5Xo2Jy/H1lKSEpFrxB5FfAi7ZuHVL
/beDUzoEQyzWDKmcn7T6efHnITzbb5F+eFr3ZqdM2L0C5JtHKUuW0gq0mgLarUcMLQi8FIAWSILF
uo96x/xV5AvUSOYIhTFkS+3i0qoVeJFjX98WfG7tNHmluvj+R5S0wSoMtzPb52hJJGVsNxtVM1Kp
iXUdvL2Rht/ZadBywquNLcjftrIQOWFXnjbn6uc4XURWrxY20e8pusW6Cesmx+8fxszp+KU5RGVW
QAhjCZL00xxULJhqpjQvqyxFRcSUb+/xbxPaMW5PfCdZbuAlhjto1N5AdQgsVvHGKwZ4A1it35VT
CGDtk32l6PJrWLOEYgf3mwJoxdMn85XC2QcoI95cc0JVndFhkC3ykLnUOzpLESo6gK50C7PO2e0B
002ovXphANIbN3CehFeTIMGzgxKeotbsLE0j/s+u6XW4/CBCCByHQj0NGYw9eD+bZTpugA0b6JXS
jzugeFZ9X4IQZDPr+SlRvsWPoP5pfEkeiUd7ml/rQ3u3HMYptj51h9ZbwNCixsE1q0raBujd5gUk
Zc4LeHtN5Tgqi1rcJ0DaLPoJ+29hhNRq/d8vaSFLy9Y9X9RdMzNAVRLBAq1st+k5Uzf5k1QUMKOO
RsjDBOG6FJXCg9akXcrXuDBuNqEUYBAEpv/vNu5T3wOXmGGT8Da68R97Ys2NIG9SMOHxBxUG0nHq
JxqLRQ5SO8lkT7igtP+wDJDTJ9vFrP0XDjGF44ILtXP1wvdmS6foQdAg+qZj6g937nWD+6GV25gF
M3nDOyopVCUhZgHDk5Q/TRwhQtA3AUBtH6GiWAgWJTFiQpog2vVKgsPH8G/2qan8niuqlWzK7H82
OSx/t9UafCVX/xChfiXXcsGeBC60vyMIY2WISDu7mf9K5yzqxC2f2To0K4CzE0xz4OZmaCX9vZ1n
yyd1PgGlJWZSQmY98aVmURFvSKZLOUXDlEcBp/QpVN6q/TZly+FFPUlDkbqQghpLJ94CF7iAtUFh
CnyRgjxW3K5hLUj2AiQUBtrZup63A1G7OU0Emiz+sDqD8qkGedVudhOwKx4/eUhTCD3OviT34o2K
cV3YCZrzjvPRre1YFS3ak9T20eomhdVtYPt8VPs3Hmz4roVPBW3j14ppaSQSrjwZ1wCUQJsXc+v3
vpL4ndNdWQiJkWGLyPLAFRjOYUKYTDSTduOqsDzRkSzIVD1jIXqFj6b7S/4Y0+VAl6MLUOst1x3e
lxWzFUXekqoXL+ApA22J/MnIhkfo1rkKvtLsX5noxBra8hihczNKAUKvAqUhtkUCkyWt7KtSPKU0
53cPNc+RCOsqsR/TUSVHuD72wUPn4+l3Bxmh1KBt9aSJ90GVD5AWG2KzhHcT/dsAK/L5lul1qDoW
fymmDKwK9Nsp2IqVLd55rHeRiyiIyA5Fx4y+f1HxfnIgbRanUsH9OdV6KMRklF9Yxv2pHrtsYRcW
4iGPps4E5hRxWDCV641gWN4VVDSnH9BEW7ud4AvmPgm5stFAPZVQHvrvovKRJfwFyFDXutD1+Cs/
Az0kBqzwLphXFR4zEcfpXDGhYfyDXjcbsQGud2jhlhFe6Qq5QN+fwYh305ki+c0mfFd0idjxfdYE
+3wKzQ9XJgqprLoYGUlk/sARiAd5qUJtjQENnl7vqLJfTjYy0w0w3BL9Ox343pQOOAOmhtrdYJ1h
hr8t8zre1wKubJJetn7A/4fP5afrv4oVW6H2wiznEl9lUWfkV1NAneg8ZZZkDLkxhExhVE3htK5B
o2IRaniCBx+M1w4qolfncWlH/dwBVDLVjAgYu6zvTvbKMsoITT1yx/jXGXtQxFAHZAKfOgjOeJSA
x5eEp9qLAGtlsf3Wx97cxGP2ORt6v16Uyp5CjwU8G44t3kKr6XWKmpY8gfKyRmzSb3b9f/dYP59Z
MwVvSeYkB1l5YWTO0NyjDVtqveRIdPYAX71WE7NvITxkxsCN3SwimLQQZYUDeIue6Z1nIZ0InXrz
GAn3xp+QfHBMl2yQlUa4gmWqvzpEI6cpzfpWpmx6sCZX8KL87A3q5SBF2jjDqTGIgXfY7H7wlLIJ
RpYGJGY5FanEyyOFDfkm73QvrZaFm+Xgo3U3RSM+kUkI9h5881urI4Yw+8EwxihSvxP3SYEvgPEe
pGotBdlS+83sOoCGNzhsB/UYU0C9iRQ53AQtcmSQyWJ+eHpm8MHcjkT0K1j5jGAaUtXo8R7Lg5p/
O8yglSippSt3qRAwoIxUQLHXy3tkyag2AeyLzeNsAB3J6MeqGqlRtlsShYwH8xotl1b3HC5fQUmR
8rx/Yb3Cz9JMXWxr5Jm3qIxvgstmdApdag9I92kAMPKQu7D3OeMJ6tF2F5dtPKFONelOgn/rwdRK
fgHqORPLgg+o7ekw2KbRi19DISG4DkrsXAqyl5cx75uYzf7KzjEFF7DHlVvbjOTcSAyieiY0TrU8
3zdWqXnaKN6jacsngpI4590W608VwvLeB5XMS51KfBb2dv4Yc1iSrGj/KULe7LOTE4+Zf/+pYn28
A5I95VfozJtH4+gcQu8EXvVhwvuf88lX1P4yGeZdsvLFF1GOsGiYxHiBCGpuBinsL5lfp033M2ER
27oPxdvYUb9wMKwaSmA1mlLxj4vOhdzRQCFNq99ncNwT8oS+/ZNRfSzYiim5HhiFKO8KJeFEcF2o
uwM1TpP8x5SLwC0ryF5RUJPglHmIk3J8OGChM3zpfI6OZI63/ep1TgrYU8W9suzSv6XPkWF9VRZK
zHDi6ooablHPemsPCbWSxv+Lui699gbA9u20FqOw0LKDzBSB6LMf7x/IklwPjcbCV/cpoiO6v1ab
wnKVf/cKxNYPqnmfIiNvIZTVYbREL4hNHaAy2mJvR6bPDyY5hIij7KT/Rp/telV88+2xPdWcXg9u
rQl0Rb6o2WXOwG5Ega9P/r37elNxCNXlVsYkIqqdl4bMKpbTkreGJ6fYlZk87lzhzbnEt9laZOej
T+Iv3plV1OEO7mmIJI5T2D4+9IqKeWn2N1ZSUmBsllLcon2V7Xu5GSmFEYe/V5WVM+60kQGmFePm
zzRRYbVwnHZwTco5Aht3C8UFb6jFTaF5oMDoTpePOsCQlrYZ1yByNld0qptE75kjtZZLw76rey9X
wt1JXR9YevieBQoYigVC4Sf7C/A7+yMXGdBE7OWqyIMQX3sXUmYVOJFGzehqgNx0IJkhbPNVr5q3
7/RdJyJ1krz3hIsTm2CE1VhCcJXpNDMMgH1vw5R6BiL/9x2Wg9jE4WmILKzWiVW/eMJ1O2vIGTm7
9IxOX/GjrWA9O+I4QBOgldpgXR6mxAFse8vEip4WMntRy7czUGmvd/rvv89ZfocpEgAaA/PR9n+p
k1bBQonegqxOpgZFexx1O5k41cmtVAES4ednvStgxCOh+CVWaCe+cpXFnmlg9rj3pVRl8jQrHYMt
xA1g4EmhDaWZNphFNjFHGFfPZEs9FxuSEaJuhdRT8pObrPXYVBHb32BmqLnZP10RuS0YeS3lX33+
o6/dQC5vYnfVkW49g1qAgc2GHU1rtWrs4+XgvfUdbfsZHSON4+9mtokx5HfrU2QxL0HwmvJSrVUj
G3gIyobdj63+eRnY3V9ZDyrkiKgVrQgDbGlJix4wpBaWhr+eCSDT/K+Hye03casbOLI3fkvGoq0o
qj66kipac/6HkqH5f7G4OML3uM81TB0zsy47tCrHJBoGHQhped+JAG3D0FAIVRhwK+SUtBlMoLmV
UDC/6Gfy9z9IpUfqSNTPftvHMQpDrPK37RWI1G0YouxHulSjwh8IhDA1B0AJ+kly2qz9DFRppHUH
EsxxoRfmTxGkwumRMrCtOjzcTIlI5Omo6sdb8wTP5wZULhUkVGuNHHFORM6g2+fOCFgCZm7R4pVN
sxC6YGIR0kn6kWRaRegli6Qy+6L78w3t/GE7ZsJrrQjNgITCXXwyXCio9/SXsfmegmvFarCX3ay9
9/p1AYzEQLgjEjeS4Yfx9TgEBEWqmHHoWb5NsSjVLhrgVx4RpvEIBe7OScTZtOU2V4CseCsD/1PJ
d+wIVTt2GqkHxCLc6IW2Bhe4FNHygUdv+wSt+UTlE3xv0XdA62xwHlm2WG7hoRdMdJmszm6PVn5y
VlIj9N0NDWwqmdh2Zf4kTd/BgYR5x2PpySZBuoHaW9/qsp5YCX+tHyrZfeqJucIJ5QZ02dKizjm2
Xf8eSbNGRGrMHYRVWS8hn80DbD3M4MJ25Xa7uDH3tYHprAQgrzPjqwphYmwGa7hcED3EE54zfDez
l/dgcCPixtA8ZauhPsLwkjPFlmo4G8SvEUockMnyhctSWY6wMlUOmlOtRUFOBqoBWXjViccPE0D/
90B+1VtpEwPeSW0FaIOAUXQJiAu75EYzH1oa6Q+1oy2H3ehGq0h7gylI9xLbw8DA82X89Tu9/oj+
QGqOI3gS29g8/gBCrm2yZai5HfRmTcQGRSI0HUuhSfa3ytn+F/iRevLbMzI9qKRntzw0lb0LnTUn
4dkKAHtnnIqnWGE00iv89UzNcNawneNzp/fKPv3xd6spDXQaHSETRZ2YYElVv6abtFmyxfBJFIG5
p/RiGVRau+2D88jB75os4YDxR7GNsWXMJp9zdFoJLkmV5RpGWKH9UncnCDMYVFScdu5WezNaVMaq
Ve0IEEjq2Zpt8SXFW2TGptW29lLgrUTm5DXtaAH2jXJ8q7hVC1Q2nbgJ4G1siAK0vgFaJMGSMSSn
xJOU9l5IHLWbUtTxMZC3GF9kOyfqGRlXEMFhEMfRgXhPTaK8dgyyEBskIwxPV3a/Xcof6Xpo6j8Y
3cEU7gpFqsmghkZmZNULwnX7b/HPIOXXF2YIQtcDyv/KuMKySTeyPmGa7PC9Wu3BGlGJ0hPJoLoJ
7anvIYQyPmyV1hngVAw/gBjLxksdI71gaysAqURYaYg0zxrjaYQmmQl1L3Izzzk3+2e/PrMvYP+M
lhB7N56P0SLot/lY+WLv3WybLX5JEl+8EuirWznx69dffkDCTX68mOdp6JWeJR1skAPGA0PqDQQR
PFtl/WuzCnP3PXNX9bJhJlF91qNcSyK8+M27ab1/gfBwrLwKMyZgAOgq2fysBPQIfc5L9/El8aAt
gGlwbzP0x18cYr5f7336MY+S7mnv4KpJSzYB9wJkrQf9+6NJzcH8hQF28/jWIPosVdwagqyrk6uy
FVwmGhY5E0XR1q3LJDOZtkp54ULX7yJD0v2rvAOg1yEuLzxt4b2PwHkLJj5+sh/5jK+kkr9WhkkV
lvnwwqngsSCDHZi4UxkTDxWOxdjLUAIzzDNOEiXZG0gLqah7LY9f1eHGlaaAbT1zW3kVMPbyuZAB
eJE0MhzbYWLtKMYPM44mt3VpZSnum+W/zdeh2vf/8aSaj1GFYSskKYsNbvicZhP0apLOtysJnR6W
ptgWthIWld0Jy8E35GKdwATHAXzw3IhtLso/U7/Nnxj0o1IMvI8hTA4jGePU5Itlgh+0+vcVAgTS
M6QlGb2YaeC7IwIBAh2A5W6nQgmGc2JI0qdbRsaTVzOL9thbmxltP7zsa2Gku8bSIgcdoUDSV01O
0liwkbhKoq+zZi9A372B2rnDR8WLHK/2P3HDpY9MxeVq7eOxPGQGjXoGy8IDe9HEVunf7bii2uUn
CR28jS1paY9TbMVkV3g/rVB5K9Xe4UYWUfeUEb50Ijf/1V9UPmeqYFeoA8azmFOJ6LCUSUbczPBe
8oegcTgrt6tOpifl+YRY6a0EB+U5fdkNxK56CUVvjks1I+k1KA0/XC1MWDgzEG6IsuJsTsU27tVp
bjhDvLy/Qh+ckQ/J6uZ6rsV5bo3P3j3OBINRWXS6pozY6d62fjHol9SBjOhtaFNQBuZ0Sb7ZhATA
HX7RvvnD0wlIYr0V09qlYiqGG3uPTZmbqJYBt+52RVVwIYZQXc9O1EoiXBcaiOljbiHc4alnMdNm
LTgE0R3YhqAQoh/gT0RRMJUWhm2vyPc2FhwVbXLoA2wpMmUARk99yNoZNt4+5bI4jJAazdcoY14O
0aTQ4w6u2j2pXG0FwhveXP7MeaMxRU8FhaK9UG0g7zQ6kZntQ5WeHgS76+/tqocxKOqA+CyakY5Z
8zP9TTenbbbIYrIQXueIazx7u2vYUYTvGJ2COjxcfWm5FpjgHRcPBJSb4yOnHZgtWyPv2y5n5e3L
nBK+FGTtEEpW+MeZTjeSVS8uIwGbufCcapox4MtMaF6g3T17TgVcP5VDKBO7Sl2UEKakoHG9IsaB
k8p3k2/GufA7BuOtkhIEIUlWJGakWI3ej2kSkxZQ8wyk5fTVImzydjVbCQyNIyth3mXvoXanoTO8
jzIArQSy8meQ00aA1qqvckJj8l2oFl2vqYHeWgXgmob+Xe/CHe3ruzh5T1qWOICM4ExShtvzulph
6/cbTTz8deTK7jApY3nrMmMLrParcBYqqh2smFKlbU7SDU3NoSmOiTQmWCI+FsZzI+b8oGK16Nub
3AeugU7mphbV9AxreGbziT+fAmnkn2b2Q6+mXrJxSP1RJ6gJMa5XoKL20P+2cOXA3+T+KD8/mYyE
UW39/55SIH6VyYQFr5ptqBLXGzI26PCPoxdhb2AMosWx9QOVaifIoDH9QS5Y2zHzkxKQgR3Bp36+
p5uEDbFDX6oiQr/OK1u2sPdlXMduO+nFLgEKaAf0HgWpmpUoClZ1l1VTBsCV3CHmaL9hy2RCdYIN
G3Tul64Ts1d7saxKH/XVauc8bN+m8JLEcguozbSiNHFoQwGmgaER+n+M0vnBNVxB2m6x5USvPbnc
4hwVTvxzRlQWBUt1E4irtVR5rAYh7Pn5MEFX5unRXkCJOjFe6sO3A19ycSGIbDonAGzIGtEpwhyW
UxlIo76qXF9zy6apiQtjZXICGfTjfauSLTULlWXuannDjjbTsB4asZfK1uzHoo+Q0h3KlgArG6Pv
X+oqNvfAVzcwzXkyOEsWY6O9JfssS5EagXAZamHTWZf1X/7fapYkL7rNqGrw/xEFb9jgVebNvFkm
dLjfWntDKzbQ2n/p3YJ3on+6EMRI+S5yT9ObDenhxNIoDw3oKL43dp45B0sERa6LX6KdGTCo66Sj
DmXzRf2+uRkhKvLjDm7uBcldQg1MmVoImB/OMWdZFJhCPuPhVYWvetppjI6xWO1guLcwS9MBIHLv
mYQywdI9apYv7E91JC2Cs+WoH6+yWRU0VFXq6+7OoivA83w6fYZeq7hIm+LIkYv9rG6v7eDRl42N
jx8xpVNebpG9Tp8zQC9flPGNQSUZqLXgNPKzQSSPmo8yhWHZ2vbrJ9IJwqEkgyAbImqM0Ap2tn8I
QttoDX1nZ/C++iUzY4zDsglq4kBvvCeImaHND0fVwmOAwWExewyOX4t2VwhcsyoL/H4zja9Sdhme
zn3L+l+5lhMh1saagd2YvpwKN5ODw87jTnGe3TcPdl3XBmg+BJK34SVDzN5A6nC/54q3Nplbo118
MA3Xn2X5+itjTbhtotQa/TfDES8dGpNGnFwMsWXZAR5/8DrJmib6g6/wms/c+VhEPHI7rBN+g/yH
zqB2c3E13QfCoQ32lmW7XBweVjjAi6ckHN0f6KKAtWNATwHYt7zr+F0VNCvB+Tw3Op+aCUYOeusV
u4W/xanqDB5Qztg8e1LLVQRH26RLaHSfg/p+99RbJAyUz7tJJfAC+J/xlj7eMFM/QqYiTWsDGUJn
reDT0CDJd72veBaKii25hrKgQhhmkkVV1wwaGj7tNYBrN7rSW0cUEmrkoDZxQuWnzum2PdwJ9aR7
eFhEKy4U0YvJJkH+HX3PXus3m7Ibf5NmtT8CUKMziXCoC8lfyDAPxvHcwRgG/ASlm3ufazC6H6nl
XipvTNI+fn7SwL5yCvbUq42WGEgzLn+u3MSw9Xu78LsX5eMNyCKnWBJJ4rgIvskWnQHwzuJrauhj
KxNDFzGTNDvBhqUXzVJ7T8jUleXRCgQFjA6vA/ZAO7oTb0AmQzKs2ZeElbbIis+0QNLEZPDUf0bz
UPsQ7nbDo9Cn0A8FBHzpcbCP0OvHZFsyQlRt+VJ+N1qMcVPobYIvF9MNfW2UY8Y/BheFJg42Rsjx
UNAL1+DzlJnC0VAFJUuZYJwdu3HCXndL5so772Nmvda+8CauBdPRDV3Ffchryn7obJ/tvGBYSPCv
tbjnBIsubr0k9p1hu+43aI9KKSemQVnJElIafyD9WdqPLy3qed0QNJm20U9h7XrMq0Ysr4k4cIsw
iyOXI62lMer9obCeStPrYD8umevPdFpMgq7x4PGH5LdGtUbac8BRzU7vXv5vnPw9HCF1ZwdkXHhw
aUo5wTso875atEMdSVvtMk5cQVXJcvr22NbfqII+SNxmTgMXjqcXgqysmBlB5toSx/5ZshmrvHlF
qDCPHLTJ4QQOHqoGlcx1O1x9evgHW3YriSFRYYYP0UPYpJqK6K9fznPL7ADQF8nZ9azAOQegdhAJ
33T0WalPuZSitIsj5tkGZkeTC1/vU2jGNSEOilvJaPgUJEampPxTOqaVMNXcsNIFdNNKUyrMYG6d
LJIzxWSZuWLAsVm1n8uTwM2Wifp6GNGbwJ31yDepp6u6q9d98h49NfLvh0OyDPmvdQsi7/+ZxJTK
qCfTd5U/gC/ug09p5DDvrnezx4YPTvTPsY+KpVZNSu4FV2zIIIGij5PnSOfrDQbxqPMrnOBXvo3C
abxEdYjLmek8u5axk6b2+Ch1LWIL3odu78GO9oF09G2ZmEBDX+G5hCf8EEjn/EmUVWDG8LOulKfj
wjaFr/RtjFedcpXEfVrAOHUXD6xFUtwqtwiEa0wJxdZRatg0i5TqAXRTjrOtGigqAHkJ8CzfrK4e
czymrK28IJaY/Ve70XVZg9CHsw+LvZaAF/nUo6GZf/LeAQt9uRPItzrJHB6ubSySfQzxmVBoJgiZ
RazSUoQDf6x0GziRxDi+HjGWU76atyWD0xJ9txLil/2JpGmo2pxBM6xJYeSQuog425QmyKFt32y7
9xlMPb+fEs/pze66UMIjLbgpIvb3K8go35nVQHEkml2Zxa4on0j+WMaIGE+joWj7k1AmSpihfm9u
48IrtSxkb+G/lOb8Dxh725wGjYzZ3vwZbgGtn10lZVwYisIimiZMQhZeCKOWNgh2ZnKHjNgZwo58
XEumW18vbVwkKuhh2xR7ltQVkksbESmH1ot1IkwqDkiThonGbxhqpSlbgyi1zTCI1nD+zUkVHZob
b2BH+XtHHQbIB8q/g+b3s+S4SqBpkbFy3588EOVCyDuDN6sqPx37YVmhiw8qoimN7toGdTgbXrWJ
O/3wJ59C7uig2fWIBA46Em0dSQU5XPxRPFn0F3/eneTLPOP2MnthGw4MxwsBg3FL3WqtPkYXzPhD
zs3f+r2LlUeG9qZO5PvnfSKipAWHUe0PgfkwJCLpNipPZHL1rVymrVGm59vjKhz9nzzHYIzEsE64
kI+UUX8AkOoH1VjxsTYUXvMsDeq2wLGMgw9yl/867R+7O/yis/APaPhQF6YLTge8AwT8jDLILGqD
OWVlrczAyLPjbM2YaNmuJKJHxfr+UY+WnjRAiCVvIoZkWwQj1rW1E8/PIiM3EXMnNiPx0KW4jsxu
Q+rp8J3Mumr2AgFCSEovBtcnRBzF9R3O/mp9PKCZvnHLv/iSRWdz+sgSV1FW0jRSXrVjFYvsNLPx
eBmoosTp87eHGs7QXOtbNh2Gr8Hef8hSQpzs1EDAHNg+SIcrRcwDnfrlT6WB4v6N6SgE2ldC1++2
hlctoTzdq20Q88Kg48XyHQ27x5i1cp+LauD48dAQwuhA2pUo3KQV1+qK95Ch0NdiH6TJr1k/iueE
wddA8OrASU2mnJQtHkUWIXed7jq+cnndQ9JpeeEWmoOlsb+9tB4GIikL0DfBPwKtFw0Ud/MthNfC
y5ccXObPAScu3kKyNKeYS+9m8E8kiWDICF0lKNbUevNLFQuf2zj0RCsKw35gFIFgr3y7fuoEPi7+
4J90bUMrJtuf5b9fEXF8Lp9YDejmoY+F64RkJeef0MF7kBop8R72lV7W0KFQX20wyVJOuNBgpP1d
iOnb8LCudSLY6lWBcXS2qoJssalcSVKpSSNcKfRqF1yS5actw5xxMrqXKW3ROTer67GDnyxi/Q4J
KjpRUyexgs8g3H+gsWoXb1aHxydvMfbgSWEXGigZVKjtT4b9FCwyLieRjD/xkyEMIyMJrRtQ7XmE
eO+CqHilL6eaNN8VsfJY7n0wjGvE2zodyE9hd3ZJDqx4zTqaH7hZGqilmGSUKz+icLMuHKnSavx/
Y3oDBuFkfPQ+eEfex1hfk0hn+C1QRpSAB2EppgB5IsRTz+9V1RXbsum8UPAexnlFXpTegvudKIo2
lYA0W8JwEfic4Pw2kAAJTMQI4DFhVZTZtPBAod1Edj//quSRxZD/VpiypQURI8+op273pmVPSdHJ
a5fZqPVWT/UEjWYZPXQbDdMwjLHWsTftp5pilMf6RDh1vPrcdFukoh6wP7T9ncU/nZfuxkGq1a0m
pPog2dE+eI/jAgfY0c3/ZheNqgObClsI+l8UWyYMxlRk9ewitikM/5zfky/VlO6kpnXd8tvptcZP
5BQyuAd3cNEwPR3SJdtfvPQqcCAIFqLR6eu7B/5khaehkhMtPRdlaeUBZZveD1+T+eD5bef7gXyI
C4okQgIZmrlRclxkadgfiAnSVbJ9J0cTDym0DmeouRmsBWavI6kb6qknlxZdr1lWJclN9jJNx/ax
cPCnVgDZi4EzjZY5cCecTM9lVLpGTH68xyxU+ghexNcX6n4fwp5BrciD6s4dLcyeWdtozYVmoVpG
tBme999a/V4+Uk3FWrTg6/2BpUa+NQ7JWp1q7QVjUMEcu6/W/iIoPLj2Fn7ryEFbdd42wG0xE11P
W1QHsj++O5ltHQO3iRZiv3eUCj06HC0b3Mma2b3PoRBzFmyqvDqjtlziFC9T+KyiMxdOltlAOjrj
Hv3X77XXZkRdMJDXHCtHLxMMImu1Ip/th+wXMJKoKHFpDMJU5o9TclRnQdP18kiUBdktwpUDIeK+
0lNJ8s1Koscsh0FDJKfAAvhaJHWWY/9Y0jhJYPGW+vmc/BOIhofiEBPr//8667M8OGPB2gc+ExxL
c0zAeADA4AqnqZn3nTzgSGAzgwsK015ezfnn+t9Wmvcf1Z+5pbSwmdh93kJI/VrT0aMtof6VqSrR
HG28qmejEC895vKku4duBnCmVWEq+Me1aIuZGrMOPXVV5Vmt/TtQATOB9wvgyOnNiSufFRrbZzjx
9GkEUTdpi8M/PuE/O0XAkhVjCas26hAy+6vxBbeh+ZSUKvMaqi8VP6a9u0YdsX6txH/mr19YY9tg
5V5rQB261HhJYd3OPQSlD1Y+9tDYWWa7A4eR1xn72kpeL/fcH8LXIiuNJQkumz1gBWHAFBQQNHBk
B6VOnYnxSsVLLH8MR2gE+CFdwS1UDJIFz7laJFSjwWydRrHai7/FHpHIOz+JYnEameGXPgYnNERW
zRdxGGfhn6SsrOd7AKbrVwX69Vftiq0g5mAUdg63DJ6yRkwKz38pI4Dqo9iyI6cN0pS4h+yK5I+z
k3Ew+viybmzRFwQ7ZDufbiCjq7nwEIEJ63yAe5Io95WmHGM9yVvwIJ9SaNCMsQTxnc/BcGjOtvOZ
g1JyKyzP29RywPhHroByGGEQg8uu6w1df3h6uH+vmXN8hKAuxLVnR8kGhwJdGal1BoMBAbfMRphJ
kMub+aw9iH8LrZvBRemYqf7ZyCJ3G+5SMDoME1h6O471h/sDEZtB97DEYoruDeR3/NlLuBCESfjS
svM7HFO8aMFJMyXpwBKSAINGqF58j55bI/oJqqRtaSt0Ercbbfo7sBPumeruV0Q27Rox4LMnyCup
4CO2bTI5vS2lOPJkBGqz6+I5YmkelFqZo9fVNcPs9p/5Rin37EJS1pX5knQlBrKV7ND7tCCq8d/k
BLW5Jys2eV1uwuktjqFX3zd46VFyXLWN3lW8v8SZc1/C4kvbO4daPQOOj7tC4qx9kjkbsFM7lJJP
vad0GeJq/oKpcUS4XqKbWmgBJocj211PM1CqQI+9zaEeKZksYGooTTifWuTPKO2EnaMsShPYA/os
h0JfaYQ2EyqQN2UGVpQOfx9Wd3DiwtADd4V+wCO90E1CDNCRk4J3V6yZ6omzkl42NuS//K/BHZAN
0/f12ZbBk7kztJCn9Arsj532Y9L+BSVVMFAi2pgC2WEP9NHi5XfaKX4Tk3BX80WNctgsjDI65hE/
ymcpV1XwtvGjjeSFJfVJUOdhd0qvZJFoiv7M/JQG7HLT2tCbQbavSFkLD+p8VLFNlAh0TM/HZWY8
JjUcqBdmQL7GCfjojstpDjCNaGLtu0AiqynaAX8jOuA6FdRf781EsAIgzRvbJfHvrqugDdZr1XDk
uAC8tXy98gCUL9xP0Izq8FUJ20tLLIRrHM1R6aMS82+xcNyivDFVjAlMEL7QyxpVRjoZK+buiaVx
pTiwLIoq0iLqJAwocSZ6jyFCYLJgEX0Dv8HDcn62rMjzvl1ZvUjSk75v/WiF+FP69WvYeOLyjpaO
cNhyPgTXnE7o3BkCsjWKR5CEtSw5kFGWO27EW3QWD915TQhxRbHrT+s8O0L4YEwycv/Zx2gI0ASX
rF5ddRP9QKEs6pakWMOvmeqM0H7AqwHymHvdo2Tpa7CFMUrRyVDkQsuPm3fUk2JPgliMIcXUR0ba
1xFgwhrzADMff3j4EYFgZILJlFmXh7wJudtlGmTm4ZMDxWE2GSLRCnWegovcTLFFOu/+xEyuyTLX
uQyBuDP4eLkVSGQ93p5jxPB+OXgi+MGkUnWP7pHtImK4Ir9cTNZAU6bPFen8iwaOseDy9KFs/0gL
QSfB+Xia06JicJl5DqDNIkCY94LOt6pZGjDfJ6lcQpt9gvmxr2Z7v5yngnyFlG1r3JuFyo3+n5Ac
R3b+Y0zdQmtGg6wxTNVfO5mLUWVPphCtIhiESc+6p1YdHjh8uBMAhn6u9KvIXXcgPtQWbhzet4Gv
D5b+av5ZfvwxEL8pLXzLz4URWr6xEWJsJfwMGL2j+vlCQRAMq6Y6mMJgbLwpVXT/RFx1AYLNPxPo
RxwAKE5E2qv7M2qjmbbshlQb1KCG5TTHsyoJn99Z4xJtPSgfPq/h6877V5t2drCeHrD4PCuSxkDz
qLoN0Mwb4ELYX+ahdbaJjGTSXKC/narqeG2H4wUDdRHwLKM2Xmyu2fjY2md0YYxF4Aal1tDzDKc3
R8xBRnD+P8z9YNJTbvlYINajWLG+5qdzRQGX1EW5nGbgc/uMvEDt/n1LZcJOaoGdC+bznKi+wVOL
Kr6LcvE+YUHNjsnsy+Xr0HrYpzxKtSx9tWFdAUTFSIH/C5E+uefqbY7vTLG3yCIN5sfwbReKKA4f
36UX+DNVNFIcrTjCRWCIoyjzYakl/Ynb6CWKsEckMrA3Ui5RdSrpOctNrGXf7xjDMFN6SfSbd4Mq
5Vz+rsU1hnTBGvn1DHAv9iXfd763OIQjF5dX4AfRXxgH/IQnb0YaFnUXaEQjSdCAbVeSUkxJm33T
t2KP/cMtO5CQRz96Q8/kUFaA0UoDNa+8S14kK6GEs5y/8Zol4bKwCfn//ahZxglOEA/piumNUijM
P4UYg6peOVGZcOH+6waJjtwUCmbHSaKnPxFR/04LIhzN06ZP++VTuaIvLT8p2hIvR6tTy3fCccBY
7Ou/oCYBbcvmQY8NzRXvIfvroT70GSauEg0cOBeEkO8k5UdXRmAMrOuOVpILPEYp3hYrFu4DLgtm
zBCgolYZ9ESajZ0WJrpns5G0f7LXx1mQ8VnXPrGL01FIfISpPEsKszylAgX3q3o9mNfhJ88cnPrC
6+6AESCrYvrEBiBys17n0Hsl+CEgFuwcCIqj15ZPRNGDF6u66u2Z9+Xan5340oC0F5VojY29AYaK
cKM13KTOn1J+ryP4ge6PbdFlFZzvhlJ+hBYch/WM4Ies2gdeCAS59Jylc/WLHQvOHJF8YlUlmRMd
EqehMuYV9FDOxnbKj/8B/ULtLusvSkm58HxY4to2f9xRkM28UUF8qEgX/ACxMT3QIQV1X8eXdJzk
GpxsPBBHu3tZBK/RQJmJjmeZ5c6CfjpkSHbAb4SGZKhzSrSlDE4RRa/Wtlqvc3XnraRfb0GxtQ68
TR62rnHb4aCZAqZjUKNAt7qQe63TmFjVKhec6ejqWjorB/Nnt7ldEmxod77z/LS9Nd4g/TW5Fpj8
/ToL2Rh27IG+2nLHJhaV/Vu/8q1GXnXMV0PpFvcAOo5UgNJKOWFxNk3FycsRd86PZLlFoqZ/Cf3B
zzRo+QbE/64VvMtJ3/f8HHwyLnXy0rmD4+UCwh66+eaXJIkUzoeBOUI+zXxf7XRO6bOVn/YdFxD9
oARC58K32w91GLJXsH7/gZQYcRzt/cNOPHjA8tTh6NuqEbQ3W1Y1xyJ0yCGsU331xjBg+UmVlbVT
VUrDd50WkNEcRANTsOAl/O806YbsM1nhVNR6eqpF0nRWrmg3mjG5ovp+pGpnXgMzh+eXaELbuk+q
fRiITw3e8oKx8vyaMQ6nSxaCLw9Ye8mxk5mbmzm8/kIrw90S9xmLgVN6a6qCYtf1b14/Eh5+sSc3
AXbRxq64BqntmDBc3do3/ZExix0kDwc6Pajp4xKNS/IKw0RE4M50dJFERB3x8FblLSrXMqLjX+ZJ
dR7QahUiPSgT0KCNTi7MPFWCuJdlqlxOe/ljqmQ1F3QzNzLZwDAuHn6h9XYCGB5CwWIji1BiDDzW
bahrc5y4L3Px2j7ZmxMMnv/5GTeeXW4r5XDgq95dkWFFCX+8xZGiFZIy/e3VTpV18aKh5LQEt8F+
DkRip3dROFNsQa5Km84TGVAmB2BR1CSOQ8BypPHpPyyqAKiIH7l+KEiNryKga0xhy6eDiIhehwTb
NsGA9g3Z194IWMbWb40WNJA3sy/2IviAYt2bJCttoEJNEM2+nu4XpwuQ7oj/h1IgbUf8v9HzLR8G
YnuaP6fXw4ChGd7Xg3gGl/mzjJjafJypTTHFz7g2socx1wYHiaIs+lXfmMofbN0X4pue4XtkoVsb
cWrgmzFd3hCV5n9I7Cyc97AaEYLL7msNM5qwJwfGA6aYA3T4547VzNGK5vgcDDxXOUD987VKkK1Y
+8T1z4YqPw8EJV5OlY+eBS7gJmroxO6LRZQ94wp/G4Y92LW6EUukLgIJOFKgKHn7zEI7fplWC1WM
yNrBlVijcEyJ6/mu2OJVDiwzHJ/XEPj8IOrcn3PWnhc+zt3UKAw3jmH2bzSF+zu6mei2iObai1F3
nMm+TiY0YAiMbUjFkHoVY7HFpO/CWV/PUR7wjrGqqLaoqhpxGBQkwmXyo4EFUuSZNI8hh17pT0lh
hkObX5Eh3SRhJnEbWjBypL7rvD6539SQ8y+QGQQ957ozlwdVXzQ7uJyHoD1KUy7ggL/1Le1ItauG
Jin25sMhyeCCUCTYdam9e+PTCO3WALRZGD1P6Is3P0HyBBgJZ6NNGXVjs70pgCdEL20RKaZnvl/z
xnZ9D1A/x4vu5t4cqo/mshRAh93vdPe4LYjmO1FqKlPkgPKmqR0Kl/o4avvGomqmhjkiqxaI50Dg
oV7SYoofq4vihtsK1jFsrBhH5RyGyiRDZlGYjJYUfBLw8DT5OVKTwsg1bvC+hmNAzBGz5qhjoff+
z4DpAhI99HZmin8W4GJP5tvda9vCv7C61hE66nml8fpdiIHoIzvWu3TEWFHsa2xQUUC6543t2DHM
F8TXapS9jLtAkaNGLAXJ9oT3vcb9PdRcpq3f4J77lbV+XVsaA+KVNJht/fpQ2Q16IukmmMN36g0t
sjTsG+ZMVjuErUdHWVCg0e/dsR/atrbZByeIRJe6JlogTHrqUgmFgN+lLXXhTikir+0xv2nizPlO
2Svdzh+O7M1Ra14bh07AM7816vylGmOSmYh8A0pnctNQKjnV6LKTZSJJZP67GPzfOfI2vwkUcHVD
fhgd7BnvApR9apPblArF8dYotjKuYpT6oAbMD/l2lwN6+Yfs2BYwu0aYTdo8AAk8fX5DNuB1oklT
jzDSYKJoZ0xLJAvXyfZ62PA999QpBOqHFiTu37e5D/jYO5wf3DXEewkGH/YNNLkcn3y8Ktah0TrP
gklKz5hMeUe5sn58Haso0nJwgmOlqzezZEurwbr4ZDsv0CdqfCaAL+B7Zc3b/RMPlM2YuJ3PO0AU
b28eo1y2wreFf5HaWQPmW7i0irKQWrctrzdQ0b+2N60ObI8ny4YQ/SuYpVWv4xNw49lOMSvfrvLc
cbs3D4B3e4Oa/Yn3pljb56m6BeDtALNF5K+P/7TXbCsob/5gXarHY+UNPgv6xI+fqaqO4iKBGKPW
GkADg93NgeAWdwTeTpUhw6lXQGsFBQTuWB7ScyMldTJRJYmpNNAFrec46rX/3jKdKV60Ob5V2BXM
HaJeMJnd4gr/Sc6SQRyASr/Fw7jUg815cz6vWhPUo2p+HydUDc+eZCvqD9Ek3WLL4uTZwJSsYUOW
79oQ83Rdz5K5/2eJpxFmo+3UadZxqncrjQU1eJo0iuHGMzaD9I53xzVmo5t3+B0b+tc7JJN+45Ej
1DM2i6zN7lL2utZrWsEXL+mbV1LsqRjJEASsmJ1zp3TGLd/Gy0pBPyYHn7JqJ0PpLSuLQqLEYwjk
X7/luYNunED+PaxHNg/SFuUEOPAhUrMiA6PmJyDO+uCtppDVfWdbZTkeYH5Qu3Q7T/hNQLSjJHN2
CwX76Xar0QEwGeDzMI49p5WY81NG3FJthjoiq5xSzz384yReSPmZV5/0oJE0B0FU9SdgE/qISzeD
Ww/KsSQZAfX4kHPQ2uRLtOgCEGi9/TFqDeXwybxMw2Y+2sqOtNKfanjp7aiM7+eHttcLKhkVzZSz
k/lWUH68ZRor8PVLKEspS0Wtx3g/2TUqYFcweC9V1nkJo4i14EZCRIrGJSCT1L9B3XygQidIb+0p
y2uFnIY7WR7H2KZgIuHRHSb2OX8PFeA6bQrduWGPXpfRQf2BMqCExZmvoi7hSyIB+67Pjf90GS4r
TuRxMOVahznZdxKHhkvcDGVY6qDUc8NtRO1qQS436Ku0SRgPwUG1zlqBfaSr2Ja89d5tUnjYLgYO
dwt9QNsgt808JI7ew4811CWWL1jyvgozwVECy4EFBNFQn+tQ/oSpg6VtGhNE2QQbrw0bMC7Nf3rp
IQeSl80CiAp7lOWpy694WbJT+9MAzvuye0Nj+ksyfCJRy9/jTpBYk1FQ/X6nI73Bn6xECVgY/pm+
7lQZZSz/mviBCNtuVvcMfCAmixWQmIH/3n/Zm8RXppNFmLycD8cvga9LRk2pq3Ce3+pwLHG5AYuf
HW5JD37od/MJ1U1Na0aXNefzKou3o61Y24y3hYwEZ/sRCIMPStF4DaoX/c7aKEj3ynpStVOnfVRH
TLA6kzufEs5IGoKO59wiKjEZMcqB4furEO9yEy4ul39Wr1U2hRbXTbdX0BmQ7Fyr52KbmtmcoDnk
ToThRuTUmkG40zJYtrMwbErBo69R0PKCQKUqFyI30QJMrJFou3m8aabMGY1MBdUamt7YFIm2YTXU
77ZrZmmV0KrX5w0t3o6tsQjZUPaVhAhNnwlyQvP0KWQfF4Cj3n9hsZn4JBI3VVEJRP9Zi4JT5j9/
X8CUzJmgIVsj3+nnuVZ7G9k5EVhJiRjvXC7jRkbQ2BFM0PXWbzzADlj+g7i4n1d5HnqIIgpFHHgk
PylwZkuaCT9BDafLqIoFfM09ADwoDUBEhyqeq16M6f/OpOkW80DmwMeuTtwHYR4efDG8CT+R2zkz
QeqIyXfgqHHjV+ASEHqLdj0NlQ02pCH0P3FBCw1+LsokukeV+mI+VNLiKOj9oQt+5LU7Q3NJlhuM
0lCFqA0KgC+LbbhvRYJY1TQCYLJvLfcOpN0sgvU5xyK5mhSI57jIWWcie38Z4beLT0DgVsdWNM7k
fnNfFe87BGS9if2hPbusCZL4bKUwZjlhZkTZAKSLZtqp9Gz9lfh/3vMPP2aF0rXJrP/FMzz2EWdp
Zn9Skuymjd++Bhaa5ifF2pDOCtBimG9SxE4BkB1VqKClHT16rrk3jWzGhUv8CWAIGueWQlWnVd9k
uxbsPZLGiXAje+q+/e1tsAnuSN1NVxPcT+TaLzLq2wScdCVvdOYLo0SHDe+PGWGxlswB3swcSrbb
INDZ/bHEKNVyqrKJV6x5YGmGdbohx+9jjCWu2QwBXA36l1vPDxvs0yHDxxvQNETTClqmILJ/H0jd
uVyh0OZmK3XGtum+P8RDLdJgZP627qQrEhIJPyWZEuxUEujTNldesEyatn+hxHqKZ1pK/WPr4jr/
B3BLxIvJQi531m+1PgJqHBrQhkJDYf8xiLSsCZh2RSb+6rxksYjCXFmrwk30OA3mMH93VTSUCoF1
1DFP1DJDHjTahLHra6gkEysV71hrI6VrYd9babNDdrf8fv4jnF5FErO5etcuNp/UdwBMuermmjVm
CFavYE6BMScT5w5c1Eiwx2fkH5QJ3WTSubF8JH7KLkzKBQ0q8ZSQ2GmZwD1DoXJKwOAZv4ZnAS8k
PP87shZLQFiCisXoAMrlSh9wu5XXJRxKxGD4qv2scFIHYEBz1UQi0P59MMNOyo5ZPDgF2jLs4ymq
S9Qs+EkeKiEdlp3gyLZHPcU3t/dyF3DGPRIexzgv9xi1hyQpVH3ZavyKMbAlkukrSB1+sUL5roI3
wcHk0xh+nNO6l1gMSNHbikcrUGwf5DF4Q2LrX62ZZ3kZftChg7mwlSZKe3DCQMD6PA82aBVfrGdZ
mb2SJOPGGImStTlRT7XQZXbWX510B5+V1PCUb3DTnijb1KGx894IxckHxYPM7Z9NkWGJpyNIPZoa
Ecofp0Ia2hvUB+D7DB438lno929EUVchl+zw9x5Wea1Px+NocYPzqOWHxQeIpA6fNBDaMw2+yLz1
bNwTmKAwGxJyXdvlw2TJc4/9LVqxmn/LFKuYsYcweB7TSk/TmjmMs0zV2m/St4Q+0NhTcJJ3KDqm
0zu9hKKaS1HArSOupBzx5Yt2bM5wzaNtzC6EUuolHpPAi63GLwMMx8qlGpono8FYLEmtuzvf97a5
QlNr8Nyylx/bx+MMS1FXTfxd8251zuiGWCUpBxYgRCMWxGpvBgIOLylOLjzGw+8rQn9kIdZae32o
3jpyCfrt4mw3d9cjXBJHkLUEwXrMbtT+WGGHOmh3zGlMnXevxvSVy6yrtQ7LPO5/siWbw663TR1F
4W181z1pD1A5tb2SzuiQIYHGs8exc43c4jmn2g5h93JoO5luteNZYv4adEQDycEadAn5H9BAoF3m
fZoMHSr/Q49Sv/TN2633FaIwe5MwpuUpTPDYkrHkYZe+MIIMiPUn0SYCIcDpqKfX6VS4FZIIILxl
dptTHIP+HrK/lUAtEv4+BU5bX9Gro01IyOeoZ+rkoIs52MHcnWyOBP8UsPWeAUVYZATvFhjw0Tzj
RH6AQUO3Z8XXEmsXo7V9SN/kYXOB2COHDd4wyF9ikV5VftcfHzUj5wV6sIN4XTXJSncyhwTRYN2W
ASIatPxMOOjHVak0EMP0BDCL86VftTcG0UhC0MaOAyT4HWEis3V2Xhv+Oth/KDOC4eoUXYsiYbDA
x0DN4SwLsSzwWe4aPBhGOqdSBOpoMC15qjdfXIhKUCWixTnlts6L4GCM8LRiAnqwU4ffEkiDyvzn
QO1pZGE14qm76eNFPaT/4uee3LkqzvKPUQ7yra7Q8spPRMNEx5EWnsaz63UAkva6aRPZ+qDwBamm
9RUWucCL3e6BiTDjfsOYb5NWFQN+z39fVeiWhUZ1UMTxKw+ZE5xyPCydBOEHQ12ft61cH9PlGke2
fBb4yEfng6uwgh9+lDwrr68VEFHZOF+UHp5dmkkrkJciBX4mleMwxNNyrS4E/DEj+r9tf5qb1xWT
HEoWvAiP47OwhFWriZwHrSSqxxjDlHEPH1xtMEEm0y10VJkXzxreLaZ33rYWrMuLnvTAjzTGKUd3
ca6Y1e3m+PhhRPoVRrwv9Xa0NwgtS9Lzx7zTWrvKDYR5cSWGfc6Mtbw8gF1+hLH4q5QZKHGoZPYz
4OH49TdGn4sPLoWx4+boQYBZiLNwEoWqdhcThSFCRruO3cOJiYEebpqUCoynKJpTKzV0yXV0b5fy
eU0J7MNv2q+lAWKT9JsDntu4wqnE5Xsk7QTs069tJ8pKqebvO/eLOcvGs5HZa7uxikjHxwnuH6Ud
Fiyg9GLT5t37cpmH6WoHZnu2Z79rIwzPLwHd71X2xuH+YSQ3vPmMhcZSXeNA4Baw6TCvyrhzZsC6
bg4C3mqhYIIixS5Lp+aJX/TZ4KUNOnzCGFmkNZBP5A9hYHAuyGLRvyyrtpc3XU6hFPms5b1iC9Xo
XTL37Ks2MPE9jdC2K6Idojjgobi1zXN1EBcoE+ARCjcB9zCocW1yCqDMA6trQTLHy4IOcAASpSZt
lugkBXGs40RVNVVaY+mdmZvJGoWESwKd19CuB93tjH8uNH3JxfKjiEoxPlohTMlhxY3Q7nBXat50
OuGZaDLR4aDcseCqWilaz1AcXcLsMZuNoja5zcgiJ3o6Mb0uuW08I3fSid/qEKVx2xn08TOcr6m/
9Gmp3NBMGyvB5z11D6/zAg/lcdARHVgj1o6dxkbMeMhNVCW6N+vSOBAUmeT0OJu65hJBGQCZDebu
4Jh2f65yVqrJjIycCpUpnrzb5V/st8MchOvcgvFWUhRpR967ui4t1ddcfXXAkitiwosLyvfxcel1
mJZ4eCAwWwvmlV7j+XvDw2d0My9bsFl58X2mEPIRL+Cqc4rE86LBFBQKYVj8o8bzik0yMLfB2JC7
Yd8xNyzVKjZosUyCFLfTmk7EFEG/Rtp/BTEXtkMDMkQGmar7pXDwyIKybRKSfL+at0fcHwY+TMTt
yi9RumODTTiVPDoHElrl0CHWgrMC3d2OT4c4wfC45hF7QJlcxj/osZIoHO37KPXBXbCgfzwqcEUG
9lorYFFcmwxYTiVPKOLMuCzxYjZ6y0wJ3362cp4Cpr0svRVUgVevnfMUj5QxkxIFFOzaOswBO1vO
rWdTFQEdC8ApwHNYkwzNxRoMKNZEXv2hXTbCiB+g64dWVOs/B/RBlqz8xRcHLMbWbXDu3It9ELZ1
g2cUPaz3n7gmiAQBV/f1JxBb1n1F3c9rLLF+sPLpslfssZg7F9lI3FibhUpyhnKpc5YHL2EhRRti
yIf5NzDANwXsUQUaVNvmeMK4gqc1S+y31ScDTKoZtRjngCJdEkxV06yhXkAAk0ks72U1ShXs1Lj8
XhA0pATt5TnOjuiGhIgF8lSDabrV5OpjkyxbKXWfiGSzwblQbVhsE0vRgogQ13Msb+mktPpu343X
6MF+MtD+i8ZPyfPwJlYYk2jC3kuSOyfJzly8Iz8VXdMGe58bnDR5lfaeeTkWrKrBCyIDpuTuftaP
8L+xxQk3Kge7Z+75gkkgaaGATHuiS5LvqzUh79BFTBMucbe3f1lcrFvmbp0/W3Lodje7k4p8zD/W
f1d+lYcRiKxSyXpy4SvvviigvsbWp8gcnlqsksYHLOQhHKcUSx/30YQNVQcfx9fWnEjTzCSG5wKI
IZ9ddlGW/rTP9QODbUVXlgxV1ury7K7YhYinySoKROHn5D2H8k46R4P3Jv7yYoxXCu6tIqyJJTb9
qlMLkKs91S2KY6CuUqQp47h2Li8yD/pOzZNoqpkaXoXE3/NH8xXww0As+e4i+tUqJ2NmYcrE5VpN
bRZUGh8c7VoVWxH4PdGwDVtzGcXTkVhm+YAAb3DJVp+Amq+5oATNfBjceeFEohFhD8cDLiko/URr
AvaIjzpeCF7rhQpACASfSONoG2xpuylWGTcfJEK1W8PnB3DGP3U1kY3s7EtpMkETDqiwPRusr3Ft
BPYsP55S0h2Oi6Ssj2U6EDPgvimYQIvKrkxWrDVw1QhPVUTf+qgNiHIXlCxPOrymePcb3Vp0i2Nk
mOvfi3H/7FdWQ9//FZtFRW2C3XwxGvtlw945fkQg+Pk6S+rpeUWEqeBGTAoDkDdnDbJRIva6IVx7
7H4e2JgPTK0/UvVY4p4bOxT8yFDLyM223MvlW//aaB4vlGZPM1JEVMRuKSN0IGJsuj+tcqcCEBBL
Eez/lJcK2kw9Nckr5DbedFGil6yXxBWvQzFU4YJJGylz/CQ+be2kftYekwIWWL5O4I6v7FEHjDgd
ucrob+t60BgXv3c/N24poJ5Zak5hxpiuOHQSv3owOlJVxyj4VvpQ4RZY2QMdZKkon+eyORNWfuQA
BxGg5sVEv81W+mpWYZQ8qeWm+Ut2kBBb0ISZjU2pkf/MzFS4kJ2KDuCoW5js+21SwScB0SkHPKoH
kLqLanKGB+sEv5mRjH+CP/gVYq7g7wJfNGw2TMXNxa3wxpb27gJ0xBvRIjijUIvcgP1s6CIe8QIe
2x9+h9EO9Rps/RkzEBU+6JPUrEbj4hvmHBhbW5IN7K3HbgR0u6olWYoi0Yp225Ae5QYc1mmg2z82
v18FoQKk1NI3IPs2wTcGRTaD6BqyymgGjHRmB/eB2K+5Y2LqX1DK1nslJbh1rTzlebMOyw7Kneat
5vAbzNQnj6E4NNYSTahuAuGIYojj95XtWihNKjW1JSpJcomsvRbOWEUoSdDHo1fzeM6J6dY7AbyB
igfYZ5OHWLoPFxSdtPA5nZRZhDMmnyitzc90XbqMtvRBSu7fHCUitEe8a/aBfczkVhvBpvGgFjn7
Bs0HxInw08e8Ou1r62ZUkqsTJdsz/TVHb02DhiUXVrdMVnZv0wEA0KiC6Vz7RPyTohJ1ipmyZdXu
1faVtiKHAkYf3mJkYCSlSmYl9PxnBuYQvw9Q+qIR4jM3N0F0aU9SWGAcurgJUo6x5KXPOxiQnxOx
1g+O+7i5hr3LhVkLT3W9LHdPR6OeHDKRCDTSFHjDWWNG6TwdXV7LpYOGuSa8B+O3FTTowuUap/N+
7R2C/VW3myhK9gmQKsAMEY4eaAOfgjSRGCkcZx/KC1FaT+Yn0/R8w98ReOkR0+qVFOAmthWMLQ7e
44thpJVAjKo0jxoiaJEFXbtcvaroYIo7Z+jotSYYnsf4XC8wsDDmIR0HT+lwxa6H1dtqBUwYiozw
pYcvD5Bqq6uGtJb0t/MAKCRHLpFrHXMHUIp8h0YL5Le2P+yyCQMSqLdWK49Y240Ef5EnabqVdHYF
kIOM8S7wpbMuL6f0xIk2bBETE6wERt8E1vVs3HaN/LD2r/C8QVKCMdKl0Y9O1JrYmADglFbI00R1
z9ShEwZtJyuaeJz7AiHyHoTMuPwzvSUj0xWngUEZsbzA6YAzABsCN4raAek/PxmcnR6o0s+mpVd6
rlRN6TMAncPt2CTGsQJ3XdHjHx4yrHLdWZfadOe4PMNwDtrt5r9TeRm3NW5TaQjGc/dIat9fwAq6
sGWpbE1am0+cIr6GtSzYwdOeMDfIHmNAE4tX2qmUTteLUX6HNgo1fyDnXxotzzcJ0+y/avGD2cco
+R6bxbDvyFGx5Ex06Q7Qqjns8e6SjXsYEaDgZ8pxo3i9NoN0uFg1DtPVeXe3SVA1+GDdR4uWi3sJ
8M9+TDrZvA3lwNMy91Pc347fDq6rYT6Zzf80vobzVb8Ubq05vSVtr08yvstgJBJMpC5xsjwVf3vP
gnIoirC6YmvHgQqTyBWgYlq9cdRFrPK0KopEIXtwPXOWc6fo9FDFzFxHlAkPRgItzB/xfJE5V4cA
xZSEAuhcnxLrR/lpUG2UU3gqwgTZo8AXyz6o15e6p6T1d6eDZPlokZvaLe2cRNnO8vtgC6QbCv91
77+8TfGy5khiYj4XLP0mn+wJwAz8zeD49yxcmVx6L+XqH+aXV5IDOPOEreiRLZubemARQKHRWQIw
1Caai8WrIJIF7ccU35maAx7y+G2C27Stkq4O4hAHQfNUD9eQ6KmvAEGqVZrkx7E/qzwlFzUaA5W7
MOEnjKdDXj929czgs0qnuC0NfRWQ/s9O91fsKa1i/mToqWV3v0Xrpk1m4SproeDvuhM+FLLC05H2
vYqyd8FeHwgl9Wr7UbjTYafm/v33aEAewTGV5dmIPr0rRg5DwE8xb+mH+4O1h4eKp4JaePNTRbS8
sOJiT20BJEfSxlcj15V4r20JFju3kkltNs8r4CU5jI1tfWC4U9mme8wa+LJ0LwgWsjRP8Fw4HosF
fzxYWaWXRNF6sA78jFmw30EZYUNjVQDyeLaOSISQ83DwFAjx4hd4hbjEcwVVEu/mCfLV6DQjjgBP
M8Cdw6JKq+LZBGodb2VyHZcN+pS2skJVGMIZlhyt6iqbkvTYdRmM7VXMeKMESLexqCGnWhzMDFhK
ltmzmX9MXz5Z2KXHOvoAk3nCxhIWj9N0QNhV/4wPkuMWrZJw470HpGK8N6+g++d87LbAMQSTJxX/
8pAUSjdrgriYv1D41R7OwUoTuxvkwG3RB9W/iWiGRxOFBEG4gyUCDBm/Y4qe5VZCxG+BVJe8c8+F
Xmf2vyl0yHGSmoZyU/6joQsb1l+Fb4mjmXHZ6H9PO1x+N28vAW8z9So5McAQQc8iaQOBetyGY24T
1AmE1Iy99vPHEIvSsam0OjGYVxo5eiuXFFj20FwIBCMryjAqvjpdIeXmhwcVijyWg5W76bfe3BUv
qBxe5AYzcrGrkkpIoHiCy9pGHhg7S3rOkXRyvgBT92jfaR8QUNjx+i+fU2KyVASnIjX2+aKChty1
vnvTeu0l2wL7n1dHqycWILKYeORJxtkrWEspiZ6DpzCFk4xw1YBqwgRKpWexs+4F6etG6R6yaX10
powAGBSnP49Gxl4yjXs6M0aw4pp8B6yI/ZyYxt7JiuYToK/WH0vpI9/0JhCL/u1qzxoz0skQhXJI
TQdlQy+z/tHLVBRW3AFG4cIuIG1G+49j+7yMf8n2/n/NqZH+o3YX27tG8zr3SfYL+3YHPjM2qlyB
gcLQmw7r1ZM1m6Jh8n9XKV9SKuWh7lckqz7OxFtmFH/9RsACw+iYSyH32HGA6l2McKc7E/UvTTKH
XaKC63BZ1DZ114Rsqm/AUEGGgB1h/4VNCT1OuFb/7IfBWzs4Ye3k/YYk5qG7d3dASxG3ef7wmEic
xIKUK5vPKeImGTkUAZUGOaLLapPAMsU/RMC1l/slq04HLc4p4iwdomlHs9WiHFCKQ6dl+mSe9dm3
X7ZOBrrFRsZjLZceXRwlbvU1CLXlyaKTaloJRUS3xhgEquRrOhZ+nThwMUh/pmbiqN9WlwJyULC/
2VnA6hzyTySA2e0BONTFrNFnJJ2m8GzvHYNuldkT+PJr1V0220ga2EF7btknlpjuVWxHwBrmSJwM
mJa105Xmt/qJywdg2PGAztgzQUJpav1ytNCpBcfJiJYP9AfEfAjNdtns6V5SAtt5XMZRPQWbTbNE
aJiTfBFi+T5XFeoRF4DcBVcP3BFFPlz5xOVXS5yjM9BrnrC9+ORcbKu+PsTrIui6OuWC0eDGWtir
4r+TI71yCALX1znRLubEZYANdWR62dhEjsI4CtdZ/jVnksZvYA86v/6s2BVG/tUfxevh8LIHiHJi
PieKMnaNTKqne7FX0gbfJGViZIth6KL5UPbH0p5qyBD7ALbJvw90R1w2CyTkr6i2X4hmpWzVJYYA
9sfLbndXJrokicBn/cL+HPZytTKl3OlKL9RdBDRPcmV2V0xF++jj+1ZNqM+d17KOSCSrg3LispOg
VCN+WXgPohztXgiJaayYhV/6j/ztw4EQR+MgihN/ZHPbwDLC9750onbKwXakTlTxohNKGFEkcGM1
5FkEItxk452QkcACkvQ7vNNDgQZwlTgu6ErlG1P9apBgfOnt/HkJK7GMJ3AiUBMqCuenj0zbTuO6
CjVy5yvzN1UF3RoQigguq87ORiWyLtkFGV0+3EKHaRfQpr5N3ULOLzCpUTWOuGhElisQQ04Xa+OC
iZC3G0WhGJPiFX69gkPCxpDfZcDFbY1RpGgd+9CcSJuoJfE3zVUpRF23278OPmk7SvdzalrgF/hT
fNtxkh/3faCFTPDOft4VB3E53zSOF37r0atTr8je5ncuVbd34hMAR8laRj/sySdIuGF2Ih5WD0PW
3cwOPDxdUpTTF611bTApda9cRCYYF007/NC6X8GKYbMAHraDnmL8vDsU7aZqvUpxmXlx+fFC4N8t
QJVM7ax17BDtrUAy6jk4lVTgn0c0e+FIpG0WBt5UuExD2fn3N0T9Te18h1dLu79tLpYsyQTKYn6N
zeR829xlzo0eq+J01ooBS/RfYNvjcN/EWvHMe4uXRAazmxuKPC+4BVuRJ63akqyw0k3W3Idntk5M
krDKZqBtgWJYDIVNcK5mzyDFsR2Ay0NNuMoXBfAGTY5h5nCi+sjsQaYfjZDwXlDG4+bvhQm7tk6c
0k8tPfCuvXRJwVfsJUiqY5DWDL8fUnRAbPvUe2mSKDZtQd06T6GmEC/bXRxfde0NTay9RD+5TUAQ
mDWsvVEn1PsFy8f9P9FlfUwGsm0eJpkEZwVBVDJyjjVWGrBCUQbDqCOcG/mtr6IJqu0xQWQYLnE5
y6V0lGru3rvnaqc/hyPucp5FUXRDTkbDf0YMWxDgH7q7FCDPqnOIIHX9XByh4L9ll1Vl8uwPkm20
szRgU4tPh6XD+PUM0Y219v9lCs6vcYXjMdIzmAKjffHxjNwZRVoyKZLfZETHUVPVZEPWyo6HWa8i
XmrDlyhkmeKC9OlNBhkyTZnibxNm86cFW40WZY9c0RRaxSce2WMT7v/pbJnBGFqrFOVgyVeg9dSy
e4tbGSHdMtXPzTP4k6DoeDvIrMWRJhHPPfH46eDK8koP2LqJkjDKxRTPHgQN6OtAELi4QkFZnwJG
ebm199o7N3eb21X71TnEwnLHuujf5ntnPQkOeGoaHqBDi9r1WD7YvZDijqykPHVfuwqLX0qaaiDS
oPiknz0DlgyYmmdgGv2RhF/zdFSyL57IjdjJlXAytNt336r+Cpar8HEZ9UrJslkEuB4oLNXeoLUT
JuK2Dj4mLmpUUxOxE16Hu1uLpnyvcyk1S1gd7ETk+hT5aLw2oQRA4LJ2tF+WtRb01d0Wlz+IjgTM
MlzpusMTOidr9KnI/RlAACKN5UUM6rKb1F6fA+4W1IvqPJ0o1GA8kiOWk+HPo7fkkTq/p6MF4duW
aXUcOVkEfky7HHLC6N1KSU+0B/LuFIOAMZfODLWnOql+3EyT4rGIQ27d7ayYUL83jFfk5YTipG7A
fLd5gQR6yZEJSdN6Z60t8Tm2+9SRz4cQ4Sg69HWmhCMLTealtdB3VtaVS/zQ9o9B0XOGh/2oucr4
V9ps9LkCvs8VUOebLgROjLfLHuK20+/5NJpohAQy65PtI9LYByoR4lrU71NIMVCpTiEqgt4Me1A0
WErMYIQwjLoXbNJQBPo7h/lmueoTiY1Ecb2Cbqh2cCutDPaX8/bb7lEXaWyqF5NkVJYNPVZDXTDa
+zx3ku/pm+MUXpOU8lx4VWmd1L8Vgq3j8R1n7eKsLYUVrvh9wnBXfinx2fx9aRAGDstM57JBmZpA
5suU/2UUhCftM0U3nAyNtTsqVAVnUmfWjXe2GVCizS5DDb4ZbxB9do+lOBy8SMBxvEEHAZlWPT1k
EI2cFPxGnaC+15IC4ta1jozbqhc17y0WqdjaZjrGUiCuFE8tpZeWavfS0spfCBp5w5QOTO+4UINo
mDrhH8+pKDKZ36Pk1lx6rxJcjVI1JbiCcut/PrvjmPEASUWzKPUfe4oyNE4qW0EgFi+vS+1P7wxL
Qxn9v3jkvgm/Qod8JtIVA0s/Oy9UTawlCBWl7xfXlqw091Vie/eRprxl7XPa3m23ePF5F/xW4bF0
0CU+bozvddVDjXwcYZQLv5rpGAwHK7234/lv1XIpwJFp/c2AxuIuhhFoqdzxeuA0MOfPZqZgUTNo
hmSqz6vN2SQLrQerIc+C56c8C3AyglefOrp5hi+onqutMPcgF1IHVp3Y/nxlBtq4kWL4WJtYe/TW
nVoEcXcFrbkoGXAt4l5FeivWozJG8iYNSh/urDhq+DQE1KsEd+OkTaL/SCNHjbWjwz4wQsS0w+Gp
RSxfgiDlWMqcPCvCQBiPuv4Tc/WgPSAN8p/cKKJDrOE1UVzFpzOQI4m9eqvbXr7uayhWavVav4HU
aYHgA8xazVqlDmpSJJ0qFZDgQoGeVl6ujoBp1D0jtGarGosI0mdS3WT7+UMiY94WV/oYnsE+K3GH
ntvTTMTrkGGqCY2tyM2/knb/P65h/UC+aRhGOG7bsjUTZ+eqkAJbS+pY/EVpl116Dm+/Za4uqnQh
dcgLh11axPSeP/eCsDXbnAwpRHqbD3JtEuhsXUxc55V86t7gyAR58avFKvPR6Tj4DIS7BZkPegFr
odMTUVo0o5l1xkaKR0uBu4QcbE8/Exi1hE0AaEe7Wk5GvyEjyWXhFsyr8MNk8c4lPejeGEH8Iitj
+IfuxZ5/kU2efoRIUfJNq7cY4c64HxVYzxb6Ri6F8KzX7w72jP4Mxh+Mxk/QO0L3Jo3AQaBlQkY6
4h77VLgZMlyEFdoKl2j0GJidcIH1Y39YOJeTxEyPMwApM61Y7/J4HG4zFABA5FquxUVY8Ps7TH04
+SDxJGMkouWFdD/77sYl8L50VW+UIZ4elTZK9FmkUCDuQEx0m6/EcANvcqqd5GJ7c90G+a9cueVO
NOpIe1+GSoHJGRF3Zfh7YcSIPIQTGp/9DJWIPYMoC8XTjC33VrZqT+er9lv8kRtuHnQ4Bsw8Zd6/
br9JOLlEGtvMaz40MaxuQRsAnFwJ6DudSE2rXdyNooeyolRxYKhSr5wXJRE6LFncy3eChs0yeMvm
Qttj94gSUUSqArT80/CETiNxt0oQ/DRyfjrW34U8IKAwiBwz6VDGYGnhsK9OOh+6wrou+I3JnIBD
UQAWw5QoTMUH1nNyK7aa30s+YXcMjw0DsZCddcNMVvE+C1KgqTwC+EKupOTccE/deWsY+A+roQUd
fAS8nsbakVZQCPKhXg7Xv9z40/clhTSVFQq4QRYWlPu1k2toLZsNesEI1mrAKMQhpc2a+e4gAJ0e
6g4HQDIZPu+3Ue2DnfQ9MMHeJJ/elN+ckYMZbkcBerWbdWUGONIKVhv+NcBMjsclvc7ZikZl0M2F
AKVoiZwkV0KczE4AsfNZF2c21XWqd6DMc0x9vNzVGtisAcRQ5FMbhcIQo/sD/GQORpd/PbMjIuDH
nU1yWZG6xp2t4mhdK8kXNDliZ5mfbFZv7kbtJTlBJuT4Hl4wKFfg6WRzNoIafd9REind7nJzOU/M
nQYLFtP9Eia0ogtFO3j0sb9akk/oNjRCVCVZjKZVPUi0am3JYR/X3czcApdsCI9rW2AgJx299oRM
ikN/p+NaVMoV6QbPKq1FuprxItmOsDoKgu4o/28H9VtqQopa5Lov+o1mrcruLFGRx5bJjleJmH/D
eNHiTIZ0A4Hri7pu7UYDF7S2FruCOUTWKyuDKlzebNW+uUyVICls6wtPe362u+XheJGZz70Po1hi
dF5WtK4jOy9hWNB+xtDQfyyBDMVFGCxYMsYxhTCoxuwUc+4UX8ikBcGVIVAIOdywHteGknuNSDIi
zN2ANdXz0klrzZ0BE/LMZfk7jMmqdQzMKEkep3tJnt6NSsqhsTeEYgVc+0bxl0WCTvGd/a0/ujAx
iYdUEsh4JAWc2tYx+D0nkTntPqTaQIlUkwt1iqRzyZTc2G6ipSAvawawxW6Kpdj86egUtn3yU1HC
U5d+JCC5MM2R6PMj9R+NBBfPZc2tsoOIF7lHVPVDI5XC8AtmVPabX6YJzIDUSID0zrYT4vE62Ovw
RAhuNbHkJKnkBPtkxzKJ1mMBz0DTznmPu4JkjGs7JTjSStDekQAuqaxPrI6vdv/pPwWFN4iJsnll
UsuJ2cx0DBCW5uvtsqfskRm1iOSNlwiwsy87oCBxolrH7w4Gsw7vzTq4d+sd3gekjshtLbyMFZMs
QvUqeqdbXTzMpVjUTuF/aOCppF+FoCwI9flrMMOzbm5d/XMJG1hPCPTQ9jt/s/tFlUG9ogryl98o
2zRH6vr0n9m8jOqVZtpkddJQXdb0NMoy1jHzFpxqBz3qB+zUj7Tj35sgJ2Cl8LTqYnGU/N0h0DiP
Ze430EGuwRRLyJiSTAEVh0UuSOXGgihECgCiJI2rLewsElfzz1U4xK8qPX/AHQwr4BPtXxw04hHw
gDhlTZGi4q6lL15UxMBuVPErujrQEbpxCesJQ1L6zKd1PBrC8zp4dsQh0c9AFT/s86lAVN0u56fc
e7ybOna6IyliX+3Ff3gKmflSNunlv3gf9OZf7o/AAduhFspziX56L9W0Eltyci7INqzcl0YoER7I
xCpsQ0QRZO4mDdkof9137qtbM1Wtq4Zsdg7DdVyiZPhbOz+7yhj0IoKfwS0SahwJxrcoeOyKRfAx
e/WbdyLXuseTalhOrZ8RlJEX9W6PrHQK73sFY1qM1gaaxx2KTQgD3e+PEfhv4OUED+vIBVnjO2vv
zMCIQjPWrK8FINfBSS0DpvoxaoJCNZSCoYgJi020xD1iKMkYIqqFF4uiAXW0wYW2lu1VnbHQDGzA
4a/MJ3Npa2NY0Rk+huTG3FSPm3LG9OJDdpeujGcDAT6P0s/BymZiYXvU3cY/JZnLjOCmD4zCImd6
7IqJsjWhihudg0t9xgdrfcJf5C0zrUdJdxUphJFBf0KmRWzVd+1ysAwRT9NtM/IpgOhbucdGeRel
sKMdIKv9HBp342LWS5oB9ha2eb673xteuVF8pe0o4n8nU4ISLiqrblKjUlliRFc2duOp2rBMwgaH
zQM85grv4nYsiYyaZNN1mdgvZl7MoswFJ1HkvSdM3lsnwmr4kuxVGBbWUIp1ksR8Bd/S56wmI9NW
i9eZ7EXKOjdhy3v/rc/McGOxXrBVGodLZ5Ml9UAa/h+fs4LDgdg01pzFSNwCVUtXBKHGGofRVjVz
SQ+ZkaCDni9PB1HCN9QY+PUc2Y//C902Wsrb6zKG+Cy6SiEWjfckM3Sq8BY5lEzrFm7QC21o2SID
XIYVjMRQqmU0dFm1q3A0WeTEXuU/ofkxjIzdlcD4iZayz49l15BMAmWk8acPPhQ90azTHGQN/JXf
jaPZEEqMXSa1sgrwzkl71MHA975MzonacF+Z/AlRv5JG6a21I58WNz2oAT55lQb+BM1l3MHjWlDy
RVRPIdQy5uGcD8RQcszmz0RJrZqGISDEQRPUSxOi8F3bvu0agBX2WtQDhZNPu0ja4/q260U+BXJQ
Va1YKGT6FmZL1pdB27pUlIkoQwbj4F7bEbtXDbnxaEL0gZpUAbozmTho0IeCqxHbNT0D+WfsedRm
rFnmhccx6WCx5lB+9sYJvem/N79j6ARnCUF4OpSixUCmfq/c4hhfeC2Hqow8BoiPwYhlwItMfaGY
CRp9btI+4dT9ZTV/4+wHBv+PooaFJ81fRWe4jwIqtdsuP6f8gUPTIuyP/OHlursUWFIXXAJZ4Rt6
CSltBPRdhUa5b5N6SMstIlMcSd9ZdoPYZBlJ3GJ1kVTrqqEEHor5mggYGvjcfb2DJSsG3Nw8SkFP
d9Bbkzy/N6X7uZ6nGHWFHhlcAqVFT3WoniuBDwG2ed8vpcG17U6MEiRn/2aHPyC7AYd3oDCZw+er
Y9XMxqDBHDBLxyXco/WetYFA899TthPOkOIvarwQ7K7SoYQjc2EuteqKC63f9S2yWFFLjNgdwV2A
H3CmLB38HGhUrzh8BeV451PAoVrn3IIrJxfaqNYTNTkHhFcJYkuQ8jvSIephNPgPn1PgxZbfT0/o
3TIfN1vDJfaAvMLYVwZIJ5vdIyKpUG48Lnm0hcLbYLV2CGgwLEot2Ki9Q9pmlnIhiplaiRvK42N5
2KpU20aw55wzOijEFS0puUFlFDgYqoMMfsmfRWrU5m21ng8RAsFFH1n7/PKjRt1DG+PQQ1Ay5AFo
33n3X5yfzCStaD1f+ajzJDdQJT0L0SYMWHxphoCwrAyXyjT0SlfMa4IFZr5Z/NBRGOce/j+rsZOI
OvQXu9+dC3TqmA+IKyhENrTb6ePoGE1By5i+0TQ0U5e/D6K65LyvF0ObUnUKOa4MCyPDULt29JNE
AAmzpdxiFVIGkdoVdmxlSlOqnvSg2Pwm/ug3RqWAcD0XTb9wYlB0c7pqh8aOc8LPeFYwhVibllDU
1oVUVkpzyJrS3pJ74wAaFOlV0ilNNqaJkQ3wRMgP7w2HsqN+iSHUcQLZWJ/GN2dbdRc022R2UsuI
wQLVO9kMtT7amDjoM0ir7w0yZolwPHuQbDkV8Yoq5K0pnfC3CSKhCHIq+UL9/bvGzhdHSv5tawgX
xgka8xR2NJKJk8xlaYbBtc83Z7qvUL4XxROCMBm161YxnfG+o1Lfr/VumaYlRVC1uf6r3V1s0iNE
Asbp0a/Y5jBEcHvZP/WekLQoiLtQ7VbEj458YAG9TdwTBogHZxFkOg3NaHi03n/4IDlE/QnTM7N4
lJY2ATQKV1+aqj/JbAM2ylZtpDTyDKHpPDtXPLddl2NzbyhqPDKktClxTlkWY4YUi5G9dYG3536/
WEeUrbVL/kMq04BXh07vkAYOAzi/JBYCuk/sLzpTEvagyeJT9ow21OY2FWSeV+pRPjWyhbSxLUFo
bodZXVR7tXaOW4I5LG/dxod7JeOrtcs0JP7fas7bGHaf8uQ/fUgkLS6eyxNrgyrWQZqDkMWTBMka
p6lYKYJA0IN6s0vq96QuakPzupwbkPltjMmEiUHKEMU8CJDqtHwk+rybshJ65vAb1rS9vswgJuXB
7oy8Zz+uU9/1qpSyaqKaCe+/RnNZ+FbqB25riA6Jgm0QdiBMHB8/Gxc7C7cOhyBkC7IVrzX6quKD
gDIdKSuQZsXAQgBKqVdcVLf780hI2vfRCAlkV5omulvArdF+aTqKUHTdAKUxeZkEWHRU9wDhb/iI
LcGGvankUAoZx0kQcVBGvmDZZ5KfZ+Ke0NTmJbrulUWTylEdDcWVt8a92quQBtGoRB88DWe+Lgoq
sO4gxJYLlxYsV5YI4Gn5LPmqv4ngoMprjOR7vkwftCFLt4V/suFwBKdME2y6peuVqGipQjtZrjAn
LyxRlsrusHiNLx6VT1Z82xpUWfY+njsvkMzFuV8jZHSmLb+WRQmJQ6nEL/gxUfKf3jWJjQOR+Zfn
z9jmKdRanEuNSaRnbluTzz7VhsbMkRrJlRQzxXX521KAUcj+t07QvtGjgYB+gUw+LHoxmAV5xXDG
zipv7unYTPE/TT7esbXEkYYhKsGj7Bv63X/utEundoI1AZ8/glj5XdA3VqCyKzsMzsvQL97WlkVi
zaAFat4Zi/gZ6lKeusidgHxQJ+IQiEbG9BruVxK7LTd7MhFo/tGTcwGLToM8K/4xwbYlkeL9awtr
+WjKKUUqYGJx4a6dlrvDd6xOY1wNK2NPCstxpAYXI/Wcv2OeZXX3JzHXe5V1zH0iIkCPkeFLDviX
n5VNYBZrYKFAjtGSofedPj4mNi8i3tsTYC9kmGqBGpKPsCU9rKvCQxp1LnVSLpELS+kriicCJq7c
TyNUaSYW9ohspu/q0u/c0BeMbUIbhXDOg14AGCWGaxdmEtej3rWk3nxWDGFgB7UWMWWBewpudIhx
AjiFS/Cs9zkn/jsReXjdpyCy2trFhgJ8UAM16bq1O5ykgK+xDbs0HfVuWTRuhSvIgRdIMge9If+u
3Ks5b4Q+K0wRjVbxTDrdgXUMZ+fEMvnT/vDaDVlt1bTeFeHSaE6KO09zqOWS4Mm0SO5LALZHYb9a
jXfrFfA8Y/ZITkZCLJwtu539zn3w84rSzaasjneX7r/3/F2eWYAeLKNaIloTFogWu0dx8EZ5i2In
ezOQpp1+daJp8lsH9fRwnLdBK+y9Cttkrk/Ki5+7cwtz6ukNxCNiB/eW2oacN2MgXSG43gE1cBMa
8xomYT3Obl3FF+NelbdLgf5YMPf9k3w34FhNWb57vq0eS4V3gcIGeMkHCjQxnxZZWY7/lxNkd4e3
AhNGabu0yFtW3QHp5vuGjwbUMppsl0tdYQShfXvmgcGEO8dyGF4Le+SvwNAzeztEomUNF96QsNQs
V140gF5i32uzjJdq21j3HtK+zSOhEdSTnJ7dWFwlSS2UQ+qqu+fdM476/qmBQp6SJMqTkKhm7fuO
VQBOvBOjVbmsNQFOwseeElGYmoB01Yp2lifJj3Rki3FRNanSOJs/2e3rm/Y88Fz1hAKxeyoTSWPD
5AE5Ov1THlhhNppqNFMwyjYJEWInIH04TUCzuUet96O1BSZHnzbUUNRdosn5Pz6i7rLvaSDD5Z0v
aClTxnoj8CY73A5xNaYf4weTDAua+uJnmLpi4u0ZO7sw6NrPA9vD8XjyR2xmJlwCaykXzYkRcmTu
55/L4GRfcrvmFGTp0FtxOWgtR0GEz6ktkGS0cEm0CcipIRwDazHO9iwWFv+KY9K/NHNUUpROAkN5
LMa0EArZIchvFClz6vtjG1yiKXoZRW1YYOs+vOYyiRNQOYeUXQYB5oXlun5RuT1mE1FZ6N/gdtTX
TSjgDuupTfwwN8UN6VUrNa1BQGRoEseL5Ou9EC+5nZhbOKEBk3jgJfP+GX7WiXcM1qam4w70YIL5
NEPGjdouodIjmG9lo4eMzGcErbAP8Pfe+sElxRXz3gwK8kesBX7FChErFY6TxJ1BQueKz0MMeWV6
p+GbNweIfXwGBV6OtAtCn62ndjjUTcdGpvdyKA5uv0+OgsxG5rZp9gJSJCy6QCqTGTjilAqKtHPd
2QY9lQd4tIGnZW3DwQ1YgyNt4/c+IeI41Rncj81G5EbRyNaCvt1uM+NiSh0YDZXntMFlqcbsAWpB
nh48t1r+P/A0UL3kz3+YwlR5Q+q/wDAlt3BBbm6jfhAp47xZOaRL2Chbbm1MyF213CVJT2aY+TPM
FDHt2vBrpun29QP9FTKwsVrHGJrAIj9YKFdvM8xCNwuArvrYszNuG2UZNxSJAHF8fcPx3xZlNyb8
UgorPu29tggxl2RSiHRlOg5mlo/HsyoslezO61Cc6gyaeUd7EXXboH1cxaLVy9Cgww37KQQIYO32
+IgOC5VyErqQBWO2YAtW5Z3/eU1zOTsnzsxWI6O4WNJKBSh0ROdWLbSC9E2p3rFsIq+L0vWf0cix
C3wpUPTAUzA9DCdpI7yVlbTN3PfnWUWEEtloog6S3re5JCzPqkJkvCmAk62cbs5PQnBCn7mmJi7e
31onPfngV1aS/wiKUgC1nqMV83Ppk7RaCJulx5mDpk/dxYzJDHKEHshPq6aCsRsfcud+7QFJN/8n
fS4JDLRM9OwLSCigtuttvzx9S+2EBUmFTETs6Kl5t6+kry5JQxY5u9evY3HBtMhnRHMuX+TrMLC2
vmqy3ayRC8GGvfAvOj5bBVdsWQgxBaGwAgWsmWQvSYNUgfa9kiAoz4ojmE+iazodqCKCmRILW5pw
0uqfs3unEUFzMC2bXYXr+DAm6WXcUDY50yohan0heJzrcUW9fXXD0/XfWy2LBRpa2yqa3OPnqBQ+
ljCkUxCotHbb3m1mS58yPbU+RdycXWSmb1hQgmbSmcQwjBXN2iZ+j6YFOd/GYOqpx5i9WIceI8+i
7ZotuXMSWUZbGeSy58Doyah+PfoyzZoSq9l7jwrBY5Mj6oSgOcmgFg/0mdfr/MBiSLLsA1oiOMBY
Dk+sIVL+VCguc6qooXojE8+nZgKkotS+SJgjAwsDsIzBvXQnMsQEqKAgvQBkNmeNDS453kF0XWYe
aMfEF3Xo8I20lbA7KEFBI/x4MyveR6lKYKJVaT93VsENDmNAbYsAFxqUibzcNbRK4a5F/ta/8pcB
JZJ0urt5/TETy6T4OMbsAsR0yaf96PGUQOy6jg5qB4yMiMV73gmXow0Bu3/tLWvIZOd1fp33OkNk
By+QbHvlCHzEnml/XqUZOkXaajDYelR4StMnER5+UytahoKMvguvGglRx7wObq6IWxopj5FIoYqW
bggcJxABRTWMnxqnEMROqkp8rEaEFaxQe9vVd8eLZwsrvbJ/BRTSQCyD0gvF+t51F6matZvhBPsq
zEEembw2VyzR6KY0nYxdKhw97KxsjRHZW+UZEYQKISXMy02jnrFblBFz7jXUbYc0MFFA+f4lFVBH
samTCuMuec6I58LruhsF8l8jaksOevlCKyIdFYjI88SnfuO+Gkov/uPjAcbx0cUNQ6lF0AiTzodB
kJGrrdQc4F4I5kPPkXGnG4jvPmJtin7MVLqikEpeZC31zioc5Dwkx9qKnl92/DPquB4/6XVQ1rXH
xTKR7OhEO8pJJUm8gIJJMqNO7TxbChHEgH/8i/FWT4IEF6d34A5TCyCi668rG0I3He2NqY9LKG4d
BjNC/ns1Ebq0MAhu96L9NLrLb9PAGg1miBwIof+W18jiwnfBiHFqCldbF9L3A6BzlVBjB7wV+rds
2aVWlEV36VGKT4BZhouw/dT42hetkBeNoY+OXVHmaXfwtSGPfwYw2qf70XQgYFj2447DEGq5amyl
BOmD6RrALdGmnlSqwI1g1jwNO2Y5h7uvcXZT8H5vjxF8KUrhWuXeW0K92HZXReSGyT4nvcV4W2g8
f9pp/Fem+4RiEQziyESTLwnqb8anQCP5hk+S43q9YEH1b/qwz8sobvB+I8//rmUyDQUNzzoltvMg
BQlSM4gvotgVWlonJd1Yarodwk1QY2IAum66icrfr4USvbr/tE+XekAkJx8c9LXcRQvBS+BgHKtn
P2Pnm8e26eFDGi6bxvPGzCiWQA4sN5vth1L62z3pwt5+H7Iz6glBP6/oPwaVlMtNam6mFVnAVRSX
VVPbaD4Aj4HiY1tqQgRBmZM9neT6yFi0/gFJ3dik7fZR+EeiFmj60nKsxApqLH80HE/CUuuhwG6B
kDla1YkwanKYsDgS4PXpRX5BBRfV2S776aglqgLQobd+xSzl3fZ3neXp67ftKDUWZF+TPVXEGUg6
7XdryOtGdffug+AJau1fJuwgMntlYJa1MJU/gCrnXCjv4o3YwjLf5e2qi+TX1bXwSPw8hvh1Betu
5RLtABc2dX2dG7JKCQpZcvrDLvSNcRzXpWzQJoMWHASIi85XOGFkKmnDryTgxXR5nP60jBzG02Rt
9G+K0JgCfhqlBJjMRh9TnFLSeUHo1Zp3dQjAW5DjR8xKQlFEMM4mt0mgyU8onHSo4S1cehdHDjK0
l5fgNhNq1Z+jaBW/TYpMT4YIsBNmh3sI+G15BkSoO67Tfzz4GRStQTmCKo4PwCva+VvL8WNAd6Nz
xV3qbWunfMzKW8NRIoJKYgltTIn78wPI0sVzavhrGo54tVCdQjKMqGEjsIIU1qlztcqp1uKHUtkE
/+n75L13Ya96fEhts6I6aoJ9nGIHji+25+CQDt0I5R8BDz3rzjmG2zOIibWFaWH6iOGRXrj3oN1i
l+XxJcSVM3slZFGNSaGCkkFL7DQ5Ptmqep8vBcQr6H4bPsM5cjBDkD19htamPJ1rvUa5Wzn1noZx
24T0/sYplpcLYYWLLmTCig/lj8zIAD0DV/A0iwEl6fakli8jdr12Rj1YZ3Xo2Xp00sDjqnV19o3+
qlz2oShgJsF6TUHa4cyUIneLS4dcrQeEijcfCk94XNIft7gNYL3DmHRknIEPsyOF9sPtD6mbAy6M
+iM/ZSVLrmMOaQ1Cm5vfc0EMQAC+w20WM9xrpE8syB+Q668MJVPjeXjM2DrsvYcSO7zfFzZAk9oB
NbpVYrEFc59rV+4gIjObY0G7ukHUVBu2zalTGDORyUJ3OSESTieWp48cVh37br1Cf97h4sieKH4A
ntLnp2+8IclNZ61qxqi3mYZoXgpb+Hduy27HsJZzLOrQgscWxoAQrQqhQvJob3cTunVO8a6vfz08
9lOojV+ZE1mw2kkyz3rthlJ1vqIykuA0OYyF2S4ccZsZXV12jfCIhqQKaDfxHNJXnXXZK5nwYMRR
+qFQsvleN04OhLl/zdqMlPxihETvKJWtih3XoBsMDQnsl+zxx7onQiaVBIbvEcZr59rbea4ufrqH
oTY8qAv1ZhQMfTrLfHOGoKrqCPfP2YpKcIk0yYxVOuu2QAnkPycZCCrK+Novda8DgpTHs1Hs92DD
qLlgMgQcVAjB5znWz1MKO/PCi2trJJEQ+FdHFm/7Pd9ls3CYGc0oa1KRtk7qCpOycRmoLsfLtgvR
QTUHvZ2mRIedYAREVJRPrm+/ofVlL1GBRvfgh3EBMNnYVCK+cBxYmVP8FbvjNR/LyZQ3BfeVOf4s
E5JfgqfML5KzVvO+FscrHMOHB3lCSYyrF+/YRDk0ByNQmdG20YL0HbOXXsNeMikC17G5nVNB4rVa
IQ5lwJhI8FrDYXz6V5n2stjNrR5uLOiX9u3T8LIE3RxapE914rk+gy1+/1kAttcrfyvmKsE+dfoN
5FfDRnvzMP+GYPp1W+mDp36yYUHGzQm5F8cmI/pqtH/HFjvAUWiEaqPvkdizS2E4kWHLiLawYB0l
rMK60TcbPphhQz4DNSvpfNh60ldtVMq6bYx1Dl8excrtmXQBzVgcLB6bGxs0xvgf8RKOOZ1tNXDW
NIrIHT5hK9msj2Ma5olXU8Ezj5C//1TPSCM+U7ao7hnJL6UXKCU3QOJCAJDjmiE3ANgsZ5SrupoA
V5VioW6Q9rZqFSNcEi98AxjGGMGmc08VwFXaDa/eXB4cbo5zlodLSuba0t/maSXKuUn4rJMHkfwJ
+R+OhpgW2o+ox043Fud4Aed9mXbJ7eW9qaqJz/oP1yP+PT2QLItHTN9elsT6fCnSJXbzHk+XQWlp
9/F1Cq61dQokSMJofPSArOT9GZub5MKqXNm7dFJVo1MDpKn5fVhOIrK4TyymCgSsmtatOEOpGpAi
Az5TMnCzwpBLZm0jBX/Y8M0FUz3dHy8QiPTY8HLlv1sOtDVpNHoOGCULqViMdjw1B+IAQLyPZC5K
+x/cWHiqmsgVkb55BCIoVXe2H7Uza2RlsHSq1DsfhCnVHze7TkQQv1CHHtcArz0aX/My9I/bv1uM
rvImNLQXiesEoln4DPXUXP4CoOsZpOa3ClNd/oHYwQf6a2SdbbkrNmpoisurc4CoyrrznpQjQPa4
N3shzMzz6b6W9sgbxAEzTkfAt3wa/p3p83aNOzNK3nTBwUBPd6b3dwHX1Ss9Eh2m8PvFx12leSbX
id4Dw5kyr6xTiy5b+VY9zARwfFdTeSnLbhh+8q58xG2u/J3C6ixzVb53vJXP3uPuLMXkyap1pLib
xkycQQXedjEdyEX4Hp/SDkx7Y5nnfbPrnBhx6Szle2ydhT21iEjSn6ngR43W267fwIsJdSo2UqK0
NfaVyVHUQ+JbqjOJZYN35XQjRHdaOTxLE4WxwDHDFgYy+ZxbpV45Ar93+9Ol3I6LLayATIw+mr28
hcTyWUMhNTmmAyOhRL+d7cXuOjPr00hnA3+ww34y3+5wgH+V7GW5a1I8AP4hrqu0rSSZguF+hzFR
dOcifHImFlg6Ki/5xDOnXJjqt0JDkDJ1kehNeB8i4CBZRZG9cyCKxUTF5zstH420YmpA6d9W4uIT
M5RNC04qltYSPrdYv/yLp9y1lZs2E0O511uWedmLQ63Q9utS9XDiv/CdagmQnh/a5z5MNtWnGeAH
kWa3Y6bKRekCgFLlWXS3U6KW0oJLtShQUPGuNBaUXQUHmp0NOwcB5/wM7AcHzKGJZBK8gWXR8miE
/v7GYmu3sKPy7PBGC/LDoov2TMcxjbOzwtIpDwaIiolDam/gZJOdzlY3t+QsGBN9lqKD+m4DnL7e
053w7HDzOFb3unmVuYRHowhyyaowXfkt8P9DEBN64XaakTXzjgpfzdZ4/M4vLUDTxMGvTw2M525k
7WCzPKapDG48e9etPZQdZ7OOMcW0t+xxJaYMczqAFwdFQ21QIddsKCw/Lo7VpoFlS5oVdWhwYaRU
67y55eMHZidxeWbbiPcL4QPN3gzX5t7E31ulzS2XuxoKcezFR1cgHe+KGZbekgXZjijzooamLcxU
1B3sD7SAUa55CXrpYD573tsEfUbugavQLhNL1vffenSj9slmTSxS+AJr+g0rVrf3itbwe29vFk8S
eVWyMNx75mFET5+v5NozN/eByUkCbIIbbX9um+veGrU5RQkPojdcOoV+NKZfTT6BGL3gEZ8G8L18
O+cxPYkoOkHTV/SzNHCLSgMb6EjX6UV/g1QFtj8l9L+Ah5Gys0Z4WDm7WykBomEpu1Nruhsp3ccK
uHaJCNdnLdDHToKYqFfvbRl4aMgJIFinS4jJwt66O5RZj4LFtez8+DtPNq4NYRqYAo10Kur185ZO
SMT2tPznEyfmdQzydbfpwE08q+pfEfq2EvfZa7gKiz8F546Rqq0FnbtjGYwE2tSXcSJy0yHee6v9
2XKXi1cCm15aS8gUI0BUjYS7jWN/6vzCERVBxYZGExiZvpqnvjJWZ4II9KOMNU4AgfNRwVRwde75
cv1UWJ5OJ7UjWMPogznSmSwJt4NHsNuJx27QEHtjRyqRgxb5LHJuOU6JONUwBxJvgSvMz7mApMBM
vKbHtsZuebrx+dquL/UTuoIBVCxEKLHstrctEK8N3FQ7piTNy1+q3oYq+EL70T0V9wuqPilNBFZk
k7erQ609HXiyg7vqvVaFiYwXB3RHMSF9p9sI/gnyZkxqShEPdTL8gnOEE9Vrv4pZN7HkWb9GwKTD
VNf8riNgWAS/ICbfnM1pTtDH8gzWLMWGQsIo+ZCgKhzbLxNKVFtATFocjfnyhhIWbzlz7Y1cddet
7WiemXlkI/zclr3+nmZVmuXkvDYa7E1k09irOEFK+TBOlAExlbNeTBFxsbjnDgMvimoqZwivbbT1
n9TEjUz0LBhj8We6BhsWM8nWcDj+T1rg6j+1VqZ/us1VgFg2F651Yd00dA+t41zpoeUemiU/ei66
fiNwW4PEgGEjSoZ96wE/VnDtXImZpWQ/39a+ZkOboVcu7DnjqWdw6dyRFpphvRr32niX8R76Uv4/
Jv6wsLIq7sdiG5KAnJcKE4RWy8ntzm+EBRwjt3gIY4vE8K0+jeAOWt32jRs28SfyD3GW4nx0fR2e
NVsiDnXtEZvaVyWbowsZ7rUsUgZz9yCcQyxsYXTplkKWGldfSgf3eZdzBPxJ8GkIVV+6MIQKrIPQ
PZxXkIAtGinpgr7YFLZ8LG07E/XNupU7iFw95GTIdIhodW1NpjBNjYfxXa8U8XvZ30PH2MycGNQH
0AknIWRj7MBhGYqaWX+qYzJJIGKPKc2N9ko+OPgNX4Yi3TfMypYQ7UQHjxgfh0UaclzBrn2q8Gil
OrfKOQTn55rVh9+M1U1vyyDHlDn7L2hGJsh34u56U6rDQbqdqzwv3ONf4T11y8p45Y01ExJG61r/
QuQcZb9/b8pmYFg4FX4mFzElzmbPs7UwMZIy6r6OHd3lx+C/UxDWBWqGLUwFmW8Sd1kP+Uo36XHu
KHtbxboWhKm1s1Ru0XT9PgqTnP9dAjHtKtQfQVFn3UxhIHqTEtzEcK6yz6gP0G0xRJYr/xY/719B
F6kchSzyGKxMPre7waZCR+rLJE91bKQJDKJwiYpFnqLJcW74tVkzsaCzjDjYjFXG58QFtpI3uOMD
xGVrqPTzLOEKw/E3ZkMuJfX0GS/G0zOjHaEoRUpnMOeRpF4NR9CJlNv4pvdrzOkrE/x3P0bcZXk/
480x+3jHk/ZzjBrcx7z2tobhkfabhpJ3Q83lvmuJKN5bcs7yKEHS+Ee2Y1P0RpRJlF+obCwnEQ9m
+CO/zw7JlmtMRXG33JTG6vwDTPXa9qr7MGEiyQwNJZCNzC1Jue19SiafK8hZs0HzfPbr947K+/bU
ft2GvDCpS/7EHA+8Y3hlHBd+rG6+ZwwYjZRFKs0wa9tKhHVJwieUc9yaq1bAwHQ44GtXi+NECpJW
ViTZSwzqaIswp0gEhqFjZAqHxKqAtIPchdwfdc7AqM+whEkCVQyLo/5xeNgwxIbayL0PVLiDbycL
kQh3CE+4EryQIkaSOAV1rDw4hWsWEsKq7TDq90KN2mPY5bLMW8YSBV1/peVDv0Et2tT0K3AKgjT/
CqyYr/Nwc0Zq/1Cgf5KxSYXJyYzsxlXRfPzvSxWYn4pOqvZJLwEpXaDHN0an1HkpiBoDt2qbexHV
HQtcYPxz2AnFZ1900GcVPaMdtMJcDndKkiZm+3hqWZICxzCU3+qMTUP8L3PBMvpV9dXWN/9ip/Yd
9x5XaGyAWjDOMbyTiWpODwpqFAiJn7vrThuwJYmeicafyabjTp89I+IekwOJZ253eunKDY43NR9N
VjHR4Iyaea9vvgwh7gSH1zS65nVzRS3W7oatUDsJWo/fwIMwOGxsk9Ddrr3SxGk1u+WO8cdKJ91m
kdfBbRu5mvqJsAQfbnISwMQVBUJ/LNMGqf7iykOPRn2oDu+ka1HeXJu00symdu9qP+JkdzuJYwEt
wR6gV41FGNdD2KlotT5nOCA8/pqr55Y7mFVY4Y2Dq4SX8EJpGa7Obltd7psF2klz0bnw6OR+wkWW
LJN71dcQod8/Qan6ZQh84XIk6pwzgGsLTYoL9f/LqrBdvCkUpkoxyr0lMrQ+bNGV5lU+cP83AWee
7z2uBGGjV9Q8vWf4Kc6eiD3GyJezLVpjmb5jGx/o8BK1f3dcFTibfNRMTfXOb2OGz6KOizNOsAdF
GBAV2BDtvg2Q3ouRARxF1w4HtO8NYVEHEY6/ztUKykHoDXWZ5MktLfgZli2FpMLaWllzD57F3s0X
UMLpgrqjiwNxApOAXcINEbRE33DCPazaWhWGbhxjR2WhKV9kc+wawzAOvpEKVTVVM/AI6iMAlIGs
W3TEChMjPPoSeEN0AGy+bQsB0jtIHf3nhpTj0JLnnoU0W0oI3MWJQ1akUKTqqXafS4LIi96cTrg1
iAZklT0c8TBlMPmrXLPcdg90mW/qPYMgZFHGdW2b1RUAXpKVoncZxggCzPvy+BjGDDuiemNp9oK8
ehL5RS1ikRMwaDIRFrmGln7QfyzniyzEC80MqZ+NbAAJkgxSergODxWaUBAmqGlmm1KzIyr25Pjc
jJGD7qU7qx/XZkA/IRVc9nOnlhnz/QBNKIlGWaj77mjXpmvgmNUi7AAWdunicbKlj7GJbmM5MpAJ
YcJCJZBssdnWuG4h91uCn+MeEWLZmji3RJarWfqo4THrx4dQ4QqJLRGrWapLX88L46R8JV6Tr9GP
AE98kdtuqJxLp7hFE7QibrK3YPkQ6AsmF7FCvTMv1G0GOOjlF2qfSjzp6O3UusCXDq4c+prYrzFp
Abk7hAmwTDHMtoJR7jL0qC7jg3LO1fMPZiUK9XDWE/pfH7sFmfqWXrLVtWrqBucqugngYZDsLhQw
2O44yJNVZ8xwNT6z+FwaRVySBmJODPt53OHlgz2hlYTzYaQMsvenOZBmYB98P89MSvpwfSPFtdxH
X2+j10pIMgYzAt/RA+9eLEHY0Jwy3toN6kgUlP6VgAjMzvfaCEs56xQW+vDCrdWzAVnT9IBSUsMA
+MpUOlnZQCBrjpwxbUetOwKyvZsbdeqCJ8Qu3VCv3bl/Gz60YejaS8PbdeJjo2cLdfBTqEgsRI0Z
l721gWW1dDg06jTKmiFVtjuI3uZnRnuzLGf14M8pD0nLI5SQzBT8uB4EuvMU6BHxluamiwcw2f6U
QUvyvjOnA54GjHuKPukN+xXABduTEXrNl7Y9yJ24bz5IusyyP9H1dvhtqQBovQcWQISFdWRKUNgQ
INsX/5dcCP5fzbLMJsAdWEiVJvBmTJE/LjVwK5i5lQ6tVFUbJA5BMYPANnK0LHIoUcHnZGZaBRHs
AguxEvozkVwTLOIjSAJT+ItHcTLOAfedUfZBf6DXZCxOPS/aCkyTyE7zl4cPp0SbSMz0gi6XbrOY
0NY4kZ9oWKXyTkGUxBZQ6Ba88uZSRaK0mZ/RizKd4wC8RDhk3vXIGKH2fYBRklcYHaCPQJZ9/xmf
w0qjkO+ejUpMU3LWV7y4YN3moSiLk2nhkK22Mpc+9dDOgvBsVBC4kTt1Q1DyeWePqGE+mBjdqedq
k2Kyhq39A7OM9pOmca/ZwBhFENaqCvUtEKUfWU8a95Dfk09Ipjpy7E+K3nk3mhckxfVwBZ56PWhv
kIbpupT6a+ZZU/kTH00mGVOo22uBS7jI1DNRmEWGsDegnFL+le+9pKo3R59eagCitQB2+o5ajvSG
rUI/vZU3NnfRc9m0IyZI452DlypxfrSTLuoOYk9kUUp9uGX990pm008Dk365TBzTfjDEp3x9Z7tY
iRS8bvjJMeVa79e8R/iyyCw1rCH+/K+1dNCSJUOIkVR6LdGTOWjrxttAsEaeIfzN2Y33TTHxFRIa
PXAebiIHJG0qClJ7QLZQ2e19W7Kl0nDHIP3fb+ENIjizW7AJligZN6XEJdvgixcqcHAQZZkpND8M
2vC8vJRvqTxXNrQ6MJvWZTz8fPQ6yXoE1K0/+PL2L2G5INogL9Tbw9AdpdIi3EVmV98a+ks812UA
VANkD6/1udQ9W9oy30x3ocxZRZqE3CFCYNm+3SycrjGqzQpXew68dcykm056ddQAybmfSwx1GHyN
IknwBxI88cE+1/hEum2VtA5snnq8RtrCW2Dq9RKsISFpDgeanQwh4oq68nZDUcUq2a5nXujJrPxj
Xw4K81N/2kHIdNhx7TI6WJeGhjGK29zHHBQG80CSkkv93hrjj6SSM4g1+885gFaOVFx71FfA8JXN
EXw4h8Mdm83C23GphAMK37vGzO7q8U1r4lMJDHDEEmYBg2a8XqNtTY8/qlzNLZ2/3hQzrxKT7QOB
j/9aNXwGNyA66dgqw4cuAY5nxD1SMdhPcaROxVXAuNgaU5OuRvOSwTY2rrBW3wCgfEDdrAsBOtYv
+5LP0UJwBQNFNP4EqjtVM8+u183iqR4hjjObdg/P1kzQX4F6odH9SHH0+RX1U60x3m9SrjEaH7Gb
hGQYGKqjb9kxSWU8K/VsOaAPQtuo5nTZA1DinlwDVfQGlpTxL1DLz3oGCU3ptoGVvHMmdpsMOij4
0P1Ui3v1OlNA7fAtFyjm0c0jzE1rz3HlL/o/00Z+uGmYtrhL7taKwe4EQcim3JtZtuivUREtDNML
zuEtxuLMDK7n+L3blNfnj2i9jdyMSepzU1/JOjceqAwxzdcK7X24boVaXoe4LrYwVbSq3RRZHoMg
WQSKZDnMO9WRIKlBmKSeSVHZMUG7ZpjukE2cQoLnSFzamSmHC9OwmtlVafFMLsmhmTlE1aXypJZQ
Z+ZYIvTdWjdP0i7V6nGMD9ZMADKgLcozGiaO1/2+mBPzKBSv1E5J48rW69fOouDm2U8MJRcKayK8
GcjJlUqPpbrD6PPMD6vF5DrGT6V80iaKLbDQQ+AZsVAR1wOwaWEu3MWHHhYcj4pflmfNCVWGi5Md
ZAUitX648qeCUjkwMmhJsEUxPn3GY3d5j96CzcmybvTxiYBxfxXsw1b1aDfnOjLddh1Uy0C7kwnu
lo5iH+GlINbLcGJmLNVQ76BEHXv1SWj1YaouCDIJAqTnn7GkIKYZF/u51nXlzg2VhRyBnpX6MNvg
Uq58iIALe5vhWwC/CUZnmiehb+BKDIovaDdVsa20BrPbT4K0W/amZVhYpuL1WHuwYeFoUKhY1lly
fOYi3Ob119+ha5NNftBY6B5GzD6jtDEIrBYMRdKW+mje8LvxZ6xYOFkewRKTIP36piGZgqeGSkZf
3UKYmlvKk5qPDON+Auu6D9EbLMPQp0lXHjL/TLPJf0wY6nmxT+16YfXaeyB5fl4pSch00stgnnAY
hHN7Rqbew0+mDEVJLSV6l3imRelPRrrEgoV8ftlT8vMeysx7mJr9Q8DwHk1z0oV36IrWJ9Wg6eDm
VnnGQy5eFLbwWS6SUoqa+XEKPdSWkSHvClruSgJrXj2AbKTe9PEJL4lZjRPaLbKxIxowQx9nTS0T
EeNpQ1M69mI2zVa2qmo4ClHJ0PC5CRV1fOhlm1XKzEC/HSiONjR2jJ3rqEpnhH74qs+n3f17haja
vN+ECOzDLWg+GLFcamnnXEjuVVCTNbttNyZ5wbGhj3EBdzeRDHbzpqqPrfqwJDXt9LJABhQfuVEK
SZPhis87GmhFwnWyxlPciocLpHEsYbsqTgfjNx3bg821npQbViSojECED3HOMTCXfi72eK65NIzZ
tTq9eHDChmqdVKAl8IVYFy0Nz/JSOT9ZVN0Z5nUr0kS4x2jATEC51Z5RyuShxzCuQI3HZz7IbGam
xg9K1i8s+I9gSniaUtHTAKdoK/+9V5V2VPxQsf9rB8nhFIO1/JeW2cJjlHLqDqnkaMfmm/qzLezc
AG39ddToPiMWhESHFpbzGgtN3sPfXMepPeD2d5SeKaWewf/q1Rm9m+3fi8olZ/Gs9cwl215jWo1I
MFA2HHIZJWie1XfbpOENxLrxsIHUnitJDk0JXH6Fqce+3tGwQBuAN7LEKXgCo9WPbteMFBmzmJwT
0qqMGRT/Ww1UbS+dAlZUVFhAwQcfPLCoH+GLPVIiy3Tard1PYIEjyZn2lVNWjfmJT85zVD2BhEsm
0pvZ4a2T0HESCktzkYbscTP5HCkquq7fwxhu4EAulrym0H+ozfDAYMk3F8duVGklY05in3RjMpbs
+UapbGDCVkpuAjR6BMOW5UhMa8dxscuW3Qb4uZbPDoNqveMZ7Kx2rsgsc2aEq1pEKc5q0tFNXH/P
TbYqG3lzNFXL1CsGaeoNSc065bO2xrgf+VYJdtdp+G7+BAMF8LWujGfr5IXI+f092aHa9JDlWTxz
ihtMJBnbYjZ+t0SVzrDxeKap6t0VeTXgMXTWzRq/D6ixJZ+8xHQRScVZ/qwgE94+EigRncxJMOSn
HYTi84ZXD/xKMcG7B8KFpbh0am/0oVDpg5lQHZeFVQW1QPgSDYcz//yo6pNqmHjQ1YYIFYrRykIw
xCdrLYHrV9J7rBgd4HlNrNEqQ597m+T4831Jvs3Og7Rkk30afB6BmEih/6pBrwHqUzFiz5+7Vmbp
2n2xA3rGIWZUWUyFZGi12kyEDMRRfYj0cQJobmODkCyJ06l3GMRCcKfTrlLmcCaIWr3pNJTGSjsh
VtsFcG6GXP4/FJxar8bPIeP4LHx3GxrWBSoWhVZJ4cCRF2lobsz9njJp6jQAS8+9SP93l+LgzSA8
Dz8P/wsH/gAm7/EZKPOLaQyNAmzZYhfVVyoa04GFFh+A2DWa5cAMtIU8KFSGVaN2he6qRZ7i3mR5
bSumXmPrOzVU33nJoO6kJp2oUwENbLBEATiKN95H9OIGoZMO2tHa3cV+g4tM2ZvqEAj9g2dvnehA
PcmYnkB5+/ES+tOPBJMivEmEF1+JrErslYbxHoAI/g+ySMyPZtwHIODmtvRKPgUay05TCdQYchwV
w+WmMfSjPnBH8UWBj7euDFPHf3rIDsko/yvIyrs7nhUbt0ptsKoZ+1L9if3QxlBmllDg88n3+Btf
jRg4r6+9Ym15xP5N3+SumrHTg3nLN0j1lUv9bJELi9iCUMfoSfu2ZMfzaD8ZvJDzcU3+U2yzip40
5l2kqpANQDw6ZsmxdNdub/A/n2Al4HrRhKV2ZrtI2te9e1j75e2oxV7nfMWV8iQqRMGfx1slL9jr
bO0IF9vqw2i+ZiXmXRzaOCeb7+LbBcWbDvzLgCcNkVhVGlG4r70Rrh8Rh1+Zt3Bfclrlu6VodLPF
dMvqeQ6TTwVKosrrsy3wYwNINa+uHWRi0rasRb3NAOiSYGk2MiE+KpXO9W5yof24D5VdBnqgOg/l
/tyHo5IwqwKYfEsEDxnFss2324iWSfyJNRxiuIHbKSKKR7+jcwvDOmj+LxLENvIRUPaED1iP6BiR
tlc9EqrlfvsOQsJeNaK5Fcu6yVKSvKU2s3/zsDFSl6fKDZ0hgkhbHdYxCGj0+dcJuytztaWM8/b6
3MScj95QnreThKX2v3GQu8mmYHLZcdYxVl+RB4UXwcUKvP86laP0IscKfbK0f8hrIbqNcs+0CrLu
TIx3gmEfVI0bDnS/v15pnhhk63S1gRaPhpBbE+rWK8Jt53H+sJKxCClsjtynZnvyAwUlXubKKvb+
mBaE9w1NsIstY5Tr2pbEwaAGR9TmbhcNkSWGQKsa6wYUi8Yb5pIOiC6CSyd9Xi2JLl0ClG/E2ktN
64WpKg0L3TpHy2IUw2dzAjpDk4sQQovwDQx0oDpKcj5vVPJDfq1AqKfQix0dpA2o41NdXnx+vQtS
FzTV75ERnjLEjDmj6+Rul8aWCt0GESoNWVP6PMqeUieeMKG6xZ48m4Lft4qnIlz32ETeRiAuoNKd
TtoO1OpmOD+FEpuT2C2UKNQdq5hYt2H0tZEoAhECVFfY72zJQUe4eUYW3ctDmHp18p0hAUFicWNx
pmCHHYckO8VbL+sezHGZ+vEi0QZVXezTp1ec7o+mq3FPR1QXciJhfvxEkHRk3iVd3Qw+G1OzXUbw
QrqEVm0Vn9aUgua2QQCV2u8pWBXvGwbjRMi7ftU9EaJvCCwIKGUzODF0h+retWE3Ivbu1bLOsLfv
Xv7Lsl6U3Hwruaiy2AXIgKlX3iK+qvLqoC55AhQmaA5zTU1YaeSw40+y5MAqnnL2b3IUUzifMvDH
TXbUDb6YdkErShk/LZ4JNftzUsqxXrRisvU8BZG/2hMWnj1AL78jQcZS/wW0RJ20lC+X3wkEVAUf
5IELYMadBuPRGop9pdJG7+BqwTn3C6EzIQlz54mZKNhSKFm0IDm6WMyp067GI0+/NPKHl9L/VkLv
e3yi+rMU2zgLNN/FHr7XEG5EiR5DR5Ua4cFD9zYqWSoEPptY6j9aq0Jny/OCU00mioZ1A0+5pmuk
y2lDHmSyhAOZjw8fKo4hWno5719Ghvdu9+S0ig5F7Dl0HsGC2wqC1lilBe7tDFzIExDEYoDHgdOl
7no6KyQDIrOTxUVlbq4N93FYZ5zFOQbNWHiqdYR5e+ChxgsaC80xrGMdBX59Xw6ccmzFaX9mOs/1
upd8wDxxiYWXtrWhi0hSmJoro+6UzZ0r9OIvLQ5Zx8oPLcdvsNj3csCkw/l83q+E+F/igS0gTtF0
xkt1Du8T/3+M0cRQFGZz2/I25tbw6uKOnIhXkpG3PNLH7wpzNn441p/nfdEpF6EU2m6GgLC9crEk
pYJOWjEPo+OGpVMGXtkJd+HMx1V4dlGBkjAnBKJ/lYa/DWIuSa4CtwUOZgd7ed7wHh72UZ9FzmgS
doCj4a/CJSeW8tkRUikR8V1g6v45Htn4oM3TKK7YlPIGgOkqXbMTTJk0L5yb5zA0qhb5iVbDk82I
+J88vQphhc//aqxdDJ5ICIJw9fFPrHRG0Xpdk+DlIQ/kDAj/DAI55b7MXYF6tXVjHzKVvgHBDLqt
eado3hkqMnbD1E45Y5jPqlt8wwA2MsWfuxf/kogg5aizwGPrmWZrtLjKprMSE4aWmtTi61MjKeul
Dhq5y5E3yRUIZv1J0g9SE1TXvPqu7UQklGfUYeZIfz54e/FpFaAAFSxr+SBYH6pO9RzRb6NwuLTJ
tkb9TCRWmiih8hIuo8MB+rJ0gus99KEven/NEE7ykvjz7iVvd3BDYU+1ZyiP4dbxXQgLvlg4qrNx
wcjt4Q/QW1RxDxpimk3caG+Z5s7WXj6UXh+sH9O3OXrHz2IG50cVu3nXYe6L31HXEiPEZA45Igjd
e/G5HhWmMf3oekRzTK6O/iVBoMWdkWRQeGnIczdmEjK0iOwdWk53aRrA2q42boPCLVi7q87CoiUA
+ywc/69mbMqnHwQQKg2OP1cZE4iz47q3DvL3u/lyyvwajyi42F/4bZtE31R4gIXx75JxQ8Cjs85M
1egc/3Aj/PDwnrX/GD+QWv79ePAVrJW1Mu+NTn4aAgfQ4Ooh9vn7B8seMVrvLGrMRaDdifohKaq5
MCAH0Jfwo//om5spzyWeNp1LLn+zPCN5RvE+Oi40DQvN9ywpE5joYU2bnJESWXcL3DVYMS8doWza
OHQs91aog5NncJ3N9HQ6YFJJoB6HWZeDV4nHbWTFTQ/hkBn2tgNXBgtpuXUQwMwGe9C4dG2L7tRe
KPbVrMHFKUiFdf5XvBB4oTrTzN3uocjpXRYXInQy0DHmXuRWY+60Cpy79FYqLYMfgu+zvAZRwvcu
JcxetJ2N7765SCAEpb0NROKkPY9DIaNQuoWdIXaT6z5odti8l5jxKYvtjP6Z+JYizVT4kQBpLw05
3qDimePsHXv00CKan1TpvpbZtjuVEMwoiuBwzFTTYLfcR3RhoAt0mmqrEhnjamLRDfJb23r3TOSv
IW6+RGIiUVJWl7h/1Kc3o0gwR9tZf8ERS77C2oWPDiCUDOUtTG1JQIuhWFuHUQosR5gWHBnELuG5
mieH3NPetUx9uLzUvwfM9tSe/S3xR7A8xmioV0we+4gZqIsFYwybqQMg83YaeDgml61QEs4ZlHDM
EQuJvOZmjeCV+5jjGsx9xqXxqC2Dt2kg1zc56SJ820gkaPQNP7A06j/0LUwKrBguteFYjuv1JC5p
2KjAa8+P0FnJ13kdJJ0ZG6HmxobIrLNWzRclWM1nRh+sOmHlP3asoBQ3nvgp0i+c1/Fx4Q26z7X8
trc+hmjVwBAOrixV5ts+jVHpqH6jdIU3RxYlZNOgIhuPSV9hS/rkHa0IMdJj553KzMvYq4UdHo6R
BvDBrZ7YpRznRbNdQKt+mo65xnbtMKauxrxcVfzZjf8TKcW3UakSp6m5kv65ev3VXJn2gCLO86bQ
a+7Z/V3ti+BEW3vBlR9VUKZw1nNMogwOmw8QiIyqfVovyQ1O9XTDVzez56X/UslgG0lySJ6pb1PQ
LvKL7ARd6/PPjhovBV3LRGE+NiygnQXFMYz27XWv8ZbSDmKEdsrVL3rrsCBgZ+O3eN0UhoR+75ax
xJSjRG6c3dijCCVRVjdHvtZkjITmiAtukWtvTFX/TSuoAWHMgz1U7r6PnEiX3B82+v/ef73Botgf
5eDn9aXEQL88aMY9BIopNDUddz8/jYSCHmwYVMjKxt38LiS4nYJa4Em1VuKEOWkb8x6j5c7zCBST
QnS5D0h7gdHgPmyKPtLo2EDjTwgsUfV31euxuwugLZp3+gGLCkL7A7LFNCD5rGlyfayl6XR7eyyZ
/UnpLim27C0YKp8vmMtghaZCGJmpeu6KOSvSicwws7E64+O5baE7M7HVRPha+YFOlyG5gzk8whIC
NoNGkenXaoa0I7IrkfDHuk+4sfnL54+UT1GwLKs4JWsfIKQidkzKHmAMaR02eC4rMNBdt0kFttX7
0eYMU4d8Of4CW07L19MfNKrTka8zqg5aOuWXhjo2dVX5v+ubQp+IvjuSBoN0KW7mDR4JVrb9oxRh
q36cEkM3TbcuOFAap5oSIrAGIWUs8QNZxo8SCxNZ9sI7ytt8Ox0Q0ZLQcR6tGWsib+jKxuLQLMF7
ASvu4ji03L+urWJdaMDoM+DyC+TNrOd9dAgTNMRnU/tnDkDWdHIHL9O0dh4aB1F6rBcEtbkqhegW
p7zy/yHL2QM8wm3w1GJlZwUp3t1VQtHJ62fgOa9wnhS8Kp1ZJrVONLIa5Q8enGWDusLLvlDjJ2l8
2obU5pTMRWC8LzcaJtavkVoBrnsOQTrZY1IulXA/9NWaroOkquUuChS+5F6pHIZvnbDZtDlSFC/O
wVP8g7kY+/1xlsvwZI5hDdBpu3Bw+YdhC1YePIscJsNj2NXgxy4podo9sldF7a5TBHkOJqGdATUg
ezyzKgVBFx+Lvr0JROsvdYcBuFbrykGD8FQtUi0blbqoRMhVOONtiA7Nfo6LV5ITtBOAFlqYia0V
JCCjHvZzlKAOQng6KXS6lBWJL74YTkLH2oWhx0blT02UmCN/qho+dj/JTro8/uFW05g2uaK8qwjI
+U2dOoF4a86Xs/z3pKqiKCedF5jNst9+DQm90iAsXo/Dd5wRPl6rW0zBfOdInxesEUyVSJhu7A8F
ynUJRn3IQGUo5vXHCy1tMDcd9TcWAqkLVrgBK+IcwSSIXHB5l1zZSwIZGEQRXsAK7+Ffpb33bU4M
pwrsIYJbXBvDrzdFLr+1OaMclFzU2Gl+2ntdRhiXP1Q2gvE+LA6GmiqeD6IEmt6SyfrJyBsbnI8B
gI+5Ulh0t/5V16MoDwogQffhzXo/xbwjUxFeBPhm8c/90vLwpdKYP37Gh4aL1NRLa2O8KFrhooie
uMMStTXAhoTe/vCNa0XNu8IOdnKgnC1jRlDsq5GU/VxCmCXOY/Ug5uoZLrmetYgXXPBkCBvgVEYN
M5uMkc4a5xtIwV6q0lVkusOj1xrF+UknzdNhj+beg183zvz9tbgK4rnlU0Adr6x5dm3MkhrKlDhb
gFhOvZzGANA5/aKhiUOUhRc1EyrJCLv6wcd/Z9IGFgoPbU0P54axRYsRv8PRP1t6g81FwP/NaaLF
N9KqV9Mrk5kPGA8NGBBHX+oB3JcvnHjQP5bBZy/TZqUZRTfl9jV0rKwqX8AQ8GVYux3pYDRz4Ibq
LGDlmxoQGd43ryOZX1caUM+BLvNLXKN/DuXsFuM8BTNcRMc5ooju8nmGvQrvZP7D8HQpACL9SoM0
A48S3gYtE9AUvRtr5TtDZPcyKpvcMKw24iPZ7cp8J0KkQmoXCBghkupYDL0JPWhHBj7yCu26ObZ3
FFgqxE5nmL5yVgQ4pRkR6ZEWapAPussMMIx3Xqg5uRnr9BoV6Mo22jqqn5VBJs6sQ21GD760cv1M
wUhZs6IYP/jOMDXjhPuIWPLEErsNYtrw8pb9JQww1kSXC7zuaIiIQuJ5aB2TN/CME2KqBk1diqY1
6j51ELXB3V2mSgAHPOWK4haXXrw9dqnGpKeFuE8EidP1R9mudd3LI4I84Qdb9+RowDhw93xswALe
tTiKXx2LM+ZSkZ638dVHqm+l/WbNYRqqgnKv82HahEzLe9AkifIlIQNhMmWWVrdmMqGemQ0ZzMg1
ZeQMtBnp/8051SeM32ANKNtOSfomGMS9mosJg2mB2Qqy3imDNSe0FY2N63LpB/kuzwDwSSU37Qxz
CVCY5EZc/W40kwQTHol6kJ4u0Jo9ND+ueIOw26I4G89BOwsiHc7OB3hQcScYNzsn2XijQ2A4A/mB
+X8wZLRoNMkV1b2QGgRpY2Lk/K3GbnLAe1IgbhjTAuytz6Gci6bISyk3N8vwHZjvhUgN7s5ycRzN
QpOrNMjwv0fLYo8hqcgx6Wb4hA+wAr8qhw6iDAraufjS5tp8suNrNq2VaLPhK8GJmlgWvQ4hjBWk
MRrdOoDH8k2yH9z1t3s75/LC2K15YKQE1xGDoz5WFhIkNR9NG7vwn+TOFY2wVGafYZK0VoLekE1n
XjTbg6X588W7hVsX9BR3KBgDcyOmsBilZdsB15iSJ8TO9hZjIk8IxE4brVhIxP3uPIpNs+DI0iWc
TyvdVbfo2fHGOPP2Ro4bw0lTrUBgjEtxP+f0HSBECdbVyk5hR77Jpq+bT53lmcXOfeEAWSnP7TWd
fkIuVKFIh6PUM8oRRPfx84pO3aI+Z4M8Czyx1lXOLPYpaBu7zr6MAMSYeu+mi/z7ClnZ0uV0CP3I
hXUpZweFUqFyvv/sqZ8+PuZODJeJ5k+M9ooZbr7EhYKTFqGwDUTxSc/+VkX+SynHM3gLUlnxdZXf
ezNEuD1TPYKFR43UtrhCNiLTrcimWRyHlm5G0vfIeOU0+5xkbJbSuxGvS8007aL1IpfQhxxgwtNn
hnm3TAnJQ71pvso6oBT9Ny4nzKOsuSW/a44T1xScJwtqPYWTGwA/88+h0B3AjQdT33yIdp+dPw07
B8oHjCw1Hji3EJhkn64vZSQsohFlvfmG7vG1OxsGrLPJ8wSCdbUqJb+oDN9yeJAv6/KhXNPuApJq
vWvjAdJR5ZRmgHN/2HPlcWxhV23sYlOP+tjSXIOHeiATyRKJlV0F/g45sVKBFc+IHDOsHTucuP6p
qdb8zLHRGjnoepqXcuIQFMr7wJAnXyrDtWR/olTqEjrrF0+KBxBtg7Jy10zvdCDS+fmjF2A4UvtM
5oVRqdm86vuHUMv1EOFSuWRyHh/tWuOWh2nYD2n29ZJTxJg5Q0goEidpq000sNUXTC4mTtdVcexO
/kCCtDf/9LFK+olEHKtqK+SWHXYe82j1NX2YPK9pe90h8BdTYaxjK4U9mNTQUAPUqLCy9+zVZscR
9U/QaV7c+Padt/OLBz+F/vytbTvoFg/W0jAC0CioBiM6XbYWlVKyob2gRhWnvpsQdnG8Qzk4bHZY
TwLFogwVsmMmma9P0xDT74DTDCNnmEoIPHN7HGDLhgzZGwGif3Xmf1cuf1WwW7HpsG+TZCYhXLR7
p3eXDbeWpI/dy7rTSBOBZEgdcxiV41ik4WpRraJY3SXfEpMilnihApIWP164/oa+WTvRFM/DcnFO
A9iyvEfVJONJTRTYk63OqszGVJaiTLoGrs4nT8qgA647hcoHsDLZyVGyR4mhQIkPYFVy6LDT0iCN
Yvc3+bZDIthkaNhDBjBpOU289V65D1E5tAII96bu8aK78ZSVFgIDKu2acfhC/t6rOdKGf7ZssdoZ
TQW4UD9iGh+edF2VaFaeRl0HvjKPiYJ7iIQdoyN1d2nkVh3HCSL9nUeJYZlZp062TbUJ8GOlFCAz
APJc7ur558Eh8hOHjkmqKtA5wyII6kZdkuLe3u8VdlFUtE1TgAGTCmP4iiFyhpRvmlDrMAWYSNcw
k5HFs3waovPixd7zU1JGbZsh69blgp25x5qsg+KqLM26GnweBIB2MiXx7iIqAEXqzo2SIh6DjOtL
OcevHckH98dIqjkUkTmHHjw+xaRrhXVbYvzg2+Fv3rd8ri3Ji9JVqiSPJn+uuhXuT22ECh2m/tl7
pk/ijK9omwMvoY1Bs62PAcqqSXB3iL0cw/fUV71eFuwy9HglIntdUCBKmJ8j2TDqM8JsnxkGK54h
CVZuj3nUGaC8EbfPgkSFuyI6zm3ChELZRsFgdQWgwAEalFacI6zWXKk1xvB10LVziirxBPZWNbhP
lpK3WW9H7fRT0MZU+IPyJB/w+dAB5oU3W+qUCcdAhO7ndTEumWbag5BAXtqJvsWfHLCvXbVw8xu/
L2XHDTwCn5Isbna45XpbwAwrOEKaIDI5PTDmOD2bn8U3wKKk1uTt3pw8E7cpMaTgsL2atTprKi6L
8RY7Gri6z574iEA5QkCHnDVKubTApRM+dJY7m73VD+H/rN1czbr5sSL5A1r1WWPqQJSFeH7i17rI
o1Bu9skJHi9dNuECAD4n2eh53c1XCu2EsiHpHs2Xu5iGZNAYq9uEW9KK6hAKMAakEz3VI4TArXVa
Z3N1xG0cBZUs3WGeCH6799YbZ5ngG7fbYdg6iMfxphTYQzgjizktgQjDQZVJeS4jZS0kVcLuYaFh
yMaNUrytiQxIYN732840GdTkDZNTH+PIK9NKV9wSghEtAWvnnwHS2FT7JHrlUxHSFaxhgyTAsiTx
XeDAi7eK4+jc4bTAo71prUBzJ4v9yCLIk3xB+LOEm3BHw/vv6tSpg1/ZjXuj+PazQop3djm2cMN1
imUSlDnhgLZb5sNYcA98yPxmSAS6gRLNAXcPXMPckgIt3mwlZGFREnJk6vUy0w+BNWPD0WqXV10d
X7UOgYflRSxDjkNA2jAMW4fxII2ZuItRgHYl4HayxREPToynTlsaLdlIhLFHFrtb611JArc+xPHG
IBWcUF4hsLrBK2OTnSy/wG6IJMvAKGmecOmNB0cIQAmcG9c3EVbSRZFowWYiAmrMWOP2jj7StpBz
PRm8WnXG5vn6nKRQiUBNQG9aplYujkAOExIpr7ycMUbLDV0V9tw8gi0vQ/U+utIBz84bdAAHNck5
QVDZqkTDbrL+Rf+D022HjbLZ6oZ2XsIfL8JFY2B3w4gHnkWNVMcH3TSf+SSdK3bA878FIm9vHpNd
5lJbE1uKfrkC1VmOiLYL7C6vmsPUc05blAok/RquGTTZea4mB/EdlXnmaGSkG57nSmwtSINnYmUW
Mv8X0defgN1w0+DTZzJS5xli/eXeavwG736q4nWdCSAhcDQQ+BqxUqGQk4k6vCzJyRaV9fQ0Geqn
cGWVYk6WtXW3mbeQ9ISfyopwv8zQK3jfs9d+qT9G4WKM0xunjLXVlrSGHc2+CK10aPGeEg0dMVf7
/MBccBeQg+t5CelwGIYtOltPV0bKROYsnJVVLdZrHhRiysOW03N/A72Hoc4wB0ylPtIICyOD/Lo+
wYWuDYGvP4FG98cGjdlesNn9D7YDeZv8vIG5HOsjFdu6qvFperrDHWVqIicxspg22hAhO1dya3+p
laJMVy+UsiJGxIeYYBS80AYFoNxeTNJHr6ZuetoVTiUJyUfV07as6td9pUcoGslouwgMqGk5zu7x
R/pzuhyx1mFEpDpUstBG60zVI9InPVQeSaEQnjsCdK38Sgw5Q/GeKqzVooriv16zzNzepzREBIjr
5xkHajaSeVqQXCADg4iW6JHgjOHphR4WjpfY542AJNmuXT6UlQ7yzZFlbYs2Y8cisq+A+2qyBbkz
O6GcmTG4OklRMQrUk6KLGuyPAooVyUnV6jYJ/L/DWTB8b4F6wIL0m+lH9Do3WBoCsQVBe+yACver
2NRRkf33Gia+KUktKaGkTnYOZwYm35RjV5seOncXLdX4lchBKjQLg20b7oaG9wf+ZyFpvVjmLk+H
eT8731kIXqEe//SA7uy0yYkeim0FpwZedT2wS+NOv+7f8S/DZL4eACST6+7MxOz+lCfAG4QqFpWx
S/sULonBBdT3+k+6G9w8Kt0JPhyTuiX47tF+bDxj4ZkEtE9OsgnYJAMASLmLyqlFN/nBPpTQnKIt
yJ2qeWKb1vf+07W9lFErOFxjdll5zMBP0X2bIa8U4TOln5zZGdklj5tYkh8tvH+N46zukMu/YznV
vC80yW/vxJp2XgymVl+bf6x3omdNGnY39u8feIAQ3KeD26200WjRncPNZ+RkWtjkZ6WMWqWv9J6M
PO1Ns2PJBMZu6gSyBjBEftt/SvlkJhskpgbADFz3sl5iZ/wNvLFIBZsklti8vK/oU/iEUScXd4aW
LGkQbYR/Agm0Tu+mWpXrVQbOqjXHjH1D0xRg7/kpp0ABQ6mvQ/W3SS9ES0fcqA5kFUOjHVK0nLAX
Os/eiFAoPJB/zhsNWNCbPhp/9zS+0p8/jq64UTK7ogxdLhWDdvsEn1/YWg5kSje3SyhLey1Cwuzd
pyQb+IEPx6MD/kCTy515FhEU6QN1DU/cVN3GIZQRm1jbZVAYyRtPYUSwgt0SghT/K+KDYGevvOg1
iSN/fGobebDP8fQ2FY0/00zX386tpZjjxcIDSrzfC0Qv2SRoIVPXXjMbbiX6mvl2Azx3apWYgi16
1BgRzzMQLIUlBFXmOZ52kgiz7onbkqxHZLD6Drf05hosla1TFqvxGy8KXznbpt8lA6l7+DbipA2W
cu6rFjkZxosRwJHmZoYokXDC9uKLjqpGcqhx2kf6pIggVQsz4c+YIb152xO3FViCYhcAhGqg6s7D
oRKzPC4onGeU7A2uePmffVHjyBThsJ7cERbp8Y6vFE5Hp8J6Qy7SdZP/4GFrycs3jv6kZptUR/BD
fZ9zGhN7V3VEcsuE5xpdb9VDgv5w5DGXVVHCuW2/EkfvM95rsaWBGfWcxHzfuNV0UGHWBhr7hWcH
mxTxeqxrJ9Lwnko4XvqTyHwbldcWjqrgm4h1UTIlQJl2RNTXytUd6lvavpaXimTU/93GpDy2td64
EtGO6prtnPFhjzw3FW4oNfx7VmXd9ZKS9oB1esIoevHt/HdLFisvAn8qXUl9IbMSxSrN1R4hEgTJ
05EqtLL6gu1KsgeZLUdRizcDeCtm2I5SQGSnnOHgw5mWTkD63tvEzEuKkG+jUAH+V48zFD0MLfsi
s9+knvHlFU0H1O2y9G/SoXtstMW1EjmCX7Jm7XSsk6GL4oGnF5QSCu8GTkfF/2un+I3s0NlWmeeT
J3o9vkyFkL0s4f8/ZqbZNwvj3P/z7tZOCBUH4HoC/utQIbLq2Ng1eKJH9d+hNmg4rdBLz2+bRKxM
IDW21fwPMLbZO4oBdgT152HVrYBIokVEzpbAoKZV8GtxGnj5artVL9AquhSrV/k4zHrctPxDPt0I
e9nugb8q8rU49e1w9yFuHCl2I5+QahHB0FfVTWQfZfo1PyaVd/ERB8p83tDxq25ghxLJNc2EVFB0
EByOO72ifdt97HKRGCfsyqk6NPfRAR+aj0iO80Ez1M+Km3nOEwOUvWPIvVznJXHp9yN835y5Zsn2
AGtVWiqlNmttYkffzlpcYKXhR3tDYrJf5CMhNwo3RZqynB6E6oz4pyMvgkj9ZWy8+EqHogdGTAUM
BzSh14FBnUetCbIb62vJsDPtoYkvbjISDDcR3Ydj/DRIvou+3GrW3z2HkZHcOeNqsGkHABOPKelS
b53RfcKPkhcUg49ydTSw3iVp533Y9FMu6r2OuxONDLAxdgy5LrawBxWaMhQK0wIB6udi7taq0yQz
7vF6xqq/fNQDJKsJASq3QCo0RWsO8FvQ3sTXbfYyAb7mLXJOIumzJr8gMMBb2s3ZxFMqN74+ap24
SHhJRmJpRiu2hYN4mdC1exsHs7PfYz2giGHz5EabVgP1fOJlTxzPV4pjkYLmkg+FVlHQN1lbAm37
6zwMipIrBX4aYlZj9VvETaAQ/PekEmLnoWmD6FjH7ZcA58Cn6fpcRei7FUdBaMPN6jVju7WGysD1
+Cl9oSrD6U8cjrbi79MvhI9Nd7zP76LPTytAW2lNSsZP+13s7hPnC1x2u64NILzUUsaYk8/PiI8t
MdYV8kdyvIBMkr7CDx/oeHwV9biPELnvmmgA4FNWin2nap7EJuvkeIub7N1NasW+4URogTD1Izi2
yv7l0kvD83OaIhhmuhqKqGc6dY0WT5IMWfUdXPESFsVhyN6BDC/yoUUy/jsw2IA9gd1So935wGp5
yMo0RZyefCd4NXTLGZx7lgLZ5h0g6n4sQl52aHRSzGfBB02ZFLrrAK0LRaagTMbmxNce5hgLQdff
g7BwZZp/Kl8lec3GHa6llgdUOvTbaY6RI/KNyr+3afAzkQNH7esNwJh4XrReE0mcMwHW9FCosWM/
lbM8daii2cCtfJalV3S1y0/o1nnErlItf6s5EquH1kYFoFTl6f7oPz4V6wK7cOnOkmxi8TB2W7S9
q1/WXnkTEBC+IwRm2Tjmh+fAuqB/Ncp+ZFPItu45jGAh/olF6obNbwqda4va2pSq/FL/eVWlqO9H
gBIKyfwyMPM/E0dE5n27uYzOz6nA9tqxOIrL/iwiXdl6tvpGWqk0AwYvXW097oZFsuP5XxK4hw7v
b9NiuqNXFiFOTcw7jNCdestgwpvU9VpryQh2GBNVFcx++kdq5IbTT80RNV0rN7XdM+9/JiPaRr7y
XBuPtvRvV/nN8pmo3j4ZFuVFj2d327X5uLYy0dj8r5d8Ep141m2TWB+d7Br+HvKsRGdjKV8g7RRC
W7yI5iz2dRApjMtL/uUgyECr6HMOY9gTGh4+dxvbBA0/Bml5ZMWTJn8o+3eiPPBRcOtDka9N2ww9
Ap1gLvhcZ2DDdQ4uugvWqsKUz2pBcRql06tE83zXYZ1aDa8uc+uA/RPJwuJkqW7HA6y96E6xWMSR
LA+ALIHlD3czfzSrJJFsX3ZyxywGl1ueSA39zJtpWQekcebEXXar2Z1r3bml/b0Z3kKR5/6v2ptV
zXaN19NFL9T3F4SGrQPYVq+eDCxNA8uovBzMVfOZZGrpFzZ078Uo+UiYo13GRxfEDzcvE5cA9wg7
jTyPKRONLHPxc7388opo9xtqMeeWyUfTeI9WF3hhMi3DhfJQ8yIiInRqMhNM1WYyUEVHAtWjLmRx
2KdVVQhc2ZV4TN0WuOwW+XfcL92HchR+UW9uWAgMM1DjJS6Els68dqWp5FCpWrNHYRuCUX9UchXM
3NwgWQvLBcqK+/QCjjoNUED7B/z8BA0HYqXqIwv9YfE7FDkH0LBnrOlDwhcmdFtzFoBuEoy07HVh
YhQpuMClN9eoYgijGWRQi0sNpqetmyZmmtefoeqv3Lvx/I9Yc6uUznaY3UId4TewMcDmTcw09jYt
9meKssEqxQWOctxEhQIXjzoRBq7MJb3lJU4UeySYr6x/u9IkGL6Vbl3/tgjvJ8RK1nLr80NxB27t
FWYBW861QeCW/sUGu0bcSxvPm7OCSKCGLUoe8LyImLadQrccXofAcWNWZ337EooWgQ+JwYBpz4UI
Nz7+WOs1J4B5pErTuysHSp3/tPRO6Cb15CuK++zw7cmNMdqyF5lpSVqWuORoC8bAaQKeMw1RLZMh
X1qVZXU7uGRzMiiKDTAdzrkG8tCLwpi5XZztKGhMn9QqTSlFofK9sJf6G8qrfjWpf1sdsLsI+g7u
lJ3sl4NKtMNVxAiFcMlCk8AyvgV8PaKTwo2SLbtaxWJ+QLoPEm3p03pCaHvM9COtC7jgNXt6f3kH
rEZ4xSXu2Md0E0+2gLnkLFA3kF21gW9XM3y5Bdtg/6wJbJhfJX/8fG5XKpDcFD+kqTm14I6U09ji
+rlfNklr3iSz19nPg0KLRhzgCBmjU7mm33htcokkbYwJQ/WKT3GI24m6hLDixuaNhssy/2Uil2LI
cio6IRUBqL+PH4+l6uareW/EwSYGgB1oBLpml3njuL6mIKvy+Bu7Clb+1pq0LSmQswZYhHN3fYuQ
q4NUSp4iqAEMdTF87Cl37+6/s8x2mwl6s8TI6xPtQW+EZbbNSiaLfE8gE3GYeRoKkkRiz8ALwpFK
5iEwqxWOnEbXWiyraQ8ru5MBdjeOVDxbBqRI4jjlpmkljjjPFWSln02c52z+QZaJrcj863qYI591
+h+VK4OjEYY4bDEpD3qdFPDC6stckBiwJ/hITLiiyNDbPYHiS075EhekXCXU/N2xbec2l6J4RvPV
pUJtH2aJkSPL10fRg6FJwVZTH/4x9x+p/B5sfa1uhsxTirDJWy1ivhDZ+S2luvTFJXmQ3+l2YAAq
zAY2l1PAcaBdQnuDt/3ZgbRb+l7njU3KWtwW4Btb9ETC5QhPsUP0K4USMgHw10tpvJRqTWBYsbBt
Bf2Tf32uPVaLIUYCETZ1OrmdEn5fq4tSVeuXhA7B9JSLjKqw21VavZnSKPLo2p9S61nhFXJR2XJb
DaX6WzAAPyv2y1VVmimbp6gOhXyfJQoQWq8J6AYZabrOhovHsJ1LTNewlfNQ59Bi2Od6NpWzPY5X
Ak41Tupkucdhtr1mshZMXoZkW1IoHaW9WSH/KoqrxFwQox5VNjzBOeXUXT+jFfYvt8/60sTJiBXW
ry2YvFwjFLqwOjJHJfA6qczt2/0ictNQimQauTWBRw9iVeP/znplVmAYh0k7YUlNqGmmy9+GU2Bz
coCsabu843q+4ZHEwbTOqBBTlKVOPU3BRQtIevMQKEk+odazLpA0BjWwz6PpY4PETLHezOh9i76i
H4TS+NGbtsrkZnd1A7LUDAqaG42tG79Skhsh0bNaOvttqxOUTIZWvHQdtii+/VoVSIYfwojOxkpN
gPF3dFuMcfvc5kdu//4KYHD699Wk23ISHzMeX0OOJg0Off6nKlQ+dSTPT+QyogJljkZFbf0xvlHD
eSAtv91w+rZe3L4n0Uv7LyQdOSIIT2Luv8cFYE54E/2Hzjcap07V2EwaPqikJt3yfzXcwmtDaYXC
h7My8fIRisQL07yn3jhsUyGWcQ+oJe9v9eYcc+bPciBRm/UItsURjQxPepHZ0hfFPb1mYWs4/8J8
yMn0GDypckGOytRZWcY+0q7jbfCuYKTB0cwMGg3cy06rdGV/9aVgsYng7gMeR0DVeW8poaJmkO5k
m4ekeTFK0KGbef/2BkCU8j1STUxQGDSYAXnhl9FmQKbET9BuAlp/P2FZqv17kMiywcxUStrG72+M
r5Djfcrpjq+UqS+Vu0bf9QP5n9LkgrKLGSpOSYHs0A1l9NoAvgJY4VZIw7T5en+B2aoOa2Xwejz0
B6NcQ4KNWB6u1GFTnT/+lZHkY07hY6XeagsOqXhrBCSVA7brfHN+S9nKfparPXQoPFD7rf3YXlTU
h71GOs3mXTJlWd60wb7YlL0PvUKcKgZXxbhdI/GBa/KU8jaEqCK0TSjJSOa5YEa+TnAAPU6o6z5k
FN4XLqojZ3gpM4njelwSL1i3jRvw9gdDRM8gpftFRcFKvKOGidFZ/i6GvYVoZg5CT9m3feE28dZS
f/i814P4prac5ubtkVRLFUTGJOvaK2czXzV3KDb+p0B1WP/j+x6oAtk4SpHOoJ8E0ax9JOgN1dCp
4nDpYz9X48VTQifXHVr3iEQf5xOUFpxBQmfWP4iMEQ9DCKCiKFWENptg0lVoXEPgMlzV0QRig6HP
ysouTr9ryhIHVtwfj6RFG8vVwt0f2bxNTc8A4xmApK3Fkd4qiiDWsXesodT7w1dKeN6G7S0SOHeD
bzVRZ9w5bxzsaAf3d6enb87id0zgXlQ/pXyVfKFIRqlH0npxcW14WaBZO5PIysZCfFEOYUESniRp
8IuUHd5t1ojnlQXpEn8milz1OI/pF9T5QAiTGXXRSg6uygNDeLGk+tPjniVp9oaKx2CONCeKxjBL
g7oxD7ti4TfWq/7Gsc/BS4byN7MzUgta3aMvW6Yn0KxEOZECYQiKJZQAjVFqOVWrVcihORilBKb8
VGckzjj8KPcBvDBX+uEAUOYU7qimz/9Gysun2snT/wtDsE9Dn7GFrAJTs4WU2M3jbwwCzPjDosDa
2v0SPMnpyAw6lF2fUKTTGA5FkW3O2KDgV+cFIMGPeyNX+rzEWA6clnef56ZRf1q9w6x/5J+qnO66
31NiXOueL83pctlWmZ/1G2QkhhwvFCkYiUTnu2ghs/NbrltKumkjGUMmXm+QfvIRd4P6E1qZtV3z
k4jFNyfrqZpM0Oak/DzhdhCl5iCBDQnTF/GPNZ0NdGdY+Ijwis09adv69n899TNYc+OKMy5jpxYD
e9UR5gy4YSTnVWUZSQhdSgps5E5ZLKOu4OKHrCa1qsYI9tZPp4yGMMc+IahI/x+THy+Z/cE/SAgU
rk55oD2OUtv+sJJW45lQvgDth5C5C5AiNm1oqRxsNPNf9gz0UjFPYNA6Rcbntg4OP/pgkt7y0FbB
Dp9HnrhI/kFyUp/lIy2z3Q31rpzGhe1iytpLTNmKu3a+3WG/alPe9uRQTrWS0Hy9ZX+jWuz78//0
0ExiE2g5l5AA4aFHReXufMmnbeAq0Yy/d+pn1LeslfN2wq7+0Ekb796rQc/9OtM8w6L4KVT3Uro2
Al2NfgLNnhHFK76wDzoX7pGKahf7bKulFbO64u887MCutEmiWsqp/tIeewE6DBaCWX/kOYrd7XEu
R6QUCqX5E0lVuj6K1f1wK9klMrmohL/LFSSOtw2j3kkk+3uWB3n/ea07OQL50PonKFQIvfFwdyHO
lImAxYRsqkeLNv5a64dMuwvhI7zwDCRFCkP0lTpYJLjKHDhzQPn33m/TsOXPeyKOGeh2DoBB/SSs
qwAJsqWXN7xaOJr0mxsOnTppfiRGz2jx+guYImw3eFVvOQm+RnCJ0EH47X/vrCH9X+s7fMHX8qGD
+2JdLgxvs+cclJQJKcmAlCCy7Faox/4pUSf3HP+eCfe0qwNuQQ7WhzOKHgI4xxi1g3V+Qw0CLJH9
Vqq9lVn0JXWdytho8SZfEw3ZfLGY/VQ6kxjxCnRqySqNHeBVZhrcfzqTxrlvy9O2GNSWU9ailx6I
PoDsHH0rrh7Js1DVQKOjW7bTbBoCzjjvl0Eeu6dOQOEVICNDuXm7JuEcvmPvunehJfzxvzL1F/N3
VenDuY6yPOPPNCfhpADjGE3gH5Qhqzm91fH5IucXqDOboYMY+IxXETDENPjQj8AiPgi78APBSxfs
A2E9bNiv/zhW5vKWaVzmB/drer7eE4+R2kblNTpOTc4LXPdiVKFMhJbasCEjfaBtkKcoG5Vqubrj
lDuJhIJaHQ33+zSvssjbPPra/guVsbhiP8ryD40z7Ix1/UpLZR9Lt5SaGV/XmQb8K+oKWZNu7j4N
NMi9bYboMG6De4uwPRprJAykoviXEs6KeQA1dmXNfFIFRo87Yh9qPUunJmantyQm98n09lKJwCv4
iLj0+LmYA2zqzSbE0nzNu05yogYs+vwADkQEx60kOSUPArWfmQ21sMTxMLZHdDtslq2+HKS0gGv0
8SaHGKaEyEaOMrQhmMXBi4XUUPurPgHgQlausx3S7rvSTzWztTTq2716WakQKBYoo8MGxWhldxDV
y/MhzT26dHt1rT3Yzq9myrfRrvWD2rQoO81A5ZExrA3Owml/iLe0yKVbKwFtCFY5tHa2RaZgS5/E
CuuDGjItxKqaR3otZAFCLQijrOtjTHoC3zRquvYjOyxp53tWAJjop3f2p1HA7WNV7m7hHFsNEkWf
PGdStM+ia9rnX8sq4WiaQkeBGUvW9JoKzzSCTtQ+W3ZcYgdj19CrqkU2OKoPRb82m2Gh+uGiI8lO
m2/JN1DS1pvsrVEnd5tgmDSY3YQOVXjRXelwur8kbRNib06Xcib00hMkTHRMzNWETVnk9YoQuVyZ
PQbRCHpE5sJCydkCx2IyQXIdruBK3k5bg6ISpkOM2Wvy2h/PmsmUm4UxmtQFGjOT/g5MYe6cVWWY
X5Zs6IQGp9TJ3zn+5FnXCE6OMbBszybS5uZXEN8uJGDPWGeMT0b3pkNF5i2bR6YgebptlN+U6liS
nB9SloXHzXmaBOXsjr5J2A3yvh8Zp9qoGjHS42/BMe6/JL/A7exL204CV/rU3rWNWq0C0IEuI48i
xY+Yct9hIT6YOmHLTSg0PoqJMN5bQ8kLC48CQbWfqKrMJqw0Fome8vQl7Fo3i2lX7a2IjfHUyYiM
51MgqvcUk7nu6nsHQJLeXGQMqVWNTM5PedljWbFeZ9xIJ9dX2svKqWVwnyKkuCAjjJhXieEtlbBD
zBd8uiqhkZdL9s8EkYdxO/ls5719ZyFwzXLhsk/fmtPoxwPHEvR9xwrc2VUero9omHO/Ibv8IPHe
EEpXA7z15nZhTRk3S1AXh5xF+XitxZZjtGgfNG69TvX/HLcg3ny2VjvN0RgA1IOPkY5zLo/m2A2t
8/tox2BY/mPxOX0VZeoxj4XliuB66+7MInx4SwgHTeyqfhT2P0UUPcYUFgnorliJ5b1MezaXf73A
WNCG3ObGxLv0rraKJZHRQLBNhKQ41ruLZiMq1kyXouH8bqBY7OKofqwdtw0OsKPh+KPE9nLIz72S
abbJ31As7QaWkg49hkFmMa58YZWq5f8ur2SReVsZYBCX8+WTCXRFobO4H3sDFLAFQjI/9IOI/DQq
feN3Dw2AGyGVsaYVp2TLqvb0OVZqAJidR3SBbOVcBeyvvyd+o/q/7Y3WHx3cOBu5yzGdB27NN/e/
dicI9xA8bqe5wP8+vM3Y1jyc6CiV/H7KGi5oyEsoZKRddvtQ1kuQP2OUJx0Y4EZKHtoHiJQaroUT
JaXgHmQFLhDiNagj/3Ag80NKFTRYuae0ooOw2le+C/fQgPppl2ILKzDDhAfWaJ6EVgSgKaZWgFp+
ifHXuBhyDLk3Sk0dGL5tlXSgGgWipFSKkfT7Evik6LorKPA9y6EkdRjZ1/4f7zVGYq/3UEmYSf+p
YFOgzo3YVYG0CDJyWyEozbkmArm0681kbEn7LTuJBCd+EjlZATO9nZZGKuU65UO7O12ltoeZKR4+
XQLyICGiRhX9hL310CsGSUortgPXekppGCNDG5w1egvUYL7klrghF/DbKFZZgnhDEMaVCZcff2VC
HuG5hJkduclSHbd4nDeFxrAD9bqU/t3qZbdTsjvjpjGF3AQzWBMgWpEcHXSQN3nyAqrL/iLtzplM
CLxM4ZDQc9PrIPU9r+S6VGliN9g0z+b8rM+HrO48dz6AA/piBFpSrq5tnP/21vygaG6mrHA6qbmW
rhdcQ6GUIKDtuYWDk4DRIrES9mi/jEo95rtTSjZv087sSLOiA+SWYPlxH9sOnOi/I9yfxx/Y0O0b
poMldYlzcD70ac/65wNIvYqvhaq+eCFXZKOkCzWBHqkTyaCeU7PjE5unshW8PMwxTwuOvbWcaPXH
FDDPQNwE8UeeOHDzJbzKc2wlSUb/RN1WypddelIrlfpBrf0SqXRVEbBYDfU7gVjmWzTpWsA2M/YV
go0t7KWFTOiWm4oVjsQxezv27wvTKNaH0KRMXllhxzLQD7Rv7kI7Tbv1Qr6/lDAw2JjQ6br5i2n7
z/2DKxbZApQYpSEkwL3CvD6niSNFsjT0XiKIB60klvDpg0R0UEqXsHLohC9e9PdDIcFBQPvKciR9
M73kAW9gMFjSNSQslKveNTcXa6A2ZkbyS2zJ/FfcJj2wCEgolCVWr6RTQUpP0t6+WIZYqNbG9P9G
MnImKDeBWjBkuzshJLvZfcKpUr+mvvTndIkkRZamp9zi5BaAmJt7CtHHwlJqTtDDfvWq4xKbFbCv
0l3TTPSt4Ru4tBo9k9kM0G6qRtLBYlamVBnKkqK1JOnRLOkDUxPE3x8z8JN/LvmybNGdjUhJlcOS
tByyKVO6tt3o62vYjo1XOFUGvODss6GYczwHicda0ApZhXDGJeH7OoWvHBkfVVjIydVNNEzHlQFS
W0C7aI6JdngCw1K5hD750+fAT32k8odq53Tfn5Fn5S/W0omm721S6ulbBYkhxf3zGvYIOMA9G/DK
VnOhuywA8o5tsguCsRfWdGfksXtyKDrHlS4EOAm/ajqKA7frWVVNYYN/p69kHdLNs3zXOkD5BHYR
2MU4Mo7gsCL0w9Sl9apHU4xqwvASzKT8qphmfTR8s0amcVcCweinO+MYyjJrcYto+7fNX+i3k8N7
RF7rygOTBThm6O7Uoe0bqbYho3k4Ly52LJTU3pDFSfTobQgduWjNn91ldV7efzLTJYgsyLLJIDj1
fefi4x5nzNLu4XAJldp5K/ApKuHIX3PVkHD2gbbk+xprebGDk8okfWDLbCpKy0t37Mg/WlkRUd5n
zje49HT/UP8Pm1WdUXY4n24z4/gmDP67YadWKFtJGbQhyyrhQF5/Y1TXFcNtES3FmDvIv3PKJdm0
3QtCv9z4rXiWhhvEWoVV4T/bHQrvq9r1AsmCoh7XQtfiTZ2t8xxiDmoQsl80wTm2v9uvXuB92n0z
seOQQoepecwxaH9Huo2bOLVClC0Wmchor9tYSTc65d1r/2c285kSsjKJgNxXYrEM4H3QxjpaRfwo
PqBy8j7VbNP0XRXFBNCe3AVq0O88bwGXrmC+hSq90qMHLOscHmmJVxXuybSZVEz+YVocUWJixwxE
QgXNY5QCbRiAKMCdZc1ddK8Eowgg1aA4sT3UuEVdDoCHSuW4uZaxRn9atEcUaMZpHxuxfsuywyWI
JsP0fJsh3RqL+yHDvyfqFswcP40sGqxXAhNtI7O1JtsujszWIaetau5kF6gYiTYahtbJXFiMcmxE
RKqIQITJC1ZovleiX57qGpVZmwMGPsUvaFx4MC3iiw3PY9MAM4h0iPWHX92St8jES6rdP4Q1TTaC
n8qW5bSiXoDCUAPOvwWQZB+43gdtUIzAjLCVDzUZ1PggFAXyJiLaXrqo+ddDBHHY0ilooD86mHsE
q8U7ym1BRRwjomJQKA1cyW+K5siMqjC4VOvyoXaJs+f7Dm5+p8h5lBDbCDl8ezK6OpUYnBw2VyHV
V7qWIbg5AMB3GrCgD2QITS/bcWrCil3RXusiT+hrcasNhBl+qpuqduDBtKb3lNn4H4sx1+/4xccu
U4WmxuSbhmmj1WXQS4fXr+Ak1Da5ZPKd/3fehC/XS4PlpAaXm3Px7De1eK24rbMYYaABIidMwL6H
thpHxfcE09DzH9YjvHfYHxI/GMyx/9an8zCy46cFJjoHH/Pxl5hEIQ9q1kMAvnL5oL/s/2u6WSWO
jYlPZOBUyb9u7BOl6OLSPF5TsjTXzeVdFrOMzKqUQXjmjFfZmadN5L4oXtwRG7eqP3dMr05Y3c/g
HNoJZNo3QLzCXZKDy8EDsKnleHFGFKQ/R6kgAcm4dnx/fLEdfeiRDEVoC14JxfXAf5hOR2X9vcng
TT2U6N05ATfdqxkXV0tXC7V95Kzocb93Ce0FrNBIA74Rmc5a8xJR1GvQoL4z6b8oQ77krWOcGV9G
fnpAECyDNDdnp3Aa/FRme9y88c45SUcAKFKIzZTu/NlvfAJ8Lw/ICMYU9biyrrMh3igVC9/y7JBs
BZd9mO20t37BSaZYE/zYgNpsq5ir00fDp6RB8rMymBC9dYIO1JJQtEqWJ7+Mws6dUWeSTX6LtgEZ
OrfSpsMxrmj3kbBPf5dBN9RZFgGfj06Vh9d6DPE24BsNF1PbzguqXI1SldNcZvGvx35QEPuHLatg
tI0BrziwDqLg87C3FNCCz8ReGMJb4LcsE03vPGxXneVMy50E2nmn3sOgtHqDfcajaTSU3b01ZWjP
g6/R4Gfglh6NN7kdqB32o8C05qT8PhIOm52kzg6+NGkVZ4mSm5+TvRcbMiinzakz+IGPSDn0XVsy
RifvqRRLVvIeuwnIz685uRs/RsGNmrd8FgtkDWqfbJ2CDdz3zDrFqgurNvU+GU/i6D5QkIr1Fr/s
hHGu0nqU4vXwoFF5cxiQwK2hAMWhvutpgSYLkI/v7zTt4P8+KDBChZ53K0DnogKl09tIOMLyFIm7
yuaUG6soE+o+bjQRFCIay6MTLRsbcAhOp8KGWdz3hPp70wxhI5R+S/hUXwvE7/oU7NoKJGBa6G+x
hYSr4/XoyKF4RfD77wrweznLoh1H+ZzqAIjbHee4clOfKjmhXHj4cnS08insOgk8SonCJJAiq88H
VlBO8MwSZOUOc0/o4xdC0PE6c0jh+JaGUTcLm2sfNzS/zcZ8RiHyMPgJLws9zjRvFyPsKhY8a7VT
PaZBfHFnuhu5LCJaetRHtmrDa+Mg8vBXoreBy//byakOnApbQhMcRZcBsc/a8PNsXjIyD7q/OPYA
sZdJEotMLaztzVVG98F40kLZy2HyVyTc1qnkleJWuGnL/GwkIonuiqCH7s5fmJVlk8zvQ4krH6JH
GJdxW7By6VxvO5dlhfGenRd7U3+MBUST9mKmsnKaAo7WRxcLy5inFzJjAjxeb/3aEyBw02aN8DOj
1t6+Wp+TFULYa5zy7K7t9XhbIdkrXw9M8lRzTVE9cinMQyVzs2GiTcf817CxIGn6Js0OeFJ8PxaC
XYf5knFOs/S7AOdOzsAYUXc6tFbdN4Lv7GxEa7yguBz4vcos09TEPFStu+vW7XBFYaYEyItyJWa8
Do7G3xRMiffy8QGpD4BYhmnW5cyYehHkR8izhn3dWanuhjZYw4mWsHv7nS7AJUjx0aEWxbmokLDS
F4JFl0RtdvnYHJGddpKi9YAJUTvZetUv0iR3JEsTtLYZvJBcz6FhjWA2CP8fStNN04qd3iDa7/X+
eTeTU2VRjQwaGFHIA3EA9I7xWdvZc1kSL+wQHRnoUIQHXy/H+bxzx9D7aDlwKfWeT0Da8Pz5YPBb
i/62WutAEIe25BSzabiC+Ky8SkW2FG1q2xv5a/X8UfuB5gHgQic/jCLZBO980vfopiCNGtAFdS4I
d6RfrMgZliOIKE2jsMeEIodL0dMmY1pjljGBe8ub9og0eJLXNZ0MjvJ2WYgesZdm5lH1OgHns/Dy
Eg45X38gH0OYY8MTa2vAV+VOc5Chc+1OG7YexHq579LoJxtAZl/jX/qh7meYszKxhYgZkzhJKyhO
lbGGfy7bN/cIRFYC7wPnj9SlrHDx7xVegcbgvGQQ+oaQPjxs/WwgZMUveXLZXAM/c7MbSHyWZyR5
mOP69t/GEK9Qogbvpg+SKGtc9TyDEJvGW2KCgHzmFUzu5HrTUK+ofdHpelbwb84ZPy/q/fcgaGjv
JhA1yF22M8tan083YqXg2/jjTCNNuCj18DMBKj/aWVtTIMpb/YzIRk6XizPHLCkAIvdPp+o88Ap4
17veKtpt/5X9IKIZpUOXobX223YJwyo8YSUNwAn+ZlUjcwHXOUe8TlFGVXmGOpD5bg9fKt2zE75B
AE+pkf+bgZ4SBU3nIf9w8+kAVSmLHuAeZWCiAo6iS6NtnGbZ9BQ+UX9GYR618RPHmypsLscYzNqX
w8R0o7YAUKXJ3A4vDqgcerK6PDE19ChhcSwtTFihN12A6SBADKUmc1ep5rqz7e8FMgYffRcgzjG9
JQlu5ylN7KM+DDeXLcyfODko+5r3UXqSKdNiVWTaEG+LrzJK2YjGGhfzSgYTgun4HVrM8EcKZj1F
g1dEBjxWmxOz0asvLeEo8Qk2vSSdBZKuWdHQNAQBplepzzvk+PH6rOlBR4RrZhEWq5T66VNLUGap
fCbTe3HU8mX+kojB4sjiV/sLtcduOLKbLmu5TJkjDKGYhCTVZRi4eavqlKX0xoNNj3Ad8cBrtTRM
ytoAsqR5V4nOGo1KAV/D3+BLkZ2G7F8km0hGNH7WKifyJjnhKyG0x7hfndtlzqIFDcyvsRTkQfql
y2jrNVhXDp+zoNrKHJmNNtSlBwocnHvmKeFc4yUdKs5SHwCHSMu0XQTQ1ZNjSQdsNuayYnd0VYaj
VZTYOCdRk7727/Eo6hV7a2RbT0FUDBS3h4xQZ2J2Oak2QPee7wgJbTN0kBrsDp/IcOt+gaSAMJJQ
xLh2ts9LCp2fvWwy++3wbH9YIgyEvHaWfnBMP4VPkJk02d/Laa/9bCI7V0hhhgjjf1v0VNsQ2gV8
BXebt6oAgMSFuo9vqZmuB3OxmM3DAr7kASkqX2H7PyHMQfkut8jphzKGREUkRnVZ1+HfxUwIJDZU
CK9668k2Lmn8Ij1Tf5OranOgUYMEpzl++jRPhZkGDu2GdQHchZS7NiuygB16ebdmVNN13+RrXYSM
StwmUH26208464Za6WGHoI2nRJGLb/mBB0xv1RAib7vWyvwPylpV/YYIAGsDvyC0ovNcaqHJkngj
8I8cQre4oAA2glngONp49N/YlFWpO1JBmNhxqSERX2O7RzMY/No3tK7i4jyPwiT786GdwsqogEeK
ysMs2uoueksLsG4rERWwHdFc3Nm+WJ1r9YZgXonIx8GSSnky2s0dBFRXH8zXC0uSJ6H4DlZID+ZT
PgLshqd6Ehc9jRVrt+bw7/b3mTNoYTT+UAIaaFh9RRI8z6nhN+8dUBWXhEr76NrCpZIC/5S8vSkW
CVWAu4y4pxhd8fHWavhU+kppWDRotbAsakm+I9MsFcJeczHWK5lLpdP3g6yMbl0cEwzwc28IE6KH
ICEaXk2lTJGqJzcvtnGVk9QqxdEp8tCt+zNTiI7d7fEmee6TsnY5P5JY3S5GmdQPyTM+MelNdj0Q
y5plRzab++6PlEjGx90a6DSFwc7frgZBur9EIgQt2KhRaZ0hzIcXQvaff3JRNqCzUVYFrF6qTTI4
tarV7Ic7sknPdNb1nzWfWpC5nhsRfCA+01gKIECsYRV1f4Y5f8KwBogNJMZd/sEuBr+vwl+MOOz1
O4pgMwKcmt3M/f+OTIBCXAOR4sUiNuWoBvTr4mcXmZcfvMmONiy4p0MCklKRgD0sw+cB4fEgSuJo
X5r/LRmT5weNsYYqz7hIYWT4lsOJlV/KoyUGMUEDV7XDXLDjwLPNkEdADEu/4s9f3eUe+QFg0hci
9RalUsc+3TYjtHlsCe4YBXejlC5dq4O7Jf0Ee2+MXahHGUr/WaJzQ85zJFf3gyNjCQaYzLQdzRKn
U99eugBdkeP0VamEnbtlmmKSqL57sXshkvTiE4hCcWEVo+3M9U6YZhwoeGI/oV4uZhnAdqfBMUVX
J1qU707BlZR7jUvfWgnFZPh/ohY/qTaWDZhiWcppR4OLJsLd6EtoDWZZCFO3J3LcBqKXO0eRk8I9
2npVlNXYuBu5bmIhva0aWgE8NI7l0NoloZ2KFWQgG29ENdww2tvmEuzwTcefMvx+hs/RPgraSInj
f23S16NuMh7dKsye/P6h04kC24MH9X+wL22HbKDfhL9n8Gdja/0HbEbaK4ZtQTr8CXLBAQaT2fEo
asIq3qP3Q5iiVvp1Cf/k99ccvqOZ9/e5cHu9y9icA9HQ1WXQtb6Qq2BDEvVX64YkOy72Z0g7BKrj
Kp3EsQZ6M9UghOMSKF5OWc6c9YJnMwvyLbidEbEEa72awLEAbN30AdXmAHSAhXYsQSSXejE1Sj9w
dbH0xFwuMBS9XfnJvKTedJwE1KzfB/RWgr5d0yKmgFIXFekLDfh5Z9RMwMXWAbw/yRBWFyrzcAxJ
uvk6nXT9Phl/UZHmcjN5loCJ2m32Y5Qyio4OL5l069dCmhqg6u8iylJFqC6xoGN0jlX492xLn8mB
rLa2ElRiRBldNsDcc/8O7KrGTrL/2933KKcO+am83FwLaNiuL0rITUJ8eIgKrMIYh8gzfkHtN/qg
GscorUmXHnDpNmpt2YV3rD3P0qBKKTYls4qww/nPjNbtvOhxlG0jpFlXwww4uPIhRrtN6r++E8nr
4jKLlKkSh2znO/sMmdBS+kyv91i//F2ae1x8f0fhRCDjis3eL7KPnqRD6CWMdL+5g+HuO8D4fJoY
kXbKmuorJfoYiB/cJ5YS210totGZWAOWkRHkLT0l/vMhvWON3U5AMI/OpsjdIJgWh8+qzqy7U7cU
9PWnFXy933lUoc+WEw0U0Z8+MP2OMK9blzV6qi6Pvm/n8b3XCQQ+qKHtXMTy6LiVbr5vWJO3CTGq
B6DjY/ZlY6pt6CDg9hcJk+vKDmcFa0v26MrkjAaY58m84XfAnmZk31D0J4ctPLW7rQDZqZ3B/mxY
kbStDDwIQRlLkUa/Di6vgtV+fXcm37hSli+lgTIzTYIeGzGnQH9B9kQWQZ9Lfl5ix6f88mfE2o8c
5ozx44yKNHMYlpi0F755DxyE1GlEdNSLF+/wG14V1WaUEcku62bALQPcKaFHWK+33qHnX/Mp9TxJ
muUXvl4AjLeIVl5i4sYiXuNidOLibj4hKm4HC7Cdp7JSaskDD3uWYTTTnQ7nS1Kb1+wthIXQsNVd
8exrlhpLBcGQItDgs7frgCwyEfbCJzCoB+DbptNZkZhM9hBeKtLBfhIgr++GnnZYVx9+DW9mRTUg
ujdBW7DwPErH7Dst/WeRId+hNxNyE3mOPMGx+sUsZBw0pHrQY83ze7WQS0C+zG2YsbPbWhgBwQds
RUtrTTLSzjMtSao4XbHAilnrZ+XtLXDPmShxmc/TMRBvjS5Usk//2iESJwVonzWinJBH4gpkq1h9
aSEvSPfeE4Bys2kMa+Eo4bebH4MEL3XzncmqeMTJDfsg91SpxZZUj1BwKHMory+o8cI4jBmsxVWL
ZQQtdQrszQT6Yomz9F495U5rpwXDNgB6N4B6Quuq7viXbvDtXgKzxX/iKXaVtEiesQCtuohH0O4A
QhvBLR20qpYWz7w+IJzseHyuHCBb1UMc+z83XA5zqnpYzq4SZboT/zNiyZqEaXXCr8RPdKaDHIuP
M5lvabanseOLzdTY8xltkdwiSJhJQMq+jlA+++AWHHszTll6EsIX3UhB/o2JMUaPzeFhLDFuDB6+
NzEZSYwCe0YBM1oPyPiNkBEHVLEIm1k5RWSLl2JShIt+XtKz9WHr+AtrRo4Af/SdIB2V4XFheKvP
bnBvZzknex1rI4M0TplHYtcF1PqEHbfnQV5cyC+N9QgbjnOqX82J02lPi3QPUTv1Q401EFJithZb
R1nsTB4kJ/QQzGvqaf6DO65+MDGECbEHPjV/+GDcP5DmOjqYEEaEN9oakVUwETKXhRa5tHQyc//J
SxemIJ1ZWOtK+qrfo6LcJ6Ut9rYpfYTYccQdp5KbmMNbusibvzgjbrTE0y3GmnLAZBC55zLG16N4
U0/ipyoyGqWfjbNOzdn7EGdsJ6CzmrnlPK2q1SpOmSqEUykJfIvU8O3yWSHUvfFOX8TtrMkkXTtf
5PO+vcNWaRhJtCvywYNSnbhxJrULmZnA75HJrMuQ8BElmoFTO7ddmJW3xU7asGDdNHJD1lYdIUhK
1cpzgeMwkABSTxU6YASr91gLJS6K11TnzAVQg2i6xwJwumXSK87m6E83/4A/ft+nya8S5s+O8yzh
zRMQxKGkW/TqSc2CBDvBpJl9bDfhuyeQPWLOk8SUUayIKN378yHVqx+FBNywFBRZUpMdHllwNToB
60aKOdUxVaz007JViXQ+NzrddfJlWQiSFGzHyCbuUx6NLclCPyMzoCjV2LeqbHsUiRVZr4tzUcde
lZALcFdf1mBdwpcYAfOKNsVDBj+mCMFm4fWIa/IJGI1jDSvqOaJOKfHMOmW0LPiHb+wmbTSUmyrz
cJtMXajsbGFo7Xo9VBkPRHA/N/Ufq8t72m8DCJT8lu9cXUG8DqiMZvfzEALY5p2w6lacrspjLUcq
TQtYGdP3qeoYIntDcQOJCACLzNaFF5POvPU+f+7hovtgTSkGrD6rDSSd2Cd+XluoOvrT0Gsn0RrQ
xxfOGpcJdHLZpFGQN9gl0Q2waIodJohIn0AHaIW3GainAO4dBwHZs94P8BAeVef534RljQsTIP8p
hlEepJLelE6/KDucAWwy6sRdTsJ33Gqdp+WxBGE4ShUK4VcsVbzk0dqFRe65PiQ92GiKBJnS8Yef
HxwSHUjX2AEgu5YlJeSyolUc/htkgv+a9GHSBOnUf+7QI72zQsTgFoDi0+eMULdRQBqlpuODU2UC
3uZi3yb+U9qnX9zZcNWi7fUmrctj5FH+Ia8uHluRZ4obAgo5M/xHBN61yevsPw/zO8cGXuS4u3vB
syrT1xXsb3yXqyS4OfedevfTzAqMOLkwGndPeKmDh8K/5Y2TNiE1KY/BxChyPPvbY6qP9MM0K1h+
4UcQ7pctpC9AyVYWcNzf+0VpXEMu4ezEFlCVqzmoMm4ndKv2lcY8Px+FOeES1dn1BoN0T4XsVS52
ekLv4S4CtC9HAu2m11TLMjhcu9TkJ8hjUN822KomGWnWs6VWvVJU3EWAZa8qQRT70HMZsIHCLtLd
Xy43rDOwMHTzqNwrhVwVpNK4beiIbab+KZ45QzE5/a3CDbPg/QGcGMNA1VCRS0ydtSYm2MHf0pBr
xX/4FTRLiBHp2ZkAD1kHqTbzBLq3lc4+MK8V/Sg9riarye9kqargOQ3AX1N4CgZgspvHs/3enApT
L/kMR0K4R5isSaLASNVuYvDJCg3vK4KyqNY06qLCsQucIj9mbMykIU+/gx3DXd3SKeaFFBsUxbO6
NHqZXw6m5EmulhZQxYHlbxQSDcd8RYcS7wjjivIIaparlFrjtAvUz7O2iasA0xjvsRQloRUe2nej
cebeGTqlLyQ1isP65FUHuIEfwQdmPoSgIDn5djX6wgNe5SmTEe5K8SuKckPXuNWSSVD7gWCLm52y
YiNWhTj0WDvUjranxixjcJARlmDWjmbRsvgfS0Pe6AHwPmwf6hnyTRCKAY1nmAyIHWG+jercUkGV
/dol3+9VOpYrnjqudOZmRD4VAliuKJLf8aVy8Y0WTcHi8hG265/I2KsYr9QK3SpYhPppxrJvInIs
clyW0714GXVbBPtx801GSArvDfmFfG2lW5wFRwwy9cwk3D4SItY2ZxaQteIIl6dPQeUVGh5HuFNR
l2XiN8y/15rj5YdIDKfnV6AKkVEgWFlglV/fRMh6P7mMlxAQVjH05zigKVBJuSZGNCQz/aH8/QB1
LmemUOyNnhxCwpp88EeJShzs0ERnhkPpUiAEiu4dGVU3LgRyKBw2JnyoXSQ6dYpxo+iGNVs6XPaZ
lhcMfnuydJ7C44fR5vtZZC866GZtIAFa4o/B6XqekLs/vALHeaSKelErNoy+YqOkVyBlisQ/yVwh
3N+8ICi2sE95M/EeflHtOx6e2MboJxEccMdCZT0DOUxOZpTBmqsfcbCc3nvrhjZEyfAY5bLnC/Lg
1jUHl7DFhpftRYOyRblYD8Mi/VweswL9t8hV3cYOe4hz+XJncghobPzEAiqsXedc5FbDCmQ5IsLc
ICa82c/dvU3KIpS/TWhZYH9NTzswPVcPenABETlaw4zeMsNEBtsGxgAeQYzr8ICOvFCqrLScemQY
cxvV4fbw++A1kNV3rb+pwWlBt+IXS+j8+v2R/nQgYIHeRIe9VoHf9S8Ql9s6FIsRbT9rYKTn2M73
VT0LZpPjy1MGUSQ5GAIPD02P+OaoKRe7MH1GGgFpL+koEhQ2pimiBnXpq5hOH/04AOMRkC5Q5N3J
fci1lFgyUlhhJxkOILEWsoypHCApjjoGwPb6uLFe/PhZTFmlJrv80hk+C+BNa7SSypPpNuDLur8y
K0vETlNuddRZpMMA0eJOcP22au+0RZQssIm9NYZJcbeigAdXycQAtzbt5XOhAmHu4QSZgXZI7CpN
AC2emE++BO2ofrKddqxoriRh8ToXU/GDhANMvqn52mv9MHjQwCJrnWCyfXDB/KUSRA8WcY2Rxm0C
i0MAtkPix6/+GKBkg6e7ea1PBoetvkueR5/1feiig/4wloDeP0ziXIo1zNzqCs7GTDCunbg1Wyaw
JGV6omAx9S97ef1kLf8MIthcP7dF1VXyl1VVJV5KQ1U+ao39SChV6Reg+K0qeais7cukBq15iZ4W
AmjJffTJPTKn0QXKcJzi0BMIKY+EHCYjq6RqfDZDii6QLA2ywBRnvycmUaaY0jUvbsmyf6KSe9Yp
iUXGoPQEqtYd9PGglBkvPjvPaTLIPsePsfLXXU0Lbna+1UKPtf0C/wTyuQouDT+GXyK3UneioXqf
CdVoWr6NVKOlBByEZQfGguoIYmkZpIs/mUViSpeQ0CUTH7NPH2f0JziiFUKybemSTSI60E2xz60x
yYwyaMNF42iHA6nV3qFQQbmu5OpheaUPvcztplmiUF0ftHdq0b73ZwAyBy2cxjL+GG/GYn2z2DLe
OW6Xq/K8n5TrTgqXCWbhPjOTRDzpCgT/eg1mBTDxBxwJgusLhUTK9fVglOrXXLgfefGfKgnvubFd
Ql7CKclV5qLNbLfQnfalgc7mCVxQUfxSOedkYBEK7qK4xeOvBgodajorO7AJxbTvZc72JSWGy8Nk
UG2iyCbasr4nQUEk+csMmyNrl2QHjOFEVB4nSM7noCT0Etw4JXhx5TtUlwtgdD/mGCC5E4osLIe/
s2fMAZ1F0KVCDlfaskEigVQUy5q0F+aUiGYkveBwZu3/U/GWRwlUiGjw7IDoMOvifk0c3IZoVNHs
fpxddzDQNSHMHT6lJGPGh2Y6joNCj0aoWZyUS5rAc7Z9z9xlX0zRAPDgNlMWXQr8dL4PTx8JKYbH
z0gg6WmXBzSGJyuPuso2RVvRmmLPeYUYuIvRjWZhT0Rc5qNLmwt2lSsp9pfCZ/vVZ/kGMhpwfGYn
MPoITGM2DdmbFcsfOgDmtXS8sYRAID13lZFP++8dkdrmfYm9nZwcYGjw2Mn08s2foUGO6vCL7fDq
ZAsT8DT+4IRVQEalMk855005DEVyRHGkeMXCxLusAquwIN4CjeOWuYXmyCOMM08Y6EdGkm3hfcvA
o6jz2HPGjj4cvmYrsbTscgQTwjhl4FzQIgO/KS/eULNmxR5DEsUPPUoy+Lx7p5czHc2XAXX1TTcZ
LpeNRCpISkm2N1vho2Mzy7CVFhwVNL8uu4ce74dxCplaT0cXdKLLqw14Mq3pWSS+pJkE3jFgddTh
+UGXLP/9PuRQ9ZEzZf06zIuzhZvc9mnApe49oHsZYXkyCTJuuJKL+MUZTmHDkhPWcvq1fACyPVjM
DSpM/AIS2jb1BKfiCGXg/izwG474JhfLBK066A9oz7hWhuVUXKYfLpXWjIfvi+iNAdFvnoCZ1X9K
GTEEG4hSy0KtRe5wLtxpRbM0CD1cDf55EvCIaBsojiJSamkCh4LCWyHt0eXZnMs0OrFWhjnWJWnk
WBkslEFnuXmbgKoOxMjQw9MdWkfS24s1x7o2mGQ+83UkzSd0I6cH+w41rbk2ynHAQPhB9x4QX6fY
U+aJpWG7A2f/xSFER90Hx605ROFIl36NgeOAdu8sfnF1rKJ7F3lKCWU5hQNzhQ9Qmk7xrICIZ0L6
8+wOV6oWVNEg7FbJDEGgncd7+V+BlnU1ps5HWSYMQJ6xqqNOBJZRChLCm20iocqWFp/uYJ28w/ex
F0yW1/tFmz15nmhG5GTrlF+3uF4wg1k/8IW1gB0ljYPX+z67/wD3tuF8TdhISgYprGQWqP9hYZfV
6aGRM4eIKRL3sVU2ldrl7drNotSFWFPePAm5WaiDQDwZ18yHSdYPacGCvozDKfxTunvai1tpdwJd
27v1KWEkOXdEwvqTQOGRyYbruNGnUn7z791hzNUrzIY1fwIIaAdj1qCQORVxO9KiVfN1z5Rprv8a
VLzmivRIADVHdQTr3Jq6pVuJYYTE17/JJxpmsaC/jbW422+wOhiBg2rCpTPPLnkbKyy3Q29jOtFW
eS/5S9xZrRyu7EzmwctYZicd+dIKuvBJST/Fdcu+J96EONBBhaS6bQU4e2kFAMwhm6MuBFDIsZET
MlWo8P8GdtRYFwn32bS0KDt/U1/ki0NfgoRHttyv14Twh7Wxy8VnYFmvO1inrSoZgH3KNrq+Q5Ov
8e/5BINagahqbndz9DMPwtUIg55XEZCYsuo6iIK6QPSFpqKYM6yMBEDoei6ifJ2C+2dnKw3Ffcnl
NdbS5FBU06Ac/nIzeH3OZjycWm/oEdoo8wm5M92kEMsLOl3Rxc693jR0jmF/CRG+4uP+qGJo0sCn
aX24dF3l3FTzo7JqwlgsEU1biR7bNrUw0RsSCioUr5M4NqRYqMqPC7ak3Zf0vINt3IUOtff2JV4l
/6/De1eF0rPiwyRN02foUrdNbFkoh6fV+hdDBWLj+w61ZkH3PQv7oryfZUp4Zt77SEvn9pUiSwgj
/PrUS+PLfmQKXfeFrb746G4fNmAs/CJoqS6hDiCWSQV795b//96Q2qinOtJeQ4wOc+SrAUC6lf1L
NqVylF1XzW7nO3uLauelv2jo++WOSnNc3U8V6sOkLpRO2ZfPLJlaMerAUp/VdrsnLy7Qoob9w2n8
4tnidcyVOhl5k21PyyEJ+x+v0ca+ET5m32GjGUnqRGx9UWuLCLbth+WHdxFSmp91bBrrXCBbjHhR
crwqtd7IEdEfkuv9qbTJuf3lwXWp6O1aZC/MtBtL7zFJ7iCT7HbGsdT0jpRMnDNKkRHXpwPfJBJK
Ozb3NhMbfGz6gRXWz67tX2wCUJT0Kd1bVwLmaM+1Qt5KwisDdpjA6DWAMs+PTK6mKIbqwOKWXFil
dswGe6A63UgKRiDMmjuiKK57aD4QH3aMlLjyqeuurh3UML3ZDVvG5mlgJ4JmRCcJZhjiS3vsFLLk
WifXbL7dLwvnMo1HcIwvIqsWBdccvaXxuEfz+qdvjAgyN0xOh6laJigPkxanKPhuCbBx47N+ymHX
9Z9+n7/nQKGoQ5NMWN7WhoXVNYU5Ddi5BBBWbIrDkTUxCy5R2IoCt8Znx1Yp1T7ECq9AaUfEWB54
bgFj6eB0bv1VFr+ftHvX7SiyVz4bR3ymgFt18Qs9Yp9+iJGm0gw0J16fT8OImXcX1MF+F3de7lKH
XRVLm+n7xf6jumwyUizS8woCxijtoGdYqy+I0WGyH832FRpafeDOPCThagC1GYuZBhLaVmWavK7Q
eXmnNdauftf5pv3H3AyHYPDCiMSAoP5VevsKwGyF3UazXc7955RqMaSJktWVyTOcXqVf9laGccPH
njcOqBpnW4/mdriORAXfHmQ5pqrDiqWR2xZfH5u1bR4WNifdWjQXEP1dMkrQS6X5aGhU1lTmktfU
/B2q84xIZa68FdUR8D4XN5EjUyDl8sXo/M+NpWNI5TXdW78iKEgAVhBDcXxsNtXV8/q2Vt4UT6uz
aA+/fhYxBU8v5xvmXYyZklIHbbBs+ZZG0/lJm7hwH2QSGrHGCw/Ac11IVH1S1gu5o23q7ENxvSv4
A8wD0pkkIAj2peBhW9tL4X/QLEuFyAhTdfOPuHdVL6F7V1GGXHEVUidx9U8OIUFI10AY8geacZFP
mOIK5vvF5GvJXtVw2y2fEVaxHTI4VDKDvlY6/8dxjXkPp9/7plM9NxVqLFuBbZ4nre90mNrqFe7o
nhvwmObSnbzzNllg0hVaL1IW87h0ak4wiwSCVvlVvbwsZ+xz06eunTGk7psvVRCJR4jzEebpq4+A
O2+kFuZCPFqMJzcHYcu3kkr8nGNlSc0yva2R/MFrJHRzi8kee8YKTT0PZ17urE8LtWUCjpuC6MoH
ZLzFKcwR9xgbAXJzcDhHC5mrDUczcWR9AbTjGrc0P8PRbzjFX1cJVx/g6JuyAxdt/l9Qfhvnjtcc
AVEWwv4ewF785/t46GgT97MYvvu/9l2VmD4YeoLdVRAfYNhtTcM3xuv5SYmW7Coz6PIpiq6sIZzQ
mEu5waldxtjk92LwB/2A4ktpwaDZd6TkaxXHn1dZLVqCRxNafD4wVhvUMfskG63PhfsGMDlYqA6G
kH+SFxfiB2He5GfiK6cc3BekboY1h86G2FSp+ohKg3GvgFbtRFJdnvkrlfhcvZH4Pn4YqejHHYy0
NtETcnqKrDa4E5sGnAPJCUwm28ayZA2gJn+iH8mZ3LNLVl5DKS0GPG4pM6VixwqXUUKByA2sLAY8
xqNVBhqze9pE0WfURh/c5XiHi8aJkt3yn6qwjTYzH1feugVAXEK4k3TaAo8tT77mwz5W2CnuUrMx
zU2cHU/jAbbc9Y/xOYmQuhSe66STFgUDGBMKr5zdPjGts4MAcfS7gU6hNyA55rvFNL+WDi4kB4OQ
ZO0HG5PoBTorr55JpEp2xfV8OFzhgSj/iwWeoUlkyFlofe30+8fBG1/Xx8oIQG5c9DWWJMRUPjRp
8oc9639oHliht1xTfBV3jpv9/yAAIIClB7roG3YzP+3V00ayGyyWq9y+mNepcqBhBvc8X5Vqa6lx
rAc4TmrI3Vk2OfFjpQr4XUJweSfSLgWrP2kq6KDvYoyC9qD+pwwIykZGUWlLVi+9iMaD1yyPaT2f
lJEoajxajRQUHZQNgMin8JVK7mP0prNwnvB3qdn1jlT68xZcQ4GlZMJfbQcik0679Bl2vGsYIdsY
xP8MnkhJ45pIwHP8kgv9msZdBpcYG5OtOdv5Ol1egn13ws4pnd5b+RubNNVxVYz2fPV+1PkANdHQ
JolOF+RkRRVkz8Dji6r4VHt3HWdiWMHvxO10Uf18Yv6Txet44CMqw7vIZ1H/WGyRYRSwAdMvMrEf
ysakK+WtTx3Q5wf2VaWaMwxIW2nXAdYu9mAnDueIJg9s6aEFoMyDGsvPpvU64128U0lJmAybtpXb
FDcKeQrp7guJpM56ZUSiTkePgmPSe0AbNfd6aq6xy1H7VBQbwyGsYTACmdyxqpnamIj6JBaWWM4Z
I7eq6wopjPoGgLNLAzFZpn/IdJSJ1+jQH4fNvHxjn4HEOSL+KjdXu0Wzl2uRZzPZS2B51vhPWtd3
T3GeFheoSpVxJhT5igfnO3TO6s6qt0aH6dRvGIgbeA1Xc6OsPqbxPtF1ioCr5DWbIel5gruIS6q/
89RLK9eClCfqscnbBF8By+//zhlcCWoe7WE02rHY6N0kemwNWuY8QJiDkyErWDkn94FedA7IdAeI
lOjzsG7mniEfdqcr4H07ypZhMMuH3OU1k7J8NOEGc5bojyuhhseLNa56VR2GHuKvosX5Pr+d2ZmK
EGagoyv4tJ1pXbYFMYE1Eldsk62n82BcihxjcDgs6etcOwtozJ7pRLL436v0tf1hPtdeA3VZbpa2
coUijdi3cIHunKzV+PeT+KuG5cOGNDFczqbpy0oFf4CzroMlwMNn4MIJ7KlFBvSM8qgjP0cQ4ZJU
GjluoNrLqBgNfo7d7XHe4Kwtt//y+q4KkHVUtITAT8Vlk8ihsSMeHfnH0rb347Gp/e74w9O0SbXX
pps04rNmwWtCC+dJuW/ZWWpp3jIRwN0PBrQM6Xt9Xo3Es+JoJ7pevNBonIwlGoU/gnKQmnK1jd2b
xISEVPPK7Uj7EUoNye3y5xOKaezd+JMWsPIuR1moOzRrLnjN2psKVgosNlpIR3h5pkLDl6+uBgDv
pubvmUbV+JYGLn+wu+uo2+UnhGLfAG2Q7Xz7RhPsugT886pfohsV2b2BguMxPb8xEQtYSDtGCPl+
9CE29yLoIsr9mSl9gBkn1MiXY9Aq8yoreWB0d/2gb9+dYdzmImIbrGOuiWw/SgDc5aEQY3gpWLP6
rQ6tIfRXraw9kYCIyzxNQzVRdlK+hPIKJ6afIk30lnU+/LKMbJAKJDDM/yhSkC4u4xwE2E7qdPAl
7U2L9pbhm4ej3/9R2tlJNmqO9Fz7cjNWVx1DoOVMr0jZE9Xmv95yn0zVrul7WpPULhiHsR/iPKjm
GdkYo96LrB5+I5iWUPe3GRrY02HjLJh1W5xEIjbYdPtOM0b2VHVt/dmultzf9hJMxhPTwQ/Z4un5
m7WTRETK/TfQbtYBxUBth2s+xbi5xikMASgG0fIqQ8GUmu009pCIm2ayfK3omEco8SBWsbAGfsT7
qSWvfViwwexXzkffZ8znFSvXATgwlVuZYWEWS6jVmDHqlrcITWrCZVmh8U6STF/MhFLrnKcRpwXC
DdBw7oH0wmY8I9tus3DjyzFc5JahpnfqQZDxplFX68B+q8HU14H6qGxvERIOsioNwr9m5cXo+PNV
LHsBCy3bCLzAv1q4s0UzmkVgXyLFkkkRhTW7XBSbky02vsBcBgibhLeG93pdTiDcngmPUZDE9cT2
enZ9kB7y8IlVfsDJW0KJVvovyMsU/2sTgZkq+AbCqUDjUY1a8ZR4JSCfe4LNG70JZWqa9r3F1MeM
JNN4Q3KV47giQyJ5DRFoLNLfZvnxkLNqfdUT79CnVX9v471WXMttET7xDtdXpipHFnQ47nkjKPf2
h7CdV+RiSFZ0YSoWXd/xOhjmxocn3g4JwWp5qlCaHHEoQONI2a9ziFgswfiw9t9lAYasiNvC/LCw
J+p3zE1dP1pJ1BIML+XePraLURKi+AqAksthLx4mtkE5Bk1K4xHhNWflhzwoxiH29OOc3sf/+rzb
zmffgyZpEShxlIw6r2+kKRCSS35jM+/1CXiGF2pDP3P0zVxOqCXg+/GI4AEinO/yN7trWMQbXlvc
U4ubpxjsUSWLK1Gx2qg0He61dzs0/7xfdT+pcZ1L1DRTq6N3hL5PdsY8tOHUn2i5KjIPgxjm8Rgb
6JJsKAReW/c22xzPR4j+fAtoI83PtG7xs7cKAWyf8VHMHQSdLz2afu71OabtP/nksIwBgKN+YGkY
SMXyW7eTTSsADTDRpyhVrvS1AClUuVrTv5O3utwd9+UwplR4dqPC9brPpd7/CbcU2lo+BNp70byS
ptbsU+XIG6p5ovWh8VZw49U6YW/kHjlXjpV7hDaWVWRWCXOC/U6bCy6LfBhB74RrN9E4kmR+Nt5w
H2Eig8j0mg5pO34sPS67VpL9lI9hQDdwRqPoqw3yimXLtxnpyMDNVquLaY4ezxHX2LBwazEAANcG
l0wLEgLITmpMLoZwhPrG30+pHRbz6P98hsUvLnTnpNaTLZ+Xn7pBQO5tOsiRwbdjM218QuZi7IDQ
sCAyIOJspApenWu9Sgg/cWCj87Hsw+a4DYU+Bd4r1CV4k6g3ubuvuBwzsrXxo12SuR3pHBX96j6d
78WV3SCIzAgvEkB8XcBe6KQALulTJpGiA+0V5dYoaxkBpmWxZs9/R9DhZaVSsuYM52YpCn9aL14v
htZ6c06qc7q/W8drK50YIPxFQzMRx/wK+PdiCAnN891t+5PLpJC4u+5tbb+2YED7boZ19W3uPaDD
GLO0ZULjegRUlg843cLxGwPDfJSjGjNBGIsbQLOlU8W2ulsQjeb8xqfeTRTG8HmWgOjcjtKL4MRX
d4ttec65lBqA8peDG38mE1DHi/95ofHXQCFbg03OXH35KjuiJJgtaUXAPoRt/3EuAYU6ehjPJem6
9IEiXQDS5ciD9IvfTR4rDsH6z/HhX7z1ab5usoLFwQlO5Ow4Dnij4sbosTESC1CNriiKcBj20s5F
vKtio6+Nilu2U5X+2WWoFpMvzP6CCtFoTj1Ii3pjK3GpnkKOKQJk3NcqLJvLZ0js8Vh/aAa+oQJ/
WfNE/Rt2yhteae/Yy+64iD1c2bvp/yMEN7JvTD0vcFWPgMJHYDlCM2Y9ndXwTeZ9strC/ypHOhBr
6G7x+08uspMGr/Bg4gtd21unhuQ0VMzsYhDcDTPbDi35A4OJva61j3PKhDT31rBbgti+ExylGWlU
1FRFkAo9GP3KF6KHc0n3eor0SNwGOLdSycVGSzyjf/eJSC+jGBdH6PC5gtfhSNlRY/5NxqhO64uE
dg2Yh9fkWXwMk41nsv41Rlr7oDIoWqzcRMBiyHEZaiI/hcF2etwdKacPmJpi+BGuSDo2UBpOGusk
n7mj8OgqWO06BSLwdob+onIDHGe178uAzNgBwoj+pOM8BWqSIy9OQZyJuK2/qI9oZA/A9o1fi788
3uqy999jWJY3Nguap0HgHFnx/rBjrGqNlc7NQgrQdZ8gW+WgvZv0DRo4g2UNSw2iPBqV9uOw6XBU
bg1OgJtsgZGK9T5FdvTRePL8XRC9uPOqB5sJBGBlExDI/j4LuxFPfntmqxx8LvX5PB9XR03nd/XU
12Zc7eIU52xF61zKUEXZYINioGOidlFllAHGju6wCua4utaBsm6/iFTAaUElH+BY2eU0LVrdyefd
jbpjEjDsZD/dqixvdoCO+PCzujJpWOrjwZHwVqTByFPv13xJMlSMj2Pju2Ws5jf5maCRI2/6x3rn
bnNufNMGWnf+2FVz4pRGbpXvyUERp2FIHFMnIFff7Z1VkQTCzkFGMV4YPRfjnyl0XaBxERyO5Vxl
cUsPEzwxtuVEOHR/5jy5D+54VuJakwwxl21my8YksNd8Sigh5B2m/Y5omf0aOGMVQUnE8NRAGJPg
74g61Oe3lb8IE9Ntyo/BMEMJimiEZqJKxKOYoc5ZBhudEVDdDf5Sk4r8IJcoRAWJzmHb7SLw478N
WJTwHnHlUYa0I/5VeIB143Oh8gAxlOU9tk/y2JPBat+IESm+Bo18LURvmSi01e9QcmNLJ5MUbABs
CZ+KqPflp2Y6T9ASkPSh+xcjX+EJ7rXgPe9R1pW7Y9bUMviK8TGYqC34aceB67koDA/vzo6c0t+A
0VJz1gk4r0LGWQJJOEjC5/DVZ/FzMwKySbv6lm1xUl0rRO5AHYsXphPvqqMA4lJ6i5N7M7YWNe3U
HS4Ke3g8D+7P+icdAo6wV05N72UE0JgSolu37upKSxz9Wmkie4UBCB6QikbxI9qkyL6Ls3B7LMoR
IrlnaAPx6tgSg9v498GQYcoEondKZf4SnUDCEV4H3St64/tD8YoOaaD+AqteniGuO5v4RwLOX35a
oGH2YHvkb0i2izbS0rT2ggP1YlYzj5DkH1xJUA/41IKZVG0uaWIBw4d+AbQsNaaDBbGeArrrRqH+
ajtDdOmDgsjh9PTrVrdzHpoARp1+YZoEUzLp7mp+ayBFfdRlyd8sjmranF8BCIcAInFgitM3/vmw
ZEcNQuHNHjTURIyN9FHjopmR5B9w6dRLUzpNHPRM2YwFJ3V/sAioiWugRAhSiZSMbLFNRNBytBtR
43Nf4JNSMDVcBF9R+tEf9EtRrA6qjq0chI3e/fuEJ1eh0J+g0H7uM61HLaitJrqFTYExPWByGEDQ
CGYltwbAWBsjrVXl9SskE2ObAKAgepQgOePDbTeHVMlweuINxpwodV/lDDVtHxE0lf1JPJRU0p/3
8qopVl96JFmVh+QvzXbeYGPUICCR6PU2K3Lw2OgBdbIbbB6JnOTpk88zMtfUZIURbCrYF0fcYzGb
xMAJWSEHjmcnCIF/jU1VK8P/U5uTp6SvEE5/dDxDN9XaJSV+WcS2IRiDr7GtEkbcgJP+nOiXFTTR
yvA4Rcnt7wYqU7UNbMl+1xstNbvcYbhnrgtpzUCNE8DIbQFJqrzrF40UhXE50nqmahT+0ak1NUnP
w7CbG/jddmwnus81xaOAf7T2OiRddPVuvUG+hIjQXL/H3JyM9GeSwW/q1y+eh2nsWVYF5lqvjpQX
AftNsB5kCCYd6DHVX+BIYTRRX0bChGZax2UJ43kwBIOPsIo182TE0Fb+2Kn+8clhhIRw/E669eMo
fZjI5vmwSUHgpbAXWbd2EDDpRMm1y0x2FjOU5qAc78ANDjfX6/MWmBzpkMXStnUTX9J8GmMz6jbe
anYP/2Iurvf2CwUCAlbPOGFgiJA4tXuieonkZuPXhwOvdFyKmoAOAAF2+qemP5IivoPNhy7m/V/J
SasDrVwLc2mmB3P2l6dvAeTdQfZ47oDS2UkZB+6M21NX7RIJs5ryRa54TnZgFonlerL+z/B/gxpS
HEf4ONZDODPcaLivhovXPNQv8pKZXEjlJ7D3w054WhvGB34J5J+hhhxCp4W7Nw+Qekcu9j26byxg
OKg/DfpDfNUT+xmZDK7M5v9rwE4v1y6SNe/KmzmiebRnuumjzakDh6r70z4fZUn05r7UJKU6CrcK
XMQ8mPeyEUtS8mJpNxJxe1DVhUsMlI31rka8fc1TPephxe5wzQ9YyHSpUoIcKvyOtXIU23VEoWKQ
u9CwNb3hwkvPiY+iQLV4KfX2mxxPVN1M06COeIVUmsimLDnYX3btHTzKDJH68Rmqbh7ce6TQHmjt
zM6Bg1V7KSImPFotNS/cvwrB0Si0RX80DeTN1349difHDvHTlwry/YKrKukAhGwdSjevC+VyDnGo
MS69b91KjU4xFgZsMH/pSbKozaKVzQ70TGUJgnNJhz0beMEn0r8JAnD9Eoss81KS6j0IolyrCPmD
BxlbUGHl8CYByLYfYUReIiZKTjPJ4h6I+RzHWh4eCEmxQ5RXvJGpfjqTsAlyJo9zBaEg+8QSVN/Y
ntht/WgqFO0zJPkbj7o8iHmt6NkXg2Ro2i6BMaLxGETENwsz61IJFUXIM/h26+f42D3qsA9gPCxr
KW0CfkgpDfqjfkd9r94h4RTWc+6BpRdZMAMvnRSN1FhCd2zZX4yPKwfvZeRZ7orrsea64vFzM/xA
ikG9DulxX5nFsCZVW+DchuqL6cj2ShIrzKjx1HxvwvpochXWrJqH0it/Os9VT3smHMpKxmn5Lw2h
2AqrSKbnz3ZarL5YBYhw2p3rZqQjpdn0IWn8+EnSzdI4Wws5yJljjLIxRE1IagZY791B6dASuuAV
AIp8HR4iMcl0UCjqpL1IOEZAiQD8eu4KyNDXzzeb/xVhA9BFqqnQgXGz0uRyOMjHm8Kni4WIkiPt
RCQFqDq5sUhRlo+j9MX/dNxMXd9umRFLqhpwcH4Z8krWsx+1Hsm6SIM5slMxMTb/xATZO6y1cd22
OBvzvng0QKfn28/GVHwwioDxOD2jYx5hs8LeRGlPvKeTlb/1aHILLci5LY+yyWNJDtyMccsBgB0m
DJy5hbSNoji/kOY+Fuv8AZ7Ywef4xGpEAAjYw0Uv9VhzNj846Zg5pPMLV2nTD3DBOoiik/YezJJ4
1KOI6+q/rKbc2dDxzJ5/h1SrLGCTvjVsfzgVPlPxBpQG2VsYmikoXxiVC7sBo2Yr3pWvJS59cywo
CSlX4LvrY0UXziAQuohdPcMQLA0/whsBkuUOWSEGkpZCRgDCweIJv+ERfbaiVTcNWddi74f0sAMg
zuL6+PRPegJlGfjMbAThdMKuhSAyTbFUNKROJt06+XGUlg/iaXC+Plkxn05MgEbfPolNPjLNlCfh
u5oiN83SoXJ8nsmzEqETqvADqbm4MHf3a/VbJa184nN7NlCulkSa1zJRJrO0HIy6oeTxrlGpwZ9A
e/8gV7/2s6gPRvHzQ6EyP1tPpbc9rHDO6cuetGhQChyiSMVIxTj1Uwi40lgxr6r8/q6AOGOImf/5
9fjAOQnGPzk+FE5NR5UJrRZRDfpCsOPVN1FF/xjod6EwsECJpz59fO0+kfDxMzb2io5vGy65hcOH
ShBo1HFNrqgeC+xDqMpCMVh/3ju4YgBuQXpsw48fTj9eoG0j/q5Y1hwWMNclhpKIejLlID/3+PeL
O9CKZ15DdHovR0jz+jEOIGG51k0npnOt2zuHNm2AX5pRmAqDIwqcOL1OLtLftzB8vXOmk8ytSsQw
AHExkINE5+pqLMYVwCB4kbI0q7PnjHUG28WNHpZLPxKbN5DHU81N8mxFt5qw4N4SLswiceiDKNPH
AFI7jOVeOF26qztMSu3IYA/UJmdQaR4VNAJWPwlg8Npn1Xzbchgq3vGum75jQR1mt2e20GHGmQKC
ryLDGtKIQM3rvd0p8TeibgFbx2GwXG3B8e4WmvZuReV+pZPONWOXNVM82DCcw2NCDFdjn7UCNnIG
nRtXqU1sAESM8bOISTtInizuti7b02/Mtzrg+LsbzJBdEx019vqK7odmYGjMsYl7Tp0XoP6NYVwN
N3ZAaC0ZuQNm6Be1M116uULXQ3+Yr0qC6brYV7LjWrZAFme9aCTvSTpjUBY/Nh0kWA1EQwSkF/6f
WRt+u+b/7dFCUIYh3haRkSlg0dxgLMj3jv8XZni+0n+ua8pQnFlOhC0BJCm/eWZg2j1KWBs0vxcn
BwqRBjHxJIdJCLVccLn6N0G5tNDadtbaJ8c2j2/9anH74ehCfG8W3LxS+VMct3rmUOp+egvCiaBu
FxJwxRzGaagTf9j3xglTE0G8LU4Z0tLL6GvHjq4lubpXcSm07pR+mgKvar25YUHrTWnJkTuHnR9d
688KKSrQwGjy4kx+wcbteiM4Z5Mhyrf27lJWajncB+Zoc+FnB0gWjEWlvy0CCCz1Ng8n9JYMIZ9l
6cH29bFLkDmzrSSReSH0z9H35B4lKbwNc9jcAGGZ1N11gQUUltzCrNYb+j7tRoaasa45IQ1gCueI
QlO9RnhmxYVpbhwy7lxgMYdzfL4zvpJ0vcliii3MEUB6wKNtSccMlKqkEAnuBP1n/tq6q2NkZ7SE
6aojF5GIDhB1naydpcf6Ipr74dWQy95Hb0mDhi0InjEIr2k79G7xTmV7Vjc26rQ1Q12N2agf2ca7
0Xvj+8gPZ2Jlv9dxzL4zokb9kq1xluVvPwL1M1NZiAFbbsG/ytFzblsy3OYViD9bmfuhNkLbGG8H
Yh8iOF2/DZRA63GfAcIs3gaRmr/hbgwj2jKkGERpbG4+BUBz2cnZ+xrR7msvVSHh/GoqPRp7V+8R
h7nb3ndvnzYIEg/etUELVU65Tr2112o8bMvhNc3ZMHECr67ICq7wUehvrn5DiZC8JwhTT9jHT1VF
fEpSyahOSrJ9mBwPAJ4+yM9AtqLe5G5HrJeBOf2xHUYGovJzJuvsiwrOkYy3PdobIVTIGYDwsfDz
b6bOQuTi57/I+jsn/dQI7+rNcHUcQ3ZdKm5Za71HtRDXHRf6sHNPsAOeMujrnBSoyho22bu3HWDo
h+DPjRY2hZnSvNLEf3yL/lmZnzpSIzX2iHLZrCSjZIIXnET83KW5KFXPMmrL1dGPHRMN9Mu4Srb/
3tSoN1ioOZzubYXvpKwEojgvS3RLq73IBgQksD33IkD9gTl52M3pqaczvGvU3fK3VjXkiZMx6eE1
8zQbzi4UY4r0/QUIhuHH1HWMgAyQnIJ49XvlAXAdZDchl1X5leN+XuYF/4tmLV65qgJx10C/r9dC
zoxyjxkY7LQ21poSAFc0plytcz6d3VTEWYpmZt7SVyahyyx4c5vmj3cjMXSDRyKHJM6AAiGh274S
cDZuGhkxySrv5vyWDnFV2/71BumvaZRQ+YvlMLgC5zNO3HdDBiaJCkfJsldqZScmEphKc4UQ/Twh
/09jnxhm0QCEj/8UCetcL2+r5V9uwNyFgHqmMo4+jyd0MzjSujb6NZPw3n2UBCFvW1YRqu+aFQup
e9HWEc3cB3FltQZmhEThZRENfOezLwL48pchjN4B2ECDChtNOPYahKIpHC3Wg5CZtCIMVPyd2H7I
fSM1w8xtadxBHuwmCEWpirQNvbRnvpeadwl/o0994KzO6SAS5H193vTAwKWkQfJGO8eXnOCdgXNK
Y3Gi1Yo/2AYR5nSIvIsbU/ApH1QOjg/5LkIouN0ZUx5veI8LO9vhWQzR2HFaOo+FpO7VsXTLPtj7
/gYd9Iu6uo2PtaB8bF/vFGYTp0LJsdW6DAf1TqYeBJQGROyV3J9t6uPkDockliH3BPUZFyGguNda
0ceLJAcKQaq6gsKXtTRyNnRmCP1oszYsf3qOxCc80F0hbN1sXMrInLIeTdCBS8HYaAj0m0iG/Ith
sxwZBqAUOebCmKGj8AWR7uwFaxfMl6MS7UcMtxEZMCg7l9hLVPkgGFM9kFGh/KImkoamL7CavFIz
BwS+EFZU/Kffrl9ukTf6A0dmEtc3+CrV1WBTYJQUyZ5ZWOvaogZRXlYfDWnHCvXKpTivHlfXr54z
IEbNV+OdDPdSoPD6m/6fD2ttZOGnyg/XpIueQvx3lLgctiDhhhfd9HbPiaRdedbnJk7HBXCL6CuE
N1JyMSH+NwT7BbFFwZwknVewrHienZF77HpZPOhAm8DRKlqbZPqHRY4B/l4oWqhqqgASx/Ct9jno
cG6Rrc2zII4qQwpg/m8Yz60CuQ8dFwPsxagFt633tlPqcaicDq0CvPfR3UA7PMe1XfeqruRIoacL
x4JadpIcmIbggJoTPpNmb4TuVTQ810SrnRKDtkpfetJNEkEkYlg54k/MQA4C86/jAiBhTe/Dg640
47J4cIfy7sP5Ex22sb8D2fpH0A06IcUs4EqiMBL4tsfy0zv1LhrtHz20CJyxFClxg30UqTcliBhS
GtW+RIw46fy7k9pHw5hYCuzhygK7Sd/Vu2G7k3LoficKwAOdeVwq0bSIVWPiIdHZZt9pLqYcO3Ay
OPAvRzyGQN9/E9j8MkvF0NQtuZzSiHjbITSROUADpg5pN9ZBUeUE+3D9dycDMpj6jdsPT3Ox4AW8
Wtp4Znwqfj+9hNTpFz401FOEvpP9cp4lLIL9Mgy2wHHEz5sMyv9/hulCoCW08Bl+9fubKkqwzvDg
hVId1Fi/j90/eXJJq9WPaIUMkZoIDOX24k5NWTqkboqpnqmYGUNN1eISjMpVeCC5g0DO7yVp/RAl
68i6VsSHRe75sMVTR8aV7/3uM0QSFVpA5bSW0OrjA8kBO/okQhNzOCxec2tzmm/LwUVMVHbRuZn5
6YyYMymXHeSIJQXO+SwuEt7F3dmKVMHl9AKhIyzpDKO9cukM7moLTt4qROvCMveUt0UF+lLGABoQ
DDS4LlE/oyGKZJS44k1V5Uj8a98KdqUSix221ssusi1lIKNc2MHvU1JHUVTI4qRAkiosz5g4U9yx
pcNXTgLeATVCa9OeFvt8psgQkxMPOCvmaH0us0Uvskqrr24tsT48ERIQ5HAxIpJNg6u4y0m4bc8U
uw7gBoZIo+Wbb85XiWRtODM9vPfkxVjb46bw4pcIR+ffGB0jAcQyJOIMLvI3Ktj7ja6FsETc1YOp
kH8ILRICkx9f48uUti5k9cVn+2I6XhEAYxSJ06V+wOP2SYTU5nmQB7icVqmxr88uBcGuCiTeWeA6
hZOtrBPVCi/Ln6agZvZ0pMcC26mFCuw9gfEv6j8EWBHpEDJWoDCfHRXKOregPsNyVqLf78KaMDF/
N97NNfF1wC3y1LA10+4XqcCcLP6/akLctFVgV6gG/zjpyTGcxVHMFEBiFNk4uAPNBly0ThBu43E3
kN+FUB2tHizOGHV2iqqKVs1R85n5ZqLDf8D0I/knAUhH8DFfvWVp4xrYrKMhlrs7bt1t+xVOjYZr
2Fyp0GuWQHfhNUU30SD5EKg/ZEdX4VWG7iKZ2vEzhfWwppelsrOSUqVy4e2okfOcInzFGRFwr0Pd
AuuWz4tKMh1LxahyBzJawvt6ylKt1HxbXr+RJPcLA4Qegva5vPP7swJk8frTBJI2Eb+n5pOCA1SM
Tm+chSP+s25/Fa3wzCSEm76I+cFInLv1JzFjZHfc9DHQd4kWO9ZyQCXePpQs1LEfh4G+quVCiX7b
BFxZsDWLo7Np7bgovwVfJCAR+M2U+WEdLe7b8gl+gwaLd3sG7uxDaFugfqSDBQkAmTlcjRjKDJmD
akNAuYilSLzb83wRlbc0ptf+q6ul61pARNlJpiGyA1eMW/Fis4lTlR7RawqpPAe7t+nPeSo5KMRF
1Nhwiv/C5vghof1ck0lhHVxP7sbEyAlvZK5ORbOCmxdwBfp9J7+wQQKOr8tti3fj9wk08pTy3T8+
HKJJEK3vniyMtfJ891ouwozTb2duskQy9m4tbgk16Y9M+GkI97nQQtclbZK/iKRWxTf8AuDvPRLC
aA2ftpWBdNNlAqYvBET0JKlDVP6ywSxpYXLtNd77EtNDsEFU7KvDoG3N8z/Cq3wexmWIkgHBTNUe
FGQaqDrBUJioooWf29h/GCrN0q8lN3c8eQgwJ6n2S6ruRlbh6t4BEdFs5AVYvKnMsMYxEJ8Ajzj6
IHFknbyeXmA0BtKBzdzGdt5XQmIyyiW2NcB9dVeQPTU5l7Ghj3HV70Sj9nthDe9I7R9pmbNx8RYv
aSF1LmoJyp17Hpf8ycalENPUsmvKV1vJ05xgaj77pDiWheF84xFVXTgSOgpYR5cfKHefRXI8qYfN
Ieyp0X2hSCZegxpN1ML4w29ZTpJnbJTSDQibUIXlo3Fx1hmTMi55hNwsuEVVc8OFiZrl0BKiykuO
VM4SL5qdgttdMVbXZJS/TkfL2q4EUDIi124H1Y5yPa15P+DJ+mplvKGjlAlI/ihIot1hPjC9anSn
ocIcS99OOQBmPBAXfS+lvrkFDbpDbl+Bfd/mIzpAP1NwdOZGQNG4wF1g42HAIwmXFN/OeVeXFdZu
Bx2qMw8MoiRKR84QPaiTUFKmLQYNOhJRgsRWEqKidkqHR1RzoiKdik7DSycI9w7Pni3Tds0zUl4m
uDHM4cYRWvNnpQjeRseyWUr0Wg4w/F7tmVkYS40q1GYn/uMQ9K1EShY7B93a6rn4wocxGi2k7xdC
IVzlcgno84C4PMm8YtiDHDz1lKv7braEBuqDGyMHm95lt91zBsUOxEQHoAm8iz+11vdzi+4AYU/Q
5uyBhcN40Yh7iauWS3CdVxQR9OQs9skzsqf8iXmYAXYNWs6VvUB/3loKtPFB8x6NhNCVlvyvuwXS
yNKMalW2hQyyVSIUoQZONd1jLX+jhrwvGUbA8Q3t0AX3Mmoz6IKBz/M8LKWNo2YsVVLVrLWnuIpP
mvEGrkHxe5O2J6fwEBKaYOv78rFNvASYvuWHeas2dFQcPMe0XTUm2E57YEOrUPk5TIycsn9Ttfju
lU8mUdjaa+qQw3LVeuN6RYP7FVG89Mx4gEkSw4m+FWb6yXZY/MhT8sbHP+O+iABNuhiEbEf7mhHl
HiaOj3y4IR90H0VpJaXJjLtRc3duilTBMOLydsSB4fT3QXEbaoL7lQ6aqosyPLbk7RfuICHy5fJD
p/RVZMAipKAVhFlFJQG55b7TfLpTBh8bhlDh4q5fCkh4fRiACxNMB0P/42etvH2b9ano8nO5e/mx
4cqjmiRdAwZKVnxOZZY69uN4vAotsQfDsYPWKj9uSUU7A5aDhV1SH+jWOScUInXLoB1IVl6fMH0m
LXt/jxtDeXHr5Zz71Ihypa8+8UJgK8ZMTBrPThD0xht2sQinpX9ujArWrP4I3jTcSRn1HUEdAZgj
BhA5KhPrdzH1xs0hK21c5Y0zwwrpHJqdnRuRjrQQxE3yrF+RlLfO4obVF8ADZMMxvKrKDMI29oNA
Y8c7amrbsiLS+TyeDknMlwWhOrXpKALh5a96SzrM+qnSCE4QsqaHVOjeDbKjSyBgj5HWu+e/GfDE
cZUGCKj9WD6Erm1kJuKDuQ0gRyb5flj16ZzZeh7PO+WJ+TnquHWswRp+jWYAxl9UYGCT1Q5j+YLr
vXv9QBQrP4G9A8UNwQqIGJ9S4HAj9qDYVNFy+hEv3G3bFynKsH+VS4CbFqgP6LfDq+FdffputaWE
4f6r/YPcTVZn8EY7OxRdt4jTq4DbiYqbCWSU3gNLG1NhGBb/1B2oqytWxrwEw4DGsH5tzL+5A0iw
+FgxdpX4MD3GvMs8F9sT3LCztT0mVYIR1fAw6iIhRysHrZObJi5m4ILqFPU6uDCKD9wgQ4X7mcuD
XLeFOxD2uhNW+tg10O71lA69X33cj9LEyrNo8seXb4YtIU3v5+I7NR34/M3I0pOQWhXp/qfCirxY
PcYVvQ0DiFy4UJmzV1eR0XU6q0TGw3CaOCRC+VtwiBbFMGRE7cr4BuE2+kvu6yhoEJG7hrilBom0
PWzqYOvGDdIGlWLOArLtxjiAs5ZWiXO9ST4Ja8PrHYzmGl0dYLXsRLWMFMcE3xIli1Tt2L2Ly/fp
oHoD5cULdjX+nVRI3bNCfQ8LvFgVgrffb5poymCAMJc9Veo2+M8ap6/9lJAVPZYIYsBYMu1gHn/z
dVvA/+AHkeO4KivnjgeWdTO87OfezcjovI42kyv41WKuwSOBNuv6vQkbZps31T8hmYMd6uZUBmfJ
ufgdJyq9cu0r0Lj5pwqPZBxw7yyFoIYd5MgMg3qjPuV7GKyITPo1AAfFu01YCjF0rOR+x5KPFb46
XRD1c+y6clmVoxaJleSq2xF57uVFnd582k6VBdfD6vFWEflRFxVqSB1A8Ap8X6dWUmp2moBdQpqX
XFSCFsaOukOZWyNKH7qb6vSD3CoW2QEJAGyWE3nG3snexKfzOurrCgRUryizs5LsGB9Nl0f6rf6f
1p44453Xj/ewGLgq5vCIjywGUEk6iG0J9f9rifQ5whZnppb5Y/qq+oyQA5Lk5AigRT0Sfsm44ysu
obk3t9JGo7+1mevxt9jOxIKLvQXLBTdXdwFvQRWqlcgXNw8gLF7jH09ghlrVVadxuCpK4uT43ulV
Ivv46bbiumJ2uLjj2rGZZ2QxL11zVDVLtN1Pe7qWI9LVZk4JMQ78hlcCRZkhvlT0wo8+8efXHWqx
8P+uf+WHnK9fXSSqeStjc62qxnJU7q2++euSV5QVy7v1+QxZhjIkUhYbRpDY5HiN4UZ1tTJ2LIOY
DsX7dsaEz9K7jObkzsThNV2im/O4ezKl1X4JMuIndg545898OboUKBQPlYlApwbPRH9tPDdY7gec
dBl61HcvQO8I3I5bfByu7lSxaBNnpJyGCh6xhMUAsHqokDqv9CyhPLR7RG9+9QuGAYeHDgNGvauk
DupUfcgsTHDHQ6Ng8qN8zM7S1mx8sQNNP6DzDI0Uy8KZ+E2S+h2udMar77IVtWJWE/0CbL0nhrgB
QCvIEG7rHkRQSddL9vO9CJaLxh9k2E3Zwdomi+/J3uEryxBNgwsX06IG9dVWSEipbyn9uZntdUXi
aoGy7Qoo1xaV+Jw5D1025lROOFeD5WK2ytHEgF2MHYWQ8ikF6mXXCx2y3219KfSF7lS5QmTndNpZ
+JettOPrxttf78iNJu/yduFSQ7jHrkTJgpZMZ5vlaQK/K96yXKj0fEYxbIV+9CQ5IWzB4G2UtJWu
6k+CG/ueKWSToCAgbcj2BQN0u60J47vv0jF7HyBNjQjvM3xjyGefr2KtOaWEd9WIkXThWsVwaqf1
B7EA+I5EZU0eksvo1mj251AKMc/HCHuWBhp1X7sSZAmp1W/FSy5Hpy3cl+u0mdn5DRf0YS74HOqw
RvjTet+1IR6EXPEsZgk+IwTJF9qKYzR7R4fh++GRFW+vcgf0aU0WYuMZyvCXi2LardBBgR72DEo4
w/eFIHdsjdvUVXLPG13ufaLSz4WAAMmcgohrp+32BEbStZfrob6qRxvNG1LnIu5SKSvnJwHQGXbg
PZOVHjZ4R5SRhyINzh0YmmsQ640HToY+bltwZ6fwSE6ZzoT0W98vIPCAdGhAEz8l5aMcvk7ZBWzp
kGNLrW8nyqp5vWYmRu53Ti1TWD9cpcYpFEblM7d19EYQuiWKLJdLN469/w7U1673mGs4Pgqa928O
uZn//OfEGQ4ZmglF83eMmUROH1QVBuk9BlDrc9YuaQAQWHYnlKnVpMG6BinVZDFdpw7PQ1Oidr53
Qm6dPc9Jx1GTs42a57lW/jbK6vF8acRtZRam2Xta8r8z6a2W5szKyh4B8eB9bjWp5BVHovc29kN1
du7haQJ5kOWp97VAMM0XJKaoDNr0TxZ0C5yK1KAOehUd/R/y2RtitgbHQdbsIYFguGMjGyWWBYy7
TlI3c/1JmBKblW/Ga80w+f3DsLxbJ3Z2n5T8+gkvKbrD9PreKD41Xkpl2xn/xIfFxZTAS5BE6bzk
wfDQaMTDn8lIybZFl5cpzLWVBSEK1KLtAODW51RgiLUKmuZhpcYBzo6u3QGS31l4aN2DRhCl3Bma
QPMttQxL8sByMDON+8NwWsLgF5LtMpjsI2e/S5THNZQ9pSoMkcNxaQZZtvTw5HvAgw+y0jCULDwI
Z+7C3q8A+Mfw6ajFcCCYZ1kipn4/oC5gLyczI3gs0HAoGMiFxQJ6f+IQO5pvvY3pCMWhxHx+UTIO
RrNhzeAf8ofrVEl7mPzk/Kj14tl/abBaAZ5uetssaSOOXcbhihMeaZUdiXfKutH4d8GybGRLZwm3
CIFkWPUbiAhgSbhNa8XZuslrFRRQkm1c/QI8AXx2IdWT8EEsQhTaRPQZiVA+aLdy0tsC6tBZqNap
AIxW5czdGWsh3CpUVREqreuO8YHTBGRChBINOYncT9Xpgt8vmSkTKXQSD0wqeeZdyvoJQZR8/ah6
csaWc1j11z+SY+e/EtYVlSiBqCGrzp5PDegM54vqG3b5/FezHmYJ2tRDaVob7Zt4TbgMNwXT/eLq
Uc0CZB4feU7toFY8SCiH4jUXm05Ut2HHCV47utRAgcFoaqIwNyjjMkYzL1v0kzqdD5aIs05zQOUD
JV+JCqzcC/wyCRTCorCwJAH2paJMygczxevoXlmIDk3DiEFuP1QjBpWCPJBhY7CHiSARSjeuh4eJ
1QaCZJ9pdFq3+9QOtSXQSzraKe7cKMsmiYfWRQ6Xgyw2aqGPDuLqz+I9ducb2QsQkK6RE2ST+/cd
4emptX0Pd8KT+FvOJgw/KbeylCXaBH1FiM+0o6wb0JTiRKxSC+Cma89yP1cgHMoEZ55KaFUu+EF8
Wy3jojnVqKRmWl3813CbT0XhxU2AWpIef68oTIyo3WA5d4BreZ2Vt87ji6XA3R53vqUYztIBejtW
SunNw0V6PCTB43BNiwQJdRQYaqM3oNVgtXegzLTe+uFQmxiU7xJR7dDScC5MqpNQzeUDgKTqaN2X
DC8VSO/EKGtoFvMMpBWD+uMXIFVbn6yjzyB0q5exa5pAF/qgxzsH+G3R33a2eDNQMn6XNIPPVixY
SsMfCKC0naD8WO3gVmOnMO1KUYzo9KXUgQZF+S59SGCjvZHsMRDeKtWdpcrG0CKyfGmjYnuLyHU9
AtAXYaflAFDsl0eHPmbFdU2NDmUy213LYZUfGWMw7P/t562fymAbtbCb2Vnlq9rEVZ1xVq6uH+tu
4sXk9LW2ofHErfGmncYIYmg9zvO4/0y/Oe41SeHVQY+4nUPj99rwEeLsv1v6yso1FM+pkDJ1IVF8
F9pip6Jc06LxMkttTvt7X0P4+XfRUIij5OA0PJLOuG2GuJuH61IMTOBX15HR9/XztXHsc1k/HsRl
rJXI2pAcCbmzozhDOSfF6yP13Pk7vvDQkWdY2UvLGWA3BipKd0ri+qWlkrIUfdz0gu3/wI+KCimI
RXSGIp5SK2BQJIss76JovteMA4RoqS+gQnsozyE8wTlgoTtFIcKAi8muuDsaxa/4FZN3bB3oM4y/
XRdNAYgRPblHNK60pF8x3fYVE6yuGT3113S1JEB2xcyw+tPrAU/6+UPWWlLlRSxD5/rNCi5uh4uE
luyJ8eq8MgvBtBYVECl/Zjdr+zVhIsZaoNoeZFkY9Q/pd1pxwYxRdD9DTzE03e4Sy8BkaaHxw5CN
Ds6gD286limy4ifZQYY8Wb6CzRhrT/Mye0l2xg/jgGVGHmW01i0jnqYIMAHAoOzMHoDQmOGpF4ez
nrjxRMZsONjbGvaeuXzSbJIxIG5SzV4wEun7fww1+GWFalhQ84iNUjRds+B5Cd23UkwJ2Xqf4ol6
3cUnFzfMtE/GtIn7nbGLfy2JLgnuA8DqEfMtAB6K90A97oeUie+qqHmzblqXXdA3WXc316t52Xfs
m06Xg8oGUDaLhW/zXE2O0NTdVwAgeEPNlFq9O4kPgEOoLSdSbTpgfbu8vYgknuU6FVhbBdU+eQbc
aN7B8wZISjOJ2RaskCW7oVCeEtX4NcG74nWVq+iIXYLn8/JjCp0M5+AWOdGOQO8b0K3FeA6+M4o8
A4aNTy1J2RpXXXeWig8n0F5KQxdXVK9g6CNkdh+VFmRwXGFy73S41Jsk9VaoxkCIPqV49Us9roIX
Vg2hUojt43yyBGL2uvfM7zTJCQB1eDdFzEYZLuk7yH02g3TPSG20SqNOIFEd3bww4wsFww5irQ3M
8D9HMycESbk/65PMDuv4eCl6EdlMhRujN4cQSk4o/ybrodU7r5t/2QanKdN+NbP4xLbGhxj516Ve
YndRKpjsUuAN1nr+0BVnQLO5gU+pEjXHHWlOrlvfXSjTmOoALz1H56G17L3Dy0EAROvJNojAP1ZK
gG8ERwY0zp3IMD+dqJlIgjLa34XW6kM1CYeqwju5v12eOVKyA76xosYq9koEqPFFDvEFcrQQUK76
Ckhsys/1HSMyimPAQp8NQIqefPrUK6zPmpHD/xlnCPASrXULbrf2BfDQ/olH96OTxZRJ3ElFYCcM
/HkRbp72QUN7rrD0Qc2ZQ2Un55Wjul+HF7vDdL14qpx9/yCjbx1Z6xtgQ/EAzojcTLweFGHhOcP+
fHsuhW92leX2PSoIs4l8UYOW17XZ3RgWPS5LJfgzoa8xIsogIkJIQucKZBqfyHF8nKcU1zl0ZOlv
VU3zwtECvwVnwWsZa28ttJhgG7L3nwD3xfT5S9GVZEyLImCclHtJrPsPa74zWroFahvYLKw77ct0
xI6zVcumjSk7b7Tpo9dND/hTMxedkAQdXvWP+TB2AOP+jVtiJDNjJBYReQvDUqfIazHMRF5mRRIc
tU6DnbH94Mq+C+rr3UVSjLaHncljyMFobhMn9fUM9s4tNtD1S69PFqNM7maPC1UxvEQQ16lfZX9b
uybFpzsHv1ZaXa255V7nB6t+WWGZn3NAuOiA3RLxjd3xqQv5n9sgsJ7MRpUG0xaP9iu3OHDhQsFH
SuOrAm6iUJ0bAkxxG3Rsjy0VDFzQPklPoYzphPyFvAPk/2J3xCV+1feP0HAQHnJu2whRnqddeuY3
+6JPTptrLcSAHgVuijzzXFWNNMlr6B6mAytFzKr6PGjQYMhhdubvRF9r0uhbMgqUj4i3jqh8AfJG
Zk2nYj8uuMwF5vzdZJMJJ1hNMk/6ivwDaCxDgQr76R+h9KA6oN1D24vJhxc9zVB805Dp/cgdJINv
h/BXqxObmRVnuRW+WMVqoN7nS5kUGo9P0gQb47P1TNvb7+QMXz9lnVFJifQgS1gyt+5AV0nIlOD9
H+WRuIssD8BLCqkvoudGnL/Vt1BMP0DElOXcaZ2fuOrZ7X+7BTIgTxJ9I8JMkPwSLRnmVelehDVj
GmUJ34TrQ/hz9ETLXTTwj79Q9xVuBOcLM4Q/4aEYLHJTl0JsUIYMLA8DUHDAKdNNoxpOjha+vR4S
vDdwNDiRVT1NNuRoDhB770zJE4LCNPn+wIOZdEpngU0A0KY5FaVlJe0J9bgdaqJIZGSjRxYiIJWt
6HZj0ITvOpD6rH3vo8JWCd+mKzVL6ThXZ1nwdndiRcv+QdK2mJg4GNJIoBzbGv7VhTr0KrvjzzGm
dabBJxz46CyuWRWrYVFGzxQhNq4xoeYoBKgJ04FAwNxSdQGbTxU+b0vtAmcW8Brft30Mos2Q0gMt
fvqwH3kCvL48+SiKVMvnYWmONJ3SkZvg2pFi2Uea/YGB2PAruHJ+Nu0SFz8OyBNYXNHbHYH0+qnF
7LcYbPmzvfbTX2nUhAELapkIMwKQ3N9nNbuW/eBVEXD78EPMuP8LEQSwBJmEvMAOn7v86zk7VlOY
KLE1XsnE8SodwOAP1YarG/NKcZraJE6vedTa41LbvbAWoI2CXfc77CT7jgGGyhe/ZIQIug3BGdZU
ilfzyz6xwPdbyC+qez1HTXFVA3iuDtS8Kc3fcgnR3Ad9lhfto5z66KuORTxkXgNseFKWoYFK/o1s
oyawJWdHS8vrlIJV42+bMn8hF15Y6D8oV+qjKXudDi1HbNsU5inr7XZRjvoVUAenkZRvA5UvCO/r
Gu+rkIISkCVKaqlPs9QYl/4PidEXXQDJTcsg5C5RY8EuPrvGAC5TMv2qc5JDMhIgMd0Crf5e6tJf
WH924MMaRP2vu6ccDBNoiYv18AQyNaG8TAMv7edKyMOdrLLl/C2yzAhx26pxL0L6R6NL8SZTHlwy
goHn8yOHZ81FmKbVHaTZIUlq27HqCTqVfFwxm/e1xBe8tJ+8bO6taEFgF1gXZjfw2BcxqX4MZwxz
SHJW4Mx32YXH1BBne+kCRsznCppm2zrGZ2XdcDkZvF1LhqxLxVGl1hPvbIPakzwsP8KTLmC7Sn1/
oJXyR3UPN/jWxIGkzagTZu1RucqCGHdaZ0BMCi+wvqufQHwiikN0HV7L2rfXhALi/fH5gl+siuSi
8s755W7SqJ/nStG1fwIfXin6z1p8GY0c/dli+hLsOJtDmjzZvCSXpfoz/+56Il2sNV1UzE0ZHzmt
h/Q0JE9YFBRVD8r3CaLJs4B0o19M/YoLm/emIDSL75yRYrtbiG+c+PdBQmmYYrK4l21uMlpTMPAf
sxmHViuY4UY/DTb46hjbsP1MxLPdzlUNf+mzQxtRnGInkNgr3nVrmXtdAD+HovHl6v3utoHcW57O
Rb9KvZpHlkwUVE2xLp8vczIv9ObizaVSYWrZiPAlJEbRc6he5xPy7J0yOjBZXSWReVwxp9Rk5k4O
1DVYYYJwk8Hb1Cu7T48QyOOOAOjRwwJXTOQi1cDfoCypZq4xdedIjMEjjWx5E5hQHBODB88jJC62
9Z5jWJf9NHXByZVsg5r4LHKSPv6FXqzmFCwXJDp0AGgU2SfAjbFJrQHtfyGGF+o3pqErrvpObQcl
JgNLYswBW4q02R/aEU8JuOFdjBRAhwwP1i42SAyMLoBYWyCXia4R0XMnRACzbAaZ3qaIEWyyPztm
4/z6ZVZmEe88ebYWF4u+4hosjPuXWRrJVHlYGNaO474OvtwtyQb8WOmicUzmuYgU8W8r1kPSo8iH
9Xvcoz97z6Zni2Y5h19fp21nXd3R5hBWcMNGQ3JVfifpfXrq4sx9sEPf7/8WH7Ei86DTbQ+TH1ly
dZaI2MRkzRRp6SbHsevVec9Pre88pByLMa5kAEAkffGv473cJQc6DuBkRmK5vPzVtLLb1cTEyIGA
nQhxXq80w2tVd39wSG23+R1jtxZJ7OfWlFK3483InPTE9TC7e5XNQC3P69TMhrKozU+Jfa5AB26t
+i0ftoIPbDsxEwuMoL2dxlKEpZMEWZDvvA3wszRpt8ymO06RQX9QdLCLLJ+nZoBGKNrGq+a5eAwA
O4XdTgmkpyApDfaj8sTLr4cT984DFn+eaBXw3YzU/3xub2ANe+flKaSMrgXuCK5s/50i/t/5dCbe
0nhFmt4kpqlaAKzkYaFrsvn6bjxt9ptdCV3mJAkvf8x1Py5iHbXiBnK7SvXn2VnYamuGduyBBYJb
5ChhYb2G+VTr7ahhfON9zmYu9iImB/EsN3vpHBVY4TQgICZ+enMLZNx7SduR4Om5DOQpfzNXQ6mM
OZ3NZZgL7XKqzeOfXDBE2sF8k+Kty1e1iMRANRKBftR3ad+MiMbHa1O4mIDGOgj6CbWo2FjOK9tp
HZr+zW/yPyJU8BE6m8qE+HA+pN+Xj8DqGb+wgrCf9JQzNB1teqMxw8UQynJh9z9LAIw2HuzsOlb1
5K+PNtAsGVU2C2AbZNrG8m7KymjJtW95Bmydb7BoIjmspNJIahTqPzYiq/KtAxldUoxorJWt6RMQ
gvjsyShIP/2hNcj6zBl551MylDaYw6XSvo1y1OWX4YkK6wtg77Wdpf8PSIeExhFzeNuBSoTdl33l
wkGPsInGZ98UVu0NyeHcVwquaB/zoRalVuZf17eOrd1pin1pjKVj185FWZPft/Pb0HdtBUfAHYwd
pH/hsrPxR5c25tyaTexBzPlaIoxlxSvmxXcZ64EYQx8+kpRBwwNQ2CvXSGGvirmGG1rGSH4hNOtp
LPv4VFkb2H9Xa9RERf85bXGaBia0N7RMUQKCkQZwSjljitQXNiSo4Z+FBqnpGH9D1ZKfaXtOK9Ly
wacd8DPeWtVFCk1o/1uw3Gd+DiKu6W+pi7cTxTUUL1atu/rpVMnhQtXKyS7eLEmIYIVZu5q5GSt2
ijd3QmjIOOSrnfO0OqIskeCoceR+SmYYa4xFJ48UFom5+V9Bk6yaVRxNHgpp96D2XybWRJmsoMV8
ui9o7wGfJt1FxOPmAB27bER7kwF36AgrhSqHgPsCyFGtVsxIpJI1BdGLscRq2blOvys4A9zE6YH/
WQLgsJhpgSc8dtrKYAjuxklgxkVOj1XO8fTL7U0NSEQlTc9QrxhU+qVYAqibqHXjX0xQJnpkqvMm
ffTbxiNQ78R3+We0o4Dhhfo1Wfxe6dlDhqAXWq5SXRsc7v5iWPg39VPCPWR6l7k9lvE5ikRqULFJ
RurPKw2WM6thAtW9TLSzotB6N1uzUqzqiZVjo6Q7qhSIxsQVivcB1IxCIMohlT//g10FTJSWzh2h
c33a0TPWlRZuP8RXlK5mj3XT2f3PAM/DE67Z4vEa2rYvzXu0ShFsofNB5i7f/Fdiy8HJPPSrcFw1
rhIz8bjacJmx1rehIDAvTf2/D/EL8JZ17WRYW8RXTdZZdrJz9wq0piI6fHhkbu2LCURy0X92dXWi
FKne1TYHOoDXeWaQv4oYsxTkaFmd0y3ixi7MafjY+xSmfTphnS+Y0fg9U8gOiIfRjicK7LUcfu74
UAIGZEt5bqVgnWEEOGDvK3awhynHoPrlTT/sn18mZfRVBduz01k1slYOGwTXdhyisDHz3EDILJwU
kTW5g44E1FnVxJ3MT/JGVv3xAUVDe73jncMnsKQxGHGQ7b8UzyugAsCi4EFKffMDaTtbpl/W4hKA
/OXrA1DmWoseuQWMhEYQXuU0EIXL1O1Q6uJRSmd9HEHOl8cwBJypi989wqy3XvxOjbLRG2IVf/fY
5SvGGyctgszYmVxN1zaAk49d8AXzLmv7Zv2wBKhsS+IAzaG3HTH9jOqqSuXsvIsLwheiC8YcwDx7
16qY0xpnN+H7m4UFLK6wgoWmTZ42sk8o626xpUQkekQ3TCc5PyBQvAESvljgLnweUe9iPoaAFqJ4
sS5e3telRstlfCHArdau9UiI2YmmJdOOA8u/qrYTN82w+44pzDry+q4tdx19xGCXUbZpQXu8G5bQ
CxvvD6GXthoBzSRTJJTvVWtOAT8QduK0/Bk7uS+qb4dWU6w4NKpRhg/Jgqc/qt09dANH2hxYqK9c
kKyanAj5zsVFtJTwFjoLjWiLrs95yD7tBYeRp8YIooX+Y1p84ZR7Ny1y/4v3dv3AaxzukF0hKaMV
0Pn94ZxvGd3Q7gfz5OGuntX57EpkYmHMj0yNqhqHWtbCGZxV120NroOnEKmYdumXMVAw+osRJ5o2
JwUkm0ULj8UvlOCMwKY/KD0kN6UiMZxOqcP1fikIiuMqYwg2gnEfrTA1IGdESaJkPdXlhrb2/cwb
Uu03YdII29kWP9pv/PsMg1quoeyfPuS9abFm2e4Sn4UXj/v5KAMRe15imTe2V0o7hbGL6A+1Ex2/
TjXMl2OZRlhtoLAeulpLyt+0eFkX5uhE8sfVoWggk8rqyxdXLxk+32Ylo53GEhtfH4ZqfzNMabUC
KjkyGeHn7JqqTekzIp1WpmGslrF0L/mKp2cWrQZTu4f5qhwAG7gvbC3qxTONNa2NY2akSJfANMNo
o3Boz39xJz54pVJgHO1db1cZ/72+JtC+6dc9gzOSItpSsDfxoJCcntUTwRlXsSaUBdVdqf75eaSA
l+iVbNYDCKVzaist/0nG4D0297ETyjM1IP7IjqIfng9DI/4pe5qRx/nD5rjMB9t4FqGlSPUngLM7
vieJDTg+XzunqdmjwTFZlAbgJFfQg4G8p9djRRTagUPe3ML18+Y2xOFBreaC1fTR8mVJnoDTM5jT
SvxO5B7/4NrIUyn5UhYLV8EF3MrZvbb482xjsuT2ngtOrBK77bDRd0cRdPTEzteaW2BeSLG/CuGA
71fnKvrNziSaa3cMUM3VkwjQn/xPS2ybOR5/huv+RzuUu05J8It+dB7NAOpgU8i/P6d9nFuSc9G1
OhLn+NyCwe4P0BzIRrtpaV/WcMjW+9DexfQcw6UdWYChYzh0yEvVzyikWriUHIi73rZKE3w+KJd7
C36h73oPruFBUXYUvlTPWkIC2fXbUAM9ZvuQONHIzha5qrBkj/6X0PhAwYbyG3aDY0ieNK+DhGaK
6RXtjvCbfYOu9XKM3TXlERVmZ8bcjyDqcrWj8dVXidcTQ62+kv+V5bUSZH5BgsIgiMWa5Uy2R1mC
m4MCXkXm+xT3R56Nw2yD5UJROoZpgUyGbGPOQ3a04hyFNG1ri6Be+1LHqyrHxvTxXkwf5iwlcb9u
uZ+6kNJKM35TH1tvDGSf0ubNC5OaUghAoAXRAjVeNAcNrZqXtuY6ITSNAYx2XYUftDcReYeV0aYl
z9Wj8U/3PbOovCUXMSFE2trHHb9JrytoLiVfCNdZxv0R1gdDZ09oa3WIpPErLT6ema6CwV8eKRMj
ZxCarDCUty7MkXgEYunyOjqntiIuZsKI1oC6xpFB6AReJOa489JvxBXuao0BIomA3RN8C9bL8137
nXil0ML+3maXKHxhDfbXjIkX3nzvT8hKyAjW0W9HkSLAJXvwcPgk7PcQJPGziyIHqVoXCxq/v4dz
aDwg86pHWfjE4cdeMrvB58CqbYplj4FkVaW7Sl/e1ywV78RhFCnVyYVF4c7y4RxY3HR561Aaf/dg
hwtgx3H1w9iQWOx9d2SvGGi4yB2ZpjS6OsmqX0XJjYmbUbKx4R49FyA80z9zwdzBq/T5JLw4i+q8
Ejb8pXyfjp8XtToUOdtlK0OO5uADodUTVkArq5zyEjTdAnp03RjGczvlzTeeUroEQUthNdzmnQIz
/w+A6+aRqlW1xN0/e49ft58rkyEHtBX/ycb8wsW8KWMrTc3M17amjEcUzBvwVFBHs2+7dcid57h7
GsNw8I4QeVkj7HOaQzYJrmDse2702PATNJyReLlXM/GmSAGYEQK6YbKIt0Ph85vU9dQ5JLwhkohW
WxtZPTs5HLLkeSSvSQivTjUNdcr2I9ViDKvpOuWAJsKU0o36LZjwDdkLole40NoOQX9DP6q4KRHS
gyfandEoC8z6D3OpGv3Eoofe1o2A1q9xWRajus6Q8p3nByWT158V2+y6br9vjXhXQjfHuVaMjtJR
itr10+4+VWUOEWvKNQiSnv3+nhHC90odf82tuPBghgO/ixpct2Rb8AtyCPkYlD32FAd+Hmw/4gmj
z+PkPjcQZ++Nf0nVMeL/H7OQKkrxXftZ8kWdDSdGJ4UFjSPsStddzaYE+2+rVgAcDnX6OqKG3Wxj
ybCLVXzJQQYmtJ0Sghaio27s2mT66UUlG+18X2SIoKobnoGl4X8UNND2SEbaBvsmCZWqvZfS4nW4
VDpPG9LZV4iWACGuBG2tlGP4m7IgtlKVhm/0syJmQMekJ5WmmiMHWaIaH9WtrZedBKo6SPu1gXSe
P+MZFhVkYeX4u4UtLJYIP20dlQZgjnGEDXdJSo516DrM0QN/R6Nuj/sZrppDdieg9iqMJA/zjo4p
dxmFbqP1TA3x900fpoINtU4/FMhtrCExgTlit5kWc4dr9nvaYglNPFCldGx3fK/UmDEKDLqUkHn4
/U4Cr/zBsP/q12Mr0dr2zSDeGjr0eAZ+s2xspchqhR7Q2mUD9eu/z3/3dKuQOIgZi8+TG4nqwRic
DrhnXfR/8fOu8GCzNjcPBmgzlAgZzb2euTpsP/9f7E63Dj1TUm1vbwjVv6ngG/ouR0jcIRs7zJGp
iI14JY1EkXCSmW9EUqqjsflTdBWaskQFvgWa3JEXRBIwykGCAUJlbc0EeRVeveRk2eEPdoOk9j86
Bx0gH+M/Jt1q1I9pT4NCQeCimyPe1Us+e4veEgowULv2hULhk+tqnD1muxsWLgfVEeJPAxOAsE9v
T70FtnbsTXyPaL4wMVnFx4g849/RZNlKkmLX7ryVI7R8N/uqbVPYMZle0poFeHiClorf7hJmLYaF
7SOSfzkmGD13rdgLnaJigM6fniMWSVzlWG8ZxuF1/6IIM00tfFj72Gt/WRHXQCcPR4X/p1X2S9uz
YHUPbST01b+sJMibkBN5UpTR/T4A3AvoPc5lF/S4KGbxncllkoefZfg8bJ6/b7FOeDajeGFwCRkb
UpfF32B94Wo6NU2uZT19YVzof+GV4Aaaz/iht8Cy34IBTCg7CMW92VASbzqqCGYghxkvF026t4Ge
P4ZRhtERmdl8/y4AK8KjF1pMRKcM/jNb6cPNbcZjlXGNosNMEsfIoEmP2klvFp0fZ1TKAR00YPik
XrOvFsEMoU8kCrSlW2DRXDQJaAuf3IlqERQGfEY0/ixA8Lz8jt6kZ/V5i1+Soo93T8uO6gJjp25A
3RRwZ3GxIsgXuqinKuSqOjIHsgLTFo4POYftxeI6e12dVmUigSuDJ9IITfq6dcLjTreIy9ZKn+HA
to4XnyUoMDmHhv7r5W3B4B6NDbqx2AVc81Elu0ON41IrzHUI7/EiePZT9ZJCqH8qdEj3sBBM2kL0
LTx44rAkeR/LMh1EYSl0HyJ0RWzEq+7PaAytXtYcVE4sEApDm/Trk0hT7RzRNqT9j4Ke8IiB5MLL
JqGSeSnLgVvbBuXgWrZOgQxgSEtiTLNRStWtJwinITTLzu2+KxZeNs07XxHVmnckLh4feGI9uw1V
5gEUySw3PVbodnk5xN9AD/gl9KE3xxBEMV4nm7PTIcye72e8L4UD9bLeQLDuzTs98sPUfDESLLdH
7Nm269zShqYoqs1fogJXNs9kGUEoeigFGx7MpqdVQWsHelX/CL6qBA2lDiXNa9yrvBnMQliPE/1f
S4YPgnVdlyIg1IckCgpU+6mEgLU/OK/qShFAatFQIKay5FIrgUGAWlDwPbj8gQ6aO0anAsdBBoFg
t1w6MIG7A1MO+rhXXErqBAEvcIWCbfcnStyQsHDwW9jqwpXv0tfEeHl6V6JGh2Zp8wQbg/M4StHv
wdXgcQC4ww7klz32x6WbB6sblPbYjSeGQAi1XZsdueRjlEwf5GqeMqZyocfHVhIqaveV7S2mEdHz
3v7VU5yBoGT2xVYG/BS0zA71LLTU8caKrUykBfqdNsAEtRcEVIue93PIK0k2qZVG6htChLaTBy3l
T4cc+jZeojsPqnGKA2maeQbSIDpkKV4FPMHDencEbXRiYjUzunfxh163ei286AlW5f0a572fhwJg
qIpvmxpAt1HEWswjEx1LxkkZXBvBeSv1PQFIeTC0+nZOoOj389oLUmGoZHW23nn1fyDuNS2azBV5
+wSSD73CaUvNqaODIMmTSRpqXZT0BlYaIoA0W7FdG9lkpVpo2SoLUeqjp6kAgJrgXTDbkVlmyk0g
1X3FSE7UKeOF2gLpVoiDAj211gHxSY6ANyUwGA4S6NG9PPpmF3v5uPj5FA4Dq0UC8guWMWrOKYDx
Hw+kkTJnWGJX/0x90h2tC+X1QMgCbf3SP3E2R3AC729FZj02Fm60miff+1Zj21XpPnJN/VC433/G
0RLRkze/ddJfwOc5nq4vSeFVriEcxbhyStPs1s4lDfUtp+/IPTKkMlySy095Dl3GTwxwBCNXageC
45uW0xJb0bOFiyzNcN1m5PSPkBe4NcmwaVR1QIsHfKfr5sTefaaIOzlNi0fEoRzFhkafZUG8Ptcz
DWrgqOBa1FP+eyeSOF+10Duo7PK6l02lYz0rAHIFk6lRURt+kwres4+3zYTAe4X4gyh4SfNL3HZ4
UKd4LnsH0/ofcp8PYCAYr0sKFVVv1uMU/YQEbEyy62FQfD4ar0yUQnF5Tkm2E1Pw1nX512c6pzw9
YYQsm+9jQLtjYv3BiwJmYG5yj1F0ueDBH/IWunIV++ckXTAjV0aQAsPULnG/6yUBSo+BJGP3dTKz
UBCrOoCotUPu+WUa3+XI5r4MmvI6SRwpJMioauITEXAMdG2gQiCLxrdrYb81byETEeEsqiSNnzc3
9FCTxG4Qjhu4fV1rEWchAtgqN7EuxTOGfexLwLpRNU/k9lHq1jFd72PMNYQPSYyBSx0hUCIsTKlV
Wk1p85VxdMwG+jTPmiu7ZCGKM7Zubucj5oDpHDIW2UJqg01vf+YVpTnVCRLdqSvMsqFkd8i+Juv1
xoYyZlh/3JjypR4kXUFIgiM071dCBgDsTA2F9PvMOCXPZNTdGly5oQmgFe8iDVPIiCMqPDmtVq7H
CbLoSTeH5SOzhhxQmtcxLWxHKmFzlOgO2pHHIJ3e8p2iFWCMn7XbK8D3CcZVXaKinmQQ4Oc+pucb
gsBrCiRrJEoGO/e11WYweDr4Pg0cQJkLNIyKcLdP/dGBuuLPIR9OAk00uaOD/POusQFPwzuwP0e+
coi+OuYYaKhr7OmkggJoUMmZTSNaGXN796cAUF9e3H4Qd4ED4e+WG7i4dxL/1Z6o8MyTuPcoRIH6
vWR1ndv0ZjgPOBRVd/33yDBDFnN3tcbcIpa9S3RJ2skhfUZp7/Rmp8Nk0fICEKHV0/RAh5I0+B5W
FXfK/KRQm3L2coTR03umJb1ExVRNd1EO0F2hSOcGVK6mU45iUhzQU9rjABZR+zrILvJCvpw4xTIL
k+XW9qROL+82IfcfOmY2INIb4IpLjIGzXU6QEr/ckVaP3C76Pp0vf705dKkAVY93kzPbgarjo3MT
VpraPd3rByB95H59PI7esVHWe6APhYBFK/BrqwYV+A5F9pnG5R+JK1VUpznRdk7GyUuCCXYC8rw3
FMQ+V4C/+woFPlPnUG0sjXnncnNo+HqzPePgT2KXg7adh/HFrdMK/KUmQDBJ+GlCZE6ljzvn0sWY
AcylIs8ndRbxy67zXHYQ1WesXI/oj37/eJ91F7ukQKjw6U5Qz29U8nqj3HH8qd39YjGyYnoQrSC8
XzmFGvjsrVCylINAwekcdkAIDZX8959TgSdq6lQNRK92mxKzonYGY6zmVKGuG/DZplCfet8GwfYL
p5KAupVUnNz+WUzuxv8u+kMyD8gEmv1mF7xMb3mzpVDcQ8cxTEV45zyRHUT8LuB8tTFjSF7IJUep
BVSfkOX1jYQQzLQPOyd/NmbiWeJ5FlQGGDOWpMSXfBz/
`protect end_protected
