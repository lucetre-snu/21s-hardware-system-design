`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
D+9lfS59pj/VVil0GGdJ59k3DOq46v/+7whNz7wCwfYdRiJPbLItui6o/zSBZEKI9gWLjOldtur1
/rmcVBQ3GA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Al4EzSQFZknJP1zXhKNIjHP2ED06e/ds+6xnXGYdohXSo6+myvUa29WxrDQ2BRCFMopuWgRIHVKr
QIL1R/lyNoyVEM+ZIozLEHgX6l1O/zTuyjCCsopsjgqJb2Wtgn8s+TaOCOvqtDrvLzt0PvLiCx3j
UkBnJ2bYuzUoN4JusSo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GryPO/G6YUeEdMxSH6E+Cylnk/9RJIpF3DfZ8qm1ecWq6hYmaGlwqiFs0cnQCPLUX5i7YB1Zhyg7
xWXnsmJ4+UqH7C7kALbZ0VgPMoxq9qXXyR3XFKCabcHGfdH1PGZgCMUJcT1U4IAGCC0HKbpQue4v
BxJxLOKucvmUl0mdNC5jktjqlol5N3LNQ1Nqb0Bi2JUbKhDXyPAghHnYm1RA1WIG/I7KPAHJRMsn
rq61TkO0r9B2jyIUh8Re69O30QuaI8MVXArXwxoLarP1bw33bj+4nw7AKPOj3d27JIY1FecXOlD+
JrglMTs1oca4ii7DTHZWrWcZD11O8wPZrSB/hg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gIxs1xJo2g0tw3pn4+ixShAOAMuK8enzcVscdNEALwVHu56ynHRf8QNrBE9hWTm0Zrotj69ZA/BK
kwI2N0AWvjk9ACiHZ+Q82pH5keVYRtMQtsAzmOmN3YJ3UkTFHW6AIALOLN/+b1CJx2DSSbUvSJRL
vYdCMY94F9Lklx9UjVtQ7r4y14DJeU9UdmLHZEJTMZ3ahOPNz53F7Y+D2abS+pN3OTP/hfwC8SXW
Y0mKDR8Tkg+zCHqpFqHVe4sN/fDWpQUR8MUszd4ygr4o7HqUOQ1RTUGx1Mc0Wtrq0QAi8Syc7V28
2OviXFf4KLhcKYs0bZN+gsgApGWiwyRvQRkZsw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lbc8rPGs9vNVJLV1Ztd+OweNWVf1r3bbhZXmEPzls7ewmRVAwHDdCz0iBVD5zHofb2Pv1cNIx1DF
Cegpi/O809UypK5vc2xsVTWDeqgYhsqvVrROg6FOkBiX78rZZIEYF4NC0rxHw/5ixAFYsGHPS840
rFWEsubE6/eEK5KjxNY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dGaX53L9Ek9wU1QC7h+mJBxY9VRQrtTA5cLqpyZvyLoi582YqMcyFxxsOh08z/CW++CYcslxK5c2
nB76qWzDGxhrcZ2LL96TaJdxfIU2EOvAbd+35O26BL5Dr65GaDwdjrxZgGVYX9zZnupIqxn8XhmC
YxZ5OIIBnPbpGQ6ribzMzlGvFizUnWWAzae4ZJK4JY+UWbuv2xdBtaDjg/1YQkACqpob/Aq4IcN9
/z+aEP0pGhrF9aYTALhCIBKRSiEmlWYFi+Y/QtDMcgPf3kf28Jl2zN9nxRNVeqUYEwqb9cl2u01M
MuW6fdTQYP8au8BQaSrUEy47B0go0sgbZVDbwA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LEujW+ttFeLDTd6Kj02ulQ4/6kxvxmgT0K9WSqzr2nEKo8u+D1wTZSNxo1Fc+SuL6Np9NoHmXZ6a
quET05vVSiMB+lIOHpijfSVwTqZ7LgYHnhXrPB5My87wRq0b9Jyg7VUy3e0yzOlKBYa8cqDKm5vE
rKtHLezwwsG/dfHwGL5KISY7D5xkA348D53WjZT2GPECqu3z2+qFTyr2skARLi+fP7tdqXthwiZ/
w32KaI0lhDwxw9CdQ/7jGNqq5B4pDSAIRhs657DCGvaZmMrfpEV3TIblWlorFwEQ5UhHeGuVslc+
eN4r6MzOumbMdENFQgB8d3D0vFnoVsLbbL5/3w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b1YdODjbk8HFhbv22dlzSJPK8onB4y/bTVR6bwet5BZoTYdYXUmOZH419afEKigqx51IMqa6rnXU
3J62hXejiIyZsm1mV6d/ZILTIg4MvKp/nsB+nzk3mwrxlbUBSjb5Gs4KJEM3QfmnigtYMQ5rNsWx
xO1OBkWglwIieiVxJRpIzrM1m6NiWCqcL1cvpMI1IywHrEeI+DhZWAgf2c+NGLeogq0I5stGLWyl
7mUNnFVREZS2ztdL9JeVlYFnkm9YAu/rEpRnd/ZFnUmo5LDgPLxnWIoTIbnJ9ETXA3VKs5m8RjLa
Y80BwwVZ8VpAYtcyfGThAvkMUN1XkU+RBOhB0w==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jw11/jyPzYF09qKNLzRASveW80p2lDhif/7GSzkqz1ay8ziMYjGu2PXCgyziHf07D1ydjBZ2Oj+T
1TciExFJYUoS4v8yaGxNYIeVg4lCZtiWwMwIjWi5TbX5hyZCCFDUioAcm2Er0tzXe+UuWzkM8uEj
VcZMHxrNXFh3ip5Q5HwOhZJLT59ez98d86/DgXZNDnY1jAn3tjdLiP3facR+GKZ2RlNKOTvP6BNt
RMIiYfDGS6i/0a2j9G97hV2faBZ9PX1JyNer2z3gD5/XUNbE3bPLm+xmhpk1/K7GiF3yvAO1dtiL
5Mg52QRrud8v05hWjH6y7rmg+wiBc1bnMIMVaw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967968)
`protect data_block
o4SFjgK1rFnXRQcv8x34k87IKeBxiR6fYgZ0+j2L7TzA3JT0uV3YnQ3nTp9aqw15ruwklCWo0nLT
TNGfI2ofOfM2arUP3LwzYw6rigO3TxxWaLTFyx5eMGQ+/IIASHW5GYYSbWBRrIz/3m+Eb6qiG7P5
V8n3t+lynbmJa1Z9VrGWjpSpzyUgxSNKhV7H6zRYdpHJGWCx5iUIYuCDV8dNDtOAX+p+Ra7oQ0fx
jtOgM1ybGWQTYTVp8R75zJDNW65TqE83kN/OnMFimmZfYQ14rEy8vxRo7b4OkiutseJgn0MZmt5n
FjdtVpnYnDjN7TvDKfMkrjHHVtr9PhANK6oJxzYigb0zrS8KPd7qr4nEw/L6WX0hIwFItRwoUy+k
4ML6F9FsY5j+LQsOp93Jx6AIEQiVPI/pNOO+B67AJQ9FpTND8068CufCbhhlqDxymhXfJY6YHly4
0rRi8I1eS4ckpT1rgOZ1X05QMaavPxvc9L5XLztPC9Oe36EFIgAFQijzk4bC4WWZJIqVcLDrjxgc
tYZNrImUa9l+gJcLLEA0Nh9fTbD74/oCOfjpiy4xK0CV2v17wGKGJJpDH5sGFv6Lanh+s7TQgniy
99gIbkbEvCXAfHPmJofkqxTG0KwIi1RhGrNbzTG2TVEFcbg5YfL445hxi7n4dlEm03ur2LeCdgiu
exbvMJdK42yDNlnWU+oNi5EyMZg92V8HObh/eX49pyX77fnPaj3Msn2Fst8px9/RN+eb6dBsCSpS
f7HruUGDA1kvd8ct27fqGWH3lCQ4R7U8leRRhHJvkLUIdsRRzqSa5OdCBmUL8fu+oJyRt+mFQkm5
RwcLfGyZbCE51w8WjJq2sXlpqxZw0rFTsCytoi++5J5Cv605c4JjLdXYLtWjpqzG0S9PgR61oiI8
eeoWwD/kvADAT81SUuaTkWWydQKifqnKDNsws7145SStNkbL9YRP3w7B5JreAbeDdWWd9j0vPqgZ
+CNVjQm3cKyFJfqoLN6XpLxqARsVdRcVM3zE/fblA2Qdh34FVhG/7ffsU94SiEHNA0esyRR7z8O4
i7JnCVwIQ4b7YpFitJskoz0OaIxrmRPBr8DrUlJMJ+jzxfp6ZDYxv9exeEtwmuAplMOLehQ4pH2s
beYR9/hkhydk3oX8f3rubGZTtwoS3sCfHppP0WXKCd+rk19/irNgZrYrmMeIU2bGyhfnOAMw8Mtr
yvDAzlOte0QCt27+VZP+2CcNCaTVn/ncUHCNFMXktqPVXsc0In3oZcTcMiay7fPEJ18+Vtltr0vQ
7Ul8hRu9D1wtyGka07LS1T4WyUml/nm+DHWBfX22ByyFEaJfyXBP9FW2pShrZIm/lKt1rTjHah/e
8Hy88w4Got9VmpqiVb3xq/5+9Q58Ht6aZtik12eHPLOlYyb80ICzNVMxNiHZavtV6G84b1Is4QGt
Cq8j7YvVPwQksu0EFThEKHjjc5MJT3SX2wZfNym1v503GAzQe/vZmDHRqwYZIutvSKoKjd6njefh
it9udIkMH8JP6lza8tg4yrj/2GGpl4ge0An7Y4qPrQj//qhz9piu/cJcx2Rc5kco4ZiWDZ3hnyz2
wwexWfq8L0G0DYSsPFNyJSxi+Ug0hmI/QUdauhTO5BxI4VhMxmHNmTv6HoIsPmErcbF4Y+DH0noy
TW9fqOjWoaaCVMYdbahIRPSFcQi+z16VWH07GydlG1FpEnacWNufA0ZsFxn7DrMZ48NUM5MjNhIr
w41qae4vd2rPu/ib24d2ZUvxCa34RVjIDpVTrjwxglZwLSaz0lRq1edzbDGtt97wGT08j9me5YXr
M+zIWwYCGsWatpa+Ckau0Aipd3Hzh39RJmpjHbqFhRz4LhlCJ8nJ1Ks8WH28nXr2DZxkcWg3xQcV
zMK/Q7FJzAXtd5RpajMH+GHAuZhK/2aWXsgytq/7igaFUFKovACkz+N/ekbtDJjcLeYTj2C5J+QC
uVH88DwBuuI43wXsGz5/R3j/6+MNcR0sON0jelu2DNP+3FmTMEVLv2yCMg2clMTl36KlscDGw/FP
SpuPoRdFUY37s4fkKaUlMyZPuSxGAI9VVl0DTdo40j5QsvNKDRiWbH+1DNT1mh4v95r/M0fisexm
ND6lK3RMliUAOe3oue+vAExrGrIRwSuj7l0W+n0U3OQc45hVxbp+/6PHfCOjzzRBvZnkzpFogkSJ
7HyeDKAFENhQBN4+3qTb5RmJDjZapZPYSeywhJdolILCVrENbbucmV8mS/gAeVT7xVTxnxQ2CjA3
VoN/SGmugIbGIgoOYJ7V7gBd2Ld94UpdTcNjbYRKmKw6bUpyGF7/cAvY3uprVrRrqmGg7NXf9vqn
hpDpalY6/bAchPt8YQh7hEuc9ECTQ6E3SIaNBlEHMnsx/PAuFoXfBIpqQPT8IjtBXdbESZhBDNmR
/KZ8l+E+MTfqBUj8KLo7lKHUXfT219L2fSX1XbyQWK1a7xFg7ZUHjx3eMZZWwZAxf2b/Zgv0fzyN
OtJws1ZBHNRmKLqai7aBJ7vOoT5L+/XsUgZLGlyYzB4VZwgNMq3cORJALzW6KqcxcMrLJ/SE7Oci
HgKIf21+TPYTJbVVjwaTFWVnaJO+rgV1l7JRZV3snbRBjo60LDKG6vhjuR8Ny7wg7z0Jpj8KHzDm
zRVbYcANVrZ370zG9Zj4MhUypF0PEy0oTKLIgGBzkrjLle/QnZ84/478Vz/zxoKUOoiT34nWBP+C
oLDlqQJmK3/fk9q+Ar94eSPIIKxeQLNS4hznD9noyfG77UVubuAF+Ij89OU3NiMU8D5V8mbgrY1/
9dLHVprrs8MDQBmQJxU6Kbntm/xarKFHeOzR+1rMBtHY8yT/+SbLlXnuR5DRnFh7BLLKpdjckjPK
fK968hDiVLibathzLB+FJDyvwhjjnFEWDmavLBSjpcgxVm3/5EprDf3AGPzRSdZX3z+fRL2eiIq4
FOUJr8735dRkdU0pJb9gjLVNNzOvvcRMvPXefbNzdfU+LRgxS3gbFuECjm3xq5AA17trJ5E2WIpv
PE13hCO7ESz0BZjTzB8AfOyt2UNFZEDIXB+2M3xsTFuuDub2k31W16gTBkV4V8t27Lgfz+ZzwX0m
i1c73Xa3E+ApriNJYlIVDHQofoi1TjZOZgGBU8P6laE/oetx1OZarUcf/LodxFa9ijeGJIMvaUGZ
ID3NfBLC7IrJ18zsF59W9wUKT5eHuYKt6HrJZOYOHtOHMfXTSg7lhD5sGpoAsvgf0TuI1083g9Q2
Yp5MlGwsJ2dqcLwg57bXwgJkP+aT4q4Bguwn03Apg4bxCJl2O1bVNrNiOnDFZvWRJvwRPa98sAsN
BF1CjkwGrnG9E1pJVy9i6y29AxqcAEY1NJeMb+DQentEjVdffbNRRtuWlkMUYqy1DOsEokj+Ppxp
tupJA5ZJQuJMf8xoq1EyVbSlQGoOAoZH1r3zfckguLhOpdjpJgItisTGxn5QiAQy/93mycGosUOr
wg6RuMv4zZNUMSgH6UYZ5EtYZ0SnWosstZXFz24Fn8z9J9sSnfQNpu687rQwgE++1jCF0BHPB2pI
N/q4HxTj1vgE7diiqFxA5ANUHZvGsPHTqpfmpdpxFuy8uUMn9PAgUYBLGHqokUrcuTuB48fyH0uX
fJOyC6P9VPa7m5Cot0MffSocopomb+F+cEr+uXjoXxKtnyA8/2rLy4xTb0pdOEW5GqW0NTfjxSFN
mFtC2lkpyQh/Kkasp0WUFMCYaqJcnt6UV0MRaUq1IHNJhP3l6zaLA1jVaM6NnbjMawySiwYv/4mA
Vdj28mLB8Fa+GqN4gTahlrc5MA79v83TN8Ss8WtuPb9ikUTUTyiEVzEeP+JoASxwZEE5a/BdO9gg
xhRyKK0hGF0QGlZypx9QdzXUA4OYmQlXxWtxZ9Hu8Vwi0v3FXonqGx5zH7gX/Nwxw49dZhkhG1Bl
3fjniCDSjLu8BXBScqpAWCfPgxKj5e+PGIR4anedSt5UTNJsKv9qa/acKiHpqL9EmlDA9vfcUfEJ
eEcj4Q2LOWqgP3lLJP6V1a4E7rtcAeoqkw1mtO4WoihD+8ypoXUUEappPZndTRRDKI8eoX9oQJjI
MnkuWRLA9Gj9NI20N10v56Cu4T40zeIOg86rEqUgSxP9DFhAcSczj+1YVv/34uEqXJmAXEsL2dZk
1yR6E4eGodq/G3mNK1d/fj19GO3Msx2G9gCt/W4y9mPk1QxoMyFz+gJsYSJHVx60ltB+k52s1Xhm
dJH89Dh0zAadXZkqOWm9iv/nZmBa/Ax22ljy5ofyMpJz+8k/Ol/8CSR1myUz6w3Gn/tkdRcJjagK
LtFXw/M21MrwFCeiins3Hk9FdwDeME/iWIKOV7Enh6mwORjVaQmsxWKHSCQYq/KyZPjIkD15DgFG
uTuNRV2TAWLhMjbGsUG46qtUm+IUXCVI0P+RQAQj0iscBYHGxBa5JIwF9y/oMqf3uO2tvmZO4Wpt
HHdgkmIT88xGSixU8Ngm0Q2rXWADG+u4JiY4m/myxa22tIYSRH03ZgGPZrola8bBJ7U1ZfBd4TNl
zxnDVYUekQkImsG63DCxaLDV2z77kUDzYNmjput9dtbUQ7BbQMqRKRy2p2pF+6wVdq51P0pOvcjX
D3qRbwBKiU74wRDPjS6XPY54JZWRjoaxyxJbreTihIY+7E7AIBPdj6FT3iiiCt8duMhdIXPYjHQu
OgL74GhNT42rH7UQkfMv+tlhZyQ2NfG0N3VfDmBBNToXsRf6LkZB9rXLrMC6N/K2TJ2IBVwoG/FZ
U1ceT93/2WOjPOizVLQkSKKWIpKLHrbCl5zRLxIwgH15UJYr/Jt65OMlUjRAPshulHz2GVgH8884
3Lk5i8tBGagXhK+69cWQcybzjyLdyAGn89QWFuWgdh4NYRcX7k0VNaQWzprD1vA0IAaXG4yW4jT5
S3evF3PUAbzlWw+/ytx90WxnJJlrsE3ADY1DmHVqRu4hTZcMAovgQ4VnMP5YUZpEoKgDW70L8I9x
2FLTQJGLxwdlpoQghBadkIPx04kSGPs1k6cLrG8RJEYmnEPH4eQTJ5kjvqV/DNFETYA29G2vY6S4
Y0RxIRt1mcoPG5FjAwcJq/Ze07yY+ltN7AYbAhrs9T4vV0yvz6RC6XfoNntamkuDeoF0GtkM58jg
Zi6jOtZRe9hWdBrfI97Od8zeX+ZxcyYkPF3FDoxaito1UDKlaKxFl4s1ARmNYCqN+l1JNzom7KE0
qqnuBJKgU0UtQBVg06uN14LveDqxE51+pHhW1X2K5my6cixmtzzy15kVwa1F+G5ju8lgrav0We5N
W7eYynF6B0dUgAx9XYlvYt/ovt4dgTCZe5E26YrD2A5Rrh03fr1FIWqw0JhrfSoadP/Xj7diuORz
isSCYOSnOKqxhqJgsSj/zPPMLUjPSUyWo7O6rudyGMyVtF+D8QD4ryPLCCQYfkD0nNEXbkJ93xtL
fIA64cgjrpy/Iw+dfWRtcFlK+AmUqn9CYlZGWqmFbBeXyfqo4KmYokjlH8UY8KKzhQ4yy/imB6eC
eanBZikNZv0/bHBxkq5plWvsw88GtKMKuSUrLqRhgb7K9RTYpR4pE1283io70Ho8ml0MI/5DPmJx
JMm+KjicxVH84hXELWO4nIcAGY7hFN6EjQYwnt6+WOlG17/EoLhuSmUTy/NIXhOsQOrCL6IFBXni
9TnnZeR+vfxPZbEa3gfkP1mcaOXXIkq3CauKVGtINAjuHGJJTuWgIqvZ2g4vGV+aAukH6FzZwp0K
dN2oJit9TKqH63nciztmNryHUpnH3HAcYH8KVTa5XbtVMYQLiuXM5Mg+9wCPoZYqfN3SmZsTdudS
l6u3uPS3uXZS9oPinY9HJL6l8W8YgWFqpSS5lVJO4XN2EhYdGuroal8ToRpip2Do67zauKeAE9fA
p7q4iXVb0G88jhBC0KVp+eioS6EKU6TuZoKZzqlG8iaJ7+9SdkTnqoBlwfbVPRqXMJlS2yKNd4et
Ve/se6x9wizXVPL3YlVmxsTYCCssO1azOrlW8NAXxmKHyy2S9/lAxTZbXM6KcvSpEUkF86mBd9Mn
Sl0epn1N+Pvnd8gwy+tESUQLHywxNu+WyZ1f5ZU5xsHA7PocPj0m098KQOv911D6qs2CcuZXYDTs
rVsumPvKOIQ4TOsT8IS2tTs+Vhks3/y8CnAPwtoRsXk/tTbFecLyi2WuxPl/tj1Al8dVFxvju9J6
KGYnbm+1BggiFbotpBV9vFxgIN0KHIZjJg/Rc9w4NHUJxf/VhqMe7nAUvodCoOTtLb0B80EaK+F8
eWT5XtWBKsndxu4wLfJv21NL4OzQB7FKwKFBnTHxu2Z1KWdEy4y0snNOsm3xMhXxUHtj9uQRWvEd
ZysrZ8BD2gcjZP4qDoAGQEnpoAms9eDmSCHwvCFH/JNNU+SA9KNecbDcH1aWL8n4OCfbt1xQY5C3
pby8rypTXOS4xeI4HNw5o/r6VJWcylQ2entOuFwFnDA2B+2bcVWcgyVzEPspl+q9VPf59M7cLqeb
cIXy0te2X7PCkfPZLhAnP5IDSvPwpHJEYYtgAJyO0NMPU/udoKaqzefvkNdNQJnhU5Zyn8G221bG
skK1WgjbqPYYg6kG0OmDEY1v1x7d2je1GZMGPAuwymWOgmj1wzM/UriNvecLOO3WfG1D+MWdDGzE
uvfhUHVrwapk17SCIkEIMBmRNiYdH2Sk30FbUZgnMS4pHZQFNd5cCFe79saDSQpSU4eOUQuwtm0p
Gt2FoHLR86mKYyF1mJ+TaNlPhCCJWv++IwcMeUJk+XJSh9N5y61Od5ETXf09gnhdGRJd7xz0VcU9
1bdFMPaTX1WspPrNWFgpxUkAK/mwr4sWdQznINcG6RTSVT9gSRXQtteGUGlmwukM1YTq80EkL8uH
ZVkO6X6QDtPHpLJLwAKzUW5ggWIAmvLJWgtBGNcTsnMHC+4wcame3m/wzBEXFGJ6Pq7253ihM6mO
O81ipP1zjkqHPz3MSjgR3Dsd4jfn4Nk8cOie6uci3ctOO2WT+P/JixavMkqmGBwx/6q/2IGqokNA
cAzeLBLEf5+ER5xY/Gn4MS8KJoSYs/wL2hk4PG+qm9tloQg+8yfbX/YL9YB6bJ+pBQD9ae0IVU7Q
MQq8LnBIY8JnCFA5zB0Lqbqu9d6D9rHvVr6UbZrU35+xR/PE8hsD6H8M3xV5TlzWViQI8WcYl6WU
ql6LUJfIorRN6Ov5tdUe1HpSrg3vAOvQ8Ou90jsdNoc+Gd6xiGvEEKbhnPvf1gsCh/hDm6pwWY5W
X/QFnR+3Ibg0zMFbA/hj3nThmGCI7GN7p8ifZlbm/AyvLkpWLVFHNLq0cTmJRe2rjY+w3JwCd2KH
AK6FSsCroBOdNxU1NOhIjnI5iPBRhK9i+CHzcjZsHCEUwZivAiozwjUcshk5iCHv2TUrwhU3OoOn
LHuiIRDVNW6U9HgV9TAE9PgtFSFhk60RVUtMi8sKcKONBFLGWr62tx5p/58zyv+VTNzLW2i9d2l2
CcRZGBN7HbcEGFIBj8UEtIPVVllSA07LKHcwXzbcRvnXpPsxD5YrNV4Vi0kz03SrVD9JPnxVUGB9
JwISEPmgfTIVfRVLxpx+67toju11D6NDTa9Q1Q/L9F/4dz0HX+tq7NFGaCTZBqrNlIMg/9BOpTy5
8sSi3BXNATluhNLfeuqKBZ7+R/wL5e7wJhIncSohA/ur9RochAhwhITvx9qwfjdwIjsT/r3mz80U
nad0CHkzowVAeRU8xzXF6kCAJrxWxnWtzXi9QhMlYH5Q79RtInPU1npw3IAfZsCBzmikRScCsMlZ
+TpFfwbA7WTgIGqWwSXW31r30v4AggA0mISzzpLNLaYKlnSSeA5wNudqWlds5IJIJ9fWtUDAfpef
wnpnjxZb1l27U8gjgGhNkdFax5ETkKUe3pJTW5liqmVIreM7gHxc1+swu99gw6OKswD7ag1z0CFh
LeGGllHbagfeo8ER4Oyu7IWlonGSRn+KcWykKoWB1nca7MuewKXCSRzeHWHX19k57izJdYIq9ZnD
stMC+hwHULIGgDCV1Ox1pAuwKreQYJuEc10PtpcbcHpwrGTsbe/T3vQdc7jAxlKHN1iP9A1BirTb
axl1iwBjICfHOEBL39y29pfZQvk/0Qi+UVjY2c5Dja9+IOmDfgp5KmXu1tNStBWeevvRItWXQsQ7
2BtOFfULerCMPQnIGf2RdzH4iDXchGxRuX/9LV4bIMBdl3KMBTzFpe7XxwKorK62v8fOAfc4SMYu
H8Z1ADL74p4cRRQdp8CuqF55ufEbudZefJI4iX2hiJl/M6TJCnoFujLK1j2ieO+KLk3IggUELIuu
Zd7T2u47rBPW9KRPvut6smdNlhdFXPXi1p2n7kRFOjimGxMmejB5bR4ol6GCgV+M1HVcmnG6TgEC
sS/rEQlMh+xg1L7ILqcmXrXQVijV9HH+MO0vfYNWeCLjf7fClDzPtyl75lU1leNdbzSQZtzyDy2Y
fL5CCx2Xihrd7XZNuib2uwUNAyjJX8/tSBSFXV0Z9GVfrhqUCfSG762U0/IQNCBF7HhEScS2FK2P
LnZnkgWHITARmx1Gkk7MGcHGLY5JS5R0eY9JOi8z4biWL5eniNpPoeuBhbzTMtjQwuIDMe0iEjwH
bzDjSEE9k7+o/UaHfsUmE8p3kVytUkrSbaQcNGVwz3vjuRcqu8phRC2332e10zjP50DUAxrQteZg
KVNyssmqWQhDrAn1fWkB8mT4PMNyOXqO7E485Iq4gh+6w/6XJjLh+y7oIjarVheTZGl3IVkWSRVb
Fe2a9ggfG5Gs4j81q4Q95Hcmdy2+OExFsT+tGJhRNqY4YtXgZdnhVhDY4NE4pfscy8jCL6+EKsJ0
/u+wgl9Z40LqhjyjZ/slMX5HbFjA/o1KcGGTIpoCvwYvCIZlllwfUcy8AGDNWtv4EgjTooldPsO0
MezTTrU8xXRSQrLO68IC4lnnSd+GKwn+U/16JexcuUozfJc1B6Clw4ZESj0nlOt6hkxorfn6y790
mOuZtqVeT+h6bsbKwR1uPHFcgPD5LbGdmbkYqTA8MWo9Xevj2zg9s6/z+o2uX3WIUSljj2H5t/0S
TiNk0isyn+ky7/2kOrxJIOpvwEX08yxqoy7bk3kygSB/4PYf35irXPQw1mRFJ0ImcOtH8anJu5u3
CcceL0UgvNnWvgTtSXfb1nm4GcxUhC1iOOf0Og2/NBVWm79jxRG1pboPRJ5bha56eA/TM9f1ISDd
sn/FznZ7xl8lVSb1yCzt9YpCXXwDfvMkMpBZoqC+e4FpPyIyyoz6pVB1S44/FsMVE7AA07b4nfb0
Oo1p5AMu3p/CVlDJ3QF16d8jV1ibL70crwWW8MnyOciJT+KyNVV0o4XT4kpqcH3CDDjc177cq2r0
F4hbbK9WQSG64xRHOduATMWI3fqCj4xlBkhCgeExxDCH+6D39QKrilgnFBFEiw7brDFHiXZF8vH7
mqjsiXVmvN18DC8T/fJjXFz1hA46hld4jjAM2xD5wiW+eSKYZBrvgePMUv9H47WrIC7a+2aTqeeE
J9Wv0NCx8CYtWDAazXOSo3Ca4f9MY7RVptb3FsHjGtEVVPbTT7OKDk8abdeOJGDfUegCKjvpaDh7
cktqUYx7odYSLJ22qYjX33WhJ62kR9mt8mRS0icxu8syZLQTfCLDCCtDsgjpNYqdqectmL4Ty+CF
GSUL9iZCbyyh8SYYZJHLpn1e1jdJ0CsymefIK1Hx+Z3UD8PgdoHehEdzSdvIr3Ffjvg7Bj24HPnm
SkY6RLcIlMkT54NnWoF+MsJSzkmjZ7dP0noiwJpjiYsrPUfn5m+nB3n02QiqZ6CBzjmlDeNtiz7G
NXOE6Cu09ryZ8AX0Rq/UpGHCyl9UOzGNwL6zGZkrxbuml7/w1wNpl+bBtlZ9TjIOT+InbEjzRx0d
rG3vgcMqjcA/rpUAQvFVLuZg2qszvrcFudGRZDnpu90hkCRrfozSpsmpUxjLY80rWjZWOHl77UPa
fYwu2rhBsMcFOuJh8YbswS2pMnUurerAUm9a4er65RefxI0ri5THilZLTuzrYt7pc+Wlwnj+00aX
xTnIiDdJRMxnjVM2IargxQKmITXxi4fSGuE/q6kXxaHo+qJmuiSSCPFDhefUHsK2oNDmxVTiw3j8
gW8ldjTIpkYU6Ufsj/h+iBrWnWkw/6WopCjXrEu0e91hYFrE3CuOh9yzfOyPcAcS25VTOKylObWx
Ca+31QNcfZwS1aEJkU2Ps2nQSyHXUYBy065QgZOo++285R/22HL1APpo1/BW46ASJ8Au8u93JsFV
+Ehk+zR5IaZeUQk9xdFglbIS3ztrNAO8iGSf7MXMws6xmmAOZsXGS4whjwYcZJsrYr4MTgbjqzBD
M0Nh6kgvzzO7Z+j3B2+9yQHm5RLqgudL0qgFWB56sduhBRRdmzqI50HBHv0K6b2iSOHq8f34VTgI
Q74nVXNu8rGMuLfqXlCDimMfzAYnJ48C6LhYnF7oHIrYz0dLw9zylSu4avyn3v5ZuWfA4J6FhK/F
09HtNPtJ+tfNWhpjXqRhSkfjM5cHxcKdMAkUbMgi9hKJfT8feUeKwT6WWPwY2Zcgj/mGJp6A80t4
59wj1ysvJkmybC+1XoRqhNIVBIqw+16nZQti+55tXUc2nHFaHEh7eIzRZSxdHIwTJYrfYMlOwFeb
jdj6/dXLsbv33K/+/cMBAzlqUtFeDqP5GlVxyQs5N/fjCitxL6tklj/Rh0IP0js1ZQrK7NeNYfKX
GiOAWs+IlDez6LpXakK/a3j+5KiVmEunzSJlTuvRCPebJ31g6SABVCsuiyammMDu9hPxn82T21yx
dActUDg/ncALe7sPAOb3ax+do3XrXUG8XClzcip4qvwBpRm40DQiPZjALQSYsIkaVosGmrCymD5b
2dl66xtC3a8POuN1ihVR4oFHFsox2x6lqryvUxnr42yJGQSP7N9/aNjsYs29pZr++Q3xctKFrSGn
egzA6oQ1pgH/qxUrdyaU7ZoQbhbqKJFipFZg/P+maZ+jZmC8MApelaj/NHJ6NN39Ccc4+CC1lFVW
Ni+Qm/i+dPeBOXMsS9mJTGMyQXhsENpTPyphSEZdx675L2Ju5Fw7CAAzWFq1HGU2fnp6agxLOF+U
GKaUvM0TU1PY8deseqAmNj+cM+z8YAvww3QY0VjWzVp6FcaYRxCti0K/IY2KAtr0Uwiv4nlVVMLM
wCs+khmDHmHqEaVAgQ58OTsv5iYJs+x7fCppQTF6PSSdcP4M5vGAcn2V3tRg/4t8wjScqILmtCHP
VCTIvyU4p/m5+97aDu0qskiNS6+B8O7Ui2XbeYAh+LRvtroDLAClCwB50isxIVzXUwORM44UTLNg
vXSPQgsEOmdAE5iZyrWSU4T4eCyLSyo4+Ikfo6F0tnynoaIwgN9uAKZs1JSizf1BxXSDFH3laM6Q
//k3mcEY2vC3IS2/vtGD67zH2B+tJh8Q5/LUzJIuv6XjVHGA4wAdXIQTefMm8qpKfhocBsJjby07
RbJqlpb0PwQZfkN3kDUDi1tr+7vin0G5OvyTsbAcuKnw9SQighNpKgvaI1rlyTVi6z7EJM/p3o4f
Tr3Nap/6FXLuRafeQC0sypLoUd1vvcR7TDZowkuD6h8ZEk/O6VEkMs6KrFCpCwyAoag6LjZiu7kC
m52LRfpl1Ar70fNiwQvGTWmyPOezWbQQqhXcKanRq0pUn8dSPFhCEWpFZwZ06bMhR39XPgu5Nhtw
9BKAZjc/39P2xBfsswa2XhRsPQum+rw99OFJEXQlwXVDEfY5oAfaT90C9KuRxoxbGWVwKMI7PpCj
CcIRGy5hBJ/O/RlrW1Sbyo9YesevbJLpj7SFy7vjaXWtv+5VqFFPUkJKPpiaiJa0E7PsBaYKyvnT
kz/n+BnpQrCrNqz+Jb/0M4yEPm1jkutrauqEJoBE44+9olfrBdpK7t+nEb898uQIZuVJdciLTJr7
i7Tqqox3x0/hLUyESgsvqbyYGOiYyxA/WnrWyhmB9dGQ54zNMsCUbEIrRZSzgbTcqtFTSIoXIX7I
MYp4mUW6Ad9AuxFZVwQHd+RfAWyMkpZ4sild+Mj3twsG+4jVSrYf3K7Q5rfZzI/C5zccAUSlGzQL
CKQITSt9XngYlxF2QCXWtNjuD0VvwXNnNZJTIekRSq5bd7jQber27u/46ilYG99VmwTNZQRDnAth
H4d4SKfCsIg7HLu+qwYDFkeLCDeGoDq/qj37szUhvp6QIoHRQJk4TknLTdfCyM/ImQUNo91mvwJH
a1XG1zi1UNPM/gJ3MsA2HZaKA8Om7xbYb+2EojoYRzmUOaGXPuO7kZ9av4tJ+sjCBnhyVlfISraV
Oifag/AwivgwKhYqcX5uJHDvixcIGCudSuk80nqHV2lkJfpi4Gx8LnZt08VFAr7Ea9hqmmSfBaiN
ffMzXb/Oo77dvfLmTpl2vB9YBsNNf4Jy0CatZyFhOkYdjGI5iNPRI0sHn3oD+j5N8PZVNcijtSal
wTl8vKMew0XciBDmPebMTMGoPZJNIFI+aQFgveib5ygqRekMke+519X10rpRO2Fegcr+fcTAZDoO
F344+kqbOWHJwgk+ktGxxH+YILGLjZNiBNYji/Y6G8ht9c0a8phvQQBBLHtuhNojWjuDFO2LQQfn
A2yjolnbesNBom59gyGVHwjhUOFKTNb+9Qn/p8MQutClb9848iNqkCA3C2oaBOzucGoxzHJ80R7M
0MsD6UcfhaLdEHigKKLAOLLujjLqKdWKT+Ap7JRrdZDlE+q0zJqlZtwSy0lKUR2ByJR4xGMSuuzn
o2toTh5Cktku7dRyYNGzh/XVHWVDpUq+iwnnLzcKlbXAXS1Ls5JEcq69hCxFRFvSsJlv4AzGBCEr
BAtFE0ajYiPC7tBmVWAe6TgbSgcSLPa7mv/vEfh8fEVWtgkqCz6cqXbDkcDZs9Ouo5vNQ5KO7nX4
OcQIxRrBUPNHEvN4tJfB7OhicNcmYt8BP+WfD/WHrVtQXN/uRGWpfzcRiZ243HM1LcV3MMECMz8G
yiZRWH/Ui0AKN4Q0dhOfs7/Dw/QIbPoush6cR0QLfNjdtD5DeG+sOchI5iqPYcY0OdBu/9v4Io48
BPNlTmCJiYJUi9xe3cJEJjtmEDo56IVBNuZ33cW+87VIwEskDJp0XQ+PCopeqn8gLOypJlv+i6z8
4eSIxsOB0g8sIVgKkbeeATg+gYkYNdOK1lbkyRol7K7YP7AlQFbkYE+YQ2CHm1aSgPn8O1B/fPmF
TCo9Py7W+2VeqCPTGY0mmCI3WgGs3VO+8ILTPMw2EpKUeCRfX6Ehug2F2aclCGZ0UKIrQMTeXXo4
wi0P7rin+6u8ytI8n17zmi23h5ImLiE3r84ZB0xiw+9ympfWujmUG9z+sPdNP/O2Pk6Jc5Y/OUou
g930E7EBgUh6KS7JW01hjUuAbU1hbVseU4KphsrBHntcCq3RaoSDzRPGbpbuv5lJgQVnzoD3T7DJ
eMZYkbu3jrErAKbDCNwtxU5aDL5bgFV/Wt3oXJVDVsnC89ZftEMQJbxUEmzLnvJnHTKfE0QVoYC6
lmzB0olsU2/246PD9u4SIlnqTK53l0i8B0vveFvZFIGbgQkAGY9ZT0DsJwNB+d6Fx38AXy3mOD2j
Bsgm4vJtZL60Rw1dUxZYCDu8v6UZ3MaQhxIZduCPuVL/O8GlWJm/+ysg/CUZmXj1+fFKrE3wEB1l
q3MZ1RTS5J4AjRDCkBS/wPujgPtiIzzarEPGQT5O/jDJteNKDzq/bj+kidfDPH95A7LmQ1TdI8XU
ZRwe/u2Akh3YJ3DMNlYLsCHMxKe2+9lTbMTNlNrxn8KXd9j/xbRznkv/B4oAOAp4NRIHroHOJzL3
lP5bp2GWVljHKrvbp1RpJljAdIBN3PlypIUdYT+9xsso5R71V/K5R7v1K61ZrWHosaxkgur80YGB
m9SgJE452vb7EHUELWr39xINnrU4qhAhGS5EUorn6ltNPwBNF5BjUuJIwB4qo45Ry/NgOgP64Me7
+3XoWDzq57I1BNSVVAssAkGrRlgEuW1n5luB13ta278LzJs2oDMauYD8jKmusoEmP+42Z0Guh736
YJl+LeqdttbnZHDkizySdVKt7A/fRl+2J9eAP/363oFMGHlYeuxAoPszDseswOExqzJHIvOLh19q
/xXFYMuGhjqPsX2n4wjlKaHSaYbt6r5DBMDETlrofdLS7IAS8/ohYV8RcSNFhDCnIF5ExYQphsyx
HsMohWWuP0rJzvBgIRoN25mRy4kHDA2qg6ue6aY8OYQXMq8mA02PF+C8YWP+kv+ydr1M1pLG8fXN
hc+Y3BxQKbhGG78Si7ZhoEmQTAHPnmw5iA+fnXn29RhGrHFc87wOFMK3/hOhzuHyHTjYXKd79bDY
nmmrCf8faU22V79QBuldjU1IArowbPrYjYB9BgTzJQr7YA/de9Hel5eS+P6WUUoqC3sOQQJoXyp1
rCRgMEIROZWI0/EMJN7UBUF8UJxm6Q1JLVZt4lSPw46N8fzU4VsdnW2ZKXwy6wQ2/prs4TFMTPsn
WuLcuDHduyDI3JEc0pHGWU2iiu8LYK0vNYAVXpddsfEE7LGCK9Daz4mcNCKpEAVR+kXTGHrkrx0w
SolSwzM4NQcZ46gthwousxID04VeazLoGE+9cbd322JftPG+n7BQtrwiNcNlvPPIJLHxFomsnqRe
QcvZ+p/tDbhVFqvuMB3OGBjPPZ/A/JtLcfNkH2TzbCfm9VLBFGbwZ8rFFbsa2icUzaH2APIsfFr1
K2ZLkWIlSSmpM+k2ZRdymAhkbGlkEwpNZWwC+xFQCKvQBLkE893iCnSruP3FZ+cSkj2qKfRXdZku
/keKYeqoBF/IFLSJ9piAqCNzEcdGdZzf3aPPPia5x82ALIpH70MDxXPtq/9ArtO+f8fhBrz3fb5+
szrfcUyoGM+CNj5eLBiottDCLrQ9ab8sOPbz3YQ7bUkuRZbK+bKZuriHnNQ3H1eaUPCNnREDuQ8Q
y23ymJNWemHdCVEAnSsjMlV0Q0zYDclc/OPmeSMaZmx6coj0wCMdNP+UcYdn+CTkbsP5Tht7noiP
E605On9P52mxdXnlqVMTtGfiIfIQfG9E9tMWiPf1kk/KVAKFvRO1nhCG1B9ubquZ9CgZNxHglF9F
DISCWvmDKpxZAqQrwv8Wv0gpZ5tDWqdFc+2QSj8c+EFiD0n/3ndZ0RMJKXEcMyb8biLmeUDJaouY
5U+G+7vTAg1bQk1KHQaQU/YPghhOeYB/wwBpaPlCrCVLuWGLVeJAhmwSLpTRTOiSCW18X1wAYxat
jrJjUcPdmMtNg4gse+6qrKxOX2OqY+vmA/JbBJ05CTw/kOk+2SSI2CRl+7Vu92ZrdEYnkzcNxgXi
uNkrfkkXbkdntkc1/hGD+HT1uLGucO0+tMITC194Xdsr0Go8lC41tCeZ1xvxBCA/5QpQjG9olU90
Lhkpz50309m8m2O29IawHmST49uzdGcALZoOhpAVkCeJBwew71uV+iJPEt0frF6MXisH5eJPbcOJ
B0cN5NvbX0Zcdg+gkSYrKQMPwKA0UQ5/fQkNnmfGatvMBJYDo8GqfZm1b1gGyVQGEqR76tSa8DTy
ehTkDFPDMiKrCuTkn6CgMvKrGGMPXRxrSgVtu6/LRoTnq9kaBkmlVcqJ7G6QSlxMNp3v+oLE+j7I
MQp/V3nVagJjts+DAAtwo4Dmb38lrZwOmwc8xrvU/xLKteGYGSUaCou/1SxBrC8QurbKEHfCYV5G
OdrJ1Cpj7nwQxGpQDCWH+5aLl+ntGcIEuUePj2+prcgagi/B1J0SDPzZ3Ai8r2y/hIvI+y6/9Fnl
cK7u4Oedw9ZKM4OLzlmzGkhhUvhgrZK9UevZvS8yqlwHInnkPSWhlEeDN265xGZjCXmr7AaPQVvA
yBmWRFttilVQroxQ4m9ap1vY4IKeUuviygUDESbUlsiBXzeXTb+yHIBY/oafujbMfl232TLuWkPh
oPsUJwcIGc+WqSNvg7nVPwoMWv7gEmeBSTkaqgzRP6cy8++WtOyX/YQk/985/9WwAihPAor8OusV
cmNrBooWmzIYBV5hskJ735ArzBTfbf5iyvwm6uF9mKpc7qiyo0AVdlSCF/slL+ErMKQCjan1r/d9
xtRsx/ZX8smPHX99P6GKzOfQCvcKTlo0GSH22Zvj4a4WE9DwAiNj/Gbl39ryIMgTLu1HruMvLsT5
ewzjMEiLTkWUKfALqdWSMXPn7EyfwQFb//yh1jyB0JAj3ZNjSGZvrMcb1BeMwltsrGkiK4H+0a5w
KZJ7bC5bGenac8AYHx4LRS7Ta0jevtvYSgzYkf1pmfr8y8xzjoOzCIqkgz3Z5clOAmTd2KRB8iUE
lErBtKezBnBAOz+Ma/IRxCQx2vBcZnNPZQr5tFxgs4gova/ioK6ia1F+VrB5jDnJgDgyXnJPhR+A
J5mUehuwiben6Zi16z35W16vfvA5QoDor7NAxITUs2zV2UTzQd6S0uaivSnzbGhVkpZavw7I6XE6
pCjSRJo/nAkvGVlZVZ7uwEQCTXv37OHsUZVjQbQnjZDs7KN7QKgrCYulvwisPiegbc0Cyk+hXOty
blSth1NscziFQpEhGG6xzqfx2MjSbyoD7O7rGhCqa4vXJGUpaIys+9in3KNInEsIKM+b1J8fPAKq
et6LyQiZdrZy0+3oIiN/5rVj32rTVUHFoG66nqt7lBgQPJ8mKP5jmzGEArmT1Koz2Um7EOnJqYkC
ia41mn+pfNZBr+FFIyEB4GhhLh6Z9nDUcdq3HTzIz/zv+uTudwWAUccnS2UBSIYMXsBB8YWUa3Y2
my1dLpBE3aFv96UlN3W1sOtZfMNDJGn3iu/E9eeSfNSambfZPN9gUFcHdeMRgTbQq72PseJUyeAE
bRjaAQu2Zm+T3HswDlX6r1xlOtUFT6biBGDnJ4FBEqMEMUpc7miVQNVKi41DqnGJ03llVzoDBV5c
1OylfQ+fly/E/2tTwr9JFnUKnNk4TsqCq0X/0qDzN5ecIEX1KOLJNburIiRo3Fi7KVh+qxK10LE9
uWOufvKzeLP238DV/e2EubjVSbAJI3rP6aR7wAFFmpWUwXWdWTFnRvNyS/Oqwh9FD9y7/HY28WgD
Yg0Ua6Qr8q0kudln5quMiGpd8zFKrw0H3DbywpXI/eOFM7Zph1Hrlsh6uXhMNAmOhATKUNiYdaV4
Nk0CudcW33ba/5Rrl7QHSp5MqsrucgcTfsx1Pvue0GrZ5ptcMnewQpWRWcYcx6oYl/eBU53na4nU
JxwQr0AU1u73q8myxOmFGxsk1wmYrEjnFG8hL+Djvm0aYTlob0dN1AJ1CR+tz66PD3ZIf49NHd0T
TYqZxdHZnqnILgzqLtzoeFwQPXfGINqWU+JzsGwXQerv0EvSxzwL+oJpoXqmdcGAPK9T04IaFtcY
q1hcuSYJLZSzNL40WSSLwv9UiDT8X5Pk0xCrRErkG2kVsp8lPnrTO+y3Qv8bw73OSnZiY3pc6PBC
fhpMuwt5BONFi18IglWXi2QeG8lzTKyvPKiqqOggMvaMR3VSwknAUs+P6mbcJBCInjyujUsrxRSt
/NUXmaXL2aRcfeyuumOFL5BddA1DQGVC6oT2mZGC4bl/Qg76O2VYjlfOgBf8TdAwQ2U9gaWtxgax
dWDQcfY86I/0dxILosllVgqOlQZAYwATcAxFyeSEnwDKiJex5EhRhusHNnH34ZJW/+nyrdU/8VnW
52aTzWwUOQYF6vHXrHGOsrtbocaG3m6dbDN13EzBUvtqgT86IUUXPIwNMyD2LMfL4FP5He+X7gXl
MM4cm7lODDDTRXfpKXAcrhvi0mYRemZ2w6qXM88qbVnlLFdf0U7itR0iE3LuZt9HmrxFqa7Mpt84
HgwkLvnnWd2OS4OfvW3LIyK07XxxQcxW60esZxVtzY+QnVQv0RHL3oPKvDJioUoTifi9Zi0DB+Eh
61PxSHticwxhzcvIKMMB3t/+OOM43ccTPvpW6dP2ToyHjSOTdkGxFNj3ZM+1Bp12gckk9TqkUCIN
qHt0lNShvxLcqe3WI8b0+cw77CfgsFroDIbgXZOZjnQLBhGOxvgfoVl8d6Wof9TzisZWewlYLrQ4
Aprg41vHxM3YqtmqIcQTXSEYWSsdjtgR6BMYfoDDRIZ3WtyRP0up5PCKUHk2BNyEsO8h2fy1EdEr
MKHtMyBHzBBWiCBWJDZ79pqHIqXnrKH14oNsN/Nh304G0EFGeNlD543tR3MgCsiez8XEeQvCPVUT
rUY8NamKRCgygsixH5ANtytEn1uBQhp1nTAk4epUla4VxkC3GUcdv8mq+3LJr5gZOyxiXdsnzmf/
0/8gIiVfy+EOKkxjIYJxrulFUgaGWMUCBTAD8FpghT7TdzY3kUNYQYlK7qVKF4kutdbkuDGpGQe2
mhzBlW9WIWdEY9PNMrdPE+PUn6lIE6lJX/2lI0K6+4F8Ir8179CGj+JBj4Q0wIJhRgs1HVLDWduH
kq6o22GV1+A6aw61NuAe0fqj6tN/cxtoN6yYZd3AHYyO7YYV1gzrVEIz2Tp6AKRr1g/hopoLNX1P
2Wl7nzDEFFwbrDFS8YvOqzBYW3cpdJbUcZQ9yBsfV9ymn4ElVpu4/98L4V/qfb+SjZxjRYGBXbbw
iXp6o4pPlZAatJ/BsAlVB8aiqKLIPgAw+aqQMIZNo+josvU637vu9Hb4rZjLSU+dX7eTazhBaclI
7szhj6GBXyZs332A/X1u2Hhlf96gi1RAqBCnv/bjgvRB+3dypVK2IsBKhAETK0WVIiNrGtsSSxQ2
BnGD9HEwpdbkgOI9/4vzfWj+KqegQxEC7siKJL7MzRUz0zDkRhXLVFL/O42yr+JRPA7cOkN50Cly
d0hXLDO8HdKHcW8nnweNrZlF1g5QJcOtTAIrDzQpJcN0opWIm/WcNYpbokv5sfKBTGt4hVco9H7i
K5ZI4r2UjVudrHy2XOD0P9m6YRjkdJAt6R7g5qBJpmS0ygMzQIrNGmKsjsUIuh8NoWf7MHip1CS1
9AvWtOx9K2DWt27Jb1iQfVcDKJF4+TDj2kOCS89xR3uw5mkYNWpxkUOAW/U+d92TfkeXEVU4hrUu
MZ2Y8NPedtZbPARdsx28oHWNJAB1Sk7tBKHFYE3TPhDgzGI9bbdnK1CNC0H9joLFErLG7DbLyRQC
Mtc2XrSBzAjybeRqEVI1wNv8PI198ODJ1BXoUXraK3G/HNkt0OIhB9wCN3N2fUZuiOVEtBlVRARe
iSV7KnS6P570CkeTBAFS876S9vlYtnmlf7acQ9adnD9maLwIL0m9RwpLLerDk0PJelPgiDJBM4Fw
vnpwwhVMYz2b7V/Aibkcn64LWEs384bt9Qf2wX3o1oRzn9xNexROVnAioSt4PQvFxPj97ym/eoss
wIRcZ7BLyoR8TrTEN89noKeiTrSRlDb+EwsqCfMI0JwWHtcUkzb3NyXaherP/jd9M+cIA3u6Stct
qOQ1gJ/pK03aGcaPv01trHzWU2AbeAtBNBkpteZMiBgSx9K88DF3Rt0RXkWwbfMMAfK3fybgDr4M
FmYjGEIbletjB4Qnq4AgEq3fN1ZyzL4E0WcO1FqiFoHL79GtJiYfrsqwIz8F+eyOmEZlvenjwLKB
41RY8yfaHA3Ywy5vC+s7jXIddZ68bCy4b2xASaCcZEckUGxDA4hkD3P/kaejv9e0ORvFtQPEFpCe
DtCanDlr2CmEi+RwSQ2NQhD4FmsnuVL51kPeD7yOwsj0+exx2GkDb84QXl5JHg5TTnJYn+5q/OIb
RZT9sAJbYBHmxABnLWW3IluSmTibtZzYv8RiF9o9zUku+50Wx5Trt6Rrchv0CuA3llkzrXlmi7oR
xcEGqlcqHMqVozO4OeI2quACrh7KB6q11JbUX8D8n9H2k+mkvWsQNIMX6aSrB6zXCdznJ7gFijsM
VaW4v4bEyLcwTwvBrg1vBawfYvLKBeNwZ7Jed2C3RQjgO3Npw8AAQS5+bjjntXJQAnQnglj6E4tn
tor7/CbPkhcaqSW5EfLEOzvPwy9ak28iQkqB6LROQWuwq0clMHAHjLrcjH3GNr6dslIsbG2A4iFh
Qpj0q0o0x9pVSNPI7+EUFWTO9I1G2mSHBHhy/G1ohXVVyUDTFbwjYKQyX4Da2OZ0mQ86XSfvBAUW
twdW/ebf/+lV63lswbGSt/ZSo8Eal6z0un/cHx8+SP2GFR8UpYgci2VsHpR3gw/uMSEW0KJry5nQ
zBPq+8a9TSiyZ61x2B9KFBFOqZ2od1Rxqh7bph8/3tR5hCmMkWWb/4caf2aRO0hzjtz5dverlID8
OV4AG8rEOrwLoTeS7pedpyM+i8OIwLDVYir0FzNE0FaTfAdWgy54VLhW5h5oxg+mqiy9g/Zm+6BW
B3MfMLlqGnyM1LsdtoW6Cus0mCfX9SkJi/64zI75HOUYp6WzdD+nKDNa5a7w+5DfRfcvTU2u/i2G
FCRIZYonjQ8TYX1XWyuaZBN0nXIa9/C6rwaciMhrUWseNsC0BfZf6g9m4/b1umD8Z+altP9YsDA3
D1qpAHykKW0BdoGobxc3FRBEmCaxyPxfj9R4HSZ4mqGiF3Dwffzb2QyDOzwMBbuYzU3vyBps1dG9
9GgubyEiz2SMrHXgLf8CazGGSfuq2ChMg6KAdar/zo0cMTMH8cHBadrSHK7vBh/cLKt7Xf+7kzRd
M3ahSnksQZw7XeK7UAMTuQG9Ckzd9t56a9Mo5rJEh2zNNu6Vucvt+Q1m47CFnYTxf6pOOVEVFvkH
xWmESvRKUl9mkxF1fyDEOls0d5tSBC7xcLgAD8PUAOy0e56+Ez+3z5IMVFylYl829G7r2vtxJT8J
hwjcL1vG+y8GCXLS+xSPVmqTvCQNZboKDdkfQjI3rgTfC3xIUaS+0ON7FKzlTptLy5aDPsJZLeIt
PWoYYc8Mci4VxkeSI4AhPj1l4+iSdfWGB0HEFB2QjicY3leoKwsh6Radt56nKiZgAWio3McNMz3A
oWHSPFuhq2HoYxSIgf54gRHkxPB3CopuRiWOG4OYtpgjBZbg/0vvG0Lfxs1nazBGuyzau2Fipv/W
Uhe8JAmee0qxNbdVfBub/gDD7OqZDlqvCWeFJHFMcEDXcfi6vDOGET18T+SdVeQlK1oSVCZJgGJC
n3ML1f80T6vBzN4mk7skBU3zMzj19RdJWSGnC3m068zsV50RXZ5Ek77WSvaUoDl3HOYU2SI7pW1i
eu/4ZlfXSTfP1++1DkLhqsE2YaB+8J3hb8hxvgxSPfB7PuLXvAUffvCiP+wTkmduV5M3ks8cjERp
Sq+hujkoAP34o0Jfc2eC75h2/ZQ49OMlqu/6IZIWLpx6n/U02ToGn8hxIwDvc7DJs9cJTL6cotvj
gFjZo8cvbXOCRNJ695cMBEToZmi6YnpQqWL4OXEWVhEV2EP73o8ryI7CvcuRKrDoyFFWKH7uF/yR
qcQON/uSI61ZJcTIn3iBGd3BT0DxsBcph5kDAQ5xLSJ3R9uYfZzz4ZzPHoHbFiOOMrQ5YbuHoJ+y
O/Bqzd6nUpLb8vvROgaQSjN4WJCBKPtJ/ZkqM/Ak3ojm/b3A0Kzm8YikTBVntvqvbdPNW6B/ErnU
2W9s1qx2b3rV2QO1LHJpp9MotSVKGOOawJt4p+QjWJMCwsUu77AuX/tekTaVbrKAVEJF/oaFsby1
6eBO0vZnL99zE0GXkmNlp7L+R4HYvuQyDtFgd+LFon83YxsnDuqYHFWVaEz6YxMk4rnNWJdfAM1I
OhJjlg+/oSjYPxqa4qNJT2wItcI960Y8z8/z3cvalWMwLz7FX1jwyi2bCg7+HK6d/RuAg+aWQNNC
pPN7TIT6MmWqo+g+mIIFuaRCuYlLEPfxlE0pkWvlwevCnKv0FMxP73K/z6E3+46sxZv5g7a1S9S+
uyyOfW/DnmojDXqYaJ3NvMVxLVIVaUAz+u8R5bBoAK/bXbKuBCGsoKwJXZkzPcfU/lzSyFRqvjEG
F8/H1gAWOfPiPQWnUaSAiM8t+U+kKfADBVbiDSs9FgdWDap7UKCpcVvr/yGyxInBj2HHl2j3yU3D
gZLj9kk8/hhbmjowgfEC+fzO+KrKwqau8o2GW2v1HWMi6DhDFtzV6/9Z3/bymrzfRisIPN+37v1J
evE+Ya7+VHPW5uF5w+ebJvmgD5IdusZux9HXWlokxvy7V6YIDKhHExgP9pfhSHpJxFZZOOGLuinO
2Iy1oOm8bm05eXve5y4TntO8kmTMCXa9wn4GGl3r1UbLW1sn2cntbtV8tLzxwphoLhqZ8pdeRBi1
5c43sjqzL9xP1m5QFSnWMOjGEM1EZdiF/VNBsYM7RdIA5coAIcsGl+sFXjd0DcKyn8dN2WPwhPit
Ds5cLJ8lxf/I8btYtQIs+bjwzDLLb4BhzGtbsej4DjhxcyrGZmme6i1mZxznh8773zYarYKS9rd5
fzCRrzJy6MR3Mg2LgIH0X1FviCGSuiyOsS9XtLqEvAvC707RZwiuf3wH1A2L4e6loxcK1gJCt+cZ
hDzDuCNBTHlSrL38+dkrPQNhW7wkJZiuPOVrpfKRWpiTo+preBXh8KXPW2g/N9FUsZAM0YJmZkVM
ReJgg0hi5KZly54356Z/yMiMIfeCDJn9X6Kaa5xtr2TYaSC880CLxuMuf7TNMqTVX+kd8Kxc5Tyk
V6eM1PULDM1OcJYXNS1N8JymzLl5fuxXRlmXS4TSYBNu3TRRyU9sCkRl493iV98NOrVlcyvd75Im
oSeWfb3VDVovsuowxdYIAV+Hg5RUBE+I8fujoxnLp0unpPA8pNdsTOWTKfa8Isf8ZWOXnxpaOTzt
avPENBSQUFJuhWTbNaK0muEbhpwb7N+8CtUJ87F8bBAUlQ8SCsbr2S6Gpcg8GflFxBhS4Q4upULH
+rqCRn6q2tH29054nEeMAgC1fA6CQpvo51zPOkvPXCqa/bP3sK9ERIbwqXUXGCwEi4NmrdG2H+1h
UzvC72k/3yt5EM24GN7+i9HkGZyGdOlIK2b/Jk+QzAWi6bluiLr4ej6/U6i3csilmED4mD0By5Qu
cjXUChqeUrFz2wkKnYuU8BHsDs9ZKMX0ZiZo5rAGwNqFVb2pVj0ZWwyKWh+8wkRP3jHN+Fv+aOhU
oqpygfuytscwz1OUheJUxHuUzHuj8/ANjbXKwm99Mz2DfG0uo5HN7vYm2c88ns9QYFr3B1gvoa5b
LGzxWXJp2UfXdv7vkxI+4LxT2S/yE2e6bJxZZaE2FqVmRxtvIyOoNK72IZ2erYxU0aZtYGG+OyoL
7nrq7SSW1NdkbIukuNLLeHgfeitkPmZ3XbSWM+HQeTn5szLk9xGf5L2Ul/oeIsRJMZs61L2Wiak8
M3vWPPOvi+nhfgtBLhuNpuyo1T+MoQP6QE7XWMJxs6bCUgg5gGfe61UncuaOigATH0bkaTP4nJWz
pZlBu0DcFXwHBWrh8X6b15KfmVb649mKhKE48JLlDmn47a+OPRw5FzCit0+XejWVW8hyVqPZUI9G
CpP9QDc8G/B/Sx4JWIkaejiVUWbhLbqQm3NTT+SUFHE+CBqJ0KrEu4o/giZbnS/6WRRBoQHBnQ6r
F40KGC2yYL+tMoWifPjkYMb5AB9jN0VEnz5MSz3tdtgiH42FQYQXbmy24TUzDpTNqcEUssvNXL6Y
MpOmcUx2uxL/U+EAtOIwuiztMEZShjWKGeeel1NWsK90hq+hv6UYtzeEBzUUDEvLlE75Pl1Vj3e0
MXsvqll0UqOLzrqpfupmTOkALLSDjiMRJEqytjQI0Ycghkds5Jmfho/dHgWU80AnOC0lsu88K1/h
gn0FWbsfO67+ZRnYJiQlGQgKFsCHRmlqEFHa++VNtuGKOjfkTTXfEoTQEvhpDBv0ihLHd2y/AmS2
ypKvF4a9XShB9HMWLTQxuUCG+UtKnbV8egXurRt1n4CQvpkzAfj+70DLUjFpV4WLBaiG8h098CFT
gbtLKtMDQPXo7v0nqP0pYx3daOiYIh+t/OW0TmnKtAuOamf1R5Yj6WKf9qFhxrh2XieSJ9iQY2BU
eapP7PpPOMfjJ0m6ey4KYgx5vR4RdJL+F+5Kh4vHTwr5Ii/7v9ffmQP7NjsNQsQrwnRfnsCHpWRQ
Xss/tVz8vmT2DciKF01SIcBNPA0dcBG22f+EypSDjMN/7a/WlTNao6Qwd1+WdrSuhlBO/nS2Y4lM
oDa5cE12uK/TRdYyIJoVJXzifextHi2Y4v4eg5dnQlgNd3tDrnqWM+n0+tQK/5HHlmvcTLs1pKKc
iAdO5TxCJQiB7Dqe8lc0QsZPDc8HzpEYLX3eE1356wXDF3FDYFvNe7jyxFcLw2I/IYzCf1erlPnM
tMOVYJgJct66X//a7pF9KQoakxgqIlT0yrmA+bPygYewHO4C43vu7RCfMhVYJWvD/k66vH7s7bT7
g7rqVJLQoNbnNfnpgZDPXf33iqhlutYqHsC2OFxJ3l3SGIUOvXBra6pLd+cbFClSdgehSnqhV/S/
HXttCyQQzB+GsGvWnAv4Iqyj9l2Xnhu4v+XBpHdbZjnVGgCUJIIyI5Qs9T+/LBNIM/4oUdob5zj4
mvNuq/06gO6ju/I2C3Ufv+dsBx2Axhd04b2bDc8L5bapVC+5NzDZ5cBO/7IxjCl8Uiw81XDfiieV
KTc6W8ca+RJ08Io0plHvfZAuz4tkEAa9Dj21l48Pgu4b4DQ9usmBV39GlAJ5CE2JJ4MXVwwobuVI
XrqkuVPxa/xaid3XVVuJg5n811xqoH+wPY3bTlf8bMIhiJMwEtxwr2k2K56Zr+cZte2u/uR0Zu9r
Rh8b39PX10hWfldeU3KJSBudD4aTVQDtdvLM0aIeBnwMcsQsuYj4V5tdCMU2JqQYyL2/aU4MsBOL
Uyxz8d1Se0MQULL+Ne4/tsAXaQ9e3Kaw8MtnN6BsfEbmBqdJyve95exz12olYPN+mHUQA5FHXkuY
F5tbFeGO/HuXHScxGXDSTlVWutmyUdzt963oXNtKFJ57IrXKdzOjDAJ5ryvfLsVtNijPY9nrqMpo
6PmcPThco/JbxUAKgatnjG4IaNu2aH/D0uWD9K8pw/L5cCU4uQZZjS8gGFKtQ1DpYwlBk8mRavou
WqvjsuZDyAaJtTYD4QPrxzrW2SKlOOk4jHqsOGWL5V1fWtTo237yPGeQQTq8jUoFwR4gvXAFlj72
mfOsd60+hDPRpWMFZMOjg/m39aEDnExoovY/WnUXDvDj+gfiqf1727IqztrqvMvPHDljujaI49f0
tdhH9m+Sc5e9UemfuarOPt+i/USGxS+z7SeqU11clWNfjfK5WfoEEWhJ/0p3KuoueDCk8+EULPAn
+HPz+WKWZyLEq6PZp21ikuOi9MRTROAs5XOlPihYmig0ni5uN/QJOritL39Ytv8zIlFW25ibRzbb
0wd4QvEOMvOz9XPITWQjH4fFbdzRXLICeDSzDvgGFfDgG0f+wI+Bb4yrNgUKKPqVhN5SiiXxAH6b
6MkRsMgrt/elEHKzLxisOcRnq3V5xDrXNyD2dcs0TjTKFqi43bwm/PqUyxCPOaxH3Cj2hpQMzGGX
tJzsX7ZVWomKfE2Geb60Y2JeQmWQBaADq7qap3HuGywwsN59KIAj07yanovG/HJ7RvrVxh7fuECY
Ye743xwi4fSP9lUdaPFF7xNWpHbh6/icD2VPKk+s356i0CU05ffIc4yk5Tkfk8SmallFs26iAo5i
hPP9XS58MY4nvKll6wUMfqKVpq/6mp6Jm4TuNi5EyOjjqXtOXeYMlaPCQLV6aIVjpmm80XZb9Uec
ms0c7xEPJJ2QqMcbm04TelqoMrnQns+ZcwAiiWzOwUEYH4px7kdEijoFtI+kXyjTsXfZlAfbSKSN
ZSybpwMPclTdUus4/ctKvsIGmSMKwIz2tY2otEZ0a91kXVsC97SG64RUgkD2Nn00PLohGkdySHsp
y3TaemV0GMHzb8G+/heJu2RZ/qlIIu1JSo4+pJUxcJcTc69DLIJ5S0KAM9Nem64NiUISBnJ2e+OM
LBUpQsaj/bsXAmWXem27bYGhMaG+itGz/3Jcs2xu1fhmQlKG2xCdaWcYWTL22icYh1LPjntQwIsx
+evlb+TLnA71MRC94dQ3wcXnLu0jqcZfyKvZUs4UrAg5QB4rzo5NPQPInEVtO1e7+2zWWQYn/PeM
QN9aSGetdbTtRmm0L8bMdQveYJYvsoG5opEsILuQh4cRMldJpMFii+xDN/jDcxKhCgjMFaKfI5pr
wzkM0Batko2rZUNp65VY/8YosbLjPgnHmoeL0p0sZTkYFCD1ohZwm54z0rEipufNT1tY85V+k6Av
0khBrZIUL3p2A2PPiUERtUFouUybs6w+VR7SB6kMnDTkMWzBzAHu9WAkzHwzISPJP9MPrMjwpuIg
SOJUtHtPoZXyoUsCSfj0PzzBRgGnWKEd8stTP+mIomepyK/aQQ+kqWoK396mQNu/yAw9pejnAU6A
Dz5SJQ4lvYXrFKX79WHq/lFtg697m3R6gZFAtZdRkfEWyPdfRYvwGmTwCp4lwL8/+9f0OCSuFbZb
8jpC4iVG2wnH6CGfkTIIlg3B9MxV6KoPX6QidTtYOu2n800wkp/IeGqmzXfOvCDAUpr3knd7b+KD
Spo4D8FXJIwuZ2tvVSZVIW3SZDacAy/s9zJEQ7247zQAA5b3yZW5iiHfF3QqyTqu9eDHn/AnNuju
DpNp3pGNxKQw7niqidrYqnyXjss+fNSEI6WMMUBhzuS2X0e30FPLNaMZqvrdPo4PRfiYlL8BWTFN
oeCZMxsoDbl47ewbd4n8GO3/dEdNReGZ3BdQODxr3z9vfL3lxnYwEcWLLRAIngdJuEfTksUNAubG
K9MvOt3Gk5H7QWa+yG7PvPVb8bxc1qi4u4L3I0GlqYddGedMSTnDAzPa5fQOPEtBT3bMiATPofmk
twC6gCFTFonntYRGJTXuunpzeF/EWJIaZNnwwEhUV6P3bs6kmA6c1cDRlKgNDGqxu7ArJhjdqwup
m+O8ak4usinA6rXA0XVBVws701+WW72S7tlAFW86MkJ0GIeZHdF8hS4dabER+kBwRD1V3UIHOEAx
8U4R+fbC/MWmZ7qL+t+X4C9dJcvNcCqtlTyCJNObCgJWnHcSlvcW2tHFXQn8Gu3Uo6ZX/HnfwlA3
0w+aLii3a86FgpYG2lQSWeQEqAgz/z1WbgeLlaJFEi4P7e4Q/TaLMaJSqVgvYtXzMk/q5ml2Mu+Z
gn4/YmSmaQ6wb8kzi6pLWqg8m6tKQ/iHuMzY+k2UL2SLmOpdB6F2fedeqREPKmURqUUp9K8Z+j2x
ltJMUlsT/4kh1Znmx0obNMohF17JLEMlvEH4Efm4NUwrOeH52wVCA+g00CqiNsbX0kvSxmLbZZcx
J/pguo2kciDqoRKGucssHMMCR3nhEaAqwjVNsZeuQnyHJPYS94n1/Cz9SfE1buPoOBeG7T1KwG+2
OVB2FMJOSicy4hr+tnxJLZWnTMmR+7pu3uxlJ0m3CLjEUqgynnxhS2SnzfAnjUR6kcjX+HtoL3Fy
664sMce6s3TiTdcGGkC7wCOKpssNIrn6R19lN6qjinyKrImaW3wih6xHInkJ/bx+skzes4qSBGGt
ugVMrG/O2d87IxMITfqltX/vnawq+OGnKKVEh+H50ourhQf/g3dhxO1b5uiVQ7W8VeBifhYoujLe
RFLQZ0dD+nY9H+vkEWU9RuuCPG9ciaRSpTt42VNhsrf9e2xLbFgnGiEBcOHZOdiBGT0W5yzZomDd
X9YbTogwTBEj/1o97R6M2yvDARPdOpNbFMIIXdY4/UJInGXumRc2qc2bzc89I9lJmE4y1PLRpS5R
wD6dQpr8X6mOoUbzMOmORbb3MuMEvqgo6Qs9eXxz5cYVsPELtoLwzJDjdCR0jZv41VxiMamjjBxy
n3U8MZrq7MXPjtHXl4z8qFHgFtG4CiYHKjUIzO8NDEoCxfgtNvniZlenN//teods+aQ9g7f5SFW6
D+SEOy1MO+XT33R+7arY20clZ/xE3encSjq4CV5/4PJlNSR/78otDoEa3uf0IoBMRsAJxT2xXFjd
BZkgd0j7de/jDxf+bVIabjI/yPUCbFohlP1AjWAGUdJJpJSc9E+042O/ieSzCQ3E1Xwk9SdRRSa9
X8wBxjRklQniQP/GY7T5jlLC1ATU1cm7oDVyL0Vh9dzgzXbvMCDVYpkzKL+F2fwnXhvf5VEcRsGE
mLS0JYINYdU1ilpqsoJo7wPTwFVBgTgWdrlvjVwgiLtXE5vuUA0HjVJq5KwBBrBuCIXAOHRlVCoC
Nz6JqA0BQvHhlI0e5eEMEuAXAthC0zoyeQOrk1pzgPh2tf2rrurtUGyRaX3UnyhYa+iyoHFHPF47
12EO/NUQFKpNAIehl5B2Q5OokmHQ+3XJhFlqCbYIjs868A4Mc3LyrfbOGZURgEfpLiNe1bHC/K1e
vTteOD3DXU0gvr1BB7eZ1felU54R4TcuVyL0uc4fpwCzL+uEkYv3tTGa6Z59HCe2d2ueEltE/z9F
q24Bd3GNny6kbpRZ8mRAGDAhl9SAHaug1mwbaG1A/P2P+eWeBAU/iCa2UuzQjpfSetVU4EA9sqYp
xQ4gInR39iqBhH5L4OBjz5/ATDd/Q/GInVv6uHz2nJpOHoajBHnXqZh0RSYHqvPwreQxZD3EhubU
G6sTkKCNSeqbhyNNmqUTBE834xJv2S5IjdHW7P2hWvQ4exP1iCl5cRowl43cNrOwqdz01AjGp83M
Mdlpu/CLHXm0ta1NNeAJbQ2Ab8N3fWIV3gPuGW54nhcxjXrFsL0wtsB3IixQz2Dsl1X1xcM4FVu6
Bdnzxs6i8KvlXzfGIj7q6MOOS4uuVAupbRCmkMfhGOVh4Ek8/1dgAqfv9pK+PXEpL4DypaR0m4Zx
XwR7CpM0aVXDLR1PzrJFA2wY0H+u8L6rpvclhBXXEfoiSZPBTS7vvxfc6SlgWVUPOOcslCBIgFji
3mcei4qgzWF7Y1dKGPEA84vwmGfkltxoiI3tG20YriaR/p/VwjAY129BcVPozSi9M50+sK+3x7od
KgWO8IiVMo6vwr3mTX36BwEfyzGylTTaFscEJQ4u1fI09/EbT4kvAWe7lBe5MWSpgcmE846O8ARC
aB8LhzpJMCn15GRXIbmLLY4iWtwZRCiFqo/6Hyl7rfbXyDly+k5Xn0RkPzrADUrrrw7KoXeHyzz/
pEB5lq8NmzqbvOiTv8P1rlkHSbQ7zEWDilwAxxAU/jAwIScQArTvuAgnJ3qo0fbFEdiRoMGTOAQ8
sDfYnNx4mJlGEatGBusJuFTcVNJO6uSzruALTpKHtFMfJRVdiPjuNHpAOiyxnWBlWH2vsElnSrYk
nd4ML3RwoM2DWwOIjMm7lLnzMFlwfsf6GZ3Rl1y4AqNHV75llMYm/Ob+cHbUcnGvfWAEo0zSUZXB
LhGMbBMi8f6knV+xyHuJIVDYr7I8ENFCqxNCRm1L24em40L1CNXLZU79i/OwJxwi72UsKnI/srRV
lFYMiVHw7QHl78NHoQgrJnkY4Ni2m0tojutS6PfIeONfwP/MFiFBYnoMyCbQVF7NJvvUT0uAwqz6
kUp7AmbdqH4Sy0jZPbFTNsBKNkBVAHQv+7A79SmRVpIbHgaj1Hfvmni7zu2HnA9f6kF5VHqHAZz7
yo849VNeNg85YRKvJHmMo24+z7MbtuNws/ZIqWNHQAyGbi2LZkbh53n6WxPTCbRwx9+bYuS2URLj
ACl4AToflSAKy8cmHfRRNIL8M8d3LHoZ06X6qeuwiY9f3F3gYZOHCYKGmRjwy0AFglL5K7DGJMDy
ZE7GrIYIXP3qur+2ByRtyUcm8Em7ZT8rp5xsgd/yILwW3uAQBqJIfkCrNu908YHvLDO3QGF6aoS3
H0YRBzc7bo+7/SIrlG27EAbe6q4yR7miC0ubF1QsJqApjbUMaf8+iZY0BCRC/vS3YimpcXN3dNEt
pCWjkK2o9buuGz6hhKbL30dI+FXi+7WNHfZ9s2WfsFhNfoQI3e6eXK8oyHkU7NDoged5KC+yNZ6p
9EBi+ISjjDalXKcyo/iQXwnU73fuSxKNBn8cUMc2Ny45eFjQ4cMjwEqW9AuRUtR7MimYCSsocHYr
26aVONd9eEsbvRkvEYPjgF+azzOyhz8oiGSuvYJUUBmtqkTZAmNr7uXprQLuQzgI54vEcYLH9tQ2
pCaYdy5CxuPWU3a9LjJbszlEQpc404GFmat7UO0s5kdgbI9tUP00WLKGRuaQCD8+TM0bMuy3mDbE
mfK2uK6mKISC8W35SHVXEizs/lPLZ6+c3it9egv0jpqvnEF+go+RMN4mrCkIPK7Q0XylV9IC2W3D
iqH0XbB7m5Bxm6L+IS8IiQbwF+GZ6YLjlz4Oe/mVATRmGarqv//HMFNRcnEUPL8VodTutpiCzR5C
WvFHR0S88fpeFZm7iqPjzmcyNOd4tQaP+mdGEhV1tTl5gNgc6hVyydbpuu8/aFV4d5hu3z8EgpMV
yVeCYi3Br/hrJY+TnIpDDT/HaE0mpcrupYZpSjHMN6RZ6r8gf0hA78PqAcp8qPXtn4vZoOuxQkcM
+dCYtaHGe6cBQj7VIzSBj81z4smqW5LjB/d6lCARL0ZCpHpLx8R1O7h7ipFC0YdNU1OzUdVRSz+x
Ri/vCo9LU7Op6MucQ8LWpQLr6F/mZwqz+/UMgYvKPkzxlwjcvc7rg2UT04mGORXRxgsNNM6OzLUT
58DMaPJqH6nbbK2bEw22gTB145dLrIeHCmjR6IqfcIA9rD0llSgQGOSSbSDJCUvkzd7Q9IMxT14K
Rp59h5npQi5waKM1GegJHU5dEdboLy9AhJBZMuIWhw8SSkrA1GznWfTmT1ITzLo7ZOWp1fFPfFoq
m8QQwvhTrkvOkpC1wkmg7WblIXY7nYJpTi9IBBa87NFl4ABVT3lT9ctHuj0A/eg6UzUNyq1gQxju
yeoFCDOyWhoz2mQU7rFf5Jiq2oVaXJTAvrMCEQpRIaZDGEE1ouImlm3S7XL8m5yj2jZW40uonagx
RTYA37jxCG+D2UueSMXWeBxAfxAiwPszH2KtH1hEk0oicNHhDQbfyBAfLWk9eXIZl7+/hXHsivo4
h4CmMpKuhlKgQbiIYd4a6FOBS1zCvNdjIhGQPde8ltY2u9Oj1vGyBCI7UBol65KHRoG06QW+WFqv
5WeOF4eJHMLQ+NIe4r2J11yb4amlJvmmIFHpnGyUP4Tl0zD+xG5NhJdkEUXDSS+A3BEFLvCRUfSH
Qp21P20J7neGhcz1z0wnW0j5PLZc9xfFUCdtaUaSco5kqyV+PrvCiRpgk2yEVBj9TunJ9X19VobO
WyJ76K/yeKgPZbsPjzcAvnzv1KOLsuIkKlZ1IbxfZjyT6Ox4GuQEDf4nB1FnzthGx8DPH6orpawV
UXaDxJcVNmrkw/GVrxd2pfR/Nj96PY+E+2FVC0/b7UhOYyBcSvSPmM3ibhiH8Wi8Zqjh62LwwX6D
lwp0g+Z0o7TqbRJ/sKZEdxYdz0mqmXyMJa121heRPlRfHJW0rmxnhVFR+QfSD/z//VjzXwfNRgTB
liH2rTtm3aNR2wSOL0ZAD7AcJtTKxd007F3dzp42MkZ5y8v2pIKVn098NZaqku47hLNLsOZuj438
+yr9mqHdWqmpxY7fF21kMyfvZV97FRRuZ3q8fZb1f3xgRBfviUvySVx5PiCbQtnx7He2J+mpTrzu
8kpfRnOj7nKRpAr2nrYbn/GZGbstB4TjlgzuCMDlImHO0KH9kEix2cbedy5Dv3BWvDIssZxA1uTw
iPVs3InkXead3k93SUHkCw1QQ/ZE/76icZUJCjdQ8CEXccP9Hr7XRO95fzoIxOHOiFjZx7k9zrHv
TJMNTgOPA7Y2taNcuMFO5UOmy6FW1QzHgLbUDSTTEZxVUy6X+90cF2a3PWRm4Bg+0aE4HTjiimHW
DQVscpZycdq6foov5TPPkkY4fTDciOCDfhKko1vuJFRPNxLayyGQD7BtXpetheb0TfYwsn22Tce0
LuK1pkaOO9UiISkuQ+aiIIXGKP9Hd2F4K9XqTNruo7bu0+KgbYMWL236TbHXYLk3MqCEVDuAcfAT
9KPk5tVJKXjx9jhpjCrDS6fAJkS9hvbwzSSgZ4zYT+XOKXYoPOtvZDRTH5Eb/FLEzn82aVzKaLpd
njGnjFN29jF42K1RH8VpBVEC1m5ijkG9VXbeWOG7TdiEAueXbAQE+RgP/BjRloBFAaayBtjw/Fdv
iLwtRvB0RYvGD6qSyemGErdWXgt6iHxpDy/wlSDTnRZfp68fH71DhHcabHDBTLU77PT/zd7xbD3f
eApguh6vAHsqrd35U1zNAXaZQBqwY6sMbkprE7cNvAvMbrQXoqGVFJq+CyyuOAYwIwHVa9gG++Ya
J0mQ71PvOzkCwoDEHBOi++pUj5U3NminX0UrN0j8wKE47uIDGAytA8kZKGzd7Mcd+M3setj99NVE
XeoaL7mFeuO2BdLKga1TJBpz5BXWjYyACq4D2BEkgEsaoONFTDw0LMdYpCd52soXbnoPbkPwhRop
cYcsZKd9WKexGguGn2JYbTCx/dUyV+urXBWPfYAB9Px2KLSoWat3MqEHsISzBeWs+JBhMw1PQVND
T0AJj8EfucbZgyWGD40z9rGRe2X0Cw1e0916lOcO/bC7pn28e7xuF2oP06Q0bvU7w1d7YP3IL3YO
8aKq+aFksp6VHGcWWHjkydHm6iQ4Y2BaLVWQbVbRnGGWbzF5j6PXMRJwxoq6+WVGfVHSSv6ez3pb
wBs4DaI2hXxD92MJl5pIxTP9qY/MoEPy5/cbWMS/q/RVjEKifwAzxo5ThvbvxMbsvw3JPOqCSptM
5C943tQlb9nERShh7kz+iLkuw6kHSVy4KkyX0LWw12XTqFdI/h0WtYJ/YPPNanRhNDqxlnJ4liIT
REFbKnDyiK2x5dbGGsSjH1jxkYtG5GcbEJHIbBjZRmFaqMoNnaBS6ZvpVedXS6XR0RrcH7z5+G9O
xNKL1dxXuxg9q8TDQ5/sa5V9zihiX0ejmH2v59T81P7yWl2JisD0R8QTZkF4YngbWitL+B41hq9M
evulXaCYbP5ZNKGt5Qb3JBuMGQ+ZiRE5+EpbNq7wBVmM/tt/kBsCpy34/pRMcF4MnBtiWVsUtuhG
PjHXFLaX/FoRk8PfWoMV8yORLAPgBB2ltRu2j/pL5uGyCkc466x3rFOjK9YgrLjMKttFVtyjAW+e
tY6ZB1pxZuju9EYlLXodXNuXkqSA+RbihDmjph6kSZwviCL4MpOFAyaFt8xcHZAxgN8d2vJTOYWK
2qITPDUq2YZ3+RXQbvmSpX9sqTfmQ7PKLwtKleyHKKbPJgffEjvLnHTGTyI2CxWQEaJDEDJ5N+Rv
XwkRu/Aqld+Nj7wQWgJN8RXFFWZdZ9f395PCd9+9PBpkPtJrfZLgdEow4tluL6AiVL0GNV60RI0c
HV8cYVdlJTDCmijQ6h+iO1WysMP0S+vo8rwI7cSqmr3Zuy82wNee7m1eJT9IgmSWDLOkC+5jERHE
qwywRjqN2HtYlBIc1p2kd998KIzIx6gxZS1obs4wND+ALPCJUKKG4N5Qathy0v6vQp1A2nCSeaoK
abxeYtXfXyGukKz3LNpyATR0w04hK45ONCdq0sWTU+4TZcbpzG6zR0FkJw8OUgu+1hI36hbRj5rh
anjZvGH2s92oVSy0x51sGJfW2Z3XGqcElVL6FfzanwnGnATsAR3z2TaQR43G7FUXbXUjxPAFNPpv
wkRHUSHRNuG5uD9bsVb/Hy49bNQEtQrtulA4g6HwVmO9H160tiiaEzXJS2GkzX3B7UfDuLDSHYeF
wC49PJqTGy/A7icPr18ILcrfsGLW1KZcrRJqRKSb0R0/mFL8xaStKjCi3lI4WwfJDtEQIQaRfK1z
xah3/NOgQf6xR4xxCk7NnJAw7EYqUgkFfugRzxe68NlIQB+gr6APsE85/4oUIE/7D6qeAMC6lqL0
AVlFfQ0W7qxAx6HgCUY/0OxNw/fwZCtDrZBZw6UjmX9P95/LcZqIrayyKOKHhWR9+bi1JRoofMpX
tnit8StvK/g88U38gCmT+OGSgRH73JR2OsdrjSPZly2v/b0WgiDO5+2J8HA5YOi99w9rVDj9EZ/J
1g+W8HAVadNueHkYmDT6cfCqz35061U8aQHzmK8QuTppujD66BEglR+GsgNdHpGo99UMdQimLgxd
2pF0854AM3S+lfaglKf4BFL81P7Zqp26hPHNtGqo53M+y37zzKll4Ujddu06WohRiE0k4lxn4j9d
tcOqRI7t14vj+taeqHdY7EamwHJieHCGp7qmrFpNyCAqMFzDP9Of8Zw8GV7wrfngLBAp6QiziALJ
lDLThYgalczDovs5+6KwUpr6MXOWmKD24dV+olN2S68oiKEGv4NY355TRvPlEGf6uJVFt5YaIeeM
1k8ikqenKNm4OxZVPrbTeHmyh2AE7mKc8xFWleYO5uLZfZCM0cyxZWOft/DL7CcKohsrgsM4hsJy
0/gV3V6idLfhxBy8+FAoxOBVM1J0N++gL6BnlKETthkjNMp7VaIZk07H+9J1NoBLUr936+zSSE7e
XUmFML92Em7eO9Gh/NtsTExO02ddUzRoHQgbK6Xfnrz/Ecsg3ljnn2IDd/4y15969DfsJxx8Wp81
ltwWr6aHODq6jYpOTfU/YH2NOoUiz3JEa2YqHLixwusFDeUFTCXL1QTG8GAwjsBmoXlyFhT3IK4t
D4bJVvOhy7gV2bFPGIcjPQbfTOvJGxIOE5KIsHNHQAC+iDLV5oVTmtI9KhOI5HbwBkgl2DEgUZsW
UhMxEibJSYbLtiyhn0zkIBTDoVkxrILQcDbAZ3kj787LtDVcSIhkFiPlWPcgL9Y6pdMJbaPx37Wu
NrfR0YTZJTAYoDVkntW4ThM6npw1sCOTTvV6hHQiwdxGx6PPrhxYVJtsMFEv4pPZIkMaBtxZbtHs
KuovNW8AbTiwfm6XUa/Yxjzr0Alz/9QStAVrjoZy72FKC0SVKRyVH0R6NM+3p4/H1WOOmCD+JsEh
lgyPem4YOQL6Qk9XMa8CcMNFyTPDM9mhb+KuHwfZWfsLWumaTUgOcHOD8rh/UmENVcbasHJxcnxJ
3x+PlTm20dmqtNbH8DM6H5tzzsBhAmZwJhRot+BfwRIBo5qLpiUNUm6Ys0EnwQIP6R4BsQfDHy6i
gcrZtcbFAeEuh/wVu3f0xdpaqua/uFf2EbM5OGKbKLzo0uXMKbS8IsVE/0w0NDJDidtkxr7rlc0v
NXrpxbRCDaMAdZpQTzig7IuvwwYa9x1LkK9kUhveLGNM6EtlaYlE5bC33mOg4tS8pdbi/SU14ORe
8WWIG6CltFdpxPVSU+Ox8dW5XLKQshy+mh4xcU2QB+ccHAA+kMxhFmaZ8da/vXX5BAHtkaOVgwEr
f8uAXXuQmAnY5QSyhmTXIgksRum4R5bySki3plaaYaPP5TYr/Hq+T/SX3iQ2Dg+9ix7Qfa/5UFUs
YwhNJ0tDVa1JGhmkvifA/GeILoPAKnpxBm5Riofr6D100PVqIojK8sHoSAegNb9upIHIh3kHUFCd
bblQIYQ9VJTmRdmxHphCgGpfmx5WnoGEN9ud8fxmHcX4FtP5cijwhEuwEDAkcwglX6a7D7y+LNac
4Rt4RoZfUcnRh0S7EYDsq/bCnWPUkYbZiZTjc8R8/TITLP8K3J/5yKStu4uq0jzE3H9BQuFFFKBE
ibHcM0VfrNvI+XosoZf1fEwqscPS8GDWCaWTv3k9CubICgXZhZKSo2+puTatcYTmWRpD96fLtEJm
016oL66I18SnW+H7mSmADFfr15LpEWLD6Cb7XqycRPNPWgWB2iLZqoGMqsidGB9MNJfeai+VZe3V
ExZNGZW0+42umELAcnKhHvSHvv1IQ2ovs7rLgKQGgsJrbcDneOKxlyHG2dbXMqZKuXPCLVxVFJlY
ehzl5+NIdPEQ4Vy3u3P9pf0ZZVGUSIgwdECn54KOCXcSxE7qXfFA5vSUX9ee6ZywO/n78ZwPAsTg
dzM7LSS3SXdxHixHwLPfCttMIF/X8wMGunR8Qogm7oSsWBywX2YILr0EMzKM2+b+4Eco4uzczLuL
pgpLeX0yrBaicR0orP9abS/jFRyB0MTXNxVRc7NdgStan43WHZl6RRjwzLfm/BLe7GoOmOzC6XVp
Z+xCaR8wiyDUuqHNNxfemB/zvs5SyUtPYFyJguPSiAIXhUdVK5rxpE/6Tbduh0IkQHB2fMRWOfcu
YzoNoCRKSGehxXZ0szN5FMxgN9QYDlaGRSaXIDD1yB7br418S+hvBqJ2CmkF0xBBliRMpBWbxbdp
j2cvDXUAynwzIOy7zolsHtxAF8W3xHcIjJ6SPn0LD++kqJcocCbVyw2NJv+mTlhuOMkpqkjWxfNL
B+POhdOq7upJviq2iY0HC1Wm4dmw55TmX6vsf0yQgSAV8vlHCz6XaVT0SnXi17ARJSHZAzEPbVbG
4F8ZdhtJrNhQca4jBCrQmf64JRm29jS1IRzhtYgb4tTwv5nTn729gnoVkEXzT3GIESycBMmtMKK7
5jsQazUaAPi6z7kYXJVIglnFCLyWTruPncxflDedMjXlXYW3ew8Bvifc7LqsXuIldz0aAgAIEDB/
F4lR/mM9zoYEN6FKAV2KLS4eX/I9E32Ed6NWKakXTNfzgkyQ0KHBN9C1IRyM15pPxpr94/zaK+jJ
o1SBAiGU6UOJxAG6HQPamERi81JSVtbOTccmGVDGouWWheNFwicJ8Gyphghr9vyhQUySHbIEMPrH
PdZ9JhobXaFKXXclQEiH3WPTCoXShT7MUpgqODpt39fXQuGIqC6xilDbYy2p0mKLCJQ+yBXsfd26
39cPLSM1Kz0lCBy+cWUUskDME1oemn+ZfhkbOOYHT9Fcztp+1DLeJBR0BEaZyS6cwh12q4htU6vG
cpqO0Z9B7iKWiHTvTQZDxG2iuBA0Ki7aQy27imitKVy9k5ghiX1FAPyYDfvTL5X4lZsS25ocDkCb
9DFCJyPPozwfktbO9jiY2LfAgIUP92da/ulVCK0YstpT+PCEtxFJQMeSC1Dm0oA9sMzK3uJX1WWA
y8WTPVe7CO4F8/RFYszTaxMTHR3XwZvX66o8EkixJVb4gjkERNrM5Y1/iIhdA9ySXlSf4iT1c0eY
315762HJTGKYp++XVJ0MHVc+rMEwxubalyvpxgaoEDrWLBXJIzqA51klTw6Z27Ko0P4JeKC9O5Yi
gi+4DbzlgFHBnulapXtPLW8gZB5QEgCtF4MCIBuv6vccS1XEs6TjHrvXFfKdwjkZlqZKHg1glXW7
oXuYEoxcGnz4PZG5K8tAnVTrtiYWaH8TBv7uny2VqNL61vGS/ixociYs/fhFickX9VT8YLuOxgvx
AATpDhPlXN4nDCkZm6KU3/y1N8nh0FMaDveitVaXaFFe+ohPv7pzTHe8wTE8d+n9VWy2fOveeqXr
PRa+1z854mnrkEm7oIPBauXBF2M26ezn97M2ncvI3NyQLxYlse/ivWbBdx5OajcZF9d914/GLB7u
VoqNv/UEP1R5EsN16GT7veP2yI/JDT3PosH4it8Gnp/xvr8ny36e+6GvMEQBh4ZSgHvGUU1MQQL0
yeBeglTN1Bee3H/LNdPhMUgKK2i0/v8N+0WwLIOoK3O3ntUUsXXK/7vnCEfwUxVhZiFM4OiqN0W5
5Od9faeZ1QXw53/ONo4Y+PhpC9lCcnAzu/8lkzx+wIp2ccetXa2SAu2RzEUo1mHEFqMki0aKBKsX
t9P86wjjIe91/VxVd/QdXnsZCWHQ3AsdxCmKD7uHk9E4+AyyGPwg1xE6mxH5j7wpUKLq6nmQx/yq
ViBKoHn5K6XtBV+jK6qeZgKN9AG3BOc/piQLchCYAmlYRo0FkDMmMrc51CoQMbF1Du9GaKDBgSOo
78JauxrNo8cGOBRR2yY2rSUo3VmGqwcn0RYj3OWtIXaJnx4dPnk51HG1uFnfEhMXcmstFczUBjFr
VqtbfRYY2K3k21B2vh5gJY9fgaKIV5EsJvn0A3pinTtuVM8ni1+IdLD7anxqJYawXtPOFid/EJxZ
l0nVPcEyaF+bCnIrg0A+y1WvGeKXRb9lYjEPx5nV7DXvSQ/XWWqeFtP2X4/to/GVu/9i/TLx3izK
gANiHvHojm5zieayDqMtNGpV2IoNyiPa1+dHnzkZAWb4FL68TFA1Q4IhAII3S6kAUrTJV7/Y2KDx
7MODraGBbk1TpKuiO5Z253o3MA7/rbUfiB4cyOwhxoDmaHKh14NL3vZ59ua/Zc08nqXw+VgH2VJr
RRWuhMtbGhhRi+wv5jNMLOcS3wG8Ax6wqlLgVakLdWN7y3qLLPzfJeFN/fJx/VgBMivq/EQuQP/N
uRl0KPYA6l5yG5eVPqT9iQxrZ8e0PjODUtMmLRHkPJu8QtSROnkjpPXaSBsspVr/xoiknrVtQk4L
qTOe753WNDVXpu58XC8mhjaBA2l0XM7SbVxjqCQwMzDp0I0kx9zAWyJUa6xO7nrzDZXbBAsUHtFb
vpep19KAPP1Dfwi0srpmRKpuk4GUjv8PR1FpAcklBJPWuZTQD7ZVFFtdrItv1dBcdUnNjb/PlmbL
BBvazUKXmu/2PMN5Jnh0VpIEKBEzqWxjRHT7ev+enB3G7HYxJ6GBcjf0rLaKWA7GmGOAaIuyXeM7
5gD+mzUENOyARNjR065BPags0pQ8ddWtKW+mXSXXEnVismfODrgsHo3/x6FfhOxfYfjBbOgjo6CQ
3cw0/kxToGm8C1yycBpSceKPo+oKR9fMmDCuS9njAQBHaX9e8sCwYJVIHXPKgF8IyOPhuPWjZIbC
SocOlLMzNLa2/as7GS3kuIY5XON2OcfqUhoghMsl6ck50c5ztR6qezUZrUo45wO+xeUFr1uAMauB
vmZKVZ9lGdQsYaKid3z8YP+WEjm+4RlpNmdHi/kiLST5VxePINrWwtz31aqrPXIIhfHmzT8KZYbr
1YneFGDeAayUPtNg880HiY8Jcq3oMoDJ0a8UdQTS7M1Z2nvnNr+9MTtT+8YdcZnznGoWDpaQuUNb
PEgrpxY5usCWrNLLV9BBKuUcPYpubks4JO/jCqmxLUvDUJny97IAtPTJ2Kn59hyrMSs4rOEraNhX
qblZN2ShHoxTy5sJY4pfKDwM+DsZuuG1FcHeLMXSJx1/yEbpXTLT03indWMlx/YW2zE5oNWgZfoB
DUl0Wjohz12yLENcL0QJNb2Zdvb+1jVIB3S7FyRwzoYVFqUIOJ+m9FmIhjb8+BlIi7+yfBQaMqrY
XPdmDOga0eItdh2LCYoFOFKcpT4oGU3YOKotJHsICb++YU9g1zI5Pq5zIsdBXyfSMW+WfOvLrrmR
TaaMPqEpOjgvHc922CNRWDjoGOXDxNcJcGCDEAEorkjLV0qb9dYOZc3LPAaYdjOaMEC7yNad0Hff
LUG9q8Ih14VF9UAhkV6+XbLJI9RsV5YRI34aG8T2r/tfR+pIOykuG93pG7W1JcFyTARs1z6J+M+p
Z5Ow56JwJkaajOXW2FKhNYsxZgD8ix7lAoujR/KFT6BTiLhdnPFUch1qyPiEZObCJT99wxTgm1C5
PUtip8h09C5yOzyuPNGks6hmeN+V6imtQLcSHD4Q09KhOXCQ+6zkkXOwoEXvpTDRR3xgJUJIyls5
sWDuS0sNxfksN6aLRCQH1g46A6KN2XzyuP98nGgSDriLK5dmo/H26vHs0XG2Q1lHhEzuo8a8fOrK
LmBatfkMNOyhO3rkinY2CzvCRQuJUZ/XooGc2TZQsMLR2nMuqPIDnGGw7Ud48KrCN9tkT8ONXlpN
BK5qpSW5vUCX2IC/69K8YUidLYuI+xApw+IuMPpBrh43a6rIXwUkWyU+rCRvNo51/HWipuDnusjL
niRRdz81/lTD1mlG/9ljRzWiDiFQSUGcVHTLthorrzrmwW/j4UBDv6yYZ1oAuYWow7Ja+2rxeQ0b
ZUP0KwUr9ekhAYU9x3Ca6nNGl/1QPq+HW4Pvw8KOc4z37JS8AwY2Wq9c9aViN2fF53IplJLbPzuu
YYxCNyKWqTxmU3LCdzG7CmYzEb/kNOYZFuMhNdVhwRnISolH+UhfxhHry5fqHqx8grUEDKWkwA5T
PupR47B0rXo4oFuirx7BdO4hhHckHDWgTTrS1gQzYpkrxUntBKMrr+anYE2tZjwBTcCy7qAZclaR
dBgzcknHpjAvCeNfzKilWHc2mGPxNZbtZ+T9oNaMj4QWJlF6waBQ68uPcc39XlsyqQSOoLSRHsUi
1Wnn+a6IsLJZFXQK5+dg2S7nCXJ6pcqE4AbLkV+0pFyTv9P53uEkp8avKbZJ0SwbZYomOH2Zxzfc
zaKvS4V1d2+YuNuLw5uE1rABRorp/7iLHtJebZUup2XZvzjxfoEpH4YaEwZ/3l7aThOrMZwUgR7L
qmgpej0ApH4f9YCYVPNjoScEvlR2fZ6+PPyDQ/gz4sBM8howm6Iv61P3JhjiC+ecD6OzAfKRuQiG
RYHtyHZtJntfYzl7KjGJA26DXZrIStdQHit58Ut0MgHU3NtuiytNrLbs8qKHZxUOZpfitb2y5meU
P4IdL0ZMktBjY8VWMmNmXgg8Pp3/eOGqujRigiBgKUBvxyVK4zMUzX1UYUU1SkmsOTXf80Vyy4Kz
BEFzmQDDIOHoZ6qy0RWxWYyZaPCvEVEBAyWjT+4DM4ShUeBQtS9UlDEzP3x5clQ5VPeyv5mBSHhW
LmVyjvOegLMjCz6AjEzOPx5Wi5rV9WaaERB/RaU78Ue0bL3z5lxZI0dGkKg2coFk+j9dWyl9VYbi
PAVIULOrS5YEubDn/yTesDMt0KrObs4ahBJFRIq15ngof8hwvqXxq2RhCgHowu10iyP9e7lG9LJ7
9ge/Ke0Xb0z08boWzsJfxUAfgvaTDn8/i3vogwW5VXLm2qUWkSrxQdvZ1cy9/Xl89Mp8XCFMJLRL
Q1E2IGtIciywaih5XrN/kB6sCTYjXzoE1/w73vCFGAHk5Dns+lv8qkOMPRZwqcXcr7XWEn50Z8pH
Y2yJr47L25YQcgCqNsClQV0jmBXSdCl4M1zBqm+B2dVYIs8LtokxpYOvTjO9DjwuQ87Y8ZLM5Xhg
DUrgpa4l9/KO6T6oibHGHm3UH4qPecAKfKRnNcX40bwKgiNbBwB4izIrh2/2mzk+cINeFmhjKLui
t90rQ188VRPTtcGp7o0HgqP5CazD2wCzpbk2TmVneLdYQmTvf1pp9x5qZUgQenvEKVNyoyhmlb+f
so/mO1CHJeAfLmeX50zAcbP8S9cF263e8GJHrB/eEDw2ukfuFdlQ1jMEsU05ID/JiW8EpA2zUvzg
U4HjqOsYhjzOH4a+1jG4aI4TEZs3tzI2CoPpEPqu55nIZrivDgn6TaCjX7/QhwDiVj8yI5bEYbuq
pJCiB33lOe6AXloflmnavU2m/GxPL21GUg6EVwEjHqfqjcTYY8zImMPYeJ84X74CuiO8fENI2uJE
HjAhdklsQe1L7AVxEhHHyV4lOZKXocwLfPUrpneUlOb0VMD1sQ8RY7JbezofEEhJnPY7SvbhOT/e
Tz4oPgXnA36lUz/Rx6ynQtUh0dUVxQLXYZTTDOS22J3vBCR5x4VaeUtHXpI1xTU6Ahr2sjoEA8Ky
SHLWa0v/21CCPIGuoDNdiqww16iCbRcOnLkE9M49aFPd/btu3LJ7tNLrtiFdYWKTSVO+DMDPSU7P
EH1Fti1g5ONatLVYJtMZkBRW/+jxt5q5L/qQRABJfrFgMz3rFgLjkSwsld9gU8fAlapPs7a/yS8j
iYACht5ykg3Vd/H9lOuUK/tfmzKsFvWn1qmLmWP9TvhzkSehPF/WJNxnxHybLPc6JKT/3+ccHjSI
8+bWOopKeju40KIB267bl1cG5UsbRkhgYpRWqGR8hhN+t6s5lx4YaPMIYV9GH3/Kiwir81Wgxsvj
ZWUNmCgp8EcsnoW6WPslrx9Un6LIme05LLkQSlO0iap7ogjl0jUUE85I6HBHVvAXXmaGg1P5rZFZ
ksq7g05mtXgiDkFkpo9zOBmPB8QLoOWSx/5EuHJzU6YSp1zbYK5f+OG7AizfQRppjwYrRIkF81Pd
pIEmUAlyxHvS66voSO9ajsQp/rfE0LluDI8fDFON50kVnDiIMgGCEvBCyqaVXqyX3OA0VQ1DZMZI
IkIpwcFVsAXof5WpLqhPNVI/isLhPZGhcnnx4HUHLBfXngHW0REfWCoMxrrtg8r4vujlh7u4tbph
SeXWv6YVxhpBvJhEBKKdF2blnkV4GbbLV6HIAKGunO0enzpxdidKdooEgtycqvt84D5YL+MGwXpI
oh/lYHB6WiSJuDzGDKVpvwB0Cpr2RjVNsSVNIx5MR1KiZi7SS9WzstaEEvSZj4GTLoK3eW9q60vP
GciqPWLbR55FC3AdtE5ImgUyJdAw4twHPAG3fwYsmu7xpf4MrUoq+HhMzGWu0rbxEScVf9G1YNNb
9SFydSW/AeD/UXCpZVOHMypQGaykuqUg7FfOHl4oId2sfgfVWMKgQSTPquurLG7TpRxn5v/O+JeQ
EbvQvKTXsYI7Cfl46yKRGZQG/RIKyZqTU7X68vh9oGlmGPvRzQ+fYdcLYdCSIYc4wZQscqGWnWNz
RX1dixyvLZstcQi3g72L7b7qEQLbd36MEnueyVARkqtVcO7e4M5VHktuPFEpqw7RtI7uplSDo/BD
xTYYWOrtZMYqLCjO5qkGdOaSrsT5vOZ4w2HexbsbSg7GFlfSVS3p6jfRBn3vmL2RUORCKkIt+TlW
L/INVLJVGiX/cN/TSDb7OGvqdUgQeI1sfCSH0HERDgusG/GzGWRXVM3ZRWHwl7DeqsTDLObqZEZ2
bD26vc32bCNzbHuY2kz0CyGOaWhp3YVXgHVUJiyhRq/MLhW3BcO26LUrWSaGTKT0/cHN79VKWQKG
EL2LX/Ri/Jq1GY8Z0XBoz1SOgwCk5pS1A1Q1fwRYcvxjIcpl1DDIUawUHTFjV9uFrq4fje4eyruj
qdteBjh3VazoK/ez+pALwU9YRRFY+kJYb12uupcucNlsjiCC+13uXNNkIY6/d/t2tMb+w+dQBNKu
sbenfLYuI2i+M7ZvEiVETXUFe93Ke8RA6QWXyEqSUxnbeDviu6350DS+IO+YJOuBEgLttb9EafEq
3Wj7VdolY2b7lSLSYeGDTg2/cTj2MuOyZqJWyNvaxGDvYualMp7xtoo3RE67IUw9ErN8CzyGClbA
bZalSTOWhq4IBERKnAyws8PJ25+nZOuQKUNFET38vJ7yE8iX5nf3bf0xXW353tJiOf9xbO92IUrD
7Mmr2W50Ppfd9YNSowbMz7EuAqKSRW2ozjfNauLWwevMn8CHnRqs4J94COm/lo38vQ4Rr0XQVtap
L4BG4cvFYeJg7F7KqDJs0srYD5VqNRroMuQQ5nMELMu7dlKLOYGi4Wg17SaM9+kJYJZFrApZPLJC
bip3k/EkPRuvZ/3I2VbBHEi+SuKX3bpAAwi3z7WNbakGrzMupootBUSwdH2rDdjP/AA5CwLLQdmm
89meROJ0IxZPbZP7cNBpPR65sBZHFdKc0Rsxk81/fKX5ctA924Dne2JC/bgXPRPbyApH6Nq3j+Bo
NLc8OK6iFkIWGcrwQOO08S0OiZFOCDSZSpA+XpAlBurkh6Y1bP+8f8zaYkOwF1wYqiMYKp0gwcXT
7vjVYNYAWZX34aPDqLkYfToDf4BZeOjk8h6PyjefmLrJLXd68ARkLLDKJaUwuEHV5jQaN0gico1r
qYVPI6iHM1/ZCUWGgV7qVsL+Ds6+Cp+IarLkiodaLdHrzIHmeBKKC/hrdjCFKxzZn1aRCSSPZWq2
zTyddrXmmuGVMz77tjaK6rj9WB2IQ1T6EdjiUKRE2D5UxUirDOwn6pBippygupw2oRSCyQGHKjJb
xelUQKhPRovU5cdaRilvycHtUP/f1yG8NU2pY16Ir4pslsO2BgH533CDxgURvN5q6iZDtUJ2Xxbx
GoPyQsPusybfRyvqktjZ3Nnnus6CYiUE7vzZBubKp1bD86Q/yN//vstl+61nV2TACg9Z/x28LduG
QuV2xMhXdrHJUrLNaE1b2XGd/qFKH+4brJ86cMBHiR7Gl1lr7yepLKTjao6vsoelaURDda9own6V
tqE4jzdgj4mgz3CAWbWseNDwz5LGFO3uuDgctdYx+faHp2L19pPoR0MhE/NOOH5uYSTz4sHy550t
8T/KiPd8oV3jvm4RS5xxRDSDddYdkEEQpXg5aIef6GxRZsJ/b6DyxHmWmM87t3g6AtjLpolF7pCd
uVBaxBmWxZZwKjC0AqidIxEHs6TT8m7NdNk/zV2olPDdi21G93amuLnVTnYh9gdAzOXXEpYoRoDr
m5V6Bwj2b0G80PBqcwNV1rIcmcp+8Ezq8IjGDF19CNzdmrYdtaensjVPj79ynod1PSgEQ0QlpxPn
TUCAEm/iNyEQnf/Z5x3+sMEzxBjvXlVHAz58+nXbumXiYw88FqJHMNZZEraUDvOXlbvXsOVpEAR2
yxBl2iO8vmZSnO3eRxS/1A7sjGRdigfzWnE5jIYgFmVva8z5/IdIRpdjQlDNFgAO4aPLVZJV0GtK
PrC6zm7Fxpam7eVPwVt9ckGx8mpMaSKMhVZu0Z/TfLSz3/AhXaWEzffW/K+eUQhwlW9UTeMdUtaa
B2vtUAPOQZ1DDI6xpZ+iU+9mPgdVZ72L/lbgyI8AA8wwra4ev2dkOyNRWVKBjeqN89PLotbk4dGB
p5QVKSI0ahtJhlTINGZUZriYrhPThTX7PvzqE45rb8/wD5Nxxel1mwqfNC32+1VjDqtqZKAqCUKM
StRIyIIwzpFR3V45MwxudTShBxBnDMX2+WRty037NwiEcph9AI/GsneKXdD2sJEqKaqxyVgvsETW
4HVyDw7Uh+etf2aezWfEgb5iwHlKiW2h7Qjhyi/jyeW14RJqLe+aS5R3M/uPek3IBNr4+V+UnvY1
dh9QVFzFIUC/vo2xbAGb8npeXduSk/zF3+ucIweC2+wIgAtix1GAM8zuByCE8J97yW/BbdhYBM5r
hvQW0qrp/g4IgsHqIfd53OGGth2Ix9woj5tuCXRYNJzPil5ICrTWAOgkgXLKHiU3g7L4CdCm/726
pD1YUiCpctEWoreW0ut0/3qucpJQclDiD1VMsv6j06eCcF0okJnCuzdWGIxmr7CyaYz/l6aopJ9r
yPwwmy+RWTw2qDVbseFBKOHwBdOpZB+i6u2St+ISjqawboTe4bRUf8QZyz/X0Hz/Z3gOyE2OSIVw
vEC6jyfwZXMqUCvTapFaaDdq381dJH6PwCf30gbQq9A5lU/uQ7guu4Q3MMSzH20cX1TDSButQSl5
KlFkvW3HJxRKvz9yCc33tl48jeKcHiL0BL8kqV7vgT6O3fFiyRwkPFyxV91tiZ2DfrnNxUAVXlkf
W5nFfzJ5LYwZHub1sM+z92aIkWSeKIgRYUKHr/1dAzKm+8Ob5p6lvHxHfI+xmE2aaxBfRgJ6Loci
Yiptgh+TyHTcFyK+OtSjogfn0E/hAabkz2XmlvuqladMtSBzWA33YSv/3bB+JASyvatz5c0nCrPs
lMR8zRcS6OFvZ0uePpTfbihbJ9xU86tPCAuAytIDs4/0HYWNUyVsBhMYgXr6Bc2erNRVAN+iEe/x
vNs2ikKSzBBvsuhoxBdtNb8IX4xlUapkCk1P7owpmDdWCoVJ/d65sJYudxIbPFx2TtafF96bShJl
NXe0CdGxFdeQ+bmybPZls6YzXnc0YbgcVfGyOR22WSi92cvlkJu8RtGIC2rs5dYRZiVZUMdAHtJC
dymnQ7LxaqBJUoJ2Bu/InENUV/6t8kLxBR9gP/n7XGpjJNF7J7yxYhdbWWud0NnYL7IFo4oCp2qt
UW0CelgJsFQa1qFrI5f8FbXkFAT37UOctOfMme17uE9evOOYZOXt/7N9nuzcK5QhLiGa6xnWOiNe
Rswmho0XXKf52oyCAGAAHoFj0OdidCSkJII3W9Mq4Ld5lXI2s8FmPTcA19aZxVxMEiwQHpQXiabk
cKduoPCc/3kdhqdA4+GwD2/jNrKiUtwiIgaTxErc5Cc13sO57icTekO8tPWo8wS4lG4a8JzWdvFK
DZXSbcYmEubldEs3KsD+dwlJIiBixiCadKz0mjCrWXAlt2oGrzHr/ev2hfoSNlJeP+gamDtooUx+
/DwYi0e/Ds1b53z2VWWxQ3yOdOKp79iH9T5xXNqRyPjhdvin+VCgdXAzkYr6LMu51T2XFxBeD5CS
tjN1XonP71SVjwpCirEXN6gQUsrsC1cY+KOlWkzfwzxjSz7Js6KpUDLc04VDK19rLifcIrfoTYwM
JiyVAeAW716Nq1xzeMhBvyQoJs0lJh88UWgxRIcoRC2ZLgpSXKC8d87GI/lPTu+hxPPGeUNI1yVy
5fL/+NUPu53YpHpFC+SqAIBAhJdeFaZyeVjKJ4vefyOK8quMWXGRUDTTBQQALHIdGfjfohm4rCuT
8+P5DjQHKJPbQBtM8Lawj+YrgFwJC42cvPJI/Vh7NHz75pcEB7MH1P+1Lj/On7Aa6k8j/+9R5LIa
VoAsjE6C12G9fxb6TgIQJQThP15GnIKCOge4i9CTplMO1bXJQ1Z61y/nusn/Mz7VwU7F+119m4Wu
11z3A+9PY8EvoI4GXbpBAobhbCnygig10yp31YQnTrOVdQ8k7gPLYULsUi48PHoIPDCTFG5PfV8v
uLsd0jLAJDi3ZQqpa8VKaRIVD0MGeKoCOas/HlH2ZQbd43L6hB0S2TApSCgmWYwDuiMk7G851XF5
KmRTNZ1ACrRlczPnoFYE+HVBRNZWf1//DDQT9n6PhJ4gqKcDw4Xp+WcjOUPahMIrO3an6NAlzj/2
KB1YrPWhyeY/GDCaXsEZRHJYC9vXvnbsv44qO9wAVrJmmnaNXvGX2jhdUVX6E05qYJThU7fA5tb4
3+DHh95fbnQ9kOZzJxdAP1bST7DHvPk39iixg3HOGqZ6BzzjzZnRHpKltFi2PmVAeOTfKYoDDa5Q
I3mMFzOMXT5RUEZYqgEmnoo2bbvYV+Fh89KtJDMB2RtkjmlwzbVfVZjqeJjoKF3mUQ3NSz7/Sdfm
NaddnZCuzrAllvGfWjB0J1esXnbgiIAutPp4GZ6QNEZbZQ8GBnCsmQIy4yneJi4j/vohWmEjiNNa
KwwTGKP+/Sj4zhttmFcDMDkFHt5XM0F2cHRvW8t9vtJaRJZstQvBfXjknJbMpDUmStU9PO7WA7AR
7f1bm3twDWpvrYw3iFPWiwowTlNAAZrRaubBdWXZBKa9BpzQ/fif2WA0nwi++H6NiaSWpzXMk4b5
XG2KLtCuWl3KRlMkgA3LYKZnwFLVwTjnxpg40YOvJ0LTG8cizrjRl8Z6PMlJnyglPgdZpgsP95lC
bP5XhQZy+bMy6OpejvLsxhRgosuNWrurgQmW4WsYIrWT5INRUBLiGbV93bjhNTvEFp3vZpbCdbdv
UVN0mN/K+Vi9gWmlNq7IFBoXkT0+KpqoPllWsPgG47tKXpWx8LrA7gHyeC9QG9xl8g3QYGTPOamR
Ac+j0BYM6hQACGI0orVmoQthoG8Im3JLn530KFMcSpAq5bBt/5Ubs/jVufrGGe+8C1P41/rTtW0H
ah0HG/BJAGHsjgw0YbYVACYaEMbDeHIhG4wVFPpypukiB2RqFCLpJs5BS+EusnIsPkuTf7oQ9wx2
IZW1URXbJMJHAYRuxILWA6kN4tEmob2VOXBK4h0FlLFfJaLGeuMfY/oXDaNcV8x2HPsEefn+1bCt
vvy+7gJh1uTejahf5Lhb6GSoVf1gJ7cNRCOpa5xjvouhRbRTmnHuMextRCGc4r/1VbmMLw+1CDL1
wKR9O0HJBMoWbiHU8u+OF+j7ZHOmrzztc0sHvXF7E54TYgcjYwrz120Zy7MxlDyoi/brlaHvu7aD
I7CL7vFvbHebE2D7aHwW/Wb18FgYdQZ62kvdtJH/HhV43gNDB1g1wo3ffxPVKut2rw79H+k7KzOj
rYm/1D69w9IZ3Cd0GWeZqdkouSpbNvMcRqC4Srzp3h+LgMqM97msc9IR2m85Qa8vLxQe+DJsliVD
ErnvF1ylur+wB7B0wzc5Ja53VLSFE8A9Yp1TxTCUbF8jO0uP0Tu3PY2sM2gzwzD0aeZ8AyOLAH6H
yYDzMeo0Cx6X3V8fhWmSKQKAZEFLaS2fSdJWqmg2PaiFHEoVK833Dw1HdbFoazzr0+f02gRcJnXq
JVGvPrxi/ALbio2meg/qilOZLVXZuTHJHFIfaAGTbPLnpAYunyHD/OfaItazSxeJ3eGynzZz7Lal
Qrn2AIcHSWogCb8F0S9xLDAdTsQFeU1SN/nfDQ4HaoXTPiOrixNSnE171XptrvFNBMkcSMcpkHvg
bcuxk10T8jNx7svg2dz8g3M6xgZ477y4OE6uUF3N6bu/n+xhFXYs+nbR4E13SqcQlW3hBbeZ9s1w
FkeQyTr24pUbgyaigbu+djTZOfd1pf06DTeVeAE+t8G75okhsJvWBzqcxrgJNqzr4sN4VtMkqRpC
vv0anVh6axWZF+1MJAleyMAyXye74kSVTSk/OK1SZnJ/Kllj+jwEPNXlCUH/itfLJFwtIHebLDwU
mDL5lrSOwcvAHHqTJUEYGDt+fjG105sG2/ogN8b2CJ2BKZzkwskgEjepxmTOarJxk0rWIuAhxShC
YbwYlyDi0+7spwvCX0QTOMtFCWB/ZWIPIn6xDM84jnKHrn51ECOUreyYBT/JGhJ7jBfGyq1j/MyE
5H/99km3SSwl8FHHA7G+LQ/rDh1rk3ORi3thz4+znjncpuRCYovjrqidmJCteX//YBwk9RthV4ZW
dzuSgseDjGCF/fleiXv7Pf6P3ZVKTUzMyjEKxNBQaiQJmt0AOjSbzqEh+608V4a2G+xeEJzWWGTx
GOi/UHdzWTOpKUk9unouwvWXWtOEZqFQNdCu2eHp9XV1Usy4GILFY0PsZNLzaA7g1drjNJoM+EBK
pr2/O4RKML2bJIE2ejp9Zc7XqIdrQ96hU77xiR1tEmi1Ejka62NmmfDzqZzhztw+j3LzhUCWQIK3
FPAIfF9P1dmtHatxm1kQ2MWXs08utcprWTfPwmDZMZR8ihyeWfDjdWnvYctp4HzagHUhcgkbDnDe
8cdqBBgI6EqqyzTBCfdVrykoUK2YvLRjBHzBiVwQBIO7ttQSI6W76wa5GO7CN5zDHoODdZLjOyPh
RSY5+Fy+dT1GwUq/IOj07Kn7+z/d70WRovmrwPNNWvx29ItR+UfsrTD7U6ON0RFs6kuMbztMcBJ1
bcSXXkkWzypE8KMQkukHQ3pt+UelQHaP4OZ/vliqSoRag0vaHdwgPNzlxRbj/yjwr6u6c4wr1ioh
l/l9T9dlQV5hRwsEMYh4UH39vCfaPUhmT4WOC37K5+aT/4d2SdW+B+vIuUCyhTpoaXKKLibgy6jX
V9br1mBl7V5VBPLG9LfsfPGzss/KImpenSaleq65UjynqLpiqMjOU370yFiDtH8blTasFIe7sC5a
PoNtkN5oBSL7j9RldmtHMU6ZzIPnRlOuI4Z5OtR3K/yQcqjIu93LqGGKlxg2T42rRH4vxQdmGYyz
WQLTbORrrysGegnKxebk83p+4fbKP9w5ac10IFpcCcbuxv0JRbR4mUH9DrGBTm5KPBy2pQ4W27Oa
6uzbpa6XiqtYtaC9KdrfBIPndObquiJ/ViMU3d0tS9D5Hf3QI+E2YL+fCAotbOkqsma3m/4+SwRN
aR5jQdq7m/aVkcBWq8ZgXjD9OEni6CrgIFmBxTuG8boE6bIsAKDiIRXvZeKBwuXewsu7RCr1JPHK
vZs/csr9ngJzQf+rVuWnRUjqWLQOogPTtw3r6vD/w5ts49vTes3CDksv/W3l/r9XdLs6b9LZfVfV
ELfSDOWCiHfobAnOpq2QZ17HG0SMCLEnrFKbtXGYkLsVdMcCAtoTQJolllBZbYryXe42qNBTmLtx
nQCLmXYH/wgfVxpI4Szs19Q0NwgfFeYu3asCLO6CaJehDjFM7MilkqoKMzARcRIpLBvlj5SCX8c4
lmNBecB1B0vMlPlOJ1Sy/lMtvpSBbxsyjcDC4OEV9E5FgovYT5fBStt50FSMuQF81hJm7C3ExLIb
vWxEZWzQsZwFIKasjW8MIcOkA/6Vhg8+e+1P91i78ctmn7i7RWQeXVvI9L4BwGJzljP8h4G7xkvx
/YFh1f+HqWKtUqCLzEqOryeeOJIDEQKtnokTJx3hQHWFggOD9qTBNXFV6vZ0tCPrTmlc0RAAmINj
XIrgiP1hsi4Dx3HJy6kQbj+M0+wT1+87169GukXZZRWMLAAxbNUX09Jecw8JYPcquSFhibAftg3M
LA7L7sOyHBaqbGWtrHK2Y4+pr1DUf+eOO5j40fpFAMoivH9naDKdSSwextW7HlghmdKJDSzadxna
rTsqs+VyP4Nv2qCA9xIAEp4ZKtAayrBzCscU+wNLDC7lwHrTpg6QHW62mlD7DglRA40sFlx4Snmn
J11jJ2GkoVsZoqco0g57eURAG4GNZ1M7X/lhkfrnqJO2A0zuljYtQMlQt2Oe1wqcAc1vo7cTB1yU
kIY6Hk79nNzUFV8iCCqT0zb11wpBJG3Lq/X9FQEmgLXiakl0R5co4kcU15Hzr3hAbMv5Cnv3HRrs
sc2sWs9PX9z9b7gjLy9LrAdB/VWrdH/tIdUH7BIYXaqib0Y4PLd+BO9qJ3udb/l82zJTfeQ0ctEq
f7WqV79WWKwOZjHhVl1d2I01L0OLEdV+RQ4KZi4/kwUNoErfqWFBDYSc9v9QoStBwRpI8e8nXl0a
K1YY2K2jhJKRM4qoWY/Ux/Luwg48S+o//wKzvILuL7wrkoyDEaQH9BW1Dn9QWdAB3EHIeiv+55qz
W/DRN45BBoDUANY6CBAQCLojsbmUvsEPpdHpi2MTyeJN/6eU2w88v8rnqvQ93961mQiEsaJPMILK
8Kzv64CGvhCSB0Y4VQueVmI6jhVTifm4fdUihWasc175HV8/aR7NiUg0/DIOjgL6mk+q4hgTx9W8
0IHiCNBbIWB6zfFGdEBGWq6m/GTpYHoHlb7zPNoYaDKWOUhiS85RJ08Ua1E7ZZgt24aKbucOuZR0
cP2HWnajOIN48hWwbdQJmfy1Tft9c1QlKuCO4WZalBdo7vjfH5N55jpuIQyQuH0/03QTnbQNN+q5
gGO1C0Aw7aWR50NUaEVEswc2nrcf65LzgCPx0F27nKHIZhSdtVBL0L4tk/Aq6CNpzP8O3wJ/Bm8p
LEE2dMxH82YAIR4Y5QnZW3KE8I4Ls2f6HrZP+al/XCNFEHXdOiVSQri0sJRDoZPoi8PPUz+b2/dC
VkHTq8iR5ZBzdCY7QW1caAHLa5B4wsGWL/sNpHHilZqGvaKJojakURWhGhgiqr0EeSeKIeA6QKE5
sf76R3yQcL24RLFYThCPp8Ht1ke649FWJneYkXhuoJYxYwRTI2KyEAM9AZ+qNaW+x6Aqi+khJ3Du
wFAnZVsrjXxI+Qnd6ZPuJJZ+6tMmuVAW/ZcK+z7CVVC8SqoLRGKZ6oMjFsw8cP558VszwxIBINxd
HMm/ZCGw6GRSQgkl8Ddt5wDMIDiAgY5HPtrCzfuGMf0FWR2XUvtaFkoYvvEvyE9kFYsWEqDZwVvU
tz1Hq2L306fHiY0k56nT3A9RDQXUdYL8Nnp/hh9E61rMCTyt1CIxO6Htz6xqcqP7sMf6U2g5XB60
n4HJrUGZutvRQk0sr323PUX0zpEs02x/g48CmZOPYidT/cEDcl3vdddLlQYAfDB2Gv+Wn43cdrnh
JZoxzqRoXaaGyeq5MR9iadCozVA3gKX6GK/1v41XEXP66FT3/ZWYGwgmGqjz3JYwM9/V9yEwhRkD
ObKMq1YxnOy3jYhjcV5/RsD+giJRpxv9zQGRlSlaQvvAhDiWhE2k2i5bWYTNFhPZe1nyU7QjwisU
WtuNbnvdZwfAT/7mmUfYLXFJII4OsoSqkrPVL6FHAbkI/TvWsKIuR/k92PLIL68+MBRsn2uBUZ4l
WqXvmzc39UK+jXMKUnO+t3b/qOZpRfuQJfynA8WZcPJjUYOhw7n+EUVeoe2kLzWzuSSZQ5ZI/Q4v
sShvpP4ep/OZha+ai1PrzO+6kgaySIkToJh1IzEBZQqmTuD0y+P2pJmVwvqovOcu47w6iI9sHp3s
CDgvOQ+Hggt7Lzdkn1WtPsGjKSdx8tSLGeq2TLNDYUrs1IniTS+PCPxUN6hSF3IBNpFE1sgls6l8
Fk7Hso0zFeBDFJAre0iRdmcQCFCKEOMpVBYKSZpsQ5WH7qOKR0CkBvQ9p8TQFzPdYbD0gCA5MuwM
smagqpcVeVTgv+sOso2cOPVxkAmjNlurfVPHk2NWRCLxUHQcL1smHnop2N53p9gc6PZs5SmCNk+T
0IGKNLSDTJvPK8p1D2IVcvnOw6IgqY+rMbjCIjZXjkHpUPB0b3T9uueFoc4ptx6xb300yLdzqHi8
r53IH4AYQ7a0XJFvlm+gFv+/uqVp8Q9bFyd+uWZagML/jWix68+kUwz4F1ZJBiQ1N/PTLu872yIc
vU7UytGXa/YaPtxsI2d+d6PgyFu7xIHC317EUeB8EPE9AoyON1+2KN9GFdrF6Yq5Vx59f1/UdqVb
DI4xUnUwdl01wSvfsdQneb/+hgi825Pxj1HSZiKP1eE+HoaE9O2Ta7RgzRL5OdVHdyeo2gNl0WEA
NydVeHBnJ1HPRE9AEbcFPQ4DpoMVw2lg1DQc5qdHBqSmn9dH1dOkBXHFZ9007CTo5qDNY5bBrcIN
lTtFay+sL3KcyYtQ+CDbNn8cgC+yxWXEC71OtiB0/Xo/iSFPwBUbRrgfhTGH6VLVKnJNA0ALILpg
pA3psSiQJEIGkytna+XpZCyDCbp3SG5A/jXEEOV0pg30jLoOiNul5ZU6l3NKWWY/UA3DQglr5fcp
bb9eGjSquN2m5E2Dy909uYwz8s7B8O6JcVPG+a+nhUeKGbig++T4krcySrNCsD1M7zYKV4qAMS3S
8qIoh2MTOa5sDgAthrAVJnvRrFbwfKeo1lRD7NltaKRnFRQ0MK3rZa5uJOY8H8sE942V+y8il0yR
iY1+jVouovYqT2VN470Rb2w63YOgXj1Y71IpNnozu4gNzzgb8CiPXueU3P+0tF95yD84Iyhvgfbh
qx1YrhjTqE3kyA39rVa4a9Hu1SZxQAqWeQfWoONJNhq870vZmUpkJAy2DN7DQ75hEKMCv+SU/+54
1fbvB4LQ01wKRG9+spBgpTkskC0dOe0JDLdOnN2VbNKW6T0cIMtRjPOYzZyQYhesrEZkPtSadZje
qkm040By3PYiM+3UZErWRVHn42v1rjh0TEMhYQ5IlpvMvDHxabDnopva4AHmLSGStq0Vgj7x9IY0
JPffvKAkSrInee7/JEhGwe+dFMln/smSv/0qt8C+RObBUk9GjEhUdTA5u5Cm9uVxZt0aJf/Fp1Di
v/OmCxONdohML6frr1TBJgGclrAXvspZG7flL5cHvMog/KVxNGLieiHrGZc8fGH24jitTsFFoo+3
4iVjsl1qCXBGrt7Li7j59zBx5XXQHSw+0mZgfvnAmZFysTjuX0j02suvy4AGWLWvfA5ZK1fhE+IA
p7vkjTaPQ5tEr4KZapOILJcBUklzqoRoIHFvcAV71g+GT/WLVrvQedyDbZaBESm1qfanBLz7FEgn
krP+uqM17RtjHipuW6+M4g/A383uC8y+QP3lKF9lVazq1yRiZe6oCnhc3lQIHOziwOsmfgrLb+2u
jZ9GTIWz8NVt6AXA4L8AFvlgyfpuRXf+KYw4vBDkU4nVszA8nvFpXvI3hgKA0foCWUs0AaHA6WMe
M9sxfjnWQ6sSjtjip8rAFVuvmIV3P8yCFQJDVseyE7x0VUJrCxChavD/WEkieKjrXrC/IsLAD8OO
iDpS+fnWCOqnZoWH8v86gz1dGjPRNLRDnBVyyPw+2wYtQ3b3d9/2jh4QzVJBpFKDX1KTSmtAzvMy
wuT5qo3BhstIWSWFPcdIjNrztdTY+56hXd0YV8HdkNQkq6ShdmpTIclDq/3qUJK6Pcg4tM1KYT0Z
Zp/ur3UOlns5v8oaeDgf9vYt6R5arJ+bar3zn8VLVjRLhmm+qdEHkkKyyOfrkOBQBXSfivst4RCY
6J6mLjn9fzyE1XHHLtL7rvqWXPhyszKTka4PPDZQRJ5tpxhDFe0extEzotENN/MAbYrQGM5Ky+8A
Q0WWBGeqW7Q5xGIP5UbJ8kIYQx/iBkG4Hbkaj5W23ig79mKd97TFSHp+5Ex3ceCBq09x1aOSztYe
NyzqHnMvGRHF0B1E8AYSNY7VUhozU6AnKMUabOdEgI7PLksx2yNnOD57hrzDaY80Gngwr+uqWgpG
RkEi9xziU+e3yhwc0OR4Ge87vaJ9zIa40akZh0UDd/3WT5wvfPjI0PKZj4AWeBqv3qUYM0651v13
HReXnsnGO+7wFWezP2EELCWGbQTOxU72AVBZ8X5tchAM87Muic5kOt+ObgCll0GUwPObUTez+2Zr
Q8TrdkMl3YGqr36OkxlopvSiKWF84GEOQ84DYDXj415/JM8YfjaAPzN2DVdzHVPya1Jp//GaIv/4
eCELLOEhH6a1OuQtEWQ/vGtwX76BW7+2AvPneQYUZmLUy3IWWQEcfLSipDaLc3hmjdW2HMwUYbBE
SMCdO+CDqh9VugYGzmxPnK4Xzq7/DzVuAsn3TC0ODaKSpbxaBFxhdpTqqKfTaku2nepM+vneTuCm
jQyNbIcL5C/sOM0bBDyhuh2es7MPX0USzYat62R6AXRqDpAgJ8sHmrI0G6KImr+iSNk5NKkPUGpT
6JswuZBYsdP+JzDVpRmGgAFl+0dKwH3CMOcoOJkflZh4YhNwJGG/7spnYavKjidI0jZnIqYdPxZv
exS86u/DcV7tNrf8rykvRajrEEqNkmc8CDVztM0WLqi5ROcOK9dpnmordlc0uTR43ifYVpQd9x21
TVHFeJiS1+Ru4FMf/gCC2CALimuy4LKRFXTh9Qmmw2OUN3rDTHb/03PvjzHcjw/8DhAmJKzxjxpU
6WfwdzjRv13rMVcCOmAgOJKB88AqPAcmBogXv9Q84Sw2cRaiWsjN5rxgvpzWgkNgN00vilQDqSB4
9Na8o0ZqY0gG73JhjPzaGlhrulmLH5o9nIWoAxstwtK1AzrkJhJKIcQfyOv1cdbdhvpaoWIhXvvD
2ssVATnYmbbWXBDE/QEVL4ZG/VF4mkONlYNOVUAz6qPNT2SbZr+uHbA6AB2Mz7HHDH3IwkHaEGaE
iTIpr/nQ1xiw8pIyinQawY9cqOCi3k4ViZPc/vh/kaEeLEtUoVD4h0UQK9+kdyPqFq8AiaSdgJ8q
QaeXQvDwj5tK5+HU4apqiO/b92QinmAXESntZE3c1j1BaqPQdh1nTJsKwFE+DccFqqw3iL2jaisR
hDYSXHju6XzeI5SXMpsrMjrFmsQ0xuQ952cq2MZ/bK2FlV+U5fpkQ26AxCST+1aN9I2QUENgQT0t
xM/MQbnhqmSzHqzcZVKSuuP3Du37K0tmc838ER9qIVvtNw7jC+hydThiwLk+6JF4R8D5eAY3VRnN
YYC3shkGGbSSDbhdfwQUs4pREZoAFQIwc7t8G8sOFoGF0LxfzrtoOqj5p3nVxqDkamGnEHaWM4i6
GDrhzPkJkwpsFqPZxJohSWCOrbEpiq/YMsZnhXg8Vm6NOVZ8Fh54mWzZ9rrFQbgIPvkwJ38SEYep
gwqHHJaO0kK8GWn3nTZ2gPTzRFiJqAPf4DB0f+edkpsEhl5z0YVWmrpnBXoNvPzDkh/kXqMvMUaz
uv9QWV6EO4hPtFs9H24NmH2BR5xsw7VZ1A/+gnSAeDUiJgWafXQAsBieAPmjsP/UcI9+VkRvPioS
P75/mkAaNEKSDuANhIhTejlP06A5KwTocWMBQatM9Cn+VzDmoyTDFvSCQ/Z+1gaBZWJiJYEwBcaJ
q/IuPq1WDM1LiIUzGm9nbDkfWtccvet70bpEmkAmkHd+74AT8cdTsVDSVJJ9qbxvPvuhmc6fItf2
/kaXh3sx0w0mXcLsjZy9em8GJjZzfPTvNowkIEo7zZJ13JJActSSpaf5Hj6ZLFHSJT4MDMW0AhxO
Qgp4qG8AM92ysexOSqMwULEAUbVNrDGLbR+OXwJeCUcJZmtKAglgNbRA+171pL7+zBaiG3k5XLVu
PydnT7Tat4p6Pg2MCriESroz2NF63yGrdw4bebuNGHWy7hURVL0Wx5/FePEHu4qNjB+zdzUBumzK
S0O3ywj2OoyrjU411HRLdR/W6WayBjAbumNfeeRQu2sD9z6oPzSTZUuT2v1jigI5rltJbL92SR1a
6afqmFGkMjPe6XcNcF3wfojXTxDPoktfsDm29+gHB6hpLcL38tv+bv1OqiH+HbJ+VDG5hHUUsSdc
c1oPrzHYhQDjvTYqVqCEBG+qgdg+Zr3mYGSCqj0EYZOaCVOblwKvVxfiBHY9Qp0eZHGrWTMmpK8O
5/eIeLQobA4QO1IZg1xdMquHEiT5nG5QgzZu5fWPmJCLh0bsUNehJlZ3SX9sBv2xDRr4JpPfrlZ7
wFbLZicS6+HjgBRcpV0fvnFn3lIkdS0AOMDhJ9pPxJlm/0LwSaUA0+MwjFpXfGub3B7jw8J//tqy
VwyAUJNLdkLEotS1RRC8D6Vx9/s9krT6rUy3T3NS6xVfMkfqTKBpStWvK2NjlPm8KN6GWiZrWlTM
FEhXEnx9wAsfdiPLRzL5waXf8yuPvPs9r6pi0C49Pgpk5wrMENgC1mne6u5/8R6EreSScll1AfFR
oQIA5OlXv7QkScO5Mki0Ipbsw7vQ30MAEBQCc61zfv/gKlNCfGJN3NkchKgbjSR8B4xi8sQHyXeg
OxsvetyWkXrYGGbo7g+APDf8nBIn3FuwdNwh7M+2VSe1H1+cunwEwbw67axE0grQb8s87W3PI30H
ZBHafrjxCsiNbKKyuff7lIRiyVrhgtikf9nykurjtoyQ4/ojoLOQf/P1L2LNAoKELZMucz7FbsvD
Zhs9pPEbtp1q0k5US4+nisfJd5MOh5e1dMkdql1sp8qYlTlq2VSbrTt4gnFng51BurH0xR8vqcXI
EOuzZ/3ol+4ojGoiSYyJVaGe9ewzuO6oCVEtVnoOzTlV+UA5u2JEHulGlOTR29yft+wfHgXeuNV1
P+8/Ly+deC82MOxWfBhpzf2BtFPtWoRwhJTdnP8UPMxeBmyMBzIWfTWfe/7bD194d5OhbRE3zo3D
LXQo/hh090Ns71w5E71v4b/F7dMAUv1QE13rxUyvHgFyCDFMqMp+gF+YDJ4mZVh3Wj+VzjqBKmMZ
yTKNBGlgJmOguqIIFs9HRxGRjsAcoDvDmbLQE5TBxCJc2ol1PQp3Vx8M3XGJ1fd+asMcGxfgJfx7
TXgalGEzyPAA+CaCWAxfkaNhX+J26aUtQLt59zKiv1Ha+o2QDaxl+Z/iCtvCqL5x3NOFlxYK4yv6
S+KisIqIBgsk4GNHz3/FFgSB1o174ZQnvbCDTu+Xn0dEPABtmCDN0MQDJJaZIVAkPVNel+GF+ELE
z7tSGSd2z1UM+Kl0LX5i5CBF/XBzixxBqVw5bezu8hgqjINQGmhKyl15bGTFJXVHaw1W1I15vQtx
7SB/v+KbFPVWYl4/8z+zpxXvucMzRsk6G7cwxmc2jEOuqsu3uJBmdwPrL7hZI6ksxqWgaA1GTRrn
WKaS9hj6CeEABDWFhYK4Oqa2nAUmqcVPAJA9+evV+E/TQUZhcmC1l/25axytXpk5t4kjeM89GQJB
4XK1htsZxy0T785iqRgoYcNurfIAoLzc+MzVkRpxZ/9p3qiBY5KIY2g9zEBkYjsEvNgmT8xNjDI/
r/TVBYmqO7RkF0bSMnuIcQxyhsJZIq+Oz2Il9gI/Oew7K/xywAkgzxGWPhaOlesB7VzK1U2owvYC
lzfb1YjmdV9z0fGyjENazHFjIiftbnfcnM4WUatqk9+Uk9hPKnmRaScFrJIcOE/a42Hr3IIevyoU
27LfgNMuC6afjC6MseEFvWCV9e1TcVIMbuV/yIkGAQ2Pg06WWX/wcd4cSkR09CPQ5TntG6ZKHG2t
ZwZ1TqTW7jdCG7wh9N+Yowddw/FZlbEJo0afra+6pk3rQhVEgFoLMortq7B/Gx6UHUSTe7/XViZR
+HPMCIfs3G2c2OZ4GlZD+EV8GXtEuOlOzi5jOUTc53y4lDrVXOs8jJf5sswjK3RmPCYXCWTmGvKj
peoW3ZhCXUnhn5O/iKvLP56DMPxwReUA72keDJ/O4Jpr8nL2SybvIxnFi/aP8ypYzGg8Km7KnW5v
up9qMv7JDN27bm4r6p0Z5PgA0oXK5epXd8kRTO7HzlWrmYCruhJhEOcB2A3puf+4B58F8IreB88I
OpVsDs307sNGeCZLkOq1Ze9nqquGNscZvxOzWlVNyKvo55XT5tRB0zygBHL8MckjLyQkRvEobQe7
J4cB2efpZGYaJVIZxRWqkAzbX1f1VPTbY+FaBBRj0oEBD24gzeu/OlkWA62mhniACrNBGtT1i9Qu
rJeyEy3mh0GVDSZkL/HVR4ZxEwTrZ8bhCdO+mqhCdyWhPYb4LGAg4Sro4DnCnScZLwnziG/3w1V7
G5u7VbEFIjKt1Z632WIqY0lq58mQtkxFF4/m52ioKzenBDnfDsim3Ptv0vXJjc/xpQLQRPxqavX3
Hdv7ibA9uBO8Sxe9ynI96fsCEBIx9XYjWm4IH3Z0A55vdFBTEFF47ZfxDLNWyBs/AhRdCtUYfN32
YCTyumuGY+G4hfbKd1OwRubCLjh6ggfpJEWAMZZ8drtincRZZkgFvAk6Htf5ih6tPBJ7dMsVVhVS
TmqsU/UwcAgfSQmIdu889yJyYfz3IyQiNBt8lI/MNGH+zvUu9FrotF0QLmY6Ovncg+5lXulN3qmL
IJEQIhdRpbTqPgPS+1NMUnNJETz1jMoUE7tt1bc/IlHUPM6D068gdx/R0eDCgpfPs4lL+QlA/9BL
E0MLUhWsD/+xfSgs3ScMk9qMllxXGgXbGS/0F2aMAIfFz6HFtWg6zCHuZiUJ5ie133FUscN10J+6
S0+Yrfz26ln5OxLtX/vYjf2vcMdZgNqzSXlSiIhyszLLbCul9sglEWdisy5Lz83Fsp5avi0NWu3y
1lccd3JuwMiRvXzwlvvarRkN/K6tOcDsY7L/fmAlbkmII2xrw8KkJokH+rIOUEygSMEnfNk2elX3
wFz99dSrQk/dS8ijeSI4hmH6Tvjuiq+T+0q4rKhntslOqCJXXmJBWH00cFMwL3/l/agedL1XhbSr
pP7HB4Le17+e8xI6h+JR1T67rJ0LBtyDIr2NseK22/V4PKmf/fQaCdfa+rNz+fQmu8NxApCnpEW/
NL/0KjwvyM+Q5zPbtnIv4nMI0YV0TtTyTM1IgTOL1ShfqU6veH9wDZjDP4DtK5XWfv3aJrTwKsOE
Yrod+pivdTF7KadYq7BPB9z3lVhTHbvBADY7pWgImQEG5aBuz6+VXYMHnkQH3ijTHXKQPo1WGc5p
zUOnMUroPr5keiK2COx+P4skpZZcAoZfvNAHsmVcaGAN++LL65F5bdbmHRSgQIojONZBbBhsW7xC
zHDSLbh8cx4oy86tyu0Xfog2fTM06XV7pMukqDl2tQF5YGLiFfA/c04e9dQUMqBkdrpVStw6V3rH
wuN6Y9TB/Sfml2vYinBowG9w2CmR7bFUcXrEcb4he3+lTaiwVfWuom5J3EiaXznk2bUzq3DnJeR8
FOubL8ZCgct3002YkYxQ3VVDLzvifmntijGJs1UtEtT4hppbOE+pyQ4J3lLezaYvpFu8TzoANif1
pn9QeJNx9Yb4WVam83IJ3/KquRfnn2T9eGWnw5Oa5cWds7OG2i90IRNnNPVz/kHSIt+Kz+3w9Bgl
2ccCNb31k8z6Za9iZIzV+VD+PN1cklgHBKp4GJ0pNpB7jr9+twCXYKo6FDWzgx7qsRa0eBM9YSmM
Z/z+VjBC2Fig4emvqUxqoWxWZGs7KlEvdu0GyTTxGo/1XbshfnIsuc7tzsJZwT4q9nHiQu224OrP
S110rg1hTvgzvvRxfj+p2/4RgIQ77bcfYc90VUO22oT27lhYfbvTyR1dv/KqGaG+vHuw1cIOslWK
GvxrVw7urfDFNy+WOQlWi6QQonQIwZEq6CFNJTB0e5aCvQmYxHH7gdo/hJoilY49501LCxbsBGBx
VKBDHBTPpfklElejwx+O+tQfo/AzZEIlK1Brq+lBuhIMzX1H+LroKR4SirkglOZ6pkWm+B87PRwl
KtXIwuxJtfMchINbuwK/OWEm2uGHB9LwcOKaidom2fsW0AYuY/7pWtrcDNbxKn9Z87Dx0jh3g41n
ofmtgVFXRK+cJCV0ZFbEIb5ID949ZRL7F/RMwUBk0pDIYoZ0qjHlpnn/ZW6K8FO9KrPp0Lfrz4+d
NaYNj/alw3XSZT2xO5RUQjFRsbaoTTnDunXamAyCFI9iAx2D0zLvtkiQz00qnU1SaqGOGieNBrJh
ISfzn+zhWJhg4BtSDjkrBCXq+rZOZv9SbxymLV94iXuSJGyVTO//aPhRWlwVnuwepUpQ827EdIpO
VDxnWfPQmg5+o5AGgKEVlclWe1yZZIHtKZSqfEuYcIVpiPbI+D/bJPFMEpnBoKUPCG6LwQ78sXZV
/iin/HOlrI6iXo+dixH2dqCTAGr4fJnUgWy0XeSkcHg6uTHPYBm+8CJvkznHP+02apTpMoKakGxZ
g62QLtTbR0H2Ds4Mj1juzQKx5bSkTlWIMOIqPWSB0bflPY1pyRfk+5MORbCYd+dqLzq4XblRt5qe
S2weZGa2CXX7jDcydTgwSI2kjzjlrOlqpnnN6AfwrZlUN5D2Vqt+JuNeVR0tZW4fTt7hbo7NwqMb
OPg9IM1UjEzM58fnl2ef24PZKwFm7PRCDNRCM4uQo7Ry1o0kePyHV7abP5tm6ROslAKQ+lxQSXK/
4Fx689YPMhtmJnuL9nqJhPCbwxap1dCYy/MUMUfatNbz520rG5YrrwxVp7EbUSzi+UoS3he1DAWX
HxynDtq/d38tfNbNrIzu+m8BVCI2fFwwUghWJGh89TcwOACc00wSc6nZ4DBxOTZ0sJUrkr6nZ8PE
lPj+4TeM5Gmz9oaTwW3xNW2EYQo4Frq4bDVzFMLLBAWxGPfLYhfgk4fhL4sQ/0iiACVAMSmczxeR
Yg6pLn4FhApZ3ikjnjpaJD6Vy5vQSls98LRw2/RcDq+D9Wn3XoX5dycGfjw+dTr7V20wsK5+lb8R
WAE9wVSeu9WVXJb9gx8UaCk76fB9ab4haNOIRiE0IFd6PZqEMWLZzQZIhhx+lJdnTeN0uHnjaPea
4LID0IjENItfFo2y/MqRawa2mUVRWIJOjIWG3MlJkVwFiR+61uzvauJwbiHRSIKAVur35dB5c1aJ
wUDCnt6GuXekipmG8nKdXksneTnR44koGPZcjwPJiTLsjLTyQYBBv4oPg5s2o3ee4c1TF+3hy4uJ
qrK5kaoCxx5G/7zDtAqmO1h9AEqqO0wbPat3DpTHsIStyuHfPoq/VKCQecfligYe/T+g+rHsRXrT
xq0xvBmEm7hRxPVCk3yBzzwB2rHBfrlCioumNm/7BTqIsPSjfa020Et25TiWpC8elzxXRb6LSkE4
K0rRqI1u26c4GsSdk4SkQrpiWRVkZCUXjg8nieFbm9AxbDEFZjhDvXy1FqYGauTDovkQVdpWFXoQ
ulUIFrZYTsu+B/W8a5GaZx7fki6IvPPgAOa5s5TGwASOVBFZZSdYTb4FAy/1gZ+if28lrziVXOfU
/dni4QJGwRb/MiCOd+deNnlV2tQZyHnN+quUbBKwF2+MliZiynQUDFZF6SgjFxG0hqpH6Dx5yO8B
Z27BdKL8eAiASmLsLt0Vbf8U8nDs21ujQLXE3tZUAoS95vJHOwSZXRY4XGac1MW422muycurNSmv
qB8AP5tQ53oHRKl2wruPieD3+EruLHpQ/3uKuv/MXFglsSwH5f1cP/04Q8iT63b+9AkWmmoGO4Ov
VsfR61i1COEPGFatxr3l9VDbVeDUceMUt1JFCNIpZQyl0ZIieV3+hTyYjnR7OvCr+/7K3gxzICED
eBYAUtw1Y2clidRUxEMuPSJnzoTA+kErNvf4EybVpkoG77alB65+62mTkX7SA/NKX/QFnL2KIrMF
OYNIWpn3HxEQewioKFpWS2Km/IuHuK3DT4CWyK/iSUppGKLSe2sCENeH/PKZDTN26UtuhCj4uMDP
VKOxVYI8KY2H2uBoJRxaOtlSvpzcoTxLsjrB0jAOoaNOr0Q8XwuE4sys+DolM50D32JUBDq1m8cV
j8x1V3q1y1rUc8ShUaHEHxtxqP/qldMjZojafIX05NxK+V3Ji9dE6IuDIljKd4b/RJh9zHkCp3l/
n041KtYVKt3IAauT4a6ysgdY9V7aeoze/c4On85prFN7BR+kiUz2OdtXN1Ef9ngmzclwhybzXHgC
0febo8XC8H5dLJDC4xw7vA3VY1npjoj8zMXf4AMosRAgmWgJnsX8B7zeBVnsAm+FC4dgcfLHjeYD
dbL//MnoKoLqEAlL7URaMcBVR+J0UgEQz6p5bq6YpqVbKuBRPXRK6twrfdTAs4fePoZY+ELv51aG
y8QNaJ6ZKFEw2bIXJnvuBuV3tkONvYWqSwtmn/0bbCXyOklaOA2ubBKTKLNud/WmdbQ23JSZP29d
FZxCLXJ4T3kbc8FeV19Nn4F995GvGugBb/2sMwm6ReXVfzR9ApI170jiDvUwFY5a2Kn93dz/UHs4
vwsmNg40Q6t4o6rChfQnNHIdwS0BYCmbSIsvFHme7u1sTHH452ojZxA7Wl+K9t/axu2U+/Y7MUL8
fXGnxBtdf2RyCOivb5I/rogAvGlExhwsQ1pDKWxtuHiNw9VyfM9Mtf2QdS8y/EMuzgtxmELjSAXp
Tg+qCXViQ/5oS1CGBkQTErNTwud8yTUHzmmFT/m4POsOUCqH3Z/Fb0B99VVc2ta7+af5hJlULlel
7IgMp6jdpFDnnu4kyXfyX8/i9PSXHI1MWgOfZPPFXi6qLxInDaPn97Uh6FLAE7oXo7tc+jySkXSM
wdEoQX6ik4J9MOOJqRjGKtre5HHR0ywdbTZewEQAal+VY0q6efEvg4R5X0QvASdr1Hxp00CDlXnP
gvgLScJqSTyZra9F8M60HaujjZsVpP1IU70k3HDdN5j94uXeFN1Lj9SrV3khJ4rOoJPDka8aT/Kb
glA9gi30ZTF9lsJF+oDYScsVddoLWk+GmCXMwS2IuzO+iy3E/Usfmze03EBgSkHvn9qWe3W4s5Nc
mveqtv/LgkrDsT6LyWYht6V8CWGaQ+gWLnYboCt+oVYTA/mwUKeCjzS6sPBafgTFoenZ72gRH4K1
1GXWpCPTAVPkYqVBlX1iGDyHcaaVXJ8kMIsGjvZJrNuW8fdPA4ajkt33lL3jLFN7zTLyB/jVCfCz
hLA7F6jue7iX+KRDI9M/yQOkOwyCV0i7G2KfhGLs+xJvsOTpM2BNz4Lmvpwhvuo8TE8semVO33a0
n9iiOA0aqEca/yPfr14XBNMtOIZIPx0y71oR4xOBKIBZPBnpcL/hkdjaC8fbwaCmZpo0zwHKcPGZ
zZ0jYt9p2WCO2IgjdREqkhS3LVz4HACgpEmDlYri6fd2l5wBrP82WpQm+PEIetb4947uTFW2hygO
EFs+rqRTkk2PtTXoTuJk/Su2rjrXOI1Na2cnCUyL42xmhVIRrkWpDbFzUryHDo9xAqPnHYQRWm7i
J6sjyYdyz+2q4TkGAwMBrIhmVuoVrtjt2XKceswb72MM8YC++g2CSRRpmYstecb9VUmgHmDvmMc7
OwiZ02HreKKtD9m+gnF9rUh8eWl6gJU6M7pGpsDHILUOjzpjvVU/g0YfaihSpEp8RS7ONadQl5Gr
XdaIUuMMJwYAhOxKx4sCIUNvx7yvBWi9bWCX/OpjY21JtKUcd48yVaNly3FCOHwlDlC9r8fh8Wxu
7eZMe/yhDJhQYlXAPFNuO1TzgpE+1XHYg5uJIuHfMVwagRS6UUBs/Ezizt/7yz3uPw3mVSHHvGvE
9dk8QZu5AdPW3sJ01EF40l6Cf3UF9/0t6DseI+G/dx+FfQ8fMCyrVnoVU+mlfpQLdDH3LkY6J8qK
Q5TiR5mwcLh66M5921a6ql21bk3UaAC6p8zbVOsP5JdhYh19f0GlCOd5gw2aqX1NU76AQQJcVEVL
bATjFuUAUSRTl605/hrjm0g8vG2myP6xRG/7NM0dgD6T2FZXbOstvEdz8gnlGVVM3+50k9XWDAv2
oAsJK4A7YHEdWyDf7O7GeVZr86Ui5EPfv5SHOYfEzLY+s5xniW3tZrsuy2Pdmw3pkzAPdcxPrISU
apkzfEmECNcEaEuQjHnkABG5KFGqy9f/FOS3+Iysu+EBAuMquS4lb1fWZZCsbRVtb7cEUxTwQEOw
ywOeKVELCPyRBN9ckk321I2cVAwHbj3VTk2wzOig4bIlmX9SN84RlUkt4y5/LTFHuEKCJsRfFYJs
uOjvfDYy+NVrUOwmZf737hX3lcA92RSjrBRExP0t2sXPqtym3SaBChbdQoBUkIGN6GF8QDqEfMsX
A9PRF8szPqQ4frBrJv06FWMP2wC5ZcX5X3F/P6XICsAt4jj6e/l50Xb3pO+X5paSUqex658tdTJQ
NvJzSOb+lveDM9wAznCKcvs4mvEy+ZA2XXvM8aNJjYqwOpWFGA7DhNzO1hU7kTKeF/O4wRz8GDuZ
eapQkAKJBi6isS3hDWC1l3FVpe5GrQPCoE8tP/jUvJgNvIKFNDeyrCLcyirV9hOMQsx7EO3+dqFw
WdUmlopxXEcMx+SK+rKShAO9pwLqOXEFGWIngxpwq0MhLwY7GPUNwWfQ3gLCtIc4GzW2+O4bF0zA
5RriwCoCUciaStUsmLYm+k7iGmqUH6G+pfQ8tv4hCcaQNqRo+akvGQ0QXoK7paAh0KhjCTQHzqtE
HtFK2sToSXGKEjBlEj0qvlx7CDZxmno8xs4UrdG0vgmYz/1PPA6SpSYOPkdMJjyAAgg9pac/Is3W
Or+9fzOsiYVPPCHTzhGgGYoX8/4KcgTm0nQc64QkKWzGXOSbwMfhRsVBQP5FEn4SZiswpCcC0Z9O
OMIrUpvlKLL+7u0kucB/jhL1PxmHS/A0vFtIh7RwSmH2qA5njZWDJrtfObgMKYZkR14hlTeUguJn
UmmdmyryFn56QouPz3JWpaDsvLUaNpwRJnbZpc7hqKlH2S9g68V+WmGHAd2QnmJKQSKrL2bN1IUX
dx+k1GXzTWsavyUD5+Fo6eJCY/qdtY/JPC/ouGp6vMdXIjZQ6C5eXoKK+VJil4CmYLiXAk2Esdgs
mXHNtZDL0lnx5W3Jqr5z20xcAFtMpE+IynexTaCp4bmCgZwS3ZQWusJsfMdQe4cnvkSaPnMoQVXk
kxZ0IujFCEJdN5Th0RQrWwwAJxztqU1fTbK1N0dYczgrhNqoBxIMs6RUreX319Xm+I80rXfCiFWg
y1hwP4y0bk7gS2PTMEyIX3iObp3Z9foUZaHVGwUYHppS8UdK3pLw6JlRVxRBTb1V81xjOKgOb6vQ
TmcEGEONtgu8ZYtYCLhZobGpU8C21i9z+5wcRaffNkPyMqhaxyYMA8CsBx5dQBD6FenFha3Df69s
x5nkl/BWgWUZPeJooAUvp1EnLoTPUmiSfySj6jAGsaj+aWPIJqUhpf2f1kNcnP0kPVVF0u/pH96W
ynIII6Nby3p5yd0b2LCAeV/g898gycrj+yFJL0DrhWjil6vyoJQ/KMMeEJLd4Qj+ZRce1KBBBkCk
xbk060OdM/olbkjD43KQYNnJ2sqoaemDXauehAYe+64o35AY9liUnHwgTPAHQvSKeQ3En1xyBayE
uxIz9GGyL9llztmuuG73jI7Ir8l7PS4UIQ9XL5912r8mjgSEJEtasrWILsKcRWOS86ISZDjawdUm
2Y0QDdJR/WDJCnm6A9kjl/Zv/mUbPqVAETRpGKozb+oOjf6j70gAqt/Cvfph+UyyWUfWoWSMSIkH
rG/HxNjkEugo36HRgeplGUqUp57Y5+iV0ecDFBXJp7ACHjjXgbOAD0bghuMn65ZDRThG8b2nk8X/
PRu0bzqo4Ctmod4gyys9e0Q4Dfp2HAd13wWNg9Wc+bhDqCvvqXj6BQawg41sy4OgztEmttjt6KkX
moWC8WOtr+p/OkDKirn34T7Z3Hs2lnU4zn3atze5pq1xrHUVtPe0DsD61xUnFKANa3T0hzh1OKKY
Jxd7SUEfoJgAFxV72RMFXGWyPiCYtnheeykpsHdpBnPNE77pOyDrUQLBX4KMzkkbEUUTdMxCwT5i
nhQV5kBgobkMjGCUdFdCKwzRS0vP7woPZ0YzQceYHzNp23cIPhfzIeHBekqVeDAtoHVzDEt9S9s9
8j5vfyeEKbowgbDF9xnDyq114T+ZKrAN6RTKhBHfiS2+57n5baxhP3ItA6uUW2nYeF+8DEdeLbQP
ZfF6gjMmwyIGPah6rxIvbLBSUfHcIrFnzv7jgoW6z5GFsEnp2Fy2Eonq2g47fpaMTV/NUN8kD/2i
fw2LLq5fCtjkFZbr5J9gU7gM08QktCmUXF0LjtrFt3JDxB7DmEzTiFI2GnvqAbSgFhCPLpEIsNNw
pTInEVWHZZ97PnkhSKe2pPYREuMW9G/8sIMEl78sTrI59tOzDV1SF0P9EEt3RqSGYMwA4CDF/K7E
JYIUNb65pkQnxDN88wzcnDsAHSmOLi/YUFMAJvlgEmMzpMeTAZfWwdYkFn5g7nlwdyPoDiGk665X
FY5hf80QA679cjC04YB1LAYFn3JA+NpU4po9PcbHnfOL/3b3VXvzG6pFTmbrCNm0HD98P6vllVSy
A9IeNG2RDGl1VSCG2xY5xVAwe1QC3YF++AVydj5WbyT47hrUeEt47jU65iuAMk0VGdHCWTEQakCv
mhPh1kUsMGRTWCEQIvoQixW7d8Mco/3i1EjDhTUqC1X71QqRfZl64a/jmZSBnMccR7Dcow6KqZDA
4/dJgbp5hH/h5zTanJOikVoBVIFOJ2TqySPkgVUnCdNI16GmQ6ISztCpt8o61Fpd+jRjdvhdDCz2
2ck27paRIyg/gPh2CQY1+kADjLJJGIrWV3vFm5ao/v6UKqa/VFx9iZO75/kfAjpulz5AJ9gnqYHA
zaYD1ZeMu37QIQAQFCce6VbiAZluveSvLM0xJNEZEv4vYJ3TnhPb57x/1lnOzgRWmVKmQu3zUZSp
kN/wCFLNg/mWBF+X+fw5nekwRFVt+J5P4QlVMWHD6mWCL+X1CK5+a9qF7gFVMQd3zNr8E/2LkNfD
MCf2hPlylx3IlUv0nGg3/j9IqNaEQ4niGtB/U+8A8/EYrMroACAODA+sPyjfIGGI5q1ZyU2uUQLP
+8UzIvKsrQS5BztTyzMtt7kWkq/BGq2dxqwcE1kdn3hFNFZqc1E1s8z5EV6my2googBqjoB6GQm0
23lbujc+HeenJsB1xHml33w4Z25t2OTSxblN3i8hLsjtj32pOaRRqRKCIUjxanLeEZjON6M2pV2k
7G5TABKjmodEghc2ZpmHWkTMWAbXQEhNCXG+ySdjl4uKLodpGoho7LDbP1PibBtAwP/AYRTvFN1D
199mKkVHJK4iOUaX68uDLFpXPq+vIs5Eso5JQE1UEt2cO6DGYL4W/5q6nB4bWfFstm9J9RzqES+E
Q2pQZcxzASHVYkDcq9eL6xTXkbE0EhSISaH9k4uypCPJ0W3XFUeF04ClEKoWJQ6ZFz/u67qjJMxq
1p+irINYKedOZ10Now2cb6IXPPR1wXzWENn7oPtEnxK1LqdHUZyJPDJXL++DGiotvHO0J++1Ts4G
iyelaRfXESVWlZ2oep+Fwy7ggw96F333FOZhjdNnPA+snwmCjuAoCyh1KImgDEoZoAeRJGiXpFdW
EJ02wLMFY18MLACJbKVyuYhWVLdD+QRf9zhZtRRirwSM7Ch5euOLbN02aGmWNTaCPWZVKqkxo21m
H0eB3EqJvHRN45Av8phdKTEe2b7nGPHuUUjb8RZ1dwBFv1AaX7p4bQCVqcjuf8fsB8b2ZJVW8beW
fIKzthWlxYEjeBifnYPVywmHebpXR9WV/bwm14vVYXQxEZB5hP7DlCcIeBcuO3Vzsz2+EiZNnPDZ
h7MQBos7j98qgTnd+r1O4nsH5/oDertFVz8tj9AEu1x5ZnReO07Eftswqybr9RtDTD1t+KkqnO0e
neJZjwzLj0mpG5YnQD0CGCicPGokJMOXbg2bQmg8R/oKFtLcXnZHbPhDvbdeEmHEcWWnPWQz67vJ
c4gs0CSX7XqI6lWq/+bHmG4ZddGxmH0zd1pB5misVrVdupAkwMF6efDmKgb9Lz2nrjMUgdo6Ok+g
4DIp2t25CCjnone/o0PWk7lRPqgzYdvp6uXA4wM2K4xs6GTub2QDfGypvPoVNOHxKox3NXmJIq/c
SnsrAcEAPLc9S5S2UK8AjfMRD/ihgffqaHch7Bh3PPG0P4ZiEr5MOhLq/dZpcfpjks7DtF1YtXCR
1wtsUXB9Ow7tTCNBGb+MqGqwpk6qjAqzFgFk9WlqdrGMbtXrfeqDjdW4XdCGH8vWciCJoc9wiU/c
zfOvpW0XVVvASQU4cxswKcYykECKyr0q7YMn+CbeFOC6W/sLPRPub5yz7pfSR9v1giWaeqz88kWU
Zjf58nMsEL+fcO54QXwC6mLcBNc2rctK2Fy300Kw2y/ixaiYczl5HzHi98XOyyXyn01U7fSCHBYd
lfaP2MazS3hWiovNgZ+QzuLZESG0fdn0pbNUvEn5jMMyvPDFgNecVIER7+KTpBLH5vP0iKBvOrdr
CpM1zgt68YCP5f7VVa4bO1affdAwTDUts89XfOLew80e3Sxniin7dIkC+nC1oZLcd563ElijE41R
gwfNtfwORuhcNsUSAxtDOIk2Wsjyvw4QD8wJUbx4rKyQLb3k2hRUkSAKXoaP8cmuygQl03Ed3K85
/EVr2a1y+wSz2xgKpQx2KF1oavrylQDNbAj3dJVWplfK2t63J8iuf7x4JFUcb1ZfREbjE1pvtFkk
pTl4R2UAOC/fdfgEyRM29/xFhli+zDyEzfT6ha+iTSBEII9mRu2o4phQoY420tnuiekYoGKMF3pB
UbeErcgcvfxV64uFbq7J20k7sfOW4SgLcrnQ+0P40BUviXTgyKn8O3rhf9QU6LuSnSuuss17up5L
WuGbq+s99tsUMDKzeRhXBkt1yOWctv/435rOE9vd8/VoLQrg0xGUt/nQq3BvjyN3i2UxAGjgMGoX
sWjnnlg07wq04k6ql87dssx+nwBP1qHqInIBtLDyOweV/nZMqFl7YfiCkPHzAr/4ExgSrJx34N8d
fa5mahK1daxXOloFfyUfUob6aSfC2q6/NHQLZgmAGZJsQq48vkWHJRX0kN9LulE3ZzeVbIcp+9aV
mLMkfUjIrg5k+/FJrs1tWJqNQMzn392IeuDFXATloJEzAdCSYqoSMoo+mEb1vSD6PSt5uoZpxth/
ne9Vm0F+pe9+I9exUgtZs7lcOy8ooiSgd/bpjMeYMMZ5CvQjpNO0qFyQALMJFCsAdnTn406PyHxC
Y6Rhb5V3WmZrwdzftTsynR+L1CP+T2Gga18YPyhHbeLnnXzz6NMGNyRv+o1ntYJhq+MSieLVK0fC
MuyBGFc7YCUBUx7vb7gi2Kcyd0weddQTH1DMJPbFYa3etwS74Q0cej1nzXmBPdMSPOJuzK8wVknP
eXjVk+gLulKtt+4jXvaXbqNUGA8GiKKHezLm574k+PIEnidCWen3UbQvOWwe2UnBSKatxpPwyX0q
qtfuYXqy8hAgVb58N0ap2bX2Fy04xIGBNsxR/6GA/oXif4yAhXLcgM+GGdYh8QnwitTOk/H+dYFP
t4UgN5GtMB3SOHfJPXOKdC9vbjwkj6BZjtH+slljaSEM0t97JPx/s4Qx2Jd9Vfa4AzpaOIAbUQYH
UVC4W6dA+0dW6y4bSy5/3ssY+jzpZ6/neCjuOgsy51VKHVFMKtWcN0WZWON68ANcXEyUBKhMM+sS
9Wm1DCgRpHFqjM6KDirRPwPkvzn954QkQP5jOjHZtOiE3XJAFeb02l+AILMcg5VhEbmf7p3vHykj
acQepJPPKexKzvkBUsCVT42s5rc2LGPSniW/vdhFKzZhl9sAn0JUXdLKl5pgkedmUlI+KCzi1fFR
ZGc7urE5r99kz8ZYecDJPiTNWPVKdHZQyV91CDnS0ubF35CPm/q+3dqx36pdz5U2pqnITF9nIaEb
fPcXFZCSrECJE8Np9/Hew+iOdbRtky6cWwja3h8OHxD8+/fwjy5KUmZKRQ0Az8PYsXBCqEpXrRVx
3iFhdjJAhokxlps+1YAhSAwSZHCVpvdZykcH0j2ur153nGN8uN1Q5tfVaUUbeL0m3ZtONn5Ir0l9
ig+CvqQ54ZLqctnoHqxRHdaZELZNmUboBOZ0XKKTxyUG8oYc7GhrqsvjblSYD9QdneYykNaGzAN1
B1zUI24XjSX9lw/xtYIg7T923k3fKIqcuoSg+T3RIVg/615TEjLOcrmMzpogwXDquju+F1yMj0JU
7bJ7hligMPXc2KGM68+PJIxAX+xj9rTAIcTR7BagcXa/ZE+YOfb8lewUIV5mhaxR98rJ5HxJQOnl
n59mO7S8S70pBxrydlG6K935ABNhRMPaF1MyppLmsKwSpjD7/W96wdYX3+hezOzuYuCs5s0FfJwi
mNKgE1OsHx/DBNVZ204gzXH0Bxx+y+4QLF+czlqauIWWf054ZwYe+KkY8Ospc41bemw/pFy617Mu
xj5RQzOcy3PBxYhBx+22jTm3QPSVpoPW+W5uhhZ5ubclvtL3YDHUNkba4M2szyZBS5DiJchZb6fQ
1ur0L/c7X25atQFH/t4VjL8MWvXAtz2e5bKZAp9GQ9bRmacQGe7qJiyqlH/NHXp0K3lywPjGzJs9
sm+0YriIC4Gs05JltnZQQWJDhW/xPK7FlGqj6B8dSkEDdZAUdNdDerYYRlasn1ehZf5UcEct+ITo
jM0EDJu0GqzJstBTJ+ge/DdQq2QpaErayszfHAd4Vu/UzIlvFIbhczn+bDk3vupVFn+wmk2cuRjV
yxZQzOVE87AskpwiJYxtOoGrh8ra3W2ORzug9XCOp5epxsmkCQWBnBqvzt9X9/K1fsKJumAUeWN1
xCgX7nPARAXv40kQV0A41om3UmVkXy1CoVHMIza54OpbxSPh6g4YY9vqKHAOPuMdM6yKDMMMbPVx
Dsr019eGn72OiVDU1UQlF+8c5DPWe30FJdlZ+u3iS9zwJ2T5tSc+SFQ6L6Agfd2/lxQmgY8Fowsv
aZATNbBzgeMlVWM3OZADbLNw23/zz6Tqm8MeeTCdbGYjVAYhSQMMKUN2p5ng9jcugztELniXLyKM
yHDrr1NXdrkGr5jbKMdogQnP5nEDinxVQ++gQi4tUy/NJ3VAgCtH/L6DMo2M3Z133W8s4XWoz/NY
j4yexydRWdOWRQPTF1R4qa9yHuJMtEnHpnvSzBUMPKAcJY+lj4H4u23tENn1eP5ZerPrjXmMYSiP
cEyhFY68FjilwSRFsCZNowysFX0GWs6boLWP1ooCTF7rgtSX8mYlKnY/LEUQwyoytiRPUrwplOLd
mao4LptWYr8aFVpBmkW6XXP4/4Xm5+2gcvmGQrQyskGNMFoLlIMVB1NI+S4jamVOzz3q2YRQaRYi
iHzgdOLePsGneXdgYxKSQuo2k5FXH2Ys3qhzM7h2o8bHqi0y8zVerGeH19LWa9E5bcAXXT/9GS+h
EoI67ruTb1mGaPZ3Do1cdr0jpaZk1HPNHDSWHXttY6QgToa/tlW9VeLIFFF7N2m+Jmm91+0c26BU
p8uSnkX1p0kxrY8gyeI9JAKgo67WCWrLADj51jzkawOI6tLtbpGmjsJYhxGlrCenruGDc5uiOuaM
JjMacwtP8hmMc6IrxXh2f9eSCQTtvGhG1MYFkoq+IzK5bTOtUHK6oXMLYbDxONE4GzO2ipI6ZECR
qCR8GulcCjbG3QAfCE210190w8l1Fuxuna1oemVr+y69T4MxEvyrLWNDf+/abck+1MbCTd78xOcx
SULNJqsdYvGp2X1dZNmwAPfwdim2nxr4K7J0dfPjUmksyCxzV9LgD5YBUImUV5gQP5zEEVbXFg9x
NjTCRS3fshoHQxeVZrg5sJQdTraYuhDzi1eM8z8TePMP4aF81LpoEDNWHzbQuoL0YdEEismmDN5o
8KkL/DgY2NpsMDhqdYu63vAqQcTMi7ShYNlP9fjc5ghveXoEGknyqvB8GqDKd9dW9YAi3XQ30Hwx
6cyLov2WKQJFhKRw40P8TfKtGNSkHC5NCM4LXiZBgAsfYtTGZMqcRHh7JNs2rjK5HlonkodX4Hp+
foy8JvJqtdN+UPe4/sd0dhP+2zqjh+C7RUpraEobf1glr5wvYWX7pUwY2XVTH8qnIP62MjsKHV2R
+6odeCGItIP287tHs7LnBR/nTDTbzZ2ynbFojpAV0W1c4QbY+w6vNGo7ibmuTGXTXd6eHFDoKS7/
fbl8Vrm1WGUM4t+MIL8M51TTwV253iY7NJk4xufNWy9Y6whsojZzHbhafzMHG2zxMGGr85G/Lkrv
6idasSn32tfaisxMOqngo24z+fqnp6fafLG/RrjQ7PjEkA9hMVVQHgLNe9DLe++URYKeMn0E9vpd
tcxPBNtpMpJrn8HK81sH8aXvByFAZk8tfz3T00R+hJY+bOddK3A08DGBAf3dU1WF9lG7oXdDIXZU
Ofa4ZSPsygeWXSWJorD55gGv2FhnuTqlmr8QiOdYJQPBl8IdK9ONeX5yl2lEAVbdg84KhUrluwcI
qFNmB4tO4Fm70RzUf+y5LUhkGtHEO9pBl8ZN4fLGBti7Gk7g7vf8T8y9sqYdlYfXGRWM2EfrNsMC
pvqQgSY6vvDniD2FAS+XufmLjQF1//urEwBFp9oCbYpGGDhRoLDKm4d2M0VskpL6HNcvn34CiXte
XKGfjuYQQtE6CL9KZACZ62HHUWRR+sD6Bed2qRkxy1uQUPwR1Ev/n2mI9Tda3vdV0epQtrrRip0q
kGyc3utk0bK08+cvLi308j78h2czyZBFxE1SVYNdOtJxSwR4+iDVJii4M6WCshYu1RVW83Tw12mI
zHcd+vPRpX5wrAZHKu2Kpny2PVPlmYHVMD6r1ikRuMzAPKYfM1o3fdrn9ptwWRKygqtvU44Xyjav
oylHZZ+v/+UNTPQKWrA42JqOZLkE/D5acYyXk/1AwqIs726AdAWwgaj+AqDImdt29gRjuRPgefxL
0fgaxPRMREU9/Xoj8BzEuKUbUuq4XOgPMxzeg/mgdPMO2WuGsD/a0aDN8afWyKsZc5MXy5S87w6u
ivZeZ9j+kCuITFO/iNwPAx/PArpS/Qpg+GIZGOB0yN95J/aweMrQPcPzWGQK6lsU7W8vxY9tPJtw
EC9PZqpwwLVvmQPDGnX9E5xs9MPFRe64kJ2LotkCbiio1xzNYFHs5rAlWVACQ4CqVmy/m0AU5ypq
0jLmXCtGciCRF3NoytA59jdxBPBgnWgENYXUsJr2ZeN/90ni5WYfqllhJKpiXLYTvG9QCeuhwdo+
5kDA9jg28zubf7heTMRJOjFEBKYG2R0ZPQiE5BpjAD1/pDVkBghP5Z+qKmhl7ipa6dO+JRMI/Mwx
5Cnm7hIkD7lxYvQbc1IXJXe3JVZJNwf4rrqGPKu4Nmv3A+h5ZUMAdHCUhJE0lzDmlSxbV31vG30A
Ql5N017C4tSNv2y0/GvB1kkT64vJ+n2YfVPamqx5xxxD+NPWYN8+SCINEkDnJroIDQTvOP9Cs6gd
waMK1geSoDargXMHpkNQJb61953l+79J5nHkkhmZ6rVFZf3pLFeK3Gg6QPSB00O1MW29lhM1acko
cUcMwx1y/TPduataCEwU3BpOdyE5JxkAcnaOfZGnxcom//zNDbYnWKuLr2CeNdoV0/oGkcgQQD4v
Ft3xBlMXXRkK4fqh5I+Y7Hy5K/FYcpwBTYwXCFHMUSi6pD1AE0gHmlsoCpLCGeoKaFk+/4dCgvIp
PQo6pfM85lAuvMK/8P4CYPhMbqWF3Ee6pF5DocLOEeH9mV7Rd83g0Um0i38HB/NlJFgsKIUp2g6Q
ww+ulHSi03nW0bymiV5yPhi/FYQf9HhNocEALdt5z73Wd/A0wCfOsZM6ugm8/NL8LvdNsJYMtJAT
VYTGI/psZfDnfEt9Wo+fcXnR4KHehrK1iC8hqvQy2x48HRXXVkBASXMCRgi6MvrRAF9345iAuDd6
d1E/Q6H/zoeGUkX7n/3k29UgMefqzmiS1aohEguwQX0R8hnuN93HB3RoyM69X4P+GOK7lVL3d8jO
mGoRflf+z58xrZQpX0JRGz3AXH7MrM6RQXiqnu7FmN7TccJkhogqo/9H81UX+t02EeAC9SvYX/cW
N7iE6zOdkTdmQy7gpxGOBHGGvU7wrtm+bjhFpj9AOdK9NQ46Z+Sfu1uqqp+rj/s+Z/qOsx+RbjVc
wtjrH8SoZVzPJsxO1WNggJ4SLA9hyrFLqg+K/D/5/5yHO6c8ruhX1k9MJLsD9MkEuw7G+QA9rkYe
jHBQoX7WF2CCSwVoj8pQ4HxBHh83FcGh/rlSJtYO+0SLrL0Hoj7bIc0HA31U53AyRx/raCcFKL0V
zsY8yYD+g75JLxcme6NkXj4VR9Q6rdQ7zWHr3Ei1LgrKXl2itMCgm81UjE6U7mBYzBA1HhEv1AEg
c4ZxjPsXsb2kx/paHm7u1cp+Cbptu0Y5ynZFmZPcpVkVOcQ0doqyiBkPcLH3OWl5XSEgJgzAeGWR
MM7424Vh8iAh1BLdQFUusoRjUWE3jVUeoQQPMCtR1yFa4GR3NYkbF2fyENMGerYoAQJxMQHdFqYX
SLVJ0FBN8GjBAKj5Gkv8A8VFTWyNAfIhh65frmu+kg//4np7bocUHsffeQEEQDCzltOzcAw59LlW
aelDVUYhdIg9IDQEuOMZtCI/S5w3ZrwwvLoS7jqhRPT1LOGlfW5UOvhb/2URhO6Kewry/Jyt1Z7p
2tpZ83rGsyopWk2mQ3Gi1mAJ0abbLKQPAtgXETKs78FVnFYQmkatG2e5WQUhmbSddrQSC/KndxgW
oaEm0GuDrXURrz/+YfI1XdHSkmk3d4ld2U0AJPIe0qJiwx5tjgt4NuGIDFpGelyPGblWULoD7dmg
IPjTFx8gD0x07Q3nVdIoTigECS3WMuD1MyTb/QyXxy74XEkLJoGUmpaaATCljDekbRF9TCC1MVqs
vRtMC24a/NKpx2j60TUvQCHkd5geEYDDIVLash+QEtyASPjbf4LSfTp/iWPKuxFJDqS+QeL+nEf7
UtnVvF6PB+Twg7Izktn9r6hYbHvYnm+YT+H6nli3TbThqyT/AOMFm6AAlKhO2lJn5XgxLspInpWE
ernUQZG1hdJY3VOeC0dPbzdqytS4hLnPtGhoDu3OMuyodF1c4kRZZWoOZzXa/hmANsYh9xmNubPz
B+hIoMg4pWPiXzTER1OoLR6VPh/jhkUosw55FCazJBMSzacd6s+TOAGfbcLrbDuAbvYa+xVRFX5L
2xk5MI5YXsD6Ibci++LDYyLIbSCTOKaMNFWXx0XfMwuL8TD3xExe+ygMDhr+4DvfDg1Fzjr+S5Ma
U48wuYCggqnRw8sA12jiDVbLU1e087VzSOeqSa0YGlptpz8QSGaA/NRrZdXZkT/Q4JsUzBqoftEj
dbzkxXNr2KwJxFROp7JAy/7DIuTsiBo84ay672hl4dblQK+fZWCBAue/fOrDgNaJnyUDVr1b0f8y
hOUbrzffIWTtN9MtPUwL+hgozOsi8SyRYNbg6JlwfZMTOJasauvkJrmBs+47AdzsRGAPNV2fAHQe
oWAq0jgTaf2GHHLJFOOIMTxT/kw9Z+Ms8ltwV/lRCOscyXElD/kQezz9ZfIaOdeO9vt9mLIbwIFC
MuOCmqqlRrqfEIeQrKNhfmBHnQaiumuPCBHaAFthskOnfPQC1PuI9qooLmZlasYU5TqCt6hAEwC1
T41hYFgsbpw5N5etJLCHrDzaSOKOlOoB7moCiiS8+SmtBQKJIm4cu3hDMrQwd9OhdIOnC9DtKAtJ
Pz10ROGECxgC1DQ87o8uzGu0jLlw3N94ctpFk/s0n14E2JAD6KnJ/hbitCS/U/WTzdWacgXJMOIi
cfiZcBhsOEldWfwCMUJugiXHwQJ7kT4CuyMzHltsmYrltvpOvpjlFromvjnADraAKGYzSdgDjSl/
6cbSzaJBKA6EUJLHxLub7uIa10A18HnFr+WREdi+zRWDOTbvwK03AdVkQCDwrSHJ2Qsb8m8WVVJk
eMdzRFtfEps6Xh9gaFYYei83/qvX7om4JbyYiqvjZY1S0cAMs6x+RCvIYB57jc132L2MiKEY3/n8
Z0hfJhAkSmzp7bgbczM0hXikSz4o1VaEKJlo57x8pJV25N4z5SSqufm7AQyXoHydeiMHK2S/uM9F
7c8+LOwe0C9CKJ0c1juFkKe++4OgvO/WN7eouRM+5dG6dC1UfIF5vQasOIqsC8z4p1VYcqW1U4IY
YsJOj2mpjje3Mc7jyJKdEW13Lc/oVU3miYA2IsKZbXJOa6V2s9ri5zDXKwfL1WEPpARLRRMjXcCr
Lo2d3KQsH92Q7eD9rtV1yrD9+JgJIHKFSJrJMXSTc1sir2E1r1GE40hGKFRdn8npr4Zn7a9wonj3
PEtDFnGJ8IvcE1jWy9jt7O4IEWS6la+mbgRDZqu4i4MNrIlwzgiOpYh0CaERlQLqfFLHhg0EIQoL
CEZRW07W/2aQb8O7qpO5DTJEhULE7ZhB7cr3D8lQhiPHozgI95TfibqhUwWZNu+sHUW6siiP+leC
9eaiUOFTIzZWAAbM2SWEBxtgNaFstybFlCd90T8k5bcU8r5K50EUNUbEDHkx15Gty/T6fsxCne8y
Rl6tabBxlpbyqRo6dbOiIFbCPpuQqYYWzYTT39zLEY4jL7wIJnzFsFS1AljQ9R0edK4bekKxEIEo
+pOZQMOX17ImbafPjmv+vs2vhR/dOjD34RMNYkWTq616EuGcfiAX0Caj5se3+ubB3miccGmWVR+D
RmAHij3mr5Cpk1IyqMoaru74MMr6lcdfp3leraWyvtsLrYat8/LJfIOXb0371jwSSRt78FvvwJy4
T46m24DVbt7vKJUd/Bqw0Q5OJWiyAJfZrAAlJF1FU7tmZ2wG8BDYILEdOx14Z+2x++vzZ+BHGAjn
5WXn7xdLDdkYSCzhHCIGxR0puaXmqG6+2USbxfMGh1cGZXIksYaqBoJ/8R2eX8fdandFXeFubSy/
tQ9fquwo+gUNZp7M+aujJVQzWxwZuizkdinrugowY/iAdfbOpIM2tz6wvtqjYcg16NgBcpqnmEdM
czTSkiAB4xtpbAm5Ux5kGJraiO99HwfNSis29GbS509g5sffOQUZMQpvVAxKQS6Ck0vNC+NK1gzZ
kSLAN8OJjGRKovbvPxH+Lw0tXHeT3P6fi92sllzlbO2a1xRPbeq+d/f39USFkcx5wAPJQzQDOFCp
iydAVdWTRaAZLA1VbvaCu+xOaRGcSlj6aDWsqfzs/j2ktPdyodEzDw86+wKIHa9SbY2rC7jU7J9K
Y6puRZYFdwoONYSEpYMXp2r2BbBWJ+JEq8+ZU/AHVEuDyFrFeusvaiLzZYdmAqgScbaoqkznJjjf
F8MMkSoNQMrRs3cZFZkX7yZb7dYaP3F8FqHQG8tzpjxpBs0y6/kD7huGg5NXucXe+POPPTXm3ZSI
4k7sdCBWWggFYoPv6GMV+Qpne3sTVAASZeoDNnp3qUxcc5cF8a+YHoaEjhPwBAhsXmm8Ejc//lZO
oQznrxLimh4RchMvpA9yEofswhHXgjgm6v6Q4DIZyrURIG7ABlOStxlA5sMBXVLNYMQhbh7y+9WQ
gE+eoRtM9hz+Eft1g5H+cR+TDd2pgdG8c25BIX2SUsHXYXuwq5GtYvMYTefo2U0gxZdo34V8KZBo
RFIq+YxxzbFlHykV7vTC5dettg5BkQ+/hcv/www9If0hGtROSC2Qnd/7PUnpqxp5mbxygYHVXZLn
zv7EZb2elLidg+3y/233NnZk/tqUKs9mJCj3eEr3tTgxA6UPMEmbYiqBJB1uKR8yfYM02aH/CnSg
yRasCmikmYwgogQUa/5KckrlrIxRC4Wd1DpmYwo/DkrCZqNMlQ2ZEY6rX1XO9dQg2S6N63hMTpVd
DiBn30xqDqRHEb0zCysY3exk6dgOnLmTS+tkQc8qa+wJYWcBK7ROHEy8+p9CGabWmIiJ9L1h5hiZ
c7A/fCidrHUx54DSW9K13RJZYkQp/J/6sper7izCASHLZm2PZZWq2WqYyQOhlc6LFS8UtsqLJBks
TZ3em229B7JfqRRQrDIBOwEAAa1v9WwXMoPai6miLwE40Iurc1dPEfbOFouNAWfBdJvFw0Tx7Sh9
/RWBo/FfuRW2CGteh91lVdlj8XXAQyDF9ePbOwiaR5+1NEvb8/e4Rr/++T94eiwmK+RqWT8Bgszj
7FMuq58wIF58BhUjZe4TS8RNmDhpuuNbNRvNtjXcJCfN0GpsOkhzEicLIoPX9lPVcIqsnys4mfYi
MuCSqWY/GypxeO4bcPBMTZfm7ZGcoTxrXFla6IW/2y62thhWBsiWAcxRNf9CdzqdAeae1bbMkgFT
9AWUOvUmBKaKtk9xKMY/dWQnc276al18lGRf4rQmmPtGvMHyhrkX10yGiudn6Glya/1bkxDZACM7
vO2HbOp9ppaU96DOG8pc76YbyUceLR1Y0VwXXFeQNCsX8L78SNHPhiVEbZOhF7V3KXn11BUJ/6sp
sm0lJm6nhyUouKsWD2UIXUfX34MoCrUP01WA9NgfVsN+Be7oDdBh12QOjTcjmEIf/ojS6z/sbfct
BPE7btFbax8AU+xofjXOQyuyfeKZTTGVH2lRc+a2ffEnSMsL44u3za2KEzQrpOHiKDhVxLfy9PQC
DNk3XIVyjeqnXvHjkvn2qHgT4WZSmz2+3bEgy0CrMCyNwEtHTZOUAjcXFkYp5+8ZAlcrgBHbalC8
5vp8toIpdlEAfHPrE6CJ95/AtPUPG//yxegTLLwh105LfnEOGwWfEYwRbcTPaN5Ikv0dYJHdLgjc
QcNN92g6wbiH/p4CrBKmD3X1j3bkUBclD5v9NvO9WJpxWdIeOlmQ3R3jNfAhw1w/bF2VKTllB6/N
Jmq2v5vxXoeDjQsjRrSdcGffXCYFuBNq/3+mG/uhrHb0mynN8w39Ma4wrxPi1Oq2XiUenMeQQzk5
C8Y/aSy7RnrnnLsoHtZk8wfgKIMjCpqWu92fUYzDj/XNubUoJ2k4x/tpVvf6+fpQ5JK6aMjkDADk
LzQPrXPep5clTLrOmF4t3zekqv7RAl3qhfoE+MAg15Xcxl7QOubhO/kyh1x8KdJdrsTlu6EqgobB
/SNEUCAWY45vAjlNfHl8IVRvv8BVB158kgRJKcaAtdYAE9jehK0YecPbEUfEhIKUk7uGM3zTm9e3
092sRd7k7FbD6TVFs6FZLQog76cs4KuftTozo2YTou8bilPODzVvHoQrSZN4m4L3L+qvf837xR9k
jRLWbyLmDj62RgFaEg8k/oLFjPPROp/BjrQiBJKB/lkxJP1DWO47BnNxJr4SANdHJy62SWXWnnWK
2L3RoVj5BBrGZr9Owti2QDrIhDYK65VB71kcj0TP4e28BgcuD73Z7VZBs3y29yQzrOkTF3cEkwxC
vGyHwv1teGmdcfnGnMq/JcdhroQuSavESPfUDlNmts1A3YgIQ2bv91mG1T1Wp4zY/ILseFn89xvM
qFH3EPBt8mpCQ3KQXN+zRPdaGytamhH/Ji/d/mO7Wn/MU/qfCfW7o+zYdYqD0eV1t35PbsPSX56J
A/+MJRdsTsxPM0XYqjBDz+s+Zu2O41KO3lttqE8PCgJpnv79br+uxiH+Cj4wSEKQ1z9/V8bD1OGj
K5yC4mm6brhOcV1UvAj8A2yfCAKL7Qy+bfcNLLuPRM5lFC/eat1phye9JBZMBg+k4GiTOygrqwRZ
Q+9jhnxOzmq99zO44pzTsDIn1+mDuhJ7uqo7BCIxD2uTJ5razVNVfs5zxygaEa88LbP0A7U1A0ex
MUhStitN1f3uD2i4pfWnP5508SCmQMMGM+hn730FZ7SSPT7y0nbXKWoNBiV2aEAAWRV76RfWR8hE
6GVjMRC3vWW82ZvR0Re7JHudgmowMYp0b5U3jx3kTuBgRFGDt05vLKswMX1QWNF1yFyc1VK0WfXK
lsunVX61D+96U8SarGYXvSSRiU6BSpQ6bIVAhtdlfjR1LGq3RIwGlE4jpeVkRyxDSjmWzPq24zH8
KyNLl71XZRXXiHt9tGccqrftU+2irdML+UIOaXHEKguAtQEN4kim2sRO5R2NRgPQ1LKx+PX2s96X
nBuNc0oGNVhsP0ienwRzt/9T06nNfOyov7Fz29JmtKt9CZiPQnp8Kp5RlaAtXb5+7CNFWN7EhOJ5
mGWhaWEp4qX9UOH8Dlvuj4Gn0zKu6QereDXYpbPfxprkBB3AWGXv0KGAunC3PcHXIvKqNhgJ+K2Z
JT1LZjftL0ps3hUDC32WAquiV1Pb9E7bJLb8V2cAmukKG6fzu6gyS0hpZIdouPWn6SSNtI3SLiZa
x/ex1/yHpYo/yJuwW66RxwYjyZqIHM6IiflXE+a3oApR1X35w55vKefSs1wNzTuVNws6Wx5UISEC
A6eFX2elWqXQomKRMedaf06KXoRJQhYFDvXSRizp07ayDqMXcwzt/c5yEn6zsVKzxGuw/1zQ8Pak
0rWzbJA0MA2tdRKE97i2ZNJ77qBOUPEVpyJe038gmUNgMMSpn2ggBIuudlp9TbvrAY/x6lY9Tnkr
t1eaYKVW6F1Ep2lCYHZr7s3koKk1HWO8hR65RsrMK2/+4uKRZWckjzvW+tIt0v6h7j2kugZXJDNP
YUs8aCYIALrgGoUOUCjZcP4Eyw6IgQb6Q7B5MPjoja5MEDtYC6LGZ14SCaMfTVmiwghxw7ieXx7Y
GtUVYL7nIAOg4rEc8io3QyZukyClZd6Ex2KdKxT3t+bbzjzSOkA4W1IClqt3nbN8B9G60QOurTnt
MIU56HZ+im0FCCIHH8ebKIzo5VztCsQHzV2sMvKeUjlMb3yORtTsehOvvua3TLcEQbNEEtyptct/
HyA1DMtsVrljTjg0cEf8Xhn6fBYugrXDJ7H25heOXqr8DmefxiauqCB1/+80nawgVuL6tlmjpEkY
j56aBu74HanU3M6dU5GrQlvkrEu0gpXxmg3TPbR3xmcr1KwiMIAzW+eooVf3mLSJxbwaS1cgLYmd
wqXOX+ySMrQJIYoV/D9R070Cw4C5x7RSHKx0ctNlrzKrg11foWluy2Z2Kzo8WUZ15BTwTYlV3Snv
sCl+wWemu8eKz+OVOEfLnu6Eqv4NUF6T88j2L7Pj4djv09IGbY+jzK/FwOiVf5Ex+XBgXUZwe2kY
Ut2HJQLTX8K8kvb39bpwuYU8In9OJvWK5GYP0LKJ9/BAC3SRn1l5bzIuRDJAwlK6/m8BkbxsBlhA
KO8JY7HVEWcYegf8x51yjyc9oAAA8ftv5f8hVabX37W3y07VOlBz3OuoySzLu5vs+NCNF0YVmDO1
mtOrUx/5gm/NCucLVKXsBe3DSG/1TC/evnA9xpXV7ZWytXk8kVmgfSds4Bntq5Exa1jXibjahxot
fUGYBsCOovDSF/359ykya0CiBIg7OpzsT9rIZIH1l/72dwyA9gWbWbqpnFzcNZ5+Cpk9JABDcI2d
I54t+CqoC3HbHItll+BsqnxbDqOnaaxyEU89ORnnS4y85Nta8zbv2zvr2YbTJuQwcRLUEBzAPeJp
3Xxc3GTxFMTADx/u1BtbWLEOxlYmh2kO/Ih0TQWF81kpQ7JFWVLMsVMzeS0xou9yZKn1aPy0RY0A
zNrlPp8Jguo/Gbq3Z15Mf7vDGSUptvDGuEIRl41301f05Y9CJDskRLA8qq240bP22Qpgbn+2Sbnt
caMd8x8otasKP/N6s9hpjwC3AWvDe38plOepwx1Kw0YyjxBOGyG8/wG51Xd6/KRfFnj9S5DjRnVn
oz5BnWsUq29Yxn6m5GwHpFfAyAy8fBYJaQdwvBY9JU8yUqut5fNUfT2DnN4zjtXmFO/TZh0BorMl
SAcqVW8mzq4aGaTpEJJNaRgIgjuwlmG3eON8l8jv+FMKXIJNO+HW50PmsETGRRoK0iaD3LQPSiVb
EFIP6XScj90I8iyPskr9e4qvBdyCzDL04iUh2Wvgo0haiqz5L9ZjUo616xBvTPBRDeOHbU9GjkZK
XfjI9epfSoMursE+btyOO/Gepe0LOxBJK0kYjsrWjQ7vsT7mO9VzNzI36VB5T4n4U9Z4mOoRliyq
fS6mCt+wOLrOYqT9uSNrg5E8k7r7Vf+jbJmMZdaC+QzqCqnDBbNWBJmejDB0htPY/Pu0if6E3AGt
Gxash+TqQrMRbic3CO5syLew+b868ncXIRflBx/F8ylipDiQgti3gbxMr2AoeJlK+CwBt8x4Cs3R
FafIxWB/d2Zq05ZNjxzu/FQh8i9R4T/gbAkTnMsYgXCBMSNPz8yUSTBgucm6VHekm8GwPLHC5b42
IOErz8IhygcAc6mgka7xkfbSVe93QoD+oKCqolpMrl2eCnL2BJBX4lan/y1lhXSxBtEXBmaVElrU
+6C7GflHZ2ElyhA3ofmfoZKWC/Q1t1c8rPqJquWG4q0VFbgXzkABsfy6foTI5bblghCBynNzOJ1s
L9gCI9XLunGyH/pOtgcNmHxXv7FlBe9d8DTMtyolahhTtB/JX7jaWZMStfYuS8PB0KsmRc2DDHym
y68PnMUXkspwmbyJhtQCGkjrb3mvWSpGDkBtgzUcfKTArz8MDQ+8sZiBse7N6+S1qsyXNCQGelLp
4qOGOm2Ij6p1c1IlaWLJKFHhS8/QMgrqxiAE0OjiF/6ttsuk+J0h4grH3i6pK2LUuYwbKv9P4ICU
8vmQPDeGCPAFftLcxOy91Y/v1nH88HY7SeKIDFP10FfqZb42LbiRueiaGjbai4P0WZVHcp4mjOfC
MZuFjZMAMh7MeAyE81fwgvYb4BQF2LbO0l5QQaYTropBe93zfIA+YKHlMRt3U4zHOmiQemkt9zq5
hm/8ZedU8WMrdxefM8rMQO7OuK+Mg+JVkUsUzIEJRrGXovozYXJq9B1hmGehqDmzMeBQUifwwhVy
oK6a9PIzUphb9ybK4SUhQegkmkxh3jEsG+JjEaqSyuf9SMfTOc6wXwzPqEjRMjfCitR4mPauCDYF
o/XibNz9uTP9wJ6OVOhT2/j4xO4bMPeDEYI4GeWfR77DrJ/1q5deMM8bhlL0AHjSpYEyOgOeielE
t8fmzcp7bF4752El340m12fVAFk4T9FtAYtZFqLgraAlWmnVWHbrgQkm57+pI4RiJRNA+uLQNURm
VFhdHUNa/BNsnKe3zmzYQaIJn9K5qpjr7RjygY1963PRur0Cfh7zdLKfx7KzntitKCIni/ju5T0B
Qdh+ylxuYI2+TrOW5HioXKO3aWjIU9ByW1LB4ngkJEwxzJiUr9ooV9vGDb1BmxN8qnofG1J6kQMj
hWAzSRHVoqRjSNIIUAd5w6ItI5efpt8wlP9Vk5i/d5/lgJe9BhIMzQCbbYK4rtUkz2HEhpamSbKi
PSV92rPf/2xfTNn6JoumVD0QGIEuRdPt/I0+XsKthJC2tgoStio/uKDsLrV3BHPYOsz1lWuybEp7
ylUorUEkHxq9Q497qapCwROvbx99eurR8gOjRviL6Bdf35b7I83avqzJ93cBUqBHe7rS5BHj3y7g
Z77qNVphnqje/Gk9QzI95dPmM0O49adssXrdpAUWsIls3j0BZmqhBhQOpjIJPZWAmVB7fV07GsAn
QbJ7hYg6PkTKXH/th++6D3Y23yN6Inrq45fugwqvywVY27/R/k3KybZbHFKUevHh+zsr/Imvb/T0
4wXbx1RfDmjkNjIcQV7mKc6wjSC+EuFEPHrwGMOdZKDfARcTQFF1RgZyY4N3Tw9yr7UKy3TXf69g
KVRt++VKxR+5rAh4BV1PJt3BH0RGarPiP7HPWhDeJ8sfAZ5XKDxe5+u+1SEAq+OH8w5pSblYyezS
0wSVSrEkwPOrB1JoLsm5eOs2wpDh/lZPtfnmkc3iVy/Mv01qTauhx1kvEYzjcrYk+DuTR4dwbJQo
CqO6b/gbskQFaCzZdRViAai0EBVruq+WUXFLQnDSoPq+qMc9DjOiCyyPfqhMqGfhpEmn84ZmyOhQ
s5DPle90Z5d0Sr7iIsUCsaT1apP0S0/pJz3iC8aY4QyrH+MYLFlKCN2n6h7FiBFfYNN8Uldpa5WO
rJyQdZel0JB7zmx4xY0SSzfMvshqJjiQbN3YabD1JuMOnvbM75M56y3iygd02RalKSNL/wqoHXkJ
1oIPyzVEGvd7C50Z3D6D8dSiFS+b7gsMeZxVBX2RDucctbPrR6jhVqmK0YFeK+BTa9zgpwu50s+p
HFYAbdo9pxcgbgDq9Hou3fLm16WtLQmPszXLL/S5xHJF/bmErmtP26ERu2E1m+To7aysZo1xHppr
TaGrtyyZA/ixqV9XHxf/7KTJfT81CmGd+pCZ1ZjoevE1i4UkQgCpo8dmcoQpyM4O/IEwPcqrDkyU
CSyzbyj68/NifzgRJi68Ttwd6dM+GHDqNEwauwGxl+XjQl5q7Be/Dsr+AZbyvv3T8RcuY0EcJeJc
hJyfmhwFVSmUhcpoMYgM+SlZNj3I+OJXfDTMaO5Z1z8KuSQzQ6+8L99eb/TjxQXJ5jD15HWaOGw0
PqumoZFxDp0i386ekghK/skaB6UuBQG64jCAOmnTSNQ1SHVpbEx+I9W7cmpTMcDmuXa357WhJXdf
mahx7g6I9OCo1Hyj10a1m5yzqmIWXZzqFhyTY3iBxrUvTV40Qnh8Sr8jry4OjlFIMU2JG3pymvXu
thT87deSj39guE5KCSKayAycC91ZVtsgiUnZ1IbF6rELVi3e1Jj/R1BjghRp8sP1IkpUVhsgtxYc
EXn4rZRYWcWRV+8fNy6kfjDDjEfkkSs9e6VHpClPKnglMs0fcfSrlaqwveRZwrZjt4xjgCVJPHLM
Z93RW71mP0jPqzXPbIzbTUnuqs/P2U/bHB+0Z8dkTJHay73ydzCRfuWe7lm0wUaqJk1FKKhk3W2Z
E3gOrGD0Ohv+B5umdGdjkYbB35WQ6IphL56PLnE7cYdT/bhwlUWdjsn88ANiC5qLfxHFAyITWyFE
mOV8LeIBKx6vW4CU0UrgHIzQ7T6lw2rXoqfSe1rrbxh7G62n/H3v2fEf2OghiJnS5gsxPNFNTJWM
zzMndxcI8JBiBX+hMWYUKwmkbYzxattzRnm9h1TUAWKxVfHLMcgDX//JZy+w82kRc7dbvnwZggsu
QER0y/gIWLOAoYBML5OorikgQH3CN8L8FQH58Y2e1wzIfx6qZvQbMMM64TkbKZy96o7OLBhdGap4
F3INOR7W6d5N0q1BYrc9P5R7xa1Y4A9sZfDXk/14P9J+uXbWmoxXsExpWBgk7DEmQRis0htfShMr
LWyzN1VyEmQkHd9XfHWt1nqyhKwaS0/eHcdOcW8vIeumiUS5og0tL9G5fzJESd65/r2Qz2J/dQ6s
unPIbm0NJcy87tobpM0Gf2Yq+01TKCrhmkJrqGnUyAE9qYlDYJ7Zguwqzb163cXZXabkTOGMkzKU
3ijZrqZbCfla81UEyvJ2bouo/rLpP/XpxXjjQdqIJsjjjj+LQp/PZIi2zPAvJ5vufIb8zGvoomAU
KbhNojo2RB+YZmzrwQwIpB9lc4kLKh8PX+JLY1AfmLf0gcCdlUluMWI0h9vqlGYFIWp5oLVbIhpv
cpB3Yvvqn8YCTdGTA207XczS09V+Ad+KOqL5tSJYpWb92zLkq0n5NFu9CeN+kna6JmM4vtKzj2Db
yC5IgR5WJMtR16UG1a+/dYWV0u30JxXoQfOb3N3aKPSMjYnoq/XtkUWxqf3UE4JKuCAYItcm61tq
gkQ9nOyFGkKRQuMiY6b74Abp7gGYEbWcrc0uC4viCRZQYW3NdGlC4AmxyOqFCmxQ8I6kLHeSj7ra
MixAt+oNuNNygnLCi1FSlOvoEFwGrcpB3NugY1eTSHKqjO6dpwt9MEJ+TNMsgMpGDn+8I+PyD3Kc
nWHO4OIdx+Qr232XwT4pM5DdFToA/YCuaDofOsk421ENkb4q1r13IK4v1AhG/5ZxBOQdV27rq1I7
G/jX//TRshXHzbb9mtxtjq8iBoQ1J7Exqd2sfRePeXei6IVo5S56JOFEovMoGvkL8ZTggsvv760q
/HAReiWMF+OjbSYxf1WABNjey1LEoif9Dlupro4zoIqfKnWVm5AgM3J7z+34YFv2oBcfx67BuYQ/
PLZrB4ObY9w9wNR248qm5n0x3hBqlsP0RfIaiUOzDNXPX5eTDq92oduOl4y0uPxBRmiPd5+v1HVC
MCcHo2fy7/XSTIsWEz0013z5kFfzan1T/1+zU/eTtysZWWaDj+Ivkj38yOOoyAOYzO3kTpDa6zEt
MyAGxbSu06qdgvngL5Nho3IV9g9Lug20NdRaEyClwPs6dw3NE8aNI4VcK5ujBVqmZqJMWOC/Ocyz
VNEwgciWWuBhytgqxGNWZGtoE+g8bBSB5AYeh6yrEqstOlVmukIkbFNQYo0KknEaSuubNKnnbJsE
8HHnwIsZK7aEd3ttPAXPneBOMky6tV8Rehoqn99FQ7hluSEKYnH/MKzCjHuG6H0LxpTEqAw8tixc
DQ7zW0ZAmg6k5JoSY9eonZ+q6JhthkGSVOO7bl4bh8qlfN0wWP9rdZOLhwf5XTOKQkt44b5NW0hj
AOxC/2ZvtC8Iyuzzoi8kmwBkzxpi3jkyGOaRAhKiMkcMuIRiCSwr2ydwQ8lFAezx5swNJrhNh0BK
6cOiCEoEzqnAdrEdZslaDuKP6IDh7zzktNNDxWD4yYLhKaae3iVEhI9WbinqbPj2qAa3YjVvhEZT
zzAPFUCP2DRN9TaeBLwTNu8j/sC62Jt+qV7emy3EQermUYviCXY76GAE5A+A0XbbFRgGTMZIy7EY
BLMQwmgrzby7fHj0R5MheyUkOAKnS79x+8huWs4w6q/H8lI3HBg2DghfJufuZd9YybAMp+ZURSiO
1vC4di8e0r56DM/FrQfmjzFQH/hETd+++dNRcjszb726FIiUVv7WnbTyw3f+beiMJFuNaGaSkS4Z
ssq5hddo5cxYw2vzjra8bxUpqvFvXHzxz+NiwanmpSlYcFjcYo6lDqUOJ+Z1XR54oqobwfAM+8Us
NmlVGaX1PaimDsY2CZ0keerxofjG/SwzdzRiAMo4yCaPrw7pf3kJQh1n75ZLyCT1dByahB66t3ya
iAPSDARg60eC863rK9PNb7voy/KZOq9JWyPvwknzvjcROCzMBHkhXxCNv/5ZHqgBuKvVXxT5JGzk
e3kEVjhJJUjhzhes5jefBiDxkk9uHEiPNmMqpzsU5dVqC40iAYlnQjvNJavLPxCCVHXNZyb5o6oK
u1sRObBtLjTKlKYMxrFRImVMEkKnv5O83Wd/M/FdX/v4fESg+wK2rrILKHyvW0Nkfya5CvgvrAcj
aFkaXzqBktkiPb7qzayULmJlfz200k6AjYpAcy1MemFVmEClYGUcCSH0MKknjYD5hFdKC09VmEWn
mEf3oM3ixUlGuRCJFQ8pSwP3air8S+jsTWH3i6tEc+Z3Y6KElOxFJ4QvMZ0oDZPTJ3uKVr6gXdk6
Raxo+/FQzAXUtKWu07r3sjK1JCYgBElVxtO8YION8sLVIKOlKl/Qf34KQTVuXUYUvkmF8GCnTXd4
B1/5+YYQBMK3m6fdN1M5FgOObE7wwC+vCL9N1yV1G/rydRQLYnRbVeR2gn8XQtEhg+hFJQ819gXM
j5C0cHDzamsbZ+PaxVeHlLq1xAcvKYVks+CpVKY/ajfcLIVvECr3xNBjsjeALTLH2uefkbeDozy9
1/5dfLOcZWjeHahUehUdLoFLBn9eDFuGcDLawjw2fV3MZq0WzunEdU5bUPn/eeRLe//4H5VQ+C3Q
KwbhYur0O7PYLCZ6HPUG4e6WDiM4ain7Z8VYHAPAAOh2uIjtefw5BfSzmsF6bX9ZUXPZqPs/ivJ8
kh/V6zYPSlitI5rT8u031R/YQ7WsiL7f4bh3fVde6t+feQ7fli7jg03utMzvtJ0tirOSExZmYlw5
84xJQyNYzrjOX5j9jwgCLF3KLfHnNYEoMNrUQ2LEF/JZqpesxuARw9OkATXA2nlYGz/rl4hz0rWk
M/4FZowgeuCE1LORp33eH3qmSX2cCBskBzH7tDPH+pLQaN45n4Xmo6ZamdvEe2Fbi049/A6apNYc
JhbL7OMoi/MVnjX7UvcPsA63mvCOOWSoX8fCFxwUmMQxBnxXKCWl6/4b1Fs7jJBLoEDxjB2iUCta
OyGjHLj+Wqqujj07y+CCgrdBZ8k80lItRvG5EOyYRHQokbq610xE4/s8tjb145/bYp8UK6z+D68W
a3p/3DiV7b23/JoZRDz/p7BrBAfjbzaqbKy4ORctFbG19v9QNpJPfz0ZyCTB1lWnFOSpE7PZX9FB
ZDF+44ktY/6vaOu3QMk1EQfZaAFV95KfPXusXq0qcOWkBriF5e+UNGh5BrpDnKE3vLZOX/C8q19M
QDwN8FVRMM6OwClhg8OjLqE/pKYw7NOkkwglNJiDM9JN2d17ojX9jDariUVMPsmZ4u/r8rUwYgJg
5aC9cZxHx4ZYHNoJFZi/Sa+ytpMm3EXuXdVqi9JdDy0reb9i5hJtS/0UbfbMc2yHFzXLiadqf7iR
Gan2sS/TPlZ1RFXwVtiXzwmdnUjyd+g5rNACh+RUpvJUH7vQfzbEz+dPaKV81mw8nT87bON+5akJ
XxVSw8Xx7bAZbg6N0KXCaTNUP6i5866MC2PUvwiKPF7sTo3PYpbTREkl+lsiCCADc4CnWhx4Nt0o
i1SmOFcN0hR3vTwvep8pki5GcdeWJH5Bd6p3jZ9R0WiFTGnA+RoSJbTZtKDUUYQLdMLf3gzzHJtu
KkzYXp3iUktEeLSBkyMURrazOxn63WOiXT+z3626V8cUKNNBTpjD0lJmLdCSQ8R+7OrLODxlX0/z
JLt5Kej7Dx1ASA96N5qzkFOmgqRGz5VuNqfXqNM9Nat8+Fi1mJn/Duelqck6EP2oZCoyjWEbYYmS
qFlLCkc88nT4I4g0eYYUxF76zoiYbxLYlG4pBET0U8AyHjL5leV2vMFxb6fPixe4LP+CbKip2XzE
ODtzK5E97CmRrsp6lpQSVj7551JuVQsM+QUVeUnJt6dLO++QRsAR6sS1Ds1SCbmf9g5eDrkUepIX
MQxG8GsUKFNJteqrX+OLC05AC/2z5zrvrXbKJ64xym//1cWOIYUi5HcqQlSxxftjITfJpKSCeNmC
Ypuq169XlCm2zygBXI/37I7Lc7CYo9y6oB0Quot2Bba/u7wqG+F6DefHHNssJiLJEE5pR0wlN+sr
SeN9aNf1PQtG2QZWbvqORV1GcAYADuC2FlFGB/FvH8dDAYfpQbckh5VpDrMejL/TZ32/JHP/dTcx
4TGrFWJeLnFWYDJlajAUaQtqGck9wLxtBKfuxZnzU+ddHxvXq0T0Bn0+RlakwbazQXzKPmt8u5ZV
qlr51aYwL7rrQjjrYJiIHjfDjLCjPXMbxo7KeoviKkQ/xb1XdDtWqSfPi8qvfaUCPAD2U2XriIIk
fZZ5+jxWKQAwVeKDDlNNheGywkVKu3cJYtR76JZ/wA1pwED16EwkGpl1bdK4vlIllSIZgk/k2WB8
OqFijCz2WCEt9MSZWzDobQlb98dnUYsi4MvCoFjahHPC29XuUW/29QGx5X27+FIecTH7HevLGcvy
UqXMUoMMByxTxdA+exp3c41O6kPMJFUd29hCAR4lAdyPCJRofZZNnHvc1oA562QtwaMugD2CU5cN
1n/CAezmpTv92ICSvPRbyovGEBVQFJzOzzsa8Vghe8HeS31aeHGRmDOYxDCHFVit5KDuqMbPpcV+
59oRjPMHjPCcGzqkIEN9Zp4DtWgcN2Pbt4aY3/21QBygIN0cknQOF1ECBK3indq5CgrtFJiequv/
ihAgCBOXOMsFGW/wUfq/mKqLSTZzBxse960ukbhnwS3qNBF/F6RNC4Wl5+brWQH/P5c2O8oHFScn
YIc41ZGOHB29JTUixDVFg0K8l/0ncIz6WNcIEp1EsKcrMxuwTZe/U1ejvQrYm+X26vwAdPHuwtp6
wzO7KSZoNTCtLkdSSHH4OLVVTAabk+ABAs/FAcfgbd+FmwoeJR7+hZV4aLWfyhcWG3Qu/ZmyyCLT
lHceXTnfkBE0hIYsBJIv1PAKMuDSVxLx6dBSu8jtbXX4BIsjAVEDRm8OMyxQ9RexoeCwHwobp/+w
1JbubcFpIAZMxrOrNHb+L+L+DC/3Qa45MSv9c6loTNFbQbK2igrsOzM48XT1bmaIxa6siKXSvLAU
stOqOLwaQ0+/6mDinmUWExY536I8beyzlOYoUYNSlESSF+ktPBt8Lk1mXDqv8PQuMTQawx0XC72t
19lAF1h0/Z9rqbmB4AIZ8Md5zOQ9ZTgiHmmA0C/q3i1XsAJpIEiC6b2aKsMPHHv6GJDTEXcVC1Ks
xmNrlO5ImzDjlx0wh28Yc/JuVgMfPWpvz4hOpBgQciLuewXl2Qdq4rb6HS+WvIqg8805kpdPv7sv
Wd+0qh+bv7doSHHIh3THINUiF7e0tbsdYvreyzE+DAnVjpQ1+r9PQ88gq8fyrbX3TbvadIqcgoUB
aXsG8NjVMBVMgCQ05bxPG0mR3W8o0TnkTqvxTIDgqOjhNCZ0pw2h+706G8OkUZ7Ta6R4RNro0MZM
NwYDU7mXdEMcfjSzzzrbdE3LmORq1qBrzvOy8H7AiovdGphMTKP7zEysZaxn+747SSfh9Pdkmicj
by5zITmLBkvp0263f9/W33SCBpvGtA+j6t95kwqOhy99kpBBlbf2SwX5GAmNFyO4U5IH19Am+iCR
l3B2Jk0IkEgT3Gvpb/gUhSINzZ6hr0b4JS6JRh1jRZta1vmpj2jlBIHdmncKTuPKJBhH7f6P4Nt2
k2CYC1nckWdd6z/wOTkzwCRahrlka71zx0zZL4EW2+A0mbh7DysdisnRAogjFeewM9y5yaHdLlwy
sXyFeyN8ZB2J3H+OGvMIgRL3Jk+ZLL+CWEx5jwGOcPtcW1h4ALtBKgcBnFsfIGj9XfUaYK0BU8Hs
9ljgGcg2pCFcEyvoA76bJzBGKNTAqxEoDBS3kRDcNdEilZV67z23fjXcvd1aMEeLa84S1Hfb/VuT
zva3n4DwX/lfjWVQ+fLGtC67FCDTe34E5DGF08ARQmG7Fm3HVbu3zXaXuHvfpB+/iHarww9shun+
OJQLPVdoLX4iaIrLy/ZXGF0EAupruJsZmoWNln/h+/8jLPR3d3xHq+QTWy4WnZGjITSNod+FiLgt
BLEJjtgkND+oMoqFQGiNKpQ8FKxWW3mhjfQQw4Jvm+K0P15CYlT2WnJQbjtd4xMhr12yVXKe8i6s
1Y4nOSiIUddCUc/oz+afc3inTKq8uSqIiQf2VRbp0USwBpCzhm8VS7fKwi3Hyuyl2NmoJHCXmq6m
Tm434jDj6NCwxPWaMj6q7ASLtsf/uPfZPTAUHx0C4/I1RgQKtl4++HGU0yX9JWYKO4DxDevRzGJ4
qYhKDbgdLl3ij/27Xpgcxl6wjByGT3eLZWWszDwg9mxYERSMboLeXJ97q75tIAeWxCa6ojc2UyAR
Oe1LG9l2Nbxa9HoPH2ClahmgHK9ihNXf9xF0Wug3hG6xIrQYlbqQXN2ieuJKXQAGHX48D4KWvCPC
hnWFn8Hn5/0h4n5ewTBLoBmGB27/c9uWWIFh6RtvtEVCpiZf7UE6WrEOtRisCbpjNM9HTfSO3VFu
3LoN9c3Kwvpx321fGggKQT4HGFBIzfwJirfDVaFZhFZXbrEy3PF8y7IF8wQTMWGXZsuV8XVkOfI/
zy9msNk8m450mh+b/4oBuAM4ppvNkzBBvfS202swTVZJbQxHgQapnzQO1pv+N63v1mDklXKsc0Ci
DWatIsEAx+GuA9IeEeCmi0BoJuHxbVgGT+V1Z3OtXgJRcHbd+VR8oskJgJDmgK4e0Yp+nDdE4wwW
0YIC3cRH6LlToAit1gGJDGpp+Lt07UMQWhxZCIrrlhCqMshoxQ5PGjn69+RnQwIcWYGwfUut6DY/
iiC6NnyMpkiES2Bi9lrtSqFWlCp4KKjmHoApRlOpuRIRQhG9zNSBDnawNTHMNbQv2l/rqELRGZ32
hW3I+IDA4Uivc5kqlpJupgKjJbt4kpAEE1fZ6eYnv4/82BQIt+fd9FnNuS5ox/zdJhAv1UHYfvNp
z608CA2Bo0w2xzWF0IbFfP+LUSeNU8lkgkVkfG5pNRdwbm7Ab0jdwH8JEZw8WHqzmMdbYDHhC62o
WXmQIqySQYeq1Kibo1f2TV4/V6DJhuxFPBXXaf1G+D/QLCMk74JK/K95np7klnHIEBA2Ng2E7OIM
MCOjA15T0CBBWEO8/Z8cIXLfb9Yx3k0EJEPHPeSQBwA7JixHkTBQMX9hLqb2UPPyjLmqHRP7dVt7
p3cMky+C/pZfCYR8i5/oJvb12wlS9ZOKpLa8YFiYISRky0z9EF4MWdt/SC6Ucjd5Op6Kth0KSJPz
mB6jUNtxu31LJqMfgmvU6SjU4DG+LFtT8BBK7aWmyFOJ5aU6M6BBLrbIunRzsIwS994ljBE7u0Kn
fLfa6CvPNxf8LakDrII8vsY/2nfoMjjLdqzjfeFmQcf/n0XvB8cFa92Ioa4hb+uJ80kYbGnAGCSi
1uFrz3eAFAua7lo8HaiiGQGiJc5wrB1DJ+d0sBDTBP65JTQvdvCfasRuD9Cdzkk+dDsHVHLxDWl1
JHN4d621KdCDkQOA44tJWbc/XImT+A6yQjeHNwqsC51nbQIl2pCdOV8VFAcZj2d75DF54IUglkR1
K29N8kAOIgBQQ5zRWWYXgQ/DsJTxPTdKR3w14fM6nIF2x1EKGdyU7DWnAaLwuL6V5Tnv3W5v7hzO
t1c29lpKIAHhrIEZLOdbgxPD+7ZWEagPVbTtJCBFMjvwUzhFFwiHVgozOUOfKV1nVY5J/XIVfSSv
SdrDjcaPlV4RbKWkoA9C1xmxJ/SqU2yKk9KteJ4cvaLP/KqMkLFBK5fn9ichjLGmQj4OE8ON9AuC
0NNh9m/A73UpK7jR+iNgTaf6EzHHRHuDkplfwFT4zTz+ojSaaIlL/XvrEvBl7t4lQad8apyIcV1D
jgyDb0LcjOux56RFrENWk7ggosdZZXyvKjEMjt5X89JzXeCQLtSACl2WbBiJePwvsYOSMzaz4crq
coHIvZt/wQ3lWJQCCgdlAd6ynxtv5C6yY7p/pf84bJIekysZa1E46GSpgaLtFDwhHHmDs60vmoWg
iETouBK4VLEvO0jLlFy7ll2fI3wrMO7q/wbvkUKVWIsxBsD0I8EQZ8wrbVYv42Z4SXnfExtzHRWd
ubyqhBnq4KweTFX15pLwqDSb2gL4Xud/XIKHMhLAyslB6cKExHd/vsU+WLOb1w1x5qJNHSLBbdUF
8GUOGXLhsJf7VWQQyG3bUC7CXLP4cErKXKPUcm7ALgRS/SmZrvDxyhm1nrWW4wN5DDEd0QPOa+pi
glBlShUa4FPEF9dL7G29QWk1AJ2yjLep6FLiF4bTni0dMbw86PCCDx3wulqV6lAQ1z8LK8JWPH4q
q2zqVhuJH2aAJjg4wjc9kcoB4YUlJRdJdza0HQ0EbAK7q2HmF5rZSiupfAvlFN3w3lunz6RzB8Hm
OAkoZt9zbulNS5f9ZYwtuTu4qHlzi0SsktIpWvaVx3ENjEeiWzd9xDdd/Qoi7hRCy0t9riA+beoa
5p3VFIREc+fZxTPJszG53G7NU0nmaoNeSfHqvd+vIfpiGPYUI1dgt464eKpm9LhlpEtECG0X1L6t
e/Kcs9cKsut8t17AMHs8TgDHC8ND2jLiuHQEaQKf9xiSATu9bJWwMtKBjN6flTw0kl/CTtG8YXpx
uM8lPzqYUqz0tTcjRU3j+G1ER5hZkhXIPxZpcY3yYL900ETL73CXwkS3Hvs10sHxNGCgw/pD2NdI
ikSd29/GtyooH6n2/d4Uvxnb5HTru06QDaIUt4YO6GnqIY49Q6BimenStGnyVHUmhFA75vRkSDaw
kDcvxtyntHKEOqKBCgAGB/zBdG99fej97KotPaLcFa41Ofmte6m9dm45iyFpf7fO/9/+e0NdTuYk
murcCF82BXAtJ2wW90tMwp5kvJcMWt15sZQ6duynreWdvuNFAWK2bBQrHGeawZvHYGvzkWhA/lOa
gWyu8C6nVGYXlXOGYPCuG9Fewb5sNosv4MTEHQVwFvLrCa5cZBR4kU0xUm5aX4s/MJeErop0eEAx
S7SrihWkm5eMbseZHx8ZW2BqmDxEdzRXENpyIq12CffcKXHPKyAXUdotHwzpha425emRbeV5mLwt
jEO/4qtsu90pZvXUT94Y4DI4Z5TAtGnUu2l6KYQuT7gI+DpniEP1Q9AYZXFGBPuaulErTK2l/BT4
NluK8IN03avihEu+9zRrn3n6T8fNQvO43vtbLS/R1eX1/nLdZlY7C/+X8uyWqXp+L+YVxLid1rX8
0huvGNN77eAR+BuwE6uyOIn0BI0Mz0Hl3bJwWy8hVMj+l+6dcHtXbDLhfxxW1KWd9j5a/7nDBWU1
P46oKwbEnulaM4nl3iYNuHKjbkYOZDvS5wnCNsWuA7zQdfqrf4zl0dCh6PyhoW+UETjhx6tF0Xn1
9Q2KWFG7HoloBxDRwGkpIvBZRciXwcwCE9LZQz6o3cx0ELHe8peca4VIghYnfRHaBeHQY3aauIcy
lwohNhFr8yNFGgrFtZpmqgn07ISPweJ5lqJ95BY8hjfAe9GKaWU3Z39XpUAOGPQfBcc4UgXJhahb
OHk9OAc/urZ7OO64ZpysIIL1d6SvPOd81qi5+w+o0eJx/8K6mhuQiuR9W/LVlJjuub4JOpj2f5B1
PmDMDXuCxNMfy1FQC+4QwAKgB+8OClEVWljLkheJhb6u74tlZ2ZO1K/gyktbzQU76R2S1hUKemVQ
RAEi1m7D+N3Yd1wQINV3gYq7LdeLoroxXYuEQHcDAbvkDxoXV/b7LK6M38ONRrmOBBooJbUJrTb6
EI+MWDu7RfTZ4khgkayi4KafWfVetvBWlVnxe+QiQdI4NXPh+13ckkIvDuJSQP0avA1xmnmd4zJu
Tpm6Iv9SktLZ1eIfCwSrPp1BXTdbpILxXFBCjGJOJTzNvjfNAYOQPxSoJ8+8D/eNjmiRYUrweNhA
BJcNyDRUQWcg1zgtHxvTf4Kbz0vqWQ3xrv03ZvJUpidaYy41ITQBnETczP1uVMn45dY1T0EAREmV
59qau3u+5KbOPI3KA1BFVb1jNO16DRQgpjry4lX1DgKnTdNq/QworgRFdAm0MoTyzPZguxo0HqXG
ybdbWoujT3NUqflmM1XNq2HeJ66kezQjzUpPeSoo10rJ9gv2tfNjnI06ywB0ZAHHEiAxwvbio2ib
dw1iAtPyuRjxokknYesFfu/lRLM5wTCAUtCXUQLNxljmAqlyi1KFvsxRgxkOftYEGIl5BQDj8vjp
ApE7EMMD7i42tdPvMWFadWCqKjbFkR7gPQShavz1gzvzgLBtwQPtyvmfpRHpbEyZBiDlG9sZu0Ia
Zhq1R9wzkc6JGU4G/9cjCOGOS5hE35QomMPXxR4JpFvB1m7jF4dsxd8xL71OLcStk3fz7cNKm0NS
sI1l0D9ahNN5pVG+dexBwHK5GW3UCGYmMSuaRF5XLmD2Kyfm+qMtssw0U6udkyJEo7yj+056wwiA
JES6YUQG9s50shqGyoKoxHRb/hDBVdYtGAtWfihjisRyqLy7Xn0AjO/T0Nnbrt06WrJO/DDKGeCm
hVD7z6xiZx8oqSrx1Z4rwzPws8Wo1DwjSeSAZ9Uwr/AUgzYd+PS8AU9qFmZ8lnWuyth8axBjNHpT
s/qWTnNOgtogSrg4MtoYQL9/c9/hX7Xb9r+8O7WS/er7IVXE9ccyUUaOvA4Yh1hotinxqne1nIv9
yw2aJNJuNND6Jl9CtY9QR2duRJs7MWr5gBooQXs6WIaEe7j5v7nahwzKCrsdV18SA78gO62EAzZO
X2MCIVeu1QnMljbM5vzzbdZFk5IBI2puIzXzznCzYiYpWPuWgNvXcEmeKxAC2hVggku7N2DuYU+C
4nsSfxLUj7Fri6HDtldPXkFd6uzpf1g8lc6yiDRPllMoewAnfxK+v8U2EYJe2nc+prf7xNuUeZNm
GYAgpMUB0Da29eyaGA28h+R86BWWSUqM0canb0A005bgGQSZsIgJeR+UWz4+FZPtEWXDo91nxaoC
OQRJ96njdTjPi+VCabiQLf6HY1u+d3p+QuLoMTWJ35Zx3KRJCQZzlJuTOUECQH7UMmUlTj2hvb4j
KikL/A5nXhy0lU753jr6TkLk/nquVIhZ2n5bI1Bm4wD6lxqDl82GfmBckrMoeE4ifpzl2z7BqUV7
GzyRJJQslkniJlAO93hZUxwQyXQr3+Qn+r0QFwZkvCoUl83C0DIeJxciPbbmbbStkF9uFcmr4ijI
vQaL2T9Z4f1kJT+zwrWwSo3Fs/SA14QoWF7mj/M8P787FOXvZLgr4jnCH9nQXnb+nAMIPNz3Jqvm
FuBP1ws/giupPJUAjAW4UfqYLTlYjOy9buooC0A7VatRv6JkwENpIOhbfLnnAMVShxPjeeLlld4E
f699+6vkD9PxQ800n8F5WGDUJhrGaglmHRgIKGKp8G06sIXx5h//GCZEIpvx1gpDkoBWDHbEVjl3
TwIX8lBBbOww5vahOeKSvgxc+bh7Egn/BpfJx08CJigfiL77+tUeJph0F+GhCT2byTTaY/6FTnwn
nvUFU3qnc+r55tZtuHrmFxfN6wmwQJm+AuK4TidxcoP72b4J9M+Ogqi+P+l6lbCg7aw75XXLnmE1
cCuJLaQvbe1hvMMg+xzVQMcPXGtVOp9RuHYqU71N+xGNCKEa7MrFEqquUqVYMHdsncGExR+d8gYj
ZaWZXAEL7I9WtC3HfV+7rLQS5e1yBHblMjlqib920YQFOnYXuQ14anDqB9C5O5vSPEB6950+Z4Y3
LrR4Us5Szy8md1lLHAgJDMYbzafaD2XPWUusoBOYJAzhyf/pNwNLNH9JSnwIWZrL/g0szLh+pL7B
Ak5lgMORQYUDuE4h/Rg56slgo6RiEcdg+SB0fYSe4RXzYy1riJzUc1xjd8A+UyP/lDdDzj2XnZ9v
oKXS3ek+UUMVEZE0IRl8m+i+n61X0RVLVMaGIPOFPSjay4EfmhXVX30AAZQvN7VwFWCnPIB8SAeS
Ttwuk+I9polQsvxAq9V54xsW8XCPxIff9PZGU+hc2f2qpgJvqY1qWMq+akf6roE5By+C/Latz0vu
paobcrBp48ARHA/KyY9o4WV5H7y2LuIT4fMEkAncfxAunPZftxHi3T4b/IcDev0ah5v3jrifX2Q9
RRDCtP+WcREl6mSqOH6DRL1YgKt3iDx0OdMqPKaS3ZMj///0ktM7+qHRBOIw9Y58j0CpsPrP63Uw
dpGknbn3UDHKHUw/fKC7OsDCXvLH8DuarO9sEGvTmng4Jtck9RVN5nLe1un646drATY2O362Lkr/
8izA99riZ+t7wVGw59W39xhQzalgrQgte/l09NTa66w7s08D1TspF4Gm8phKU6QgYZaSW+sGbKyW
Dat8Yv2i4E7DwAhrdgHwK7ydikYrnUpjKP7GKoV2H5llWPrWJJiLTxlpwe3/WV06B3zSskgJIPLO
kovUZUUc5oDPZ1HoQAXGAbAUuCu7akYCPoNb9XG7GeCllF1w/fdh0I/uslTLrPF8ty5ILhSasBA+
bDFxXq2r3mABQEU+M5na6ff7rfc/h547JTr147xFrrzAIDBevkgYA7RwXSVRG5UREHhkSkFOa1Bu
V06alD5ZO3PZGAQoLQT2ZWUuShfqfIzKfV0PlcsdWrZBnavPVSYVX0gVzYXATAd/tIS0qQqzkPS5
d94fPK+Tav4W9bGqjUoIGSFQ+MNm4RBqXcwYcjW/CCMKfVXbKoyV6OViTNVQB6ZZv2qyp5jIRTjB
XGzjGWDFkEKdVmqEvk08ic3d514+JiOQl4VrxLKZxWTN5s/PpAO474ESEznJW77Vs3d3e40AnrQH
VR3ZX1XqjzXFfqfdeo/nqy26SaMz8tvO/6G49aRzqzo18ortwrf3U9jZXusmUoM3Gu8XvZQB24in
oTjd54dXcnSblEJ2IzLqcBsTzRla9hKreeJDb9ItEMhUmbtVCWsifHNiY6rsRe8JLTu7bLQ/Qifd
q6TVDnB+BPLx6y7Qcwvcb2/Qrfqx8vx3J8RIHlmuY3MgmIBRnW84lKppMXty9IwjKgMPA4ZIRMTd
v1+H2vPFvRQLNeGuhusrQxkEOU1hiUgEyRgLMx1/sxaDZRfOf3cuwAddoMGCzzzEq40aCM8xi6qP
d/Q03T6m/tFuOOv0U6iyjmkjPp823TUq2U5ysdiktDx89DN2aWb7xycKS3uvzisWZCRswcAeYiHg
kQUK0prislXnexE0gabvo+mTwO0woIghqbE0Md5b4P0MXDjfxAgvqo5viK2QPLiEk51g9+8T+mGf
WV8QL0NHt1EEzgDHx7ogOxNq94epypIMqEaE5+Mz7gt6Hbwc4ak5NO0iJyK0o3dTrZnV6IPAlEyb
mIa9doWCpCzTeDj8TBpD63AExo/2rhx/uST6rmqGf9tV5ECOYtJ65hpAksm2jM+tmqciaoQ47iV1
DoaOwjUG9uf+UxkdmYuGkxnguvH7gV+q+aiMsgOQ2h6nopsD9sJiPJvpBpQzXXMHoFWu4tRik1IV
6XW7NmchQein/94b4FZNAAOlpiB5fkfnNxcBNhJpoLOAinyAJvBCDJoy9H1EhAinrlNwNpPnlZsh
hM4VIw0LfgpyfjG+rLbOjVXy54qI9wBDafk5sjQEXL+WTpvo9Y3QFWMTWB3jv5fgTBVyPXg/wj7z
dqpx0A5AzvT1Xp6OLoVGOlCNepEsbIXYy9GzhXRrWJzwSytqLsfu2su/81JaXE5dGrd8iCGAMFiV
DeVEcXm2j43WzuhQCsUqnyP8zvup7l0gJloOFvrVWhTowN+Z3snUxA6HdiTQ6gkAD2Du0NlUjaxU
g58+hyHfGgDCsZXCXe7YdgNUN3OfAcLCT29QaKXGoEqlAJ/aWDHGm0eH7xxUzOrrnnKHYKZwjMss
Yw8ieo8J2cNxIAxSmZJGe3ITGjFmCwvaEhIMXfxDsHn9ibolCi5F4zORkNjfojQf3Fs8aYZCFnDQ
RvEOe5v6+LQrggyGJpm1sqtmX+OIuxwPcwC+DuoQq0MW8sjf1OmQD1hvMoe02Yuz5CtfIqHqlSAR
9IFt1NrVnDDXE/c02A1sXqOJmPCb3WqqGmP8+CBp2+WIAD5O2y/YM+ixanlbZyvF9VxIiu9z5InP
j3DIjDRSMUvkIs8qftwBZn8Wk7xQZXJuvd6+pjh9uVdJ+M9IJqtp20fbaTfdZcbOc9nYHu0qJGP8
HZ4YAYWQnwUevCgCW4h4H49n8WjSZ7GMGvEogc0uyzXjmVtT6SULJpdYMSDX+vm/E3CsRTLYicA/
K1DCafgcnyKLbhpwqvSLZK+ZJzEFPhTM00o5zRO36eDKIxNfUEpdYShnfPb/kkQIYNE6rIKGHSKt
KiwsOoHQWP8CC9fFSB55x+6Tk1/KnoyxDzyzmIharkF1njyAaf5Y4kc+qbuMuFxx1ECPU7Y1FbcU
wvze8c17zLZhQ8/bYLZX5RGeV+b3dyTxby4QGZLnUgUY+xBUUt5sn03AJVENDZY6eFL+p049wgqs
odX03E2hYPY3slfq/K0GsBLOWdFPrIOAbaL7ZDpeZ4z9TBqn0S+dZ/poRD95COBNao9YyQaE8yem
NfBv1P+T7ThJDwWOo+gzgDpnYS1lhRgd4ALBtnImv5ya1aGN/vmsJAVlpbAUK6HBt1q0QAzUMoJl
h49dxsNRcoHp6J9CzVoFmvp6tlqyKY1/Q3PzRyqVF6j3DNMoVwOa+kET6+vfrWrTX5HJRqXzf1PQ
RLy5Capz662haO66OL5UupGilRlkNAgz766BUGeGcNDAyRX7LzjQUlJDMBjGCxgmgLSfILU034g5
irkPxQxSvSC4jfmulk8HoczkDkInxdRpNSQMZniXqmXilD33243BVv57MMTdq1CsPFBMABll9Q/n
aMWuHCCaNeAW/6t9wkA4qLl+KrcYWy+0JQcm+AQDMRBU/+pen1JX3vTdQhKeDmo9UC4bWObP5/Rg
/AR3/VpNoNvG13A5CflAI1LzvBM+F8+ewbIT/jjmedvOvpfdiFSzzbFiCYyyG55OTBiWPBBy2zxg
TRXw+zm6VYeaWgFpvXaEiZGz6jVpKE4xM0yU1I3lLm34Dzr3sSFNkxscpnCXClqdpX675XDeESX+
rfLIlNEA38bS+BbrLzyAiJTOrelzTAOClwx8Hsch6rka79GH97cqYm58fs+Rghom5Mke5kk42hSf
COfHLbWL82G4utM1TbqtmIY6zuO7jokypv32UfsozS8REKExWqn+JOjealnU0vb35xyeTXqs7yTK
a2T7s4iOzq8OXrw2thEqDRLsMpBBVhP39fHUBDkFbdcBztXvyH8YYGjLgj7zpQjCvkAKWDV7qt9K
HrgLS50W+q1zUIOgxYzprPuVzsNAGz98qfKaM5Wy4USsUDulB+CnCxLeh7A8OuEQllX2Kd0AduG7
3LQ1G/kObp0b66it5XZJV3mFZ1OY5PVx0nPE60rjQMOORooVPAZnpJHc2eymvMWO8owTOYcy6U7e
E3czRFzJM5J+FuzdO3PCwHRCuADT8MLVfmC9aQ2Dvg9a7WDuvb9ynbOqVRYUEck0Hk4A72l5HN01
VJd/6DCXiN6PPT6+nAXUy1+1SR+t/VhURlyC+JIcG/EvPo7rdKd+gM+6AM6xPOHLiwRYDJPVqjeN
d4mpKHvRsNKr+GDUrOhNxNOD9Xu3nzSMO1d6/ORHocWPnC+S+p5qUoAKGVCcKvJJHeV1zliAesTk
//GT2bUqU8B7jLDPd9VUnBnGvmnoYAPMHE2SVvRZPRFwxT9UlbsdBELeuKb17DTW4OfvJtD8a8Zs
qmntkbOyOqTJyIitc2ghxtJojowJqDNGm+d2OL2iwtUdf/ETFxAhL3d2A1pYcTPQPMAGQmOIl3RO
BFfuVvkA41TzZUkXaBcQXbax1Z33HhMJBJBs3BE7VY62jcoiDIxZOMODA6b/QCDkK5Tnbq4kJt1i
mp3FznoGLO3r+S59ZqB0DcQukdHkk2ZsPIdGfiQlHhtqfdocYAvL/9z/413hJsme3Ks6+zXcIh1Q
TsPIJlq4436fpFWYj/HLLqiG3QqPrqbHPRuSaXhKXc+AmsYM2QEI8kmUGyhYBo0is6oZ64XMQws+
YP2DrH9BD9RlsoPabxt7QisVwN800Bw8rbpFvdHEyjcjNPP3wLZ/bVbnONjGIqUSLdCrAOZvgfUK
4hRBTiKobzwQwuN23RpASZJsGVrA+nDE2+DFHdTvkTNzUor8mljcyrAyAOJm+xS9p5OuALihUtB7
hIv6XqMMm6XijcWYp2OwFpzISGA/WPDiHSlsBHODzbfnMWInTcxoCzNYGmXG0al7aeYtRwwXKnXR
vPktanhy6SQPyyHEJD5K3q5skyjsnj4a4PycUX0imTSWBUi3TiWP72Xd8rXwoKoyfwOJmciEu2Lm
mq+sTJ6pbjaduRxrFgEm/2QMf/VEft61HbLPYnQEEzg6RWXaQnx5tQKcXrWLLL2tUvhSHJYX+7mO
Nq8dWX/jCFFhkPEOoiAcE+LA9n4+pxUpyWedUosym4TKPfAfeL9wWvET6cOZZyk4Jz4IZBZFt2gk
cS9wy8A9gdoCEUuTDBrLNlb977l8CqHWKaK4RifrrtlCgjV2CeUwmddlWqOMc0oIlxQV/No/RFLe
290sk7A4DJ340K2vsA4idgXqQKcr0WgKrQ5oLVfnv7FzJLxiWRf+WgbTXqYtfd2NDVjfOgunoTNp
YVnofyBykD1CUoHgwQLMrzo0K+3QFZJA60STcX8POr9pJZ47m69iaIwbMn0l2eaGSE73Ipf5BgfS
podX5uCoaD67v5/caIlniMM2ErY5Dk8o9lDpAbw/st9sLz/vuEQhqsIfFJNcpCWff+4sWr7d8waO
OZO9pZvM/hK8NYm0GYbkpWZq6/wX5ON7RWWk9G6nqzGYeBb84UMnItwcQNI7cDiWuLh5vrmnArij
7ItLoxeT5hqL8jgJ6zcVCNXuztG5SxHeS1vLGGmhJCluIDT8XsanHm2sQSW+98XaPZ7qsgumup7+
5D/VeOKrRXJxX3ej9V2Obz4WjmPPguP+qxoE0GAWO5TK4qlf8xKjvUL8rc/Oggv6VghLyw3jle43
VEypiwuY8OPJ/lLWevXqzo9lj0Ua8aASBuJqeaNVVG7iPGtTSaisX6lMUo5FLecU5iQ6hWF8JRfH
DTr6Cj/3kGQsaobKrdDf6SuFzFyx4yH2dsKZVVOboZDD7bRkBkiJtxDhaATQwmhN98VHnGj83jUf
aQ1OKZ2I0R3xy5erIqQWPSFo6IrWd/KEFpiyjYSO08p10nez6C6whubowmbwg4IuPiGGvBa31P9W
y5wTQEC49cCrzpeIAGdX63/Iiw4Hw9gkJ0bisvV/87gS4G3dI+WagNqjOSKmXQvtVdcYQRyCAmBA
QTd2tXwKIO9a24BNXUbAFZ8HPinuLmOaJbEvhvX5P4FwrNAMbPMpfEDEWJuhWXmP8vt31p1xlDVe
/X0MgrU8Ln74DnHU0IiF04wXqOAJBABnvwf1qrMEoCqvHjZONqVa1QPdy99eCjv57ryBeM1EsjSq
I+sXn2XXvqGGKU/RCTWhkjQP5mrbBOqjC/lCiN/RWd+bCbaUOFz1j2Rhd2pdPgTSF4sa6/zgLCLk
5+tGauTqkn5zy3FoXbNAos2NkdAu+ovqrv1iabGAPSb66t9FSA9t3SOJXAud1RW+PZTKtfDhuGCY
2xnLveM8Dv2uop0GL736FRqSMbeK/tvwbu3jShX+m4+sJx5zqxULSE1qSVZ2MrE2WOQ7LFHU3Z4/
Inb5aW5BWB7XgAmlSvfdYUufdbUuZymopC2yo+LWo8y1tB1NNFVz9qkcwZMYAwLqqm1RSzazaxZO
Irp1sIifpzcdTSqqXh65OqWPXnmb7ex3ZHkWVTgpiPLmHTUcp9z0OvKDi9820f0Qlyba6LSr7HXf
W1pSl2YikcqDi9uUpwWDCL7vuBiCSA+3heksp8tnCMpAj3HOklm57vdlXfK5ZrR3i4Qa4CuS2ozf
hXttRfc/6db2RzgBXrV6GHlLiAtSV2fJOTUALVeKIpz0TnjZT3wCg5poJgOSxp6OyGbDQxeiFVHm
orxFGX8G2suma1rqTgP3BcPq6YaOyZEfrEJ+F6/AACu3zRkIshg7PqbKIQnMNLDI5zyubiQLkdDu
MopfgYwIp3sNVuhA5uh3zX2wfcfdwva46yUNjbjBxkj7q4eNqJanwFl9cCuz5+nOVu6O8tzbQ+AZ
hKV5KPXcapPv7Kk0x82yU3HZotNGyJH605oH1OK1AnKAgh7vFM/rxPJ0NfOs+711hptNN1W61bJP
uxlT5L4OQg8kpTugH+mdSdxWiy7/WhQR6majO+P0Vcvw/svwITRtv8qdFQeGyd2mDS1Kgjyg5fqO
3DkdXRrXS1RGoO3pGswz3R4Tz63CgtwEv+NHE7Xb0DimvwhhQjc7oknobZbyxyRDStl8gWPdTpw+
/rOg2yeyNv3pGbMpWzoaTNBBAQXdCphIgBtRIc+kHbwbkqqtCEg3Ks4xxX0tJeGad/xLFfaZFwqe
XsrT66gF/QIkg715+LQRYdn/b2fsK4Z9C9X7MLKytoR48iGN1q+sW9ufob1wsk6C8iw9xSkT6RAU
R8u0WuGzJ+PJYkJWR4kJUP3XCHdKChDHFJcC3uvhYmw/bFfk24shErCydKHuNGEc6gkcE6HyutDO
rnf/SbBB4xkdsMLc6MHAR2IPG0l6DX7Ltt7VpGTkqU1fo9x4LgPJ76NVVFUPOWKx9VzCBgWJWqRj
eulWB9ub9JkXUVW0qtRlPDLB/P1of+01pCc5d5lmVh9aSOTnQvcAfXMsaDcccGSQfz4c52lUS41t
qtnsovMns4X+2Iy5SsLoYFts/JhA8fcgxiDu9Y7eODfJoAwxTPd75zLGXy2dXfS4uZVyO13+NJ7P
lfRySYyrKJQWBcgcvgdIiC2ruON8qu9CSjETCa+8gJoucDqfgJ7AUI2vwQYs8C9ZUOm5XVs1wh7D
w7mHQCXxjGIPHwXm1jj3dFHRbuUAe4WfUzb1romAoEQ61u9qgvO2cKKE7imR//+Ufc/tfyggIPoi
VK+SchDkLXR9r0Gjl2Rs2Kq97aESGT0RkFw451pGO10sadp+7mso0Y/t3/Gf237/V9T5iQFYcKwu
RjrRfaXJvH2CV9DomZqBP1tqfOXn9C3hsABZAEto1NW5VRKQ8ajHO52ipv9ocVTDR6cO0cULHUI2
onUjHlI/9nDo/1juXwJbLIFOAQYMhk7+4P14vjr2HObwhktKl8WF3E4SY+ORN4KthrvV5vL1udzD
NDhqKMneinI4mYyd6j4dC8q7rCj/ftp4VuE2HbjDklvI48veWDDQn4EROD5pSLQnFksJc9ROPhF9
kNOzOY0MJVIPg+Er1ZKuNw0yRjj3u8wnDbGO+O4Vn2c7ELnZKlArxfLZCUCdhvWLb+PgKgjjmGwe
uG09Q3q0J+lHulyCrE2Chavkz8HfdxzVdw/euqQjQSBOHee09iBQYUlvtX/zdZnF7hqMLYPEdezk
M0DAjyIZ86k/KS3pB2HOokhjWnzgDZSdAagbaEs8e9g4TPkL6o2jyv5hlC8OzRkVf7IPzcFyGrWR
3RRuwywsZmeLTQy4RY81qSS+dWPCelLmoQqdL1PrntZym7GWtx1q+3rwZUqm+pFGeWUjuqCC4UbO
Ew6nApdpQZOO8cIhPxDlayzEOz1jwV6OnQCE+Nv+VkXIvKLNd94KRIWk8aOkHXZrxkiCdz81PUWN
FlRDWuENG++kcp3yVTNFNoR3XJ+mUlmeSvayITeq9wWG8gHpXOkGOz9F3l38QXBSyJLwdfRJx0i8
KIdwfCffhgmS1hfkR247x9zRDzivCBZMAcWksO8pai3AhvJNFOcXEeAWvUznOIijMi55hu3yHz6B
yAeDsDtdUuGlq4ROOez7ii/oRxUy87uxNiFawGNo2hMUOI+sz3SkFs9k3jeRGAacvMQ3wtv63DF1
KPZ6XKd6iYKce/m+vWZgJL4jDotmHOQXL05d2twJRYwL1AgOVzOC4U4pHWJw+PX1FEmXpZBcvot5
EyfseOba6EFPfIrV/V42BBzkopTOHa/l5hyYtYDzPjQusa6yOmD07L0I2IigmjkEpLQ0IK7q7Tug
RfP/yAzjqg/vV0enYjGe98n1nhUKqrMGpqo5dSghoP9XLYau7YMGfxRn03+zrsDSGXhZeWtaieyu
TndPWyOsu9qGSce0IyAA200XLQojZ2HnHS1r1vmHqE5X+mHGNBfHWcE3ZtHVAr4QSWyHqbNQm39k
sUyK3u7p+67emGlg1H7El1ZRj+/bw+RWw+9JZBKyBSz550DV2MlXtdEJKGJeSuW3oQpQ8QwSWOnn
hHwcGBmYi1x1vSqZEfxVEs7uyg5iw9hpynrENZacjGpt1+umTsngPGU6EWzD1EfPqrSfJtCf58M+
diY203nwzZFESith+ISYF/VfWiE4PgP98trf8VvZbEf7rPDfLLarU1rZsOKlIqu8NlM3dQifQ2mG
OqOXtx/8ZChND1uEUpxPPiSiYE7Sckhb/HEnyYqDecIDyfhu2JaT7MNrmWb9tQNoeE2QvrycZvIW
btLeJ5VV57PClcBb/LP+NE7vVdPCIXmt9OMm/MpRPkQluxtMS3ACvxsI2dlBQ5zJmVgOum8YtxWj
ZGUSR1Tm2B/4pm3Mn8dH+GYT0eu1/OJtGPI0Xuol4h8VbmdoZmRkiU5KKCZUZZ3J24V+QD3AcKqg
xIHPmQFI4exaXnnuLh3MoHbllS7FLeadZJ0G98YGpgCAq8le0o5QwKh9q8d5UPGZarODbkhIr3e6
2CSpeo6mHCYKNNPpRw3mTHHzKrhxB/tpoIajvGnamTxPsHFxL18W3CxypyuH9vNDGoYhuFYrcvnh
CbF6p2L34BxCJiMFWAF233rli0UnlmYLrA1cg7O5YQ4u6myybkf/J9G8cRaUPaRK1Z/1pqIwZZG8
OMkmpeWjsm5ezANiyyo9Y7y8ZnY9y7Ln9hkpfcM1tDas4tEMBfJrLpBj0fSlNTdv22NnkHo1A8cf
C4rbAF50Mu+Pt1aNbE532JqXXMKhLlD0vHLYst6sfIQ+W1lOedWiPdD3DN7L++EKyD7P+Qq8GdpK
79XoIoDVUOZrj1+yhxUgLHh9DVvmq06eoCJvNMNsNvlhxfY2jAmCS06vrofZM86xVB0wSm88TbYL
Yj3oRjrkKHocFWcQ99DFJpWWHwjVDhBqpvk+hwEWG3lmykFHAUCC+2Urp0gkC+49AeBfu62mDiwj
fUbjCad05W3NzDd49Z9j3xmFCmwUbyElEX6O6BwK8T211ZC8dx3yag9yukM1hqQI9dGYwQJu8JVc
wGcQ8FNiCu6WU60Mq8xk7MjIsnBNTA7uLGrp8J4QiSpRWxCg1Z/VBequbk5gvDARlfTS95uPZU9u
EwKRizVGYNruuiF/IbYcfYLn/pPiIL4QZN1MRNDptUkVhCxROZIGmxoVFoR6pswpjoDYQTTs/7D5
aP+w8PqOLaJj+hvXE/FLmHbi7e2ZRLzHrHhr+7ZvWsip2pfDhu7xgavOIoZnikY7FSCaBTU+b2oX
gEVLpskZU9/aR9x1BCVWMkAFVQFPsruMCS3L7UcnN/dQVlJfXPhCL1/nVUQYPDMIqW637KxKzy8V
QfyZ1OocdF91GrrX4Rc+5DPFpP10S7x2YU01db+4myz7/8dXDBBKMSwuGCEKSJcl9HIRjit/wDAr
pazmnV8/lUz0L9rCRpLwcPhZ4mvvOgdLoZEMHJ5F8ON9aWptGAq0IuiyQrwOgv6FQtnajcR9Au6r
MFAs1wmNPaitIKqKvCaBf3bi4P+oDnq9ATaXChW8P14G6sNfNTfNXrI3i15ypeuAbiwj6r3Xl8K/
toEmTQsS9YUNmOJl1dlLIKZgRdP6Np7P128ptCwFqJOlWUE7j/otFtkCgGiOHd7ITJo6pY6GzH9h
A1DbM1mBTjAKRDNOUKihWyW7MI20uYAk/bAVXpqjme99ivvKtDXJm4iVjAtvhbXOp9gRejFg4Qxf
RM5lSKVGwchVl1OiZGiWaOViOcUH09Q+g7B6LM8wf7BtsrJSFd3dx/4Og+zCpFYCkgVNDmTCN0l/
qLIqV1aTBe21e6nnm1vLr+yMiEyFxl+YiYmkBZ+xxMVhsq3b9esaHYDMUdDJJxB9Z3yI8VrMwCMB
4eR1bFDhMOrsB/aTfvHFCChCdB42pauLWHhq5MurcDshRoha5LnZjx2D2j2p+c/jTl/u9vd48bQj
2TqmRuYYYnLY3vqm1H/Z+nn60UQahdM9DgbdlPTYEs3ylLuRucj/uAzoAZQiwKNezAG1d2suZ6xi
JUhImLmCQiIc3Z6KUgG8f1jL/DbppyNe/VGjx5F7BAZxS+PPgVEDGcpDG4whdSKO+biko37XZcQC
mqbCbGKcKmAXY3BazpoRpoGmEen0Bdfni2P+3YpS6AIzJazmmNg89E88XjBPxFlKdym/Gz43/hIj
LpLXO0C+x/NNAnwraIjtomSN99081Hh9L0JSkA/EDM9+xtW6Rl1BeLkcdLGRAe0x3VYKTG7pH041
CLI9l114mTDMFxOQh17Nv2QAv2dbelHDvkdpBJMzDX9qCsXm7pUELjHvQ4BbbcfY7yRxsHm2/HLe
0bDKaq5RLkPiThsB/5+zRiYmoo14xZuwSqb/oxCwfj7Ny3i9y5lAjtBZDtvMsoFg97h6HFK+KKMw
KID7j27FbczmStE0iJXpxnzp0eZ2xI52hLApQo1tRbdR8JUzlilEBxLMcDpN8ILFxe28r1Y3qsP/
JXeiFoyVq4RqzRJz3BI82w6lWAWQ3jK4OrZ34+qD8/Y++hJstr1E5kFDX2bv6nTIEzScPdxVWPwZ
K/Wv0zoQZnNq1exGE1TQH2ZnBQkP8ar8+0AX88BrPy7twkgduCYaFfkJfO4ddd4oObn3JnRQM7Gz
rwrwvJWPAQuRkO0uz7o7nPnTo9a5yGnp3XSFEt2YmNnDtskvZHpqcbY+HaW98OUmW55UnHD+uSOh
/+aitSbL5tRf5QfNir0i/lZLaM2FVaY9WYaAjR2Zk5pzLZ9NZpPdKCWO/6Q67qfOfjcqX2jrcobQ
Vexs4VsCK1IQLj9Hw41lpo4poOhRNIaUGYe58WEu+zrCEcNksLALXLaKpekvbSujPzZqvXU25l/E
BAoxc3ffCdM3ds5YBcKCgHbx+TS9+kpsuhGQku/LC74AhNSK/b2hvREb0Fb5nMSitR0Ru8qpJUvn
dmzx6J6bqK0e/mjF+Mxy140QlMPuGtibzt7PyBSpLjcUfXjKCAkV5BgDHrl2x/lrFj64oBlkldQC
AeD6TF6AUPDOm5HOXRPsjMoswV5ax1dMfaHp6avolKfhy6lNXogVb0m36r5ngnVsvbet7wSuC+rP
2ifgCfldrHg1W9tHM4mWyDvsqO5GoG4msvYXAJPG8EWGHpwx1qdhCSG/ozxp4AQ8gwld92VD6Ui6
ABTWPr/39dUupPc0dxubN6trplXL64N0ww2RMnaIuBl8I2tDxSBemQVGrea9nuTZACB3kJ+eamPE
epA8xRLPElj30eNr/9uLcfrYPzY+0gxZFFmpM/qgFZTwtTFZxmPzcU0NZSa7iZ8dKwHAyCHmv0oO
f2usyOMMmPIyDDWiydx8JKLFPVIY6MqTA57bCZuvdvVNNmAPO1L3qrLjZG52K+PpJT+8Ed5OOpMd
HQGVMis7EfCzsdI/7/6xjq9gUTP2IfnsZFY1Mqx6u/QnsjmozCZo6l/uKrrh4oZ2dFiYXWlu8vsD
rDGARBOXNL/9t0UGJl33peup5WQn2GzqQb4PGGeCVQnQ2aEJRIjGrJFUt88utf/3EvnSAqoZEZ7R
nvReY9sz5BgQHWQSfHKC+zqtZLfdRH0RrwH4+GJDRhxJIaOnydjPBJuo+a1OsrB9gnL3MtIf4JRD
6vcaYAhO2YkYTtzll+rmXaD2OXwp1nUoATgsrruESHtNNAWMjKzawxwLPemVKLeaZpaxExnD8lpI
PHECWZfN/FGXKcDgd4+WD0XoJZcTj1/Dk1jTDTROwpLzq8lVfz+4KaLvC3GhoqRB/C7Elu5+Fwgm
A469Kvr7rx1eFGUdMUk60D/5bCmyPVGiFuXUY14CeeHow94by6385BMExalioJZF30TtSQgF4mVt
VNDGaIQlabjlas95V1+gK4fUfl3cxgAvFWINhG2Yj1KXRnjk+SVLBzmpliMXKpnuqVO/iPek5b1N
hVdVA+diJfT8+Y013J2wijnKa4Geouza6tHFbHpfid8ul83VEVnR74aRrlodJvFEhawCZYImqFNO
oU/7JiJ9eGB2Uop3/luq5xnQgsgc5fNVoR5f1vUWLysxyHc7kGniyjd65csccviLZTc1H1Mn7MMp
M1leETi/Oe5SUqocfdf0aWE7c3m9FdyBt/ZbkDVPX06YywzfBsdtGP+1fWr8L2vFoOI8utu1IrpR
5OToAWvTnS7L8awUko9HzAm8L8ujlqwYa4m7hyeMJoieAimfLlBgDZIV+umrIVdjNRVXFFecgZh0
+Rscf1MtYsA9OlmHJA/zQDgjT+kXxL/ellpuWSV781f98qPQ4CgSX4BzDUNpdxyry17CJbaKq2Tf
PgFHpCaRrrUOD58xILTSeznVsxs9oMLMrj9PJDsyZWZD15bcZ0Jj7Z2b15XS6mvHujY5ZqmN+6su
rHtV70QLOiHfkeeiG1c5okW52n99YosDeo25TfDgUlmXKePRqBOJQ8ZOmDqEh5jdn2DpLQno2otL
riom5HhuclfSGCDe8EQpgn0BTCB6Sy83QZfNnoNvNCAclT3Z2by6DCxNfNdmDLICsH25tuwMhHEr
74b3eYSSP9rAv8Vc9m84AUw/gQPldOc+mluJgqoMQopEuohkcaAH0EHrEB7ZtIvRLQJe4aN1gqXD
QLcq/dFxcc1Wg9tP1crgXgri9rtQBxm3NaSKxLlw/pdV+0moqThr15oxzVea/Po4GLBLt39uqwpS
yizlL4aCXFTTTGm9W6Y2SofxYJLYdreUmAceyGncSxBkCS5iv3IhHqkxu3ZEzr0/ek54wlHMisO5
ixcE6Fxumz1+LFRKUfzHUrb6Oi7EqlC2LreQqwAUycdvAVtE3ZGVllvzGUOI+X/fsSvinaA8uRAo
UfqN9QmpNWm3P/OiHM7YtNq3jeKMIHxTXr/nQNlpmBuJwQKF6y3X3wXjIA76sPmgMUZz4wsVXuQE
VIGeG6o6xIPa+qE163CZW85oW6ammcOSE+X/GO7hPqJT2g1ytB68ZNkn8OvEzq3LbwpcUSO3/yU9
TH6rspzJSyaLvYJhV7kQPmSajvUnuzHO8J/3oBTiLfKCsLU/CKJLe8M55anPNwyTpALVpZ5pq/Zr
rUfDLNPhVVInmzuTFJrjmvpI3PLLJZJQJ+1lTtIyO3QxVL8UxjdMKyJv+POVSOt21oCnfRdsY1Hw
80Xutx10/K2JcpjmjeemWni6HkMUj4TpUP8sjHMcg0n2z/MWiUlewdRBVDcMZgVU2nS+Y3ag6Jlv
T1KgWYmTup5Zpneanpb4FWmkW0lO768/HZ6ynXNYrrdASw4f6ODKFcbJymydhfwfjGdih2m0cG6j
mqJUR8LHw8Pa9f+d4GQGq+uUQHOItkki1uZTDo3xj05A0/PGUXUO2vIpUT0GZjxUucexm0idCtvr
P8Lr0DAP+7QJbERIXeE7K/snAGCFT7vU/RjAwxTokLe2EXmtJbON5wDuT4HKDVhexM6+9c/z2h4N
tx0+lq1MaaXO4TbNUSDJwe4kp4vhqfbLObi68kLzpEpWVjzqPKDlTkFfQbFvS0qhOAmbEIRmPj0g
nKQD0DrQGAxLpbNB5yI08UVuRrsmEpgXkaXOqilpM3ns6Ov4mmCsw52/2vuj/OzdZdyj47/iNCNp
8QlZmNo9+mMRkT1Ry/FQUKLDvXJ9fEWZ1TbWgYEdgCGhKu4XV8v+V4P+vBCNP4Pp7j9HyeMux9Oz
jYiqkEi4UzGD+6Lb7R1exsSzlfL+tUs54j/rU9sv2f/C5H12WBIYYNNk8KTRa6y1/2yOTH2De4QU
u9QJRn3HxBSyPoVYQLQxxGQY1fkkC6OTOaWG09g0iX9s4ImoxavWurVQolUiM7EKoC8eh0WhKXPy
t+InVdcyJLz/wLYoZ9182PP+Zjf1mWqCyEsGqg2NqoeYnHSQiVkUkrA34uHok9An8EiYuWwDZF0x
rdKhQHjMyjUldGLfV5zSsvcb/T8xsP8ootHWZKM6ENUJA87Wjj0IROo7q1K6Q0VhTyv273Myp9uv
4dvzvYZZR+LveRY5UB+bmptOueUAY49l1J855pkOYXGBOV43pL5byrhFDWhWKcmMm6W6GnwNAUlK
m81ZNwrFSz4JhNaCWKhnFLWfgBTRx3rYFwbbGu3yk+VL2zx69CJkHtNPTDAdYXNU17X9E0ZIcX4L
/m+7o9X5qg+wlXwliKdfD6JrU8HXaDnLeN4HCyEP3rwI6iR0rWbOzUR30KQLLbHp/UnHsXi/QwFy
y614XQh/4VQx0lIWZ9/bebnaOH50IPPKk5DxzAMhorw7u+d5zWTj1FGsqkE7uHEPzAbkbL+iAb+o
kYZ6s67znj3x/MkAfL/Aq59MC4sfP7jEcsWbRgju4X6smVCKCaRhRdILrdnWejCnhtkjIjz9mJhl
0L9O0jqna9WE1voVKSueEbxzvz03CIx86qY3ITFKLApZ+O22k2q1A4AVLGc7C59MsDJKEPngDIvF
myfbwHHGZpZw3INnRAsfn5uUPGY+GfVxEScEPRyXV3rVp2th75FuFW3Y7HIe5RdqgFO6wGBab8aH
08W+w2iztVGEQIOxerStuXtHOfpTCuhUZ3MaBinGGNuhgrugZmmG+FVb0IfFJWUIRVg6PlukRxJI
qGf/jFDFEqe9hBwdYR/tpUaURpxkJW3plJQASjtPjeFyKkfOHVYd1DvYtYCMzC6qJ71hyRovMvqc
hycdOShFFVVubkd9D4uqnIXiC8YI94RX/9BjssZPtnoY3ESf7h/VdkJGVfSqp6zpy0S0XZQxvjZP
/aAMDUYGR9vu7Idj6V/oWdp8TXK3mLKw7/nNxMenxTDxZvlrzTMfiag9E4lGXA6EaKlj3PeZ43/t
nyx72hhOMSx6izGrTZgIvdbukiBO1aIcdMGSbvULgQFl+UXyy0j8o7QPcVWLQdrr013L2W1ubKgA
/einZkRbVa60mDeGyNxA3r72l1XYnWDJ8j99ZGRkgfnhGnpuFG4VR+6BXlsgR/Y0EYhF5deTUj48
w57ddB6zBJ+4FTY4ilIFRshMc5l/FDSyHVGiKcJERJYOAj26L11PlKuTriO28GoloEKHXqt/nhLl
yCkZtrQpJlf/uFjw2mSwfud1unUV0gFOMk1fZdojx+Qld2H4fFOJglwjHlSSzI74b+wWs4KgOyg3
7GObxoJ3QAFgtNxmlH8kSZKeQ03bg2ipj/m2+5ErlClb8xEdqbe23EGucrfSSUnD7W0o+/qOazGk
3stEk5D6Eedowi7rlzj/GY3dfyEmRbeaRr5vTJvygstVyYcczfqXqJfguFcCOwsZEnA7wV+Cy2mz
uGezn9knO75OyY4t8luAjW0JAUhD2QCqwgo+F1qeWx+trncAr3pcwnJyicJLoi5g9sIQXVYybSXK
S4ESllC32Ri7Fp4N1BDPQ0i53EEVH1LQuGeib771uy35F2kIwo2LSeTH/3TL1xwq86kkxcAujjoh
nEQgyekwkV1sej5LN9J5GpQWJMg+Otvc3kvnARzVDCluCX0tqd8UfoO3EINxyA/VAw0iK2h6AUT8
fbnbdNbwpXGFL8a2xTYSECJcUtu6I/uuy5+2wRCJCaVDvxXXBF0L9tiAjklTJe59fprxzjMW78IQ
SRD+zKL2rA2v9xp2vWhNdrOyrMGZDiCpKMHqsUBYNK6KSzCEVeInAQTmBuEvq9YbF2xFk/02Kafo
SPnlH5jK6drN2nUxmNp3tIrpmNDFsNGAm2IZNv/Nt621YQGXITMxO7cw3CQbRhIXLwScnF49SqQD
z4FjUcBXTsYu7sHmzW1/Pr0HeD55wbulGpkwvvdGOoEd0tTy2n4gKRjv74tRg6zLQJG0JgRTS8x2
yjSXXoVs1J/98meVuuJ5mfOh/BvdsGRGvbaAbi9MUAVjJgBRrmA7eFzO9bkn03VE0X0ozbvt0ijO
EJ8X97hXe8EQ8pUJDIsdqWAM1vwHCNVAiDoBLOxTedQEaG9dqfmhYa2UvVZqu6VSFGwFGCOvZ8oH
IuApqkFn0Ng7lfaBOjnl5Lj91Dq7OCK42p/cfBsaNZ+bydi2SdioEpP0cB0OYBpLIQD6y5VZ1bEv
oeOZ+gBYMWGSXpasjj7hDXQSST8VDMboQXe3lkneoLpPn6Owmwe6iGWSmGzWSDEE0vrf65CwvAN+
KCfgTgx1RNRPTHb9lF+bbVj4RI1hXyvY60jU3lwfNUDc4csa1c8qPHebT0+TRaD57l2kEhKl+I/X
XdEdee8nIODPRhenQ6JaZpORfzpIir214VMiaGsOEZgG4S5XNWikfhNc1/n+T2iwPg95gSiypdUQ
OWqMys4G8ovEP71QkqM9AqT1eCQk3OHEByp4F7Ek+HprHgNW2PJuMgjrUAY1ILbZTJDsRD/KWfsm
at9zYY265enOsfAGiqctEF9xEEPr8Cvl0io3DuDaFRIGxHWwSEetGND1JgLWqHvL0isVFzf2iXXV
14XNSN7HA1DpdH4jNRUZWoA43udOG1KtA9bwQfUTkLmhJtKQ/dJWZcmol9E+sxIUEPUKb0lT14nB
h0QxL2XE/Fah1IbsgMq8KUebc5CnmnNQiWjwiI/hUe1RRpySBmT4qxkz71hZR8sTcZfd78YRqsOO
3Ct/3bnoj6n5E9ewH8rWxWlmSxiFSIRgVHo1pJXrMxq4Vv2VFuvTuV+b/5T6ZJ1ydKsy2IXGacZI
4vIIT7WKDPai3NHfsGpmL1CiIdMNVR6VQdQZ9b6FQvWisOHB/u5acX4nYosaClTNod7qllZ5Y1Hk
uzrAvpw8d7xsVZ8zQU/AsvFNNQVQwolIK54IU6pvk/SYqEfo5E5AyjoGhF0Hsa9+YffY/LLnpfX0
tTR9unYpUIKjo3gpVS1uCo5VkfP5l533WmaeQHZe3OH2didaoghWFge7IqaGJXqTqw3l6o2AqMRf
/UByezdz8dbtVANAWphkpEYj7Tk+1ORABI+sfe5THBcq5ek5JtCC/VefdsFalwNrAWPi/Q01mf+v
z6oxN9U/pN71CCVLcTa3UPDV7XSrC+XOqDyVBHYxYlare8AX/cDRIK/KCpzfLBs3K5nmLYiDeAQG
RK7KIxrVAZtCYK0/r2pG5tY5rcqktRXgF7Ahmqp11hN3PIXSofYhylx/coZXp7Lj69/q9sV05Byk
qv3gmQDUyA+N48MlcTulqnefYqkbXBTuZlmI992jB/g+bZdpEpZww3m0GJbCqf7++TKkGLg4ikeD
F745Cc1zOFaBrBb9bhoC0ndcGMrpQ2LfM+vP2s6JPjZrlRfGm3VoteJJi6Vlx9/PTMO6b8hoF/My
aZiFbxNsa5xEf7qAKXIaBMMRHgQYpgkWgmIkRDoNl5NJ00TituvYA/fO8WIEjpomzm/ALp1MUTv9
m2C+RIp39K/2ll9mIGXUnKEdV5T4tWPynJQEJRI8b9f56UzgCBhgsehAPn53QPcEDqqq/97g2uCI
LSdgocrcJvr3aczjBV2r6nGX3pH/PeRkanECP88l/t4V4muvYUxpp59+OTFUuuNxEPxyFyAtG9wB
RMomaS8yut2OMweprUiXqBC6+3PNJFaG+ATWdXV20x768RysK5gsFVbe85NCylD2qd/HRlce+FzP
2Cgi/iNcItuQ5hYst7KwSaS4jYGQPdxfL40FHzc0Mx8Hyxvt7WUjUV5P5OKKnX4uYyd3HbeLRinj
FUjHI/7PQxtOqfoWarU0TfdkQNkLIeSIGxA5ENQeilBIQ1KxGZfVtQXSkbvGy6hB0YkLMJU8HLVC
mIQgStKCPWVwN4C/22gfeKGOz94V0w5FpNzT8rzWuc0IyJ95Yn7W0cHX6bTawURVgwiTjNlKIciX
Po7ksQznvOsG2LdQhho2TonFCFAFxl/RadnmLYk33BE4378RewN94/5nxMeFxPIGQkeoE996CCb9
AQLM+gm8hhQ15imCmZAOEHzA2PHAlY96jkN5hVQOMAMS8D4akd0nK36pCtkaevpvKlYnhdV+Pl0a
iOswANT7mAR63Iltc7OlfCUP33ujYxH/W+vWRQzy6C+le2Bate665MccT1p/Rp78HiJb6PnjZmpM
Gwlvz7U1ZwXGA2r/lJtzVPYGRiM99rCaZllO/LFJl7hgBybq+gV/HQQQ0o3gJKSXzRz7dRfS7Jsh
jvFennI47Mt+fJfNT/FJGDGaM4wzAo7ESxKHK1qSo6K2BSDUcCE3l/PIfgPM3tn9/p/tJRvGfi9Q
gROKuM85gXMyrpgP5e+EbRwFc3WAU3HYGjosjFktbSpF4BkBkzjEBkRGMbVe+MqILeSc6EfhCch7
zd5itbsGjhhHz+shz2Yfkjo03PbgDrP28kBDuQpQWQc9eONTF7mcBN0br3xWQGpcP0jDSGsYFkLA
Z5wypOilwiy3b0TXmg6IyK0gM/rLvk/l1JMmfNamS81qhaA1d9M7G5+HdzOAgC0/xBoiL51tIXZR
UtVfKWVHuw7Knv3geFqavuKArVAr2bHPP9QS74USv3oFndCfO7hjSbeejVeOZEcfeNgbZJ8TLfly
pORxLJ4087nj4W2HdPTLnCTVsfzf03CG0Jv87wZv9I/kCn5bwd8f9/hue/PN3wyLJOIRowoQ7qtw
XKASzluRD9cqMOqnd7xIcB5BUMmtQPb4vJx+R/AeJNBBymqcMR+r7ACnF/PXoRhBjZZZFtwbkMxl
ji0YaL2iNRm9TdXiBbtkTH1p6RrgXV8sDLxBcW9s2sCQy2q/JDK8bSRMnE46aWYecovvxsA8y+1t
Ps0NtRfBPScwve7xUENSPvIgDewqNqKQMPai1QlNA8ndbKA77VcnIOaOHPeQYFTVgtdZR9vLzGDs
fXimiO8x+ESVhPhJt+BJccIy4SHJppMhYWAyt3RNxekz2iDzylq4ALRBwqGT5VQemwG4QCaxnmaY
/RHohGN9tDyO6WB9IbL2vJ1QGndDZRdpU5BZ38q8WpfBbHoWnKpUVUgNyS9TR3NsvcS5mzqR15k7
2tzfpyOs7S+PLPWeMwgv5hwpGz7P+3wv/3ydQyi8MHrJ5iOeuUzDCvN2WTDHi2yDMTI8AkrVbs/l
4w15BO4Y34ZyspcINY/8YB/xg+RxcLOH50/GvtGFMPcLJ+ys3HcypEwlLQ+zkgSgArFlm06ac7Lr
HgLwot8VYqRqt3wN5GwgqI+8ND9UvAENp8tWNP5ugXd0ojr7aggNGsmunIEsjfQH+FS+kF/TEPYm
q2ljCV6vBGVVdi6bN9ojIcllQQuyZatPZ1u+wxBzTJyH2Dcc5fPrsJE/sY/nDQb0gNJSXF8dwLuw
TJwFPXcGbnXe9MaPUG/QhabzfdEq8n7amxaBthwUUTEeDM5jqGiYxVEeyVipnyNgslc4x0UADQCv
zBRhK4RIzCVDMpE4jSYYOWbJAOjcdl8MCT1As50lQEUBkxb0goedS1m4r5UuzX4S4W7JA1VxOucv
qoEaSnLf9H/4MRV+udoZMulRImOcaN+lP6K4EbwBxl7hroAnTY7T30Y3QuzMEBxwdoKY6QNdc1tA
Lazot5GbNKUBrpfJ7h6SxuyNBD5sDB+8zKpFLzeiNynkAkulTbAwBSxJEFs1Z+wfN0yJ2Ui0t8bh
4mXTnxGDGp//u3BdcypOuj76pVaIT1EpYp7inTOlEgncoJV+uOKmHq7j1KoAkPusUFBPQCA/Du9d
WcsfRtpV+0RYSOjMA+RBu6hYQGcyPb0lOsvqQgC/Yw2T/wsbOkRAdZSWFC0D2/kKMZFfhUJhsnRX
O4Sx2Z8KXrumv2mnvZQwYFc0Cqtb4gI0XjKj6uyVswDmwL5GU0rqiv7/S6XMQtCJu60yqWSAJrPG
fcynPMKdu8FIyFmYJZvdh4qSsFsMxnLscS1tV9sijkN8BmqVuWCX7tqW0a9bFh+NSgOTrsxU35Ia
I36sWRPsY/W+4AIaeLk0fLWq+EVmBBZ4ScYAVuL/6uci8DdyV3sGMZp4E6u5IGmsnUmWwYdNJB78
x4J0/GTDqPEREvAPEUysDBFDYS55bNjkJK23x4a/phVmIV/XYu7ppG/7yBYRUBYijk+TUVl3vnmH
x4sObkqu7eukf8UkH2y3QeT8KdlqlT+2SIFevPyXMWjlUgrdty3E6L/g5CvkihhLIpfplaJrOQwl
8lrabpq3SesiKnUyJIgpxCY82LjErSsui+qkqMkB3JpPHPJ6EPjqzTdkWD1UMPDZHWIEKrp+wtrA
MAUW9nz99uRzJLqBJIP37D8VTdaJ1PXj32VvFppuRXN6/ViBOaBXzKwTQLbxguORVFE40HfaSv3h
z6NnjzVE6B4OoyJcJ/TtQmHWgY04pcTLxTsGALbf3yHoz4Ko9g9fjV9z8Kqf8W5JT72BRyaQxV+P
kXbyMzyC7FWieI+wZpoRX7IazJ2Wf4rypLQe6syrKm6Mv5WIXYGQlRDgWnM9UqrUIljLvuHl5sKb
yNqc+6Oj1EV8REinGg0eGNUWrzQScrwooyhxF+Dn2wnP1eF2TO53J27jwCFjUeaAtuk8dyAeywek
JyQ8gz5jjKwIyR0hdtHy13hRQrDUrp4V1Pa0Pr4zboP9j3+D2rgkWcCRrxIPhFlr1YTaPksHkRQq
y+9Krqu0Iz/Q/ZGh7VDg9Jr6SbGux6sLmeMWwIlMUE6MTmj+kzWIpVQLsFklOSUkt3vJoy0fGx7O
jVLxIDCym3p9vwlkgQ8RF9L8L7axh6m37zhEDMNodaG00V3rTt6TtOEaEMbo30MbNXeHsX9Z9tTd
2oTlMMuOeWmUEkWFA7Ua3fSebda1NY2FxNdMWifikPUFyLbhwhv/hip6vzH/s24Q6/or+7bWOtcC
kqRkna6SMLDK15dGjaQTZHt99EgTkmejzepkn2DSc/JlXNk/w/tGgvC+28PRhoOjQH8TOiJ+qG8J
i88/dWrvJU0fb4Zr3GesnLjnuaRP5ElizaC2vqK5wdWVXVoBBfuyVNe3R+ozKFa2V5/3W6cW4tHZ
zfrMTbof7z5tjJNxsCC0n1y4GRqcZS4A3T2M8NqUsuvaz+IiP2Mbh0sufdNeg0b6mqByDi/pMMq7
DhImRr1NlSJikpQOojXJ85w+ZHVlr8ymTU4Kv4IlrTpUVifg3grx11nwvX7sFUvtWX7FP9iCJ5et
wWToEOMiRPhqPYyi6QRKAV2rvSSF8ZPwSScaW1cK3AgTDD1ulicXYbpQFUgbSc2yWt29S03zwpX9
/xsQaZrdrDmXYXM5CHxsbjlrOz/pBCfRGukpfzLUdzgY8csj8GTGDY5B+8fYiDhb50xh5Z46dJ7d
8toy84cnRetxBvp0Yio3jlbPM3544sW2Sh7v/3RFI2g8cyxeEANelF76jFa9W1TFN3TIeAqDNJ9a
j9q+Eq6rNHm1cCewNiv5HP7GP0gefJJCsp6is9VX3gJIqZIjQSkEu6BhCoYbNCx6Xj83r8eCw6fX
D/Y/wljfctHvw60+dIcrJiiG/BS/gz30+UXPO7CztCNgi2A29Tk+lZwu9dtgdc9s5eHy8nyG5e0L
ha/v25L7asfRKMARt63l5jDtqvYEcqqMx914LTAAjX2ljhW86OqwCIAKus3SezpkUrPAIncnSqv/
zteugkJuSbI3n/1KqFvl7+e09+gxQ7eLHtCsJ2aUI4sCa38qA8JLiU5WD9pG4HWJSEw1GOeDGC4n
1I8cv6MV8Jj3Y5st/G3vfzAgbfrMdbRb/1oqE1jkV8sVxYcytxA8hJWuJ1p1DbRgpqIQHB8nhnun
LxELjAZtMRLqLCqEF/pV3jaAh3vz6V5j0YQADR/jc9s1mdSiMRWgEE/R65ISt9/oY4scq5itDPOG
kKJi+XRIueY27qYRbpQ33JTBorA4bPcHOxFpr5DZH7tPoAj4e0ZTsR8JOYE1BiPYb9aHfA3HCsu1
OrPEt2F/EHgK0s5ngeN4TkvFRPce745qUdsq4W7aRAkw7W2FHd6AQkML9Z/SMi0z/3lGBYHzv2y4
UE9vdEyOkhGhIXcOSMyiznEWJPGluMlTe3+xgu5Yn8nUQsomziWLp7VU+2EVSafexfRn6X8jwa8C
Nlnd9NJUcABaEwEXGVcIfJqba+vtMp6oiEEmqBCtfSndhH9VCaURlY6mgUyedhdZfaOssZEp/c6q
cFMY/cIgn1CiwuD+s+qzocl6FezjrRGxqEMRhIsV9azVxO8dWm8nzdCPRas7EBuHneJ8lrcc9WCM
AAi/Wk7lgkqUwvemDssWbRE2AeSERCeqZ91lZqiaQMFzLgkhWz1Gw/MtJatayx9BbtEA7aGsSyIa
8xbfI7Yq7KNiFrCbumkmmxRF6XSuRKZD0nwk6+IxUcdTCRTmDx8yMsIXCcA9PJ0mr/9LijU9IGDC
OMnaM0vFU/g9xW2Qt6UMq8Xs8TIrhYuwMx80aITggsAQ+0JxNWE0C9jNSf3tG7n9bXI3pxrxfX3L
vRbkXKaqnrDbrcs1q9PWH03OaTA4iFpU3M9D5YqEeW1LHVg9yJquHH0DOYFEXvmw6FK9pskCBoQA
NEpmG/w/CQepLVZPiD/VTFuJ0Xri8wbZQdt9U9SL1QHXaXQSDR67nmC20zgX/m/L74N8RqqEhj4T
VNdHv+W+L9xQYQSFIABSXPOyfXKHZw7I6zvlsjr4pOdLYnbM8ZVDgb60+cIPJJ7u6uaF/hRiSczl
vvzaURMCiYj+s517VEiDunNzSDC7sFjp1vQ5DjB3XTAQD1e4Kf9g+sCkP3YOWbf6F4Axc9cpv6kN
MTAL4f3rC4P0/sgR/FsVg4cWkdeYMu70tMUjTwgS80OQgdLCVnBjKXH0aA4AveVblRTqRZPkmlZW
wUk7gdOfou6V4973sEjrbj+VyN03dN27ASECFZHaiS0efT/8g87S8iNcuQ/XtpWYV4A7tPjS7A3G
0PAvp+0C0SeXBzhuGe+oF7rBKqi5jGANLqU9rnMiQf3IXkTRUPui4ju9ZMq4ZV5sf43QZroH+qkn
YWgWP17JzERt7y14Sy25clwrqe5HJXMeOj92/UGMsstLCgqyaxK/3GJioGlBoGdpDX1vwz+oUK8A
+68dSlcbHTktsXE69lo0uX2Fz4KzWBl59ChH6ruzCeqWky4Z4unCSPkksWVVduLR0v7u2zQJt0GA
URtZBvPHZCYbWRr7hs60jcYTfS7N+a7NZYhEE7auv5t4EMcShogSEevKGQqVmW3zV5J2VQssU08U
3YGIpSNiztwSpkLSYHHX/w6iE2zifEH6sW7bn+klNGW6hS2HRa02fxLVoqypOosV47+PNXt4eBPC
BIM01QS1wlh07WKy0sNp/hH1zHMeylyBI1+nGq8VM73wvgk0/RP4LGynYvFQq49YAumpnA66gz5l
MxlqLIS389pP3TNYEyaWmEX+in/pWYKYF/vaILcFh/oso8lnpgvkoXtkZV4DrLCfIWqnsIASvP4k
Vgcpv09SC+/0xcMSoAj534cYOkL5hQ5Q9D8iGiOdOrw2Mr0iFa/JIIiUU1ZPkicJbZ1IYDfKiL6M
Vd6ZM3/GhEwsUTJQMznJwNl6ZN3jUC4eHduMURmP+U7I9hpUbDhKrEuQKUns0KpQADJmvTt20FCT
WmaDwOiZy/XAz0nVXrvNYo5mVTGswYF6K3O3xHhLdiFqpfbC4z5MbZdGlpTouACbju6w6ZAshos1
vhckaU98DlwMKLsPAAcC1TpXP7OWhXk3YksNt8jhs0RBjMetk/AW/MuIOvVGhKz2Xkt4Pv5fO1+Y
RQnhmDv1juFbnUfCS5AdMht+nT3HrhyAxZzUNleixPbbX8QYj1XTfXInjZfl3kWZRiXJjt+AZ8bZ
j+iKCdgIq1ZxyXlrEfCsOj9Xwp5asQBEA/vRPaQcLVsnDHrKR1UUaPS2RT5g3CpJ+VWFd3ySSxSz
yEfXaStOET4sKcI55sdXuPsF31jgmtU0/+AD3rNG2YGubnA5B4gxide4JhCP66J2z+GwGawqKi4C
yZ3Qp7vvZNvTrz7O6ELr1Q3QzFix6r5QkAhugP5r/vnY4MoOVFfsFxTSEMVWGqq//Fuz/4kKz5py
t46f4V4pnAFx58vcwqMFeOXyVPnVe1YcOrRb9pMiOSxlMaKvaSMsBxcZ9o7mtQ/chfi6bkvmz43O
ttqQ2NX1PkLq7ORwvy6NADCxLW7tcAKaHLj8gMBYxfymg+QUhvP0hYTmGomTNPlGUSBySBDufDAG
rXiWshy4HZbU17V+V0CCDl8EcBNS1ott8TyrbZ46boe2oNFgFhZcWBnTpu0Xu9Rpdp1kOPHKckgS
0EQ/9RMhrXaVz4jS93C8hnGGKM06nBKf6pqqN6iweXVu3M+xCZ1afOyjQdaOGbiTZWVQNnoqs2DV
6JE5QK7WiMTdqhyuq2mfF62B/7algGk1MCPUVtfIy4+S8m8VjiNPi1dGqw7hU71y/WpsgIVZvuRk
TaLGep47ulJ5mZv0uA6C4Cy8XHYUO0b4HhS8EzfnNWZNhKbLS3rmMEXiR59wV4LBoCgx4MUVI6e0
9G8lD5D+VFfc5jB2lT2jpN4EGjQuvzTdrdeWD43OyvOHZNOLoiMqPkp/9qBbCLS8WW7B3BMU3uFI
ug66WBT+gXQsA6FEZo8OI5/UinotWSEte+dXRphi2gFLrBXxwCR9QsUwqJ9q6d++r2Lu8LrSjcki
CFWGGZmqJXXre1x8T5ET9/5yljRFfqO3XNm6Or9IlQ9HvW2UfFf66CvDIGKjsRg6mz/sdLlhUGJt
4x7HmINEAlfz1y7GfY00GoXDxS6I1IwXm0Aq0qorpyoM9cqGKRaO/Y1SZPOqvT5WS3Qv/JGkh8lY
owgJKSy/ofBKtv++7rhtPq9Y5y45L1RizRKANkeqZ94OsRbu4vG11wQWCxJGtNV43CoPs4fONv64
ddsUUhFunrZoaWiifsW72trudapmNd63UMB3tXdD6+0QJClusUJzqCrxQwJnpXjGyEMhd5b7VHX5
/Vu7X/KGcmm/90gHXUx4WU6Ykcxad+BuYo3vufDwB1rvzc3r1r8WLCvP7PZVfP7B9mn9X2C9gw9Z
UWYdAwuDB7NZcbZJ1nUJYmdAu8MwPqxEhyaqmaRTSUT3WoIxsYI/bb9nadJgJteDyLSaaDjxlknf
65YqFQZ2KUImzUL7MNhr23S7tL7sLU327QYziDlx0HVBZhsAnwNJwjuliPIiXlkiqrIIM9O1tAbj
Jumza54ucSo0u4g239WqhSOcdAf7dzRY/eszLNVs9BX9Wfch7v4+TyreYPKTK7IyRz7yyDvNxuzz
rUCQY8P91AWYnLxO0k6lKbJ/319BUiVsdv5IzlpTBevuPCOa0d1QwMdvBso8dxjz9ft50Bl45oRW
dZGRYqYyIEnH57TPu/LfsxLQom5SLJEBWs/dP4J50D+g9IP/ToWVuMmFMB0HhayQbo3bjv7Y2aG6
bi2cNemmAksS8GXgJHTdvbsdleTWKccFBGMvIoeW6VWgnt3Qf4yQXrWTWRNl3X2Kp723/UVUbMif
qx4GOirHP2H1KzzajPbtxWuD5CzCvDrMQetSGGvKvdbiKc7mXEf+/dlO4709umQPd0qmg3nT3d/y
57K7MyYqz+WDUg2hSTYcfnm7JkmJUIOUna3cKoljR37FLfDXOhioGZ4Vvy8vJCxXZiCBCQY3fzQn
B/KY1cUomCUkU9vQFkMU4bQjBUITFABvLAyliDP7ajzlAAQxNxpwbobFJU+nOt0cE+S1g0+nHlnv
p7042RjAevGTaA4W1cmEdFokmUNebPeVAWCZQO3bkuj/cqfrzvnqtgrfoLeleI2ULWfaRKDAu3D9
k+LsFkgA7NhkrgyZpEmNKL/HJiux5cY3me81mlWXpcI/onMIYe5VKJnkKVdDvh5nYAqoJpgujo4t
wH3HElv1FnaIp+VAFU9yUSoW9DWLmx772pcyqeRGs8ESv/oWPm4bav+k4YrajOlAGom6QXdWu9xD
LxeqES9oQjtM+I+KX22UDFu+m4gFOmIib74kzZbyDkQtypxgDMbCNUuLx3kbqqPlSq/xpQDY3zwH
o23Rap6mFj4n40R8gzHJAiE1u/c1PaV007Jjl6h3SIha6Rnq46A4QK/zt2M0PjSfe2EVOfg4nrUS
GzmOU5hJZZzkgkBSUuTaegtfKPU7zXSHcgD86WBrzEnAdJrjtWn6M0cBwNX7XStIruht7Mq8tUNX
ddT/NvL2hSXFWYaRVfe1jSQfy/YkPnOhsbNZLvHz5rYvNhSLnfvDXLpowG0GUcvzBaHsoYFM+x8u
u8qdCvmfoogS5z2c+0TgAu2AYUZbhrOy7zC6dI5TV733NjS7dKFUu+LVfv+UInpICCW1+sXKS086
nKcsFHrc98N95g5S9Qo2YUYyR+Al82Z7mN1Oxs4Pwx/wc+YFtURwHIEFCQLreQWXtebNNqkVB9Of
A4VZikjn81Qo/BZ2JWKOkAmUDHVcHnsqsHDCLeSm/8EIC19B9ChM4o0ailu5BLBxCtyqeguHRwtt
fitQU5iTlq5ZWJFu33VDaOKVbB2ACpybW3tt87l9qyohE343Sx4b4wm/wJlGSPbAWv0tiMlydPzv
1x4QaQI86N2ztAzYuZ+oBB2SBCdi2HHV4czfW45qzCMNBXTRPTiZeqatyFcHNyaY8yHYQYRxxLMU
9s3J62li7L6nAw7zIVN/tlpuoWSgGuSWUpFMcwg9DW+BEZMtcCaXc2ZzmUJgmgZkps4nYS+UhHCo
yN2y6V6IZDvl9jjLSE1yb3Nd6FxO8CSltwlyPxhUVJeP+3bPr7C1taCS5VgI6DAyMFLrctfW56qg
pk0j4XICjwchSM/ioQyNj9/Ek9ft4sn2y9QfBBpS+ffGAZjgMzlXrql1IUPB8mLklbfenGvLWqR8
RAzqdes580zYKVV1Mj7Ia/vB+jGAynIuKUMznIO07XT4FsqRWjFvdopqUgwe8fxryNomW2Fx8s9C
9VmqGF3FGLuZl4y2pscJZYEAVeyiFW7XfLdOYW2HIPLJYz5r3OuI8yXzLphbouSsRVyAKzJr43B9
veik9r2kiKxk711rv6SlWEaKdq0PDCXUD2JmL6gUfHjTgu7ATvlvZyNz+fe3ZpyKzFFKnptL4GU3
DjbAUT78/hAnMKiTxnkSqvIGnQdGCVAbYte/gTRsQL11GeEpIebjOhfO/zpcKvSnY1ApugsyOyws
CSvlSRn0l0mkSnuZlBmXBvILxI+Ky/SrqiZcv79Wqmc2Gh9Ql3nLf2eUJ9ZLcoMjYCvyl4IniKDn
kXAEcbA+2fdLyoJ59j9ciLUfmA8kruMpdBsLfFamokb8oVDcxDmb0+4WxMpF6r1q+mxPgDWMKjCn
EQHwsTE/Of1N0BSYTDDCmrzWhOgDh82leezLI1GKsIOjEez3NvueKDZXCudwUaVwS+4o5byauSjL
W20W1LgAo6jKuCPhrxwe5x6HXLU5lGPEN7CD6Eq8YRVul9DinrdkHR/vzhPOTQfpVP2yTpowUCkA
bijiep/ex675gRmAxhBN3IxnPgRPM3yrbpn9ANLSP6zRP9xs+CVhZsu1TqEuGYEw8VW9PGIuFXKr
1HAaiW7STZoRkzzmdAacT8sVwZLXGHhf6VpF4I3WigTZpAzJkbAv7aiaiC5eib0L/y6aUfRJb7wF
/ZiOWUeYXRwI6YZLJ2/N6q9yVioB/utBFT28iFGK0338f9wtM+JEl1/+wMh9ACK6/1TO6KI9wLOY
Bl0nIbsUyQ5NecGvPZVL7fSV6raFCL9qsOPwe/TKhZUQfWvlSwlh6F18Cq+Z+3KaILeeZzKItnI0
OlhGWGIbhYo7gRS3h+/QrgvLGonfOQeMIdl5jIdRrJlyWEZ7tf1j6W7rI8ETxhORI4kJ9Isr3p1A
ZwKLHNBtOWZh+8OhRq0GmxtyG6dnyqYOZlU2xFtXgsKZxe7zd4oOhv+vIIyRzV1sw3iIKUqnpdh+
kR2vYA6J0sGgEWAsvUJljBYMmNaNR9SMzONbeI2+QA6n6Ea9p46aRoO/uXeffIDoRN8PCJsFZ6/o
bR9iCYcAk+Cx0lQO8V8QlT4/UTMx7tckcMwSQfaLockkroXLsml3DLVsOHtneTOTNRAn0UFs67xD
RVH97m8UMS97QC4ZBzZc/NItT279Pd7fZAMl6FA6U7FqqtR+366NCwI7Ys6mHUN5RITGi0NVaODJ
3fC3iZPiWGHGr4zYaVRcSdST46WkyOUKZEP0D5U2OvBsDsVVGJmn2ItFODkYA+2feGVsE1x5TKIX
h+txUrCnLYQfz5Y12OIr+9UR4/5dykvL1/VuntRGNyja2EGA7oStV0oeOSCxHq2GKCyHqVP1oR5q
Q8QGc37tEAENg9998KoHMVJVYu1fXcOfQ+df5U6P3r6j5n6ijkbWL9rqoxc86c8A80btUVkQn1OE
YH+u0BGMlwtCQ/fc49H83UL9/4VU2U68HwoP/8MByi40E49WB3QHQitp+q3VW/8ZKXfsKcqel+mO
25la3pTB+Ln2ZIuMEIeUoc0XILG+dHwwNkKAawfz3mPK7q/yC6hfRbxwvA+kEpfZf3IddQ4oIDP1
itSo4064D/aD0HH9otWZT1okUiaOhjJOsVFZ7u9huDKEWxymBDz1qjJyVYWZDjyfYyqZ1rMT/QZv
TCenxiT0y7HI9zbFLqfd7LV2kxLjFk5vUmuPFzxWhjkaw02ZISAWjyuuDfkzaMc4MTePZfYXFImY
HhaKtZctihQ0ie4QyOU4Ngilm+DM5HZdENvQhB1/1leNbIY5tf6v7qWKmNOZy6AgNt+jQ5ARxUU1
jZYxMQETFlGQVvwtJH2NmAqwSKf35p+wnFMHBir7YZ66143BRBvxm2aNcqvSe0jwpZCPb/QSLTSX
lSDe57Y8JgzKeCIqyGMN7G5nLkd5pP+6Mew5PfNLuioDCj/6mHx/Y67QyFtVLpC0kZXVm+09j0DA
qVGPgaj21ZaGY5hTnkkUNpaxigAE5mL2DCH4a5j7rMX9QDHK4AmdscdlpLJTh4P2MfgJ2htUCdO0
Q4DYUOMnBB6Wdtxc/PX70jG9ZIAvduk59SfWtDi80mzSnbmFojYy8AVBD3GNHqgdc0Qzo8kzbNI3
E1D9aDiG9EV4tNqBreKy77EaO0y5xTan3KZgjZNtHE8Hvl13dzcHzVk3ZikA4Iu3K8TK2kX7w8CH
g0wvQPuroH4FxeKehk/7MMepKQYr/0AFKtmUEZn1UhuZHx6Z8Rg3mf//LKuHN+IbYY5W2p1DrE+g
ZTbwQEfuQb+zqvUH4WK/61ljRCSmNglL0tNPOpxg9InfnvpfHuqAibTYWYSWkqTyC2vUKm83GS0Y
PaRca3xBG/yhTYO9yrcSxA83/ErrKJxxIj54Amj120DIV7ua7sll4iKGC0/gbf0VGbnTSidRB8GI
MTadt+aGKoNA8TbGy6hixbjM97bBGB69fzl1PDRgsgUOfm0NKqL9DypHHgmVHzFSet7bA3UcQ7b5
FsI2UOrUqumAQaV8qQ/c7KDQug1k6jfMYwlE1XpD22FSupaj7BdV+2X07cJ1tZf6Z/O2e5T2uYlX
ilkycGaZAKwzbDX1fzNOMFHq1y5ZectIbYBVQYVOwXp/ZTtG+2zg+OuczxvwqCHwqtsaHrcv++sc
8vOPEZY0WZZqW0UV3QSaG4MHTuNayDN3X2dQ0NVRL7+Z0PqfF0qBkYAQMHqeqRqMQIqfbousr7+p
chuAm1LXcmYuJmfE6Y/4D/myDDiB4+EVCtI0r4hAnH450JdswbV0Co76Im8/zC2cuyPUGytV5oaf
slHtdVZjhxnRjAHywEYO76MzHWBrbPvesAZm6NMqFsBM+40p3Y0sdNqqVoSX04aY2hsA7Mln9RaN
gN/PVs+bEtVOzQDLjFCxnL7NyIIw5yTLv8jJ+hgtDPdxXqweZUBZzI/r7e4ebFIW7BYi0hts7kXH
bqAiiAc257Lqkjb8gkhd9g/8OHJ6nPmRZWFQaT2/2CfhlUDjoy/bkmbtRCiSaVZh9UB2y7hRRmQI
NZntEIeR0F8hKDoY4JHg2Vjfw5DnFVvbq0X9JpeN0KBx+4NY2pk4QzbehiTqOI2Oo6SDmMt/45XY
wGFCzg6lrdScLikJ97eZwXGFvjY95ftnQoz0GPeONI8qKk7ruVPz/9a7uTIGOa91HIUecFX2SDs3
M0lyc48Yt+vTQvTpxBFYgIaRLtdIPpT+QS8HK8gh0+d6NgH+IsP6P2EjoocwmswdSr3vUdrWjr3q
a4vxOMao9z7pK2q4ObAbp5MdHWOfhsi1z9un/od2/ftqyy6WDyzm9F32gYOpS9jMbwXAAxSjll9i
GI2/LlpUrS2oA7YW6EG5iIszg660mz5+ZdR85njMDg7pB5EFkuFnwikvw++RGwAMozzGIpFBBnKg
J4p3xzFIptTdYM96v+SB6J6cYpDo3caitHl0uXOFpfJNpLYKKp3Rt2R+BvpD6XfSwTR08KTWwSaU
7wfK0awMfJWl7TjRGieyzM8X+ZOEHouLkrEvdZqeR1vFxMP+WXumOu6CZraz1JciiKJRB6GVQIVB
DPvu0kpxZP5S+KIVHL6f3bmKfr/rSV9qcM63qBMax5ou3aeURFa7nPliBIgqcEr4e/PC8upEc7Q7
ePEaacigO+jSnQadlL669ypddu1HAgDQYDGTXVoFflEC3kYLeBL80AVgWMIu/JvhwRVAPZq1cSg5
xe7RPqS3eHBV2EshTtrk6ALnq1y7hNt0FvaqlOWfxI9IKO3e1SXtIZSeIaHztNn5v/hEYVfdG+ZX
RKOHnNdEbQaZRMfqzMWX9Km6wlA2WjdZLWCTQ1IuCaFMrUAaSLKIOVYHrytf/JS3UhNGKgyiCi7I
WN2LGkWOG7LYevGR1Bx+DAnRzgv14C9rV6KN4T+io9NEQY7121QOqvyVkwFCflCvsjBSiuc9s5Q+
cVii6dSpJ2SaPKfab3mT4ywvMGMHNVRYqxFxFPKdfP8cdAmnW2RNNDn02LTRw1nvE69S944T017d
bjdLBfSvDroLQuJVvsatE2PAZS7F9vI1t/azcF8kS6FalQsf6EjvhGaQMt+7rFdZQa7MzcYNeLmo
h+Mj3MKBXSt/bZ4vRaeQNj7WGWQCZxHKThVO64iIbuVrqxT9NAqFZybcMCdneUypd5858r6Wpp3B
7QEEss0ChbBdK1mGN04lRhA0Gvt3jLy7CJ4NLiW87oJ4AMeULjGZyesSGOz4F7u4V/sHum7J5E6b
wQrIqZJP/yp8RJYY7Uy2UimIvgbD6V0CZeTsV5M/NhHHIP1DzQFKWBjCQj8f0lotAcIxiDgOPXwq
uMfvjB/tubdEMaORka04u0fKneYXPNLg85IY1WGcgLXvvaTP2uxG01HEhzjmAvWQihILqk2y6t81
kcDdE8tQgUHXHm6WJODbKjOxk07UJaUasgXNFsjp9qjcOcxM0k4kgi7mLc3tb+jdJndgNL5ks9Cw
3R1SDkqMEfj7fBi1SWIImOym/DGQ1CQvz8UGiu6+0f5ZCu5dJRp03mzPgVC45eW4TpZoLt//d9hY
sHiV/sAqDm9JxL12JpZnTtUwDMnFTk7sCAkcGkftnRzKTHB2rwQiM5FLH488p/9HNjg1KWEEgEj8
EwtrGQJ3c8ZkRApR5MxtE7MnAjGApzB/RUdqwOKZZm/ckcsSIwdx5t74CQBV8sM38qxoc4T9rtQN
ToVuN34Muc8Plvc8PRQc7/550maj/ikaMrJD83J4qPMJiuj+eNUSJw7JlMu7qoKFj703tKQMYet4
Qolt3lkllt/BzPhWR4hWsdQns+wy+bC/qx9m2fZ327BHfQo/4osQpagves8VV/Kv8HUGpwKFofSZ
FlzKyJSPMFEgdY1oKsHdocOx/2Wb8Wkl0V5p/foJDSwwQSl+DzV1NJJTBqxE7HiDFTkjYRHaDURV
K+uYBnPJt6aFc/YhspYcVxCVbUVk7OL9kFMCpXJzgBAjLu3LRGdgf1S6Fv4RQuC8HNSPOQdrIHnN
o+r+UMjqlKAANRs7XZFtDAKgvvz5hwhesDvwooRaBIBlIx12vR6cp85aLK+Tdel7sAS+9TRR7Zdp
s9Aq5eR7avN/EmlBebcOboX9TrI0cdOX/pu8ZL7nEQxwHaLEnDV4EyuhOCUBmSVYlU+KXDVhESlH
dZGR41oNKI8csvXJvgWLavLxUfziz79YaQC6OCKbDCZ8Nt7hTTQeAoDbD+MLznpZpYK3Drd+RKsC
s8sOhL51Xek3WeAhecvvEPJdIAK8FM5AJGVVnpaKlwRm9hGNV1uD/j+yG73qwKoo375vwUMrU73N
qOHkLz/K9665OEetUo/IORgG+vqt4L1Mz5RnQxgmXVmH5lBJdSj4jPtntL4TKvsUBslCFoPHjo10
5KVGUkYXLDGoqIqM4U+CMO5+HamRdaaSwNjnMnP63oFowLKANnFhE8ZEaP/2xQ4vKd3fGij0JnZY
9M1y4sEcQVD9gQT9kXCko5aSV4wXLyUY45e0ZOnLAyjIqHVPU2s8BBZFWzCSs1ItS90iCzjO0jb8
mvjSGlaax2qZkY1SktuOKIwjkbpYrDuiHkjp21JKO/fZNEsZuu3e0774gr2qW6Q2LoB4c76CWO1C
/f8zEKQGoFaxtmR4zzHGm3YBq52iAa8bCOwlaLOoBMwEqL1jZdPfzVxcNw8qOx74lQo+iwZtYzYF
DwGeKpFBKvbXrMsMW0siIESoW5xxVYWBaI5oAkK5Bqq7Vc47RNyHVPKP1Mt0j3+Nj7qkjNYOeY4J
YEEoPBJnlXJDOC6OcHmcfKeCA9KlLbqieJteXzDNg1g3mb3LycFsiDbRm25kCJaVI4GbPpwI9eHx
/Se16c1gXT4/U0wQt9oQevM0dNJtwd2yeA7BTv6mkBQiWhPbJ29OS94nJgE7QVOkPSi4wmxfnxme
Hc94Bl4nqA3CbfyU4RHenf+Z0my7Ih5NPNGt9x/3ONyC9kkpQpstY5DEDZt4Rvkl8zdIid2QL1C6
0LVl5NLeCJ/ZQKqlDS9He/O82yVIBe4b0Zx78bhRcos/Wx7NehtnODMZAkm21Hzt1gV06/VBQ+S9
4Lb0Fuc5cH3K04ktkvV2sIB25xAeYkxdWPaqTKvT80ejy/37GOoHhPxTb2eYqC0YzvPjDnd1KqjA
+EZmGGFu1MNdYbwGUKYNHdaEnOO2cQ0DD6nB1BqLhztLilbentsC93sqB2/Epl2XiHqimMrCQltu
4V/NZDKzjhdhhU0eVrK+53q8lnHurtJs+DAvUaW6wCTTwMepVwJngECTqy2RpRV5fdvLUmKtiEeg
uCOCntztTyzJSEGTBfOwpPf5KXqNXLt1s2ryAbHSRff/c44Q8xIPDmKFFaxVMypkxUrWrdyv6i6t
nDHX/81ZWzKvUOGB19uMrfpym2iYNOufwA8V7kf1/2IGWdjD5wB5rAHsuXc0lictg8CCZWOtgNZD
ps69KSL0+oByw7GLPjQjlDY2RAN/A8vuaW15VZkstInIFk8aF1p8LLnQMfdqwj8zgbewgKQl+NZf
GxD5/9ER4afVrF/MAT4UDpYU6vSO7MQCmPLJ1MRP09u2/lTo8m5bk3oaelkHk841RluN1566xawa
D6MFRzC0LlX2QrLE5/FxOjE80pGXVEh7/W6Iv5mnsxHA9ol6gqhsajlbkMtud/iYvkPP5s+IXbFA
AlVIzDYjZdG44pxe/2t3VmjvSIb2Y4ABFjpLjMVQe+rOQUgU+ZW0VLczBl7b0Q9Vw5IgGXQxiqaz
rY+4WZjEv9NBKc7p8qIwWJkmMaDiXVhcSwEISdX9Cb15fQgzvqyIWe6SzpZeJScopOcBqe/V6qd/
ROztKmsKTdTKrjn95MWuJ/1BCroa/C7eNwFY3RDcjVcfYUikuiGYguitn/iq10/0k2ghUsxcsPn9
lrsElStG13d8a+gIfi3D9AD1gU95aFfPui9bn93tSqT9A0pQe3Vne8CeknZ3pVS0M6bHbIr0Xrre
idGsXuj9i4YwlQJYZ0Kdlj++RmuIOwaog1fFjS7BFW0xQ7SJRLxO0xdi8YJYWoEWgS1b5Ozmv0SS
LQpf/xF59mmbYpmMz+aFy6YkE+0r5tOTt05cUed8ihkzJCSNaoH65oXyZcn5SZc+uTjo1Ak2O4u3
WgnfOeptc1VnExWPoJZ6ISU9IyvY1HDod7aQz4k8j8BR/uKo78As8pHzFyKXL2yG/uBEJO3w6EW1
4pSWB7O9/4JGF12LVnuT6xtJHbVa3lzmvbkT2B5SDQjbKDjCbnsCNtACzG4OTr2ICfQ6DhSMHaSO
ow6f5QZxUVTj7dNSvDShYzHbhZ1rFoxVOYZ0H06e9674ksJgRPl93Ostq+UMLoEbn92TVfIKbDTr
hvGfBrBHeSjSaAAB0wZulG2ovYUvAIuwyF/IHcBSjK8ZMpZbJ6FZMEUPXjdP/KdXK4eRwXe4Pz+y
u8sEZFUclAqjmtD2WpolpXQjY69FnXcXAyv/ZI50J1ocZs86fSFuFbxeqLufqZdncy0IdYQA1HoN
VwZ1ukYlHl1pXYr4mbABdhcmeF6AfxmJHPrrE3fDwH+PO0/x36iBNCsmdQm2eoz1TdDe5KNo1Ym9
TMkmWISWCKreltrBY4htJ/yJYL/qHxIMOIha7iWtueiPZU8VITcC6GhKZm7FLTo8lzhBR5HdxW27
x2RUh+vAapFHnEbEf39Vauzk8XpqFGjmPWMe0o8xI6UZV8hBNdKJQUAHU43d4j0+Qmal08uaF+8e
8RK7s1OFJwbMTXRmMNO91wt26j6s3EFgr74kZzNL5Ksq4q7KBbQg7MXCvB7RBJ2R5Z77ZnVvO3rc
+/vobG+/gCLz7Da54IhZCL0jvb5UI6X8HCY/szmyIxeT/bn4ACOYpjgsLoLJY9TX/iniE/riiYFQ
TiUKBm3YMnyeEYCVItjHqGZHdYJdq4jKLvG6IufkjU5SmbiNyFgIYpOpHLekBXmpczrHzOjxVc+z
SAt4h0cUcAc0m7SIn43h0Q9tbH+tMIXdu6tBurLTrDiaizOe2mrPcQ7r7qPoC4MRxASmudHgMaWm
zFUNT+55Ono99tN9cs5Lqvz2atvIL8B6UNCMep7p8rnMHoN/S0z2N5jCETA3ART8fC/9ySMvDGbj
8UuB1gyks8wDDYIvZF4rPRFGXZ5DidRHivM2xcSHZpqEcH8A/M15z1jTbYXeKTobjl91B5DpR43f
OzfHhMd7w5TWKUaS6h7R6uQsCCew1Yav7iFqg4vpixjhKHI3/3vY0RhtConw6dQ2bUzBzwGAz7Hp
7VPpkZ4bRooMgNW1JS9EbWJwAGUVtoZFthUoRdptoFm/s6keUoDO8Fe7UNROIdkmujxLgmWI/OjX
LRQ/Bl8xvEGXfxgub8c25CWlU4wJRhm1zfzU71iTADL7kO7FMOWI5+yqoN+/iI9u4jf5RukrPHcT
epz7Zcd2oyL3KhdMw3RPEqtjI9YITWe3mzdCeGwYpj72sUxgZZDwr9hNuHE7r2pGYZUGTT2oWIUR
EESGkulswWNSUIZBFVVbt56uRgnJiTjMOgOSeT5noeBEl/9w+hO2w9vSKuopEbAKbZK21sywLj4l
+t78KEBSGaQ5QeYeJroJDdz9plQnjnoKRAX4XAX5FjhBT1cSVHMQGp7rwh0dostZkTXsIKTsDGpT
t+ZkYnenEbWji59yU3Fs/drBvM6eWtSzXXuwwLfMrUW70Bf7x24zI51mmCPSXoHYganR79RSbWDQ
RT9pPi1K4NPaef75HxWVsEZijuJ1+LtfkjBsLWHbElYH559HpWPLwxk+lJsASYHbhL01PUCn+1yJ
DSPAKeUZn82pJeaCRGVYz/N53QC4PT3dDY+SS894UnJz8ju3jw0w2sivUKUtudyN+sTnMauqqQT0
Y51AIqLosqtdjtBAMD2S97+e+VCeOLyLL2c30QK1knGV8JixBKbzI7HKyYfVw74MBeYLcijeusVr
Qrqom7DYCo/JdxKuVgzfa9BnUOAMihDG9iGP5WPzOOUksTtl01CNiqhuIRGt+Daja0k08YlR5F5/
pIr0GJGQr1Yr882Y3pfLdPl4cnHXzutJwHlhNVC7rmHeO62WugPfgMX9/n9jca5qnYNMTWPGtD2S
HAVAlzKHlYnK82vEQ697MFAYb13hi8GIwJSOz8IanddCKt1qNvUgenPJUI7yB9mYwiN6FPX2HCp/
Stw9U/BsLWq+t5Kkoi+49eBL+UAbxzVkY/VnO/GRL7gljt++QEWaV+1NYjimxyhVp9zBcuCvMiHL
nezvRxVunWO3a5ZFEApg5l621irqCYxzmx1mks03m9cPeJbtcCPatIJpzgDy9p/5mQTOch8zAE9p
x8HidgLhWtoHBgXZvqx71svQJwK3ZW7fE0aOZ7WDmgKwyLA0HDNCkI3nVrHhYiv/3LAs0EJsAh9v
9YI+uI5w8f2kpfrXJJaGLo2A0+gSQSoafs+AreOLh6NcEfCeSy+9MmxRWQ98mezrv+o7yfhmXKiw
qvuLNM/xwwK3g0EMo0JiZ47Oq456L/q6N9J/+7ZgRHYJhTRn07iR92+G0Dw8770ZMFpIdNcJBctJ
w/K79QkXYZTqQYNdSoOevzQ9WE6PmiCkTTyp1VTUboHPnztjDHoAfHPlT5wJ+MhywK2Kgcx3UreY
Z1lfO1DGolxp2tm8DJ5BSIq1yEI74ytJGYwSPfwwjQImUrYYKvxA1JhDnL8IaQevCqawlXYT4Tlx
N+1O4F6C6e0fFZ1hfeTcQmirQuQ2YckiglCSc9yaIu7QMXNxwpLOWxKh/c5xyMqtbD7rkZDcpcCY
z4y244fN2jXbZxRSk7lwYwlD4k92wqd2O9YrFGH00NSfZceFXBjcRnlF1M1eHHeY1T+fcUeochk8
SH8LRpI0GUg/aP9E7laAYOvjvF8zm/EOxtySq7tdjaq40RjnZuppMsDC83fah+B0j+FMbJsBWpuH
7nGy2iVb8fdZtgd5Oz6JwF5t1HsW5L+1XF875C0P0xkfV2mfljsGHA3QGRrxfXDPZnQ/DAY0GrMt
jaqnwS6po2AIEfc8KtjJM2K34LjieuRdW9mNnWQjmXTf9NISqsS4SxsNmJIeuC5nPX0PFAnNDZGq
vuKWtRSE4GbSusFTGI0JfJa98mEJDxhCzqGaJwtHfNkB6IWdibxID776kmEFntRMo8SKTTGBnbWU
XQZ+wKy8/9yg21dxyzQGq6oNDTSoEWqlYBHfc4LRui2KDzvXTIqP2dJkdbuqwV6Zrp+RRxGRP2H3
+0qIq5VbAgE5n1gXKr/c8WGvukShFEUsH3mi3Ng85zObQhMv2aSXyLQmYlwoqwZ1UPrKeJ4AKTRG
sweSHwUS4zwLFtQ6AZ2KcqBQsX6D2OkJ3RMkaZBWBiY9iphExQJ9diP0TGfjM1IPzPWdwlPHCbfi
PlbIWS71jwl3WwMOWXP7Ab6SgZ+nmv88RRCnNw4WFR+lyFkZJh/h6lt1PDTCfYzwE4lQNVaKwElx
PnNIlItJxW9XsT2plXc5Es3GdPOXoCr8ATo2pHmgcphajf6VDUCsKb7nr8uzzluspqI0d397z82j
/H5mg8//An6iOGhaeVeM2S69avrOHodli6jeOfPPZTCaxx0y7PeFJSlVK/i+zqtn4ztw83XBBuT9
1GcB+mBoA2xl4CxPI3gJzP+C93fIyW4GsNumRNnZcFKXH6usJQPEWm2H5+CoFz9SysJj7jcTdE1f
M3pag1WFGA7PEvrr0NYV+PprXIqlcOh6Rr9Lp2eVaOotbbUWxeXnN3WoBlhP70DaGp7bqFiagNlB
2NMiA7OOkcJu+h+cLPfzf+tTWG269197V8Qu6D0JRk6xqLLMzO1CFf3tdbTkR1w0/d/NgUz+EdU4
SuIPGFOka8wGAhxfSBw9fLrNWm5JUIQnX+Z+HBdqnNm8NyVjkEl67DbXs4pXYCvT12gjM9lpMX+E
FTWCdu2VKHH4C6uecjllocl51FkSmXfJsk1EluleU+J54Kw+q7QEZMXF4tVslsnFgdZ8kXBGST1y
1P/IupgfyMwelBB/rebwH1s67CvaiU+JZ/2wzKOS39YpEagdWN90j7Em5nRACsCmsCCzQXC2ksQK
HF5hPN/4MDQ1KgVDwMX9rEifQZ3oz2YJ/MkRZvScvWGtqbBT7DqQwt4pPDaCkc4fFAfGDsnTl0R2
Qk9p5DXT8n000yBcu+gl3xjdR66ChaWauqPM2mHYTw2GNwjkRfcabJv5d2ctht1kTyoUM9XAJJxB
xVgBj5XjkVn60FYlZga8bikvubhAy0k5eap3m4nnRW7W+VRf4yirYwpr0YyN8MsE0ulrcbE2+9D4
16Cm5L1TJ+rXUEQQ1ir5tRCfzLc2gg0KOqTdRW0wUaRLUM8saEnKdhCclb4ltnyIAhY4hQ28PA6a
nK2tfW3yGaqWnt0GiIsDCRbEQfZCyiDvWvhFP1XHtOtXAXIUj91ArGTQaUO6RlBC2xFWKUXpZqau
1FsGZXO8rOMJoUCh24YKCoPv3e6YZFMlkyIVijE9Ju8KFH8UZBL5C4lfeUixFU4VN2N7YPzbKtWs
vrlAyE4dQgKWwAr89LVjWXr+kYNw/AFpODEZmCOctSpK+8g5JnNzCwCT2Ab9TyL3Z0sa0vtrwZnN
nnYScyKjnt4Cgq521hoR2ohLbAg/tpDWiXgwuyRS3fSiCqXrMuqQ13mccF1XUHOhRtvkg5Tkr5kG
teXArZpvShuvTAZu2ttXnUSxbYCCeSI1O4hx1DUtPtlG3h3pu37+r1pKFehdopeqof7ZhIS3IeIV
8cy6S4H4GayqHhBo/flbtdJDbVOG4CFPKqfj24xtrPolfgv6E63W4QmbE93b/pZsOBqY59hR30lB
1srR9YNDXNoJd5uXZKW4UQARbAUdUDvYhcj5QC+W/DwJ6YTPxA30Lquk4rvgfCSc0ydPSTmI3Kzd
nrfnQuaPm1e2uMAd0Whz1HNdUD4grKxaoopMsNfi+5FzSxGfEVhxVKVs6nWUIcuaqyudqybwDRBa
XD/VcmViE3rVedqQ9lf0iDMsmoeR1kTmWxOtmmInqLMEfgfhaIElSkEEuRnsbDPV4HTqpTAtX806
ozft2XcQUuuSegDUOl35iBxe6MXNljzSj2TyQPsYSbPfSItj3fgGQzNfZZj2tyeUis4e0WOvq+/o
Azf9sDkDysDdVLegAvLb75nAjI7d2a6pCW0BlaZczud922aV2b2DZe+YJiSo8D9gKnVB0nM65qKx
IM9ekq60VnphNc4Da8D0bFssa1UhdbzU5n9oxCG5/MrizeXSzSbEFN8ndBU/bFtjY+zEzGsWgD95
hfZxljdKO565dgB+l+HdFlW6FCjDXN0/C7dmMJZ+4f/RB3QBAaxvWZPx6pHpu3tAu0/zTT9jxYQu
dE2XY6CnQUHvu+bi5nY36KcSDYvRjb3OpY5R70anzevaR+JwUW50WKHAvV7wDbwGQ2ATzSUCIcMN
xAHL26F5kWkWujszYyBj4DExp4wxjXa6a5abQPjqc4V+ZNlD5QgwLwzuecCK6VEiCW31WmPC45PJ
t+L5xKvHbSzb7oTBHJWthGaUyH93KrPrgdqhCpdxNGu+izW9yWF9eetJ9qgRpstYNCYPR9q+oafo
9+luHNsYFpMTYvZXqyBDZQsqRJSf+3YtSM89HuK5ZDAy4UaPE3kJE0lB6+pnt0k4PcCPHcB7GHH7
8ulcJBdpIkVmAmlp9cRfNyTn4SfawCfWwoaoFfb86ookPmO1Q0FU/3f4lO9ZM+CIPuFjF4T7j3aT
7guUxWgP7PoVlZJ4f6Dqq9J5kMushJVf9BjmjXgcWpOKC2Er/PgT3+HQSuE1D8nI4Jo9J3qWuWoA
juoDEw1PUyMQXwVpGCgz+g9JcxAttR8cNCh7SKM/vsBqlhWl+PxFKsUhc21RfY2LjMFRA/nP6qw8
k5CO03YgE6WbwWpTW1BB3EpZZ5KqhVbdX+A3lTj5UfkjPp0gxUqeY+T/tghX0DwnQKVakh6BNx0J
WGVNYMiEom0t4mrjOl7dsrXuYyG19X5PenQdQUmyMtJ30aaTWPJlh380NHRHRL5YIsBNDq07OOJ3
U26HxRBnAPSN268PXlmIYiwAhvaiKYfrJ+KNASzMCCxyeFt6IKFvu3J6P7D/Q6G9XVfyrbi0VwBl
1ch2V3rSe+e0IIQLO8jhF3VfeQZr7wbMjXh2ckzmFW3mTQuYSy20qMK5g1l72d23F68jIh7iMY9V
YRbjQCBdGoH0KQM1RL8O5oBsoULq5UIsFggiwaeHjQo9JiJjw7AQaZ8/5vEQUuWubVjgvU8ZejYJ
X2jKt7v9x1H7dt3Ff+fpVQdVI1MkEZWsyZjs8zzXf96PuwrvucXAXkoOWRfgCcI4Dw1qY8nSOkvH
CDm7NFldj+9Tk3l/y9rVUeoKLfnTdtn4kx6jk5dEEhWbMekfOSNCG+zcn5CSciOJSMaTMeuACBcG
zWQiGId0MYEKIiBpSTpD3Pk7fTdQbA0L8P6MH3WeVh3nzE31jQ8E5Q1l84VtO3pwPszX4kxUTaG/
E09jm8pDp0fQ8lIOfHI19e6pmOs8w07TPKZ5IeF480HRXno0z02tBDyDgB/Sz4FgUZ2rL13cvBpJ
o3IfI9ZfTNVuCm8GAMaPNzXaPKDXev6cQqAywwQ0Dt1M91aGEFvWXJwIxKpAzulI0mu2BoPDphsf
jBvk+40NY1YqNLJb7OAIPErjxm8OlayWhMIHLWyP2RvhUFaRvOSLpBn3nAtLxH1pwSkDNOUh5sXe
sH2G33Zf4iiMlyu6YZTiQEofSdeXLLqszAHFziEd4N2PK1iBoMfjhMNn2cg+Cmhg9dprX4sHKL5i
y12NCWFLG/qyZtle3S14ex82PAEcyotwELTt3FGEmfkDJJn5vHJRAYJCs6cp/2soAoQwkiUNRAxx
X5qqja/O2HGmw5rrCO51nl48oSWX1NCD2l78e1oTmo3uSID3Ra7REHkoQsfNrmoGgs1x/0la67Xb
6HB1oWjKRrGFUOX/iTWLu1R6XK8dpKTFnCRbyIw4Agcps7KGqlZKzK2XqzUQgjt7hKopEV8EJ9i9
0ryV4+bQTxFLHnAV5PeqJLiiobqNU16nHZpEmbuZVKHbh5dOmnviRAbVqOJSSFFsc18Tbeyqdu0X
vQ/e0n9pfyOc7Xh3oLCaG1Xia+MAjtnA8sGbaVHpCC71a8vjCSntU/ruifUo6H2qybw/wVlK7NXM
l3ksthzFQW6AagvQjK4y1soVk9Ty4Eu7/xk6Est/Mn+fCu6RjIyclP11uXBgDzKnrIZeZbQ5fvZp
ElcEXaidOVxhzpyTFACspalevlsSWQm1c7PcKa4S0CWmDdaya5/r77iWt1HcypBvPjy15gpE6NNL
fcWzJluhMigq3J4dq0q1hHOL8I1KD0P/oDnh7tONIA5tyGdIJ1XA0/cO/eoUOu3SMolJSpLRR3XY
2VBGpJqshZNV2V2kOjNSXK9B1dJsk+kXt+IVhRARrNYNp4HRcA7UZWzursEZZvvteFjtxENaJQxP
M9Dh0FzAImUlNGwhsjQhLqoOQo4rS4uqz+FpWinN5XXLeCdvVYXScsTQYw2NtI+H6ucbtfN8y5F/
Dvy+2x8QcZ7LyV4AEUDk7DDejr16eDTPUmnpySdbFQwHXDWj+Cg/Px5hnZnxYpdgB2H1ob8g5Jh4
rq8ZiCgvsUE0m6+gxunG+kqrqXi/0HbPTOUTfJsMbYnK5VpyoqgX++SFBRRfDQDnHaYXimnnnmY9
9V0a0xB7lAMkD53eI9ck5NVqESkexOr7RIz0NuKIKrTxGbiDnatPIGHqZKo1hu8xLy1SgYVLWQh6
2+wDShE5rRUf7Vw5C//yBe+oNcpsxRmQgvzwu5tMEzLOLA9BiKZna+fWkGNpP/cyrxrNjDvaDywU
F3fCrk68oKoBnFEnY5QWNR1d/jFn9NRs83a8dFTsYnQ4p15T+ohUQxQB8FuxLCvKQEeQS/oYuoMB
iqM1L/WcWBwtTiSs7fBLd0f+qi4SinFN3qMTs04/LtV81o+T9u6lLiyA9MhcvNPc0OipYz3KHR8u
8bIiuC374jCSYpcvP25X0qVqcws/Utyn/+niO0Wjnq8NnlKk5UKTA/vVd3qbU0ykbPSh3o1bLzMD
h+GpqkVLSLQQdNTRTVLjd6ZWjd5mr1rKUScr4USA2VL3ReC5mCDkUfEpPrCzfGolFqXhsyPaQTw0
+PaWcHfWH74wF+/+e0OznUoeGj6HdtBC8pM/IVwJgIbhUZeZ+YQm5Fa6cHfVIF+98+MiSdH8g8q5
mf+YXVXFs4Okq9LKfPUU2N5Crq4FwTUseEjKhJJAWksaJ6sgtopRNNaY25mOoHzsoBmo6uTHh+mT
NYKQm7OVBFT24MZYPy6CGKDQqmO8SsEgL1EJcglUK7RtJJdGk6c85aLA7VAniX8i+zgzDyqT2YFe
Kjy2QpdRp06f9Frn/8G7eK4XPolEbpeyV65aD00qqdDXKt2xgrhJujZIhazutN5MLGL5y6V7YSI0
IzO7jfghwhcZN2WMUMEyIEKJCndU11GJPRKFxsMiz0SWBVD2xLmAYoxGsG7v14fLYJVmx9GILM+D
YYqTAcNVCo20G+Tni3K1CMyP2djzqCgW66NFC8gdK4be7eEdu6tOkPRIA7LBRA5+HsYX8nBvRRrg
nIbHBznhtFoLUhzxfIJ2UYl65xM9VeEk5AJGi3MuGUHKjH0n+xxPZ/0VZ56reYpVCCigX03VXLst
GVO+BWZmMpWPfTvrVnemLbumZ+HN1QsSHA9sxvPqQdWI5CiiuIbUNkO38790AMH4m9K7RYl5E37Y
kTUnQ1gElJuO0V2DwK93v1CjGC5bCGUcMwcLm7ldKssx0inzLoNuhB/odvY9VC4LU33/bMrYuqDT
CbZH8BLAB+bA2vpRt5aWUzgSWluPhdrVqzlm5ZpRNZbloaE5tzMoHHCbQeHQUKFfs4QsI3w5/A+Z
6tDeOr7PMNe3z9TiRdtqSJuN8kwVWeXZ2ndd+FFBgTKnTvtD8vR10yH9Hfmtt49AWdR5pU29x7nx
Dk1PRNUtdiElRWfzkxDT/3oMfP6giVDwasso5Js9JYIr3E8oTsCd0MJ0ZSFgJv6Ewp93+CJF4b42
/stPkX8HAEQKgymDdps0lyrVyVIn7qpOpC2W0bugJqwA9R3wK5xALQao4vhHPSV0OhXxhY/rTL/+
tZBp1yOFVidcGzLnrhwjpyCBwKC9YuBc1vkHcDjt/ynRSo9Gp5oQnnJzFYJtrO0p6e+P7rAr46Pn
JfWf3MJgasAvanCxO6/HEWQv/2vwPT28HOUy/C27XLO+JJKuTCrUyi4rPhWiYTJtqTTYen5HEBOR
Y4391RddeUnZt0VYKReelnglvw3K0i5rYvrWZggQUs27iVLgSM7qyZ3i/ZsrCg7w8cSk9Oq5dogD
8w/8416JUHXroC3VliawwDxZPTZDoIC4bvsAzEkLq8ywBN+26L+pDwSDOLIKIheOtmqfEaXAdo8E
pbi8000TQb1wldvu7dCd/JJ3wejdPfKzI/JykDIRIDWeICRlfNgl8GmG4xSmfCyJk8V1TK3jgqrP
9WxPS7rY9zoxvFeH5tdiX1hzn2/NDfklMf1EF7BjXEKb99qlFG6yem3R7//OOh4116vJ7FUA+nfr
7SYFs+I1+yL+NC0QI/c4/rqopAe7Qwfc4GucFZ76QH+Lb7TwHmeexhUaQ/JyZA9G4x/oGBh1VnLo
R/4FTvyoESOfO+N6UBWtcjq+R7b9CsmtthDXtfrdBqQ6DwhUEvn4Oo2tQVl36oyUeiiskPK63SQU
0Dxt9sK8KaPW3Ii8kWYxZa7teqqFshlOntGASzyCnV9npx0qFGc3KIfzdvwhW6+F9GgZO3sgvvOM
9vAXnTHyc3Vj8EyFv7+i7wS/E2hn2/731WuLNVFUU0wKn/982GhMAf8M8ytciZpqshmcJZWy6uJo
0iJZw+sTQdfAFLe0s/XHAi93EuuKjyp7PfVTBYwUb2+312sav00KA7Kklgvgo455GVazK950la4x
BCvrY8gNNFaxeC1eAURAI8yxfXBJo8aQUh1QHycaUO85J+56NPSUKNaeLkoBlbXxAo1e9nkZcGWT
DuZrLyR4ccWfJzPo3tU3yFwp70ImSBpupPD0p5S9gxv6eKeAT8tgHjqVs2iDMGkJ/AFNV5ccRE0B
b59bxZy2IaZlsbFrYtB4MooYFNz41Gk+yjjCZhnV732gbs8Xt6oBhIPsYAnx/O2wSR8QTIwIArRb
sjLCu4C7/PTs9jlmPdkqR76vAKLZsWkq3h4NExoIc2CehwXHkzWWGYiiFiIa4gcWRVulG8jNQnCm
BM/yjIXLwfpGnZC19BoUfBQ/YsD3cPKp1gVDwozrDgT3aSeIaeduk3Yc1z1fI8BMgLa+Npt7WVsd
7G5chhbhkjwCsjLWa9kL1AYr6Y3ME0XDv58ixZgCcOcEtzIPk0OHyHgXHj5/9zaiFvRyM1DmTTxK
eAI8QO8RdH5/w7kQtgbA3YbNxuli6cFTEmqwtQfBxozFBoJPG3lQ9YbpApIyCi3yNQHmwhc5FCdQ
7xrkMXNKHB1b4hbiWJZTfqAH33hpkOdn2qTSKC8H0L5NsP3UaXuKtVwerJrdOQ7Jy4Xluc/w3MtM
C5EzTQUhkgoYSbmnPflT1kf0LlZOnbqtv2YFCFaNP14F9IhEjSl7SW0adAj+LNkDkqujr1QJIBBh
a1kFdZPHuHEsHq/dmukfdifiznpLutjUBVgjM/cPLquejERA5oOR1mE9SIiEopGy6660B7+L8f3i
AcWtkdlN0tnOWgCQtko2sGkNDHn0iBQzFbip/s2Kv4bVQvlnBAhn30+PZuEQYl8fCP/UKixPNEPo
hcZAHqNxHWQFjh2zWZO6GT6d+o8N/PXL5zA5auO7HvTznFMugp4U3y+BwFMiKn3R5GDDMSMswFRx
5y597rhJgnejAOp2rReK54NhsHLonJuvt53+i1yIVGbVv+ZhDYanv6NAZ7SCPZ8z2gMWTkMBTnlK
uSCk1eT9W8vQlIKXU++YwaamYKgWfi11sC/t7fDO73ellvWKzL5co0Y4bo1wz2+SPWCpGTPfAaiA
fPLjxLJgFWXEz1RIarYNwbnIbWFZXSPuOYjti+zbpcoJMc6Q4VEnxDJOFcvVQ3d0nfNZa5ZkyIpz
sZDDvs1RrnLC2vVtnBLaTkmvZTVrKkoBb5hu4G2h9CglNhAdS6xWE6D6vj/eo9iu9IflyRXpIg9R
s2/jzFbAbWKV4GIfJVIEmqRX3YNFFVpohHjNWhGNl4c76i9XDAji3pfwwEpKW+GadyaQadW9yFcF
D2uahtT5m65HOJ/ALuvS6p2mEBkefvmpo60vEH0vGkiGxtz+aHPco5OhnvQyK1QMVA+OT9Aq9drZ
Zc6iZYjW+4sTQebnB/f9+puBFxgYlZRzWHupsBHcj6A0Zgbz5vbe72QChSBQrvoiU1RwgPWeUZ8n
HKVrguMKMTlgc7s2ZTarW4Q8o6tjMKEoXHFXInXFBOFJY0xkrtmL/Ye7BdgAru65TaVRTEWoZwzF
+b8p6Au2aImrZrsOgb/AvP9lnWHHSnOMwBhitul9ZGc3xwqAxsiQuPVWVy9HtSMet7WLJ4EsLs9W
v1RrAVup3I4kO6Ap0UqXWgvuUbTVdZoic480HWRrOYq7riAkIv6ZhoRoH0rM10IKLNLTm7DGxdMN
bahhTVDmu/jhFiF0eopzBTiuZqDxb+8GlEraC82Swz5JZ0TbxXcvdhs/YLYSpGl0wpksx3Alp3Ye
nelkU6Zs4PTl+SB+P3PaJjw3w2+6T4HnnDi4ZVyRsemFZF///jW/IaAPRDg1I19wlsYFxabS4ysv
I9m47DIB2cVUaBOCaTze45lcN6B7ZC7zhHxm1VqxLhpzIMNqhXS20cg9/jvVHGxUI44YotDFXu81
s3yJwz56KTvX4a4OYL6vaZp1shcaglQrsVfvfMhiGZfgBuUy2+fe7zRkB855tN42jIcfTEr/ENjn
y4y2xUj1k5M+kZiwZ9CUdyb0GJEkvM13Xod7tvH1iX7WZpj0WUwEBNh2Chc+eDoPSappwCNnr/Cf
xWrNNaA+c+4KmOXk7Tw3zouQ1JvfQOpRvDzSOZigCvPu5HdBbqj45//4NCPo1rsmK5Gv6iRxSXim
ahfZLI4k+HDQqpTvTKnAifWblaNHcAh5Lfs/SGPxSCFlToMXPRoLuactGiaUsMRuu/HizP81bF3c
E24psQB3s7JbBeVTYb1DLu15U9+9PSLqTNjBkyXEnei69d6iKv+w3Dfu1aOhtQGysIIFVC3yx2o6
XAi14T4ogguKY8uIAUPodB92SqZG8KD+6Qldssrfapb2Kn8KXkEdiXngAlX9hzF769RlrptVWv6A
b8hSX9tjZpf4OJ8WLWXougKDW/QZ17IwvFkWCfTblblCoGO8r8RFltC3/dNqF5HFDW1+pGOFev0V
K4jaVwqzBJrbEoP2Z7KZXOiNCi/WlhQJBtAzcsIU9Wh0LgQ4NdJiXYlgXGXpAqcL6uiUxUN4ds/u
TARfooKwNE410wjm3spkNI/AQQ9LeK97+i82OMgrPRKIBQNVEg+asdPISVBVWWsT0IMn3P77MNLB
IEd61VuRAye8Z+vbUHEwONRouX4RE0b4QY/4lWiTQ2u9etawzUq1oOFuSrxCgcLRWvmkO16jU8jW
IC23toGXGpEYH/UBDy7hKXlRw3t21NMqz/I1hgiMX87eNtL1fZhJkTVR9AqZ/8W8hmQXLsKBZup8
1mFR7if28xpF662asE0scdOy1z39hw330WL+M7TYr3UPM1Yn+xu0ufYDCCdaLDDCLd4IREKFT12X
11JO11aSN4GWNb+uhm+8qxrm31VZd6vN5jL5J3NXTBGA76vT8b5AXKLlp8Syv5qsKjfB5R24o16U
ulqZY5jrhfIHHek3XFvgYc45NV9QDx4lYFnnNfwQeS2EHLX9heLSJrGnOLsQpYC3+4l9v07uYFXg
moIs5T542xTaKmE8gk9o0+W1L74uTxvhrdcHWjJBGvSRBByub7MSJcBERgo6yF5F8S5YZaW/31L4
J+NF43IjkTLeHCW6S/dAQubWNQOiDN2YEFICt21Zw5CHdYOP7UOdSeb6zLU8aS8Ki5QR9I1qavAK
vFHKWOQQLpvt00KT+sZFhYWK6dg96mcX70RnVicgcwQuqywue38PB5ESqrZujXb73DWJfqaWbudk
ZKq0OrluZmrvpq0SChVWLC8dy1C9ouyG52VkpvxT2ABTz0HUuYmsok+xsZTa7T5QKxeAFFkexiMG
rMdbkHRY1/Bn/pRgXhOCNhEjvb4D8/bTlV4D/Bv4lrd+sbcMOuVTCTx30wI2Ux93jk4oYautfZOH
79/PvrS/KmgX3KfXxBjn31vd+8Qd/6xRPgm62pO2CVJ+k4R+ZGKuTmPVS/yF0AxQTn7Gj1W5Cb5w
hzJRroYYSbnydru26Qs7XrqG3pOcprlIZktdQ7mv5aBHRXKmO2lmLLyvQfZJJidcdi4OI2jwQzJ3
AtY02YQMpTZGNbThsqRJKM7vo8uVwI6+lyhZtkG10QQ19zP4bu+sO8hUmF0ZXaMRCuuMpLrB1/ZY
jOWJmkwwoyS7WxI78Sg0HGeKYyt9hWNGVpg+51rh7SOm2dThhBvbmikE0E8oVat0YSYfWLD7XSue
ifWbEVOuHngLHL1kCoU2sRzI4MhM/WrC/fWseDvBYCplH24uVAa8zs6ofjMuZdWmS7ZMne3vow1X
duK0fhX/TG09LaYen9B5FY8+hpGeU1UpZ+LYN2T8f6h4cFl/sX6g7xhIHppCI3jbNeiRvjHsIPDZ
kytW66/upTKeFrf4mH2pCi2tRK4+0+7PsBi3RLct6aUkcIABfAQsNphYDBV0NsPmmM3UhkoxfD3f
gEtVyhghvXol0IGJao3IFqp4oRnjE5pIIU/ueMRn4uuDUMMdaSGzP6mBOLf8oY/uqjQu2lYJU8xP
/BNe9cj1mGw4v62HG3+mTFdEcD9kkWgofwsugMP2PZG/jiSfWRot2jjZVRQE8KIG6C2M23zQFcOt
ha5xRPXsycwek2tJkjd6OXRtBZ1DFBRZxPVCccPN/bdKjA2nvlA3DjDmCA85C3Q8/Do+wgid5of3
m9cYsX5N/d2w1MF0JbofhKFWJFskZwktH/9qmjpm0tTq74R4MqFcn1XPlM4Fxc1kfiDAqgCCNv9P
lFqK9QNCxtaEOX8Qynf7FG/S0YeGcP0B70ItMMIQGtTXnrA9YcU8btPtsRxQRDZeZhZ/4Cy7Ys0W
7r9p7N6DKtAa/MvJycEcTY4VLKadfPihIF/FTuv5crGIRNhGwY/7FDa/c88mBHBA567x2zp8VfMp
AMKamgtAR2ybDiEHTzuI/ciBy7o/r3k1CPiyl/lFF4AD69W8jWkyIZM6UsYZx9V5rx8I38aIXFO8
wYm/4rYj6fwHqIE2EiC6ec00aXuGXv8PrnTG+0U8zgiPJjsPLAByzlvkIagCjN/l++MI6rdycgEd
TU8uGh+1zY+h4xh2Q1O7nrJD797bE3WSSmVCbLsAGu5qKPNy05N3QZ8rsQ2dIXyjOQhhrYC+Ao4/
MB6WuXDxgzcBeKhiIU7GzP20+LIBdCSMDVGqZ1u6RlMPLlNbjWgc62FX5AEKDxSVakqjetmPA9HG
GBiusiXprF8LKQlQOo/xjImQNjKZUZTHrlL/ziPd9+XgKAQ77RSx7qO4l699h9/s37pesf17kyCk
Il4wl9hCV3LKXu04BtoY6+6B+LULheFSjWWXOjvX1FO8skl708W3qVICQLsbpQCl3p8VvkKFCeLz
6Vj0hhLifTNoUX3FEiuZtNNVHK6K2fo6R8iLfSuncIREIpIlq58VA+q1IGT85OnpNGBCqjbypX2G
Wjq5OZNL00dq20vub1Vcxmhan0tFpAZXMiKsdpkIX8JyTXYFO1CkvldAKDlUOC9dODrsZq+csZhz
/6WobZ34PeqrnigD86St9zpeB532z6UHQdgU1wrrC7JxKKlEpnGwMr60YTrI4/HTQaN7VptDkErD
tlHZf3hEB25zuTLN8yO2Xum3ohlavKlBog9gMiseTV6gQWdnQLR+CQzZ2/4CFfOvz+aqyGSZTRBD
Kwm5FzzeXzIr4q98J4pUm6fp30w8imimgb1ZnP8GbqRqANeJe8b63+mSyb2mVhbEqFoVWKnxm+KR
BbjHWH4NyjtwJTnK+D72UC29hCICN2/ZROmoRsYjEbgmzdLASb5UWs6fQXuuvVGRTfP6YyptxQcL
GBLZ6WDHNZtba05ulWGj2yG40eQ2LWOMVkd127Hb1PO7VxL28AD93YYkTKAugOS1/+zKK6Qy6KUV
3NQgeHrh0OJ+X50tJuqoKQL0ikgMynv5VQoJbN7KMRc6hOHLDvLPSIo7tbT0H5h5T6PvaVpA77GL
Wzst3Q/+Ey57jw4lquh727o3gT1RXrskFoqkyzEgdKIgdF02odxUe4YaqMI69wy4TcTUjHhKo341
ApDZRDKqmKC1Y9F/+8sFs75cIVz//qh6yxvWjeIT0NExnVSC2vhdfFsrr+dNPr+CmcD7mCaN2wQW
e8V+HVmopXZe1vz19wuLUE6qbFDOSJfuFkqJ98PhBGi0MjyVGoEPYYFch0nKN5ttZkYdk/so/1fd
ChfITNwuHR0YkqPuLcUr13qQ3CrMG0BGxtJIvDSiPGh9VwbEy87f9cplQxmn2cZQlEd7npcM0LQK
E3qXrw1KW2JRAhy8hIBsAx5cD7BnvZqTFN/ThTd20EVT9wg4YEf6Y3B28uJImepav8JVNKnhVSLw
R5iQloQVv3odoEocTpS3Hb6819NCByXqI2Hjpg5bN9zsjya5ROa+mgPo4j758s31y9Ikox0VdWrI
ZWNkj6cwJuf4mvpgFkSqN2L2nAoAcWO9ol6XsO39fnGGUmhAriN5p1dI16tSoObfkF5LpOTezT1p
yd2Q16iaFKFwGSLBvguM8Caa1iWBW9cHLOzbB4ZM3PBysf/QXN8TSlXLEJc2G1h05UhkRMr+QPi0
t48iqq/HFwhdJokMGc/4mU+iao96HwMkiztPpoN81wCvl/U21mCKHoS+bGklT7TpkMVcEHRo/S+a
dfsyEaBVRkEfifchWASLE7jI+cB+uGJijZC+D07jQfwex9wmxUEySWeMUerrdxyTlNkBxPLtpC0o
o7rh516tz3+SDb2vkA60Rierpz3PfDe159NHVf8bJAbVIWo7iNnHMXJur/vTNrPWhtkBjv4+3Ltc
4BBfYXpe6Zay54on+VWWBkjJlPbdcjrVPWS39t3y3zojDy5rPxd7VLXlNrOlET93I75adY+l0M4r
u4XsirEhbKdprdt4MTpbcn/agGwC3WA+Vfo7X9z9WdQB0QonC8QBvpaRCIDx0bK+x9wVyK2PlkP3
ofm9ZbbvQ0ZExydFLdYMx7BOgRbCZ8JHtM0LN1zAf0uVL835UljqfefGyCxTQebbG01KVFR7CLfT
vLtEF04Uls9PNtExN7SZbR0VJqP8AgodaYV5QLiuwVvGKTee0SMkSInDheVzZmnxPZJJtjnvwA0t
5WAInDTLpubIwJWmmu4EFy8DJdY5WAW9y9KTxOqurKnc6NnUUIjbO8oGEEaDruc92lwU/8PVar9F
lcm++BkqcsZuh8fMwl9/BHBjiZtfF2lwHjV+oKDWxjKxJLFwDIXV8gM3zB4EJY++t7ve2a8dfbhe
PszOrJ6RdrWDIWwsZ8wsOc/kX48vUJRq4lNpTUSS6lvM7+stC6UYKLpFqqMEuGV92jP0pCQSVLIM
gFQiFSCoFDqQyXg2Kf3rZmyu+PXh4xzPeULnUhvfOZOa1eNhYI8yoZCrdvydqLKoLG0Fx3dyOQPg
f2122i8lKfigu94pAxwRQe+rLtFgGa6Qtv28SWmB+/+yZ+OSqwoedrUBljSF37AuDQkX8d4VmaP5
VBmtlM9PckKebJy+0A1m+oCFtoyaInUpVvz7ugzKyH8Hg4s9yhZbaQUANfYt8agwQi3fZ/0Z3ufk
Cw129LTxi9RAP3eINLcqVsdIGQw4PxuBWuIxf5I49W9cdV3FYRgwno//FPvjXWnwZ/JHwKpfEUJx
oT216xeBNeNXNaqLGh+5DE2l9FaqgPi0OKlVH4rUKbP8LTNkPIllDV97qFuO9RnIEZsd/CbX8IHa
/KzyPQK9sZzcYJP+eyxec3shue2ixTNc48EjBrHY7IZliFtlG+X47cpvuWDsogTjLQPwXtqNYjss
AGuISUohrAw4RCLuOLJJA5npMKtsnAl5XMdKYpsqsxe85KX8ilExsXCisVKnJqFyd2wDOYTGJhtE
kbVGUCBGDxslseDTrOjxV11sr/dT9ix/UqHdLkIag4XWtw81XD9KDG5e0kJRDaxn1/3aLJXB868e
6tMaLIqyI05TQvpRFscC4mgl65N3s/aDYo2PaANXZjq96K6HgxbaFYwgwSH9MQc6+O7Wj81eLXwN
vL9brlV1vkYwQwt5Ys0GJt/ztlhRbiyU9k8bViGmTIi1tUxcO8yP8PfuiCL5+mWGmtqHKAoY4xPi
H65vNSwfp+jnyACZ8qBcWCfZc6PyqzHkomeAvZemHRvloh5Ids0gMZ4f262UN11N69eJQSOudKxK
0Dzp0URYhkxb0LrNDZC8mlhDmBobcXZBFUqE49Dtg8AAO+aMKwCKwTyoYj/dRL9b4s+qmtsCWPhR
NFLA8uyYRr9mJDpxqptTFCG0CsMSaU2U43mEtTnm8Z5fQwHpJTj4g4zLneeE2rdFVnDeEDRAbMWN
0lup+8Z5fLOLGXbilnWaAwgkFam+aZJOGnB7px4VEPFOkYr4vPDZZhTrLOIA5HWc+csoTy8QWUEB
g5zUkH8wVeW7dmj5UeyjCvil7nVWKCjfKNp0JKIouvCI2FwolQtaWbRh2w0IsfgMkAAyXQelFksc
xYQC66GKwl0fPwm3NL7pqHAksZtGKqw+XPJm8mnTVcoCnduhrin51ogD8oRA1/LlrvQe+j1cYg/l
zzNRrjLZN4actlKR9WMpCldkafyANQQx6yO+4uLuXtx2SkoTyBY00toV0zy6306AyHih5nozKpUs
XeUkqEhpOOzeTIUsaSqpftvKh+lOFpBdtRohEqZaBbWtLdV4phd9DHzgJEWjNjfTZ9Ce3YjmU/3l
AhdmIUsBYfYANMAHqoj2nuewSaAOaaHjin2IMr9lTplLe7yHpP/2pAEDoEZETpodE4UvDfLGh7A8
2O35yEOXQik642pQIVe+oCWIEsMFFzMNDW2P8dYo41Iz/Qc9w3LgnYc7ZQbna29Gnw3jsmbh9q6V
8NXc/me8ms9w+VvViLm+F6GT4qSoWz7Bn1lkkunGujuoWCyvxvJY/ar0XGUaFE/VB8Rz3jYWmiOi
tCwkt1/3EuBui9W136vOcrNXqifoGN6SXFWVAQ47cZzcFgskqJ/K3cPJr34WZDhpQDB+vi8EogxO
up4Q6fhcuZCRwLXZUjWj9yQWnLR3zdF1j4QuMutXVN+dcPZUQQNw7lKQI+YulUnul8RMoT0C0W8k
ks9g+xbwc8XDt2cx01+wOz77IJLwCPUL6glF/PaZvvAY0vnWFF0JkLPoC8E1u6w/WLum2MOanf9a
k9e3NdKioaVpSUmNTuhfbzus7q2jnr5wlWC75lSzOnCrVl6mnkzH/25yP3oqnfAIJF9XANMuJ+Hg
I3y1kCMQcHnQlOZYj+KyKuqR4TwOC8/VonOZVPDjKzRRAltJKtvaZfN+k12Uj1pd1T8OyDZqACjb
Uzq5mRms204VpexNFDTfgo+n1NDUR3d5UqGqKM1XFSDw7GcQVuX6qUjwxSSnHYcBmeJRPOYnQnPK
c7exnVl+SQAy6dYIeA7OQuKBOvhp9/Uxecr51wMUMD3QyfOMkT2KZ+xDQNUUzL1G6WOLRSy73SMx
CHGJvHIijk11mN0yQ/2+4567hCFzpaAhz+IVWLKh8kvmpewvELNyBHleCn6Yoqq45pFTL9HMKa2K
TjYAW1IELinlVebwJmidHQf+IFACo5TU3GW9LbI1Slp07+8ZrFedy2phxudosQbPVZFoKkei9LWQ
W+TRwJz9mnNP0ey72E4r3q7vcYDH0ZGzmvmT5zj72rzbweiaPsNBWhWAgpu1Q/xWbtNKCAF6zc2E
B7KtQ6uPBRa8xQjuXMwVxUlmDck4X3y632pdKSZQuRNNK6y98zdB7FNqv9flxsT63eAKoGZ5GHmO
tlvabIWYu2qh0zat4GAFsxd7a3fvQiuRqzD5ZORGujhdvkRfBiJSlv3UGJfYJIQoC3yxgkFeoYBY
UN+4TXsgfBm6+fAy+WAWYK9ZrkpSiTNvMCIKrFvuWaO4KbTO1P64xL71ckrB0VN7Kb1g57LF0Wqn
yAyh5gOw/kfv7hDxzHXk12MAhhVWS1bxbx8YTGnVNTUnRAA2Q8n9BF4xwaPnHNW+PSrmwpMJAKTA
dZNBCwScdhd1usG7yZcf9U0C57TYSM/tRa83D0oUtRhgTcdZZCGSYPpqO2HCFqRMHcln7VaABSFa
8l4lCukODAtgZVKvkBG30SgmzmgHvIUvmeSBo/bQ76nq1pSeQ2/T7yO70YOq/vfjZ7u274rzBC0z
MDr+jKXSmUlIyIhMCGmuL5MmX6Ed7gkp/wijzz9rV0/JRsRBMHi36WAEOPl2ewVGIleA3j+qb7RZ
7duDDfMoTsK9FfxtoIJ+3sNa/L5GmuChtPRDzHknbKYchmUOmcZdl/B4/vN6fKo2z8jZHauj0NKh
CORxS+JJXWm3hzF/KPwXMXTfpnWOg5EcFsK6EGMFCbXk8ZMnNyl8jHZCzAcBdxvR3AJRQzbjl1xi
kF6OZNOMamnnuz2rUTSJXYqDB///9FyqcLX0t1KcU7vKk+T/z2TacEYIIyrI+cXb7jaRjVPMcScN
tuxp2b9v30Ssik1YxYQHPfZliL4h9s5vtBNcggkQEXpt4LxEUfl+ujQGPpEFcNBhrVCGbrXhJsoG
y03hFndvzbKfpbKKcDDoDhiMOMyySU9ESwr3pCv6MKHQjrS7l/c9hBkvHTggg1KlDzv+6uxYKJ6Z
HyMFD87+U2nkAndHr+a+RH84QGEVpybyw/v9Ih1oI/qD9elv112hQoMQOCoP+yilWSeQeCR9uYwE
M8DZlcIDdBafHYL39OUv5XkehaSGdXu2z+Coi5/1JOgtxRV2C6f/BxbPh7IReGiMywLl3bTfwBjt
ARP9gV2649yN+So/OwVuBlKTeQiqHcIxlZtqbH9N/iVJWLtRSObh+VMEY1oUguvI3cCGL+xCXh6u
3YVebFbjk3+0+ZLoq+HH89U17PQJX9jaAb95NTaBmFOXHOiFqrZPS1BjqzPI+GnX2FsH1gEU0frx
vMhn2jXlCOjke4zRE1Jxe+gVrmYoTWfoYU4HcjSPGbstZjSfLujl4taMRPCxpJcGNr6svo2HYdDo
JRYhsW45g/YaNCo22UPRvFYdwEFfwIU4r+9f8GoOrn5BEpCMXTiaEIysWT/l6z8edjVDWfg0r3sb
eBftLDWb5ee/BFjqVSFUnKyHQTc/H1+4pvFYFKOHklp4o3sy8GEd4Ox92gLGFvAX1RiE1aauPU+a
ziLVd4+DBDWdOepdq29CblTJ+UpUI7VEaJD+vgabZiqJdRzF8KRBxZJ3vL7KNNpIkjWt/QXOajR3
4fT6mZY1x4iGuv4Lv5aes2jdzOCX386rgCQnVM7rGbuUdcOn6560eeQ08FNGlGibfHyH16XYLkVs
hdASoRUlJdP7tBmDJxaFRciX8EYHkKFx1YdDegA9ACWOF7GvB+64foht3UccIDM9VX/SBrADyt2x
PbtFr8ThOGFpzoOlf8c9hrJ8QFEgyV+wsWzEiwde/dMZQu0YFOlcfOrmFxAx4CEhis2+UOSfrsLo
QfWiERH6a57uA8hb5i6/o0DdlSkZWilzVRgL7OCCvzSlkP3cTUtY7iTcH0sLzvAg0h/qhQrA8aOX
Ne3ujW4LODrTJPnbdZK8K2ZGjPEis1cah4UnPQT6oyxW1d7lPJzCdAYEkdIGU7vO/6XOVPHdl8Oz
1KD/bT0kxsoUvHo0wiAgzepQOjWzisIQAmo+xZsR0hh3gVj0huvy7CLqIORDDikMCugcppzQyHC6
Lub1EWWSfnwVrG78CYlECTT7YTD9Igi6kp7nc8zCKYHRna8p7guIcFupp5rksOjxgIVFmlpPhWJx
7DzUQanFPpEM1OpI4h4Phlndf+tdApswoR8xWu8lYwIN9obsyhnPH/Ly4tf1+NS8fi88qdOF7eFF
PuwHTShQVxGqvV79dJyuBmnhb9ImLGnI2mgr2oTIWmq/T8ocrnA+chRBBoB/aszUV/cluEpmUHD9
CXXgH3hSRI9+CDmhzYDKSYUxQACTzKmByo5dvk96wsZoarViz/toWHndFDaSRAsXE8FchDGtxt44
xBRGiDwv3KVpaJpMIy9pYd4CV9NQKX9TbMDHWiaseXTlzM0bjhk1A2H6GsYIj0Lv5BBg1cjuIXG9
JQgV1Arwue64Ot0PxSaEBebtWxnCr1EehyCGEoW+XfwMuctbBysqQy9YTeMeu+ybNY0IiKeo2wt8
RNUMT6jorWJegZhTKqXLD2MITBGZN6fjEIUTmAj8qnrqUzlxp2H81O/dqzA24nNwiL9f1aDJAO7k
6Bvy+/u30z5flG5fR18xfzYlvFXR3U7hL9JXeiMoyL0gfy2VmzJxgqrJZb8OuXIsO+UykjmZGo92
nDNa/n13wI1rY7t0nepHlTL7DGIf/+us7u4qjCHryBD1bcvSKDZo1KCPWqcLebFvnC9FtigV5wAF
ULVHpxAsDB5Z6VVdeUAQaqPySyLxEtfiHSgnLsCbDuUPwAR98z0sSaxRgKJe3vgzv8HF6EpPMuE9
oAKSnlyrhymoXtpCS8w4FqeBT2jnnDktYD6IT009cDpuhvPfX8f7CbTLW1ctu5ao8wFZ0p0Up4av
jsk7LnQVBnQNm0wPUNc8rSgWOiSmVs3REkrbOc69IiNcY/yzwyky2UnaJAddVRDX1iUHkKWVnJjR
lxd1BOUAQjLlkFZjluuXJx8k+ternXVChRuFHJHIC2U3ZzUCMoNBaRkuqCDpoZtVLq2Ir4aGH93v
wfuWCo7qUNdz1HfMWRJUionGQiX8J97Ec2XSvs0O5HIKzrDcXwuqgZEyp0HBBSSA+AKTlDbgURSc
SToFxGlhS6u9ypimz4KpZi+NyCDTAv2SLbER5FYFvX9zQMG/d1xmw2AicDN3dgyOmt7KyskQA8Ve
iafK2OEKQCB/pU3C8e1kGPoZSizrKv0gut/18GH6S00VPvpCJE9Y73DP+40p5XS+SL6A+jhxemYo
4LUz0fOkDmEF/YKhEY8O0w+ta6u6b7Q/Tu8cw7zyalo1L9/HcMawRy3Qf8ts+22N8//z4eyJ2YgT
bixDHOlslZAyWWZdqRzBWm7G4lDLCOISM5V9UPoAOvNFy2qBzi0qcryI6+ZfMyuAaq9MxDz/FJZD
SqfM8ePFEFDhcn4f57zv6gVS23IXRWuYGZbJ6OhKABqAwSbYG/cPMhjLdpJocFPVuzAZSlrmDDpt
CZdl56hLoFUHaAZNBZXU+ajMcMV6mZtTBaesfWI95uiAG3f25xpmeHhcbDP9sZyjvYVhHXksASfE
gMolSbHY+7Yp1/cGJhTo7w45AQVnW5prCjsaCv5/jVd9Br6etNYXBp1kN8N7lMNTfxIicrzc4tiH
7Hj+O10d5seDswUlFypmWLmYRRq81cBlIWOC0VfQQzXqxX9GR/0bsPZ/UpTNd2D35MSlWHBuQ7TZ
pbGYjXwOh1e0RgK0WL5VwYs00NESkT8eyJXLnf/z+UZAYAMluKXhA4v4UFBFDaeF2vrMuakQQMuz
O43GtI6HyX7N3mQiTGF2XCxrkKHeYZ24GrIvQMwvmPuzg1S7HnhNAwwuwFRGccLk0xoAdSe6iNSI
EoAiaEs1F9D/xBJcxQkxnXgbuf2OnumtbOL2t3vn5dTEJx+OnVq0Q1A+wtVpleWzVcWOW2urYyX0
OO9CuPy3jIdkrpVoXmd2ek24B7jmn1EKjwqO2V2idHmU8VGXglvF45N0gJM0BrDZlrPdL+kWhN0g
9fD7dvPUGVrduWRI03UL3Rk+SxRsGm9jbSVSgz5fXwLJ4odXV5qWWqOiXwn2NR194b1q74MBHUF4
Ube1KANzemJZbBFNPkXSZtU+rnROXFXp3qRDJcFGVFMzxwDiMUdyaqLm+FWAvudDbeJ6UOoiqlts
MCPzbtbxr2Uk/Cqrzzk6L7hYv4lApqLZwG9jt5wyVHRMHvnNZb9W27S9oLKnTWNh3o0V0o/5H7Q6
HkCt/2C45qqw1w3tbbo6G7p//MCX4msNGu6AC/y/BduDANLC29G8HNsKAldQOp217WuXbiCTnR7D
U5lo7ySg08jgcU13n5QFmWWSwAxPchwZMy2Co1GrXgwtYmFGNRmc63bTBkoRSJahcRG1M4K6pE6y
iMM+mF7vUCO9aN7UzId0XnXtfNOWyE2YPd5rT8453ODZXD8cdlHdhNau0uRoGOheX+vxOXG7fWgy
h9ME2vcQWnWtpMoBCW8fl9rKfkhOmuqM4D0mMPTsL+wkH4vt8fhTEKrFI9MPKunohNxtd5IV3nZE
ygEotxp75irglNz5HhB8vrCXWitWoKvPBA4aAiYMT0SWJmP3jhCItD6CnDqfvKx6joZqAQj/BpJq
YwK8ExLxmmU17a61lUu5TkwQ9JAzeO59oU9BGw6qSPglnHUBC//o4ic+1TtuLry1Ey0/dIiCoT+B
yjOcMV6YADsRwv0t8p6QQr8m7Zef85XyhRU/GEM76EnGjLyBxIxTuyyzWMV9xHnAPwcEpL00EMXQ
0RQoYC4efQKUzSUbaQEGCNiOW5fcBTgFuY3HN9DpdG15EkwpChoIvYnbvXHA+QC+ZW5z6FLaa/1Z
OLyufzWjhlFOBF6xCJfXCnN0hIyWeNx79nKBNDTRrGl/uyDQYxT9jFX7yvQsG0xl7XUr5Ic9GmA9
uRbJKIxkEBoJjoZNgmGgF8XYbdFhYdNHpJB60cRCvmERdDlhTQKljItXFBG6xPd4UDF3f6/XORMc
luUt0P68Y2uQDhz+VUQcxFnaU/2McEA/yBg0cyGWSjPAOB1SfKh4w+LJlJLkDwu7en8dP27S3DYd
QLnheMKE50kEDmf3oosrvC+rpdOTi1yV7M7JIWLHQcSZVAls24WImvRHkiwsKx/01mdCo2+rIGuq
DfkJy2YqwuWDM7SDaxTLd8P7rdoYUHkRqin5Z5UtyNmpoXjG81BJ0rdldpkIWzijl28I4mMi8ezn
l1e84zj5g8gCwMtovdfVKHaEWmwj3x7WzEEFZ1uQPBmf/a6E/nGQryWY3rQTto/u+S7OzrfeghVR
niYBb/wv1hgJYCbTwXv3cKJe/r+vwwS6L1ePsYQT/rdLSyLetytqKgZt9mWkSnoDUY6QT28RwbI+
D5rK6VCiSNRGuTA4la+xVg5rIBd3deXNNgS7CT+1MfPvA8rn0x4MDEgxOyKFIyO1eIrXnAtTlH/K
RmowMwxogye0X9OiWidgblMta5yjUlwRDSL8EDaKiP7H7WJvQwxoOvJbsh4z6DcgLEtxK6bZcpPI
tlYt7+D9jy8xbbBFM39aCt64oB6I6X4TAJesTK/Bn09RRIrSFzgHf5xEpI9UUu+mw3m634H/45N4
zjpo1qZY7h+0L5VPgHcTudvj1qOP8URFxre8ys03+wPfCLpqCHw7blb2Ws1SVRnvYxA3HBKf1jca
rUqnXoRLpvchfB+MlzemklymxxxZsearA/davQI1EQF6oSlcNgu5YSku3g81V/JXZjo58ytlZoIn
QvmVBMw4eKmsHoMJcAMR/JLPglefNy4htSDjmbdGFXqwr73f8tuB31c+42ZM2FgjvyX4IAzDrg11
Y88Ey9zwajMTIySKC3r3XD4FyAJkbt4JvVeG5/jfds95y5cZKfBfxUSPdLlnWnZCvQOX5nqWvFBC
oJUfaVoZSzWi7YOZKs9CprYgF2mBTiQhNRnCVWASKgWcY5NOXuH8uuuT9w1GavFsTqGNB2Z+gbns
sibVlSl7Cl4j1Nem893gdcog9Ojzy3/SQmOAFaGgd2m4BRE2jMG3c6PT2KyFnDKhZsLD7cYD2HoR
8WaSK0GrFoROJ5M6yVujyNPBgmwMsiKi9Sq+wqEReqffny7pxC6tjm/oiIZ7HFVfAr/beeD+xtTx
MKI6oXZSz1qip7OBnyGTHppxKR9f/luuja2uRPb/6TuNl2vp0f6Xhul3wdctsfR45eMk0SblP6RN
iFoGN7lFJRKi2TGQeMAYRVVSyR8gB6muKeX41L3YiESfS/6CSwfDusD2aT+AA91UyChTnpKzTBYp
UDeb2kr9DsaTbeHTpl1xBMNiPKrTcfXO/EC1wVKCOMwCaW865WbEoFFv0G1MGGeOE4hnM0lZFT9E
Dyxk+HFJTsjv6eNXExfoWhnyohQLf7rIztamxY1ObbeWDaJnXQNnkuZ7w0iDGe26u4D3YXwRsb6N
MwFcl83XMv/umPX52iy5VXd9K4w4GhorIYnHzqHKNRnQxKuXTkRvCDdimPzHAqKrADqntdgQGssD
1B5kumdWWa5dyPOGsw+M3PiXApuk9C6G0NAXjP/CTPqynor+gd/R3BNU2wGHPy5g8D6Jyu3H68jV
vUB6w8Xgi+b++vAwWmdfdteHt21w43Xnzvod9F0ZQm3RaDTmE7sI+S6f/W/Jwj5iqi2eWCyh/bza
yLAyxHTagFhntfsr0grgVgXHJ9aWHJxa2VYNBzrBjoMOIiCTd13oEbTzatAutPe8HHpQ4GKIPG9O
IhrUjkHak9PV7rW3JdNiWvxnMsfYCTYCnnhumuIei4KvtIlJlUD8hOGFC+kqJrwziNVU7ts+8wvQ
tx9xWiT8qWdLbpY/4+gFOWvWYBEJff7H8cdf+dI1QHP/LU0AzUWva9AU03zo2+NPkuHTGwfo3dgo
geI2dpKfsjvE3DE28EEPjMGFiki94sqL5+rC0XTl/+IeFmMQe/xRgM23yJ5IXbmmhR84kWJ7rgvv
Y5woiJ7xvF50OnUU8GKl8xMMaME3fOv86czMmrHpHIb8h59KEWJnRMzDcvpenuRMRdzZUfCFLAjf
LID22dv+CelwStVezKbuewGUVcBesFPaeHisg2yFA0MFNd4z36K+iaI8OaB7DlmRdzv1Sx5dRUGH
wmvgo3J2sCvSdlPMu4B3S/1dYITuAHg8kINxMOwd9SCzZHO1brDEMr2wbS3/k+ziZKzbY6hNLqj9
wUQRDkJN0Vzphk0nzsJFZuLijER9BNG2+vrLpV/q6UN/5gNRbrjDPEpr7DKtuLm7yccGzJyb7dpC
+wuzej+nwaqhvsHSaDO5VuMRhcZT0LURrM1w2XxcV3D5jTYf08vWj+6aaGk+Jo9IcVxTZq2AUHJ8
ByLfNrUi4NTxQjL+3+7Ylm1QSWsmc5jNnksFuwJN4/z4Zea9IX/lRtDJkpFOQ/munZZzIIu9H7KJ
gw5EZGyj+bgYl6u37FBTXHX66XT1eoDFau1jX95pGiJKdiMc6qSQ3PkLFMYO5z6bL7NlslzLI7wu
K67ScR2D9ZE975MXbLLS0aGl17QT0g0ezcA7MI96KdhRTgwxFv+dFNSl9MYzbXdQEdHPMKjUVBNY
HyWbvne8QbX9ThJG5WSh+B9wwKD8yDO2eYcGqNFLXts0kx2FN3bGAuZOhRmAxAqhuqxs8LaK0UjT
0H77P9uN6qOmJyFIVPCM9YaQTIndMnRt1sbwHm1Z4xpEOrpAQseP0A6SzO3BIDuesdR5pg/JkI55
KGfxhlLcDx1BfUGsWvZGNmmrL5KHtHsc8a62VTbnz5+Mxn/CSbBOYGjxvdrvmm5UT2xOqOxEUccJ
s1tDbZ1iARtDm2e1mR62o5yMleQ0jQKr3m4FboRwKYgHZFEHQee1v2OJthoopWaz0mm1NxAXVKxk
C1chr0hZAsfRi0Kq+dp1xY8vO5buqbJGxfs0Hfdx3tTBaloHVN3g9UVCDqL1fAmfclK8Yr7AanRh
Ou/clSgayaNuyZQvLyFOEhCF3KdEKqRgCpGdOrTq2IrdLkYN4gu11ZFHcOQKSngIg/J4/rGhYg5u
aOaLNY0PpPeMYytDf/sTmXmvVSEqrnQ0Lh2IejNqD28IC4kHfKuNJogJCebXn3l8tTanTbTXJ/a9
7iUIg8rVwS9Y+tFroF6tPTLRsQBYyI7t4uQ2v5Cpr5YgTiin0U/NRhJ8/HNPn8QiRhacNg6vHWEB
1XII0opb6OhY2vRURYgCCy+RwtsjwDBrUMIjvzHq4ZcTf8RvXr2jErkrNXSQuqPgk58bwt2K2FpC
pWUyJG5QLN/dVaYutn9dUumS9+R9eDf1v8P25EPVzFGDMBiiA+vvCm8gwPK872t0Gdtw+k9SU80X
2KkSCbpDU/B9YQpKD4Q2cYU+6hxe6iyAfdH0MiW/aAQCOd7EWGXFCmkVAcplVNB6MQRqEC36W0TT
mBjx3IP2xCTkrQRshYzowxdNAXNuZg6L/AtLJsja581/8tlPcpZhpwrYguxITqhalqJICYZ6Doj3
40rrAbtsnBh8rW3sx+AScjcfPTPrEXOWglBSijulwrBYNMZhOY7nAqovh0EZ7j4HR/WPsGmAzTGb
LBosy78p/HquLFOEja3JVcuqHcDybZE/N//YtIMqbyDyVYPcgZHyvJVcC6f7NspBmqwKWWc25btz
jVhXgu8vI9+JikLrABXEausnmhqwFGBUol24/M0p3ISRv7amy2tA1oVXPFvWiHJ356m9W/hLLwHY
lg5VP0KPXbEoVQ9J4JbXmkYvF/fyFI9QzFiu2XmaEEhavEKWJGbH0YZ/nsNmM6tPuo3JaBFDdIac
TzDK+GalCyEdSMa7LR5DisUxlicXOYFNlNNtF3tBi2W5s5zd656qclOUbGtynzc8wNbx0kUxowTX
hguk82MpIUeGp69EmSdBQQTeeUZM2vgXoTFguYtf8fjCeDGUPawT651RRxE+hA11C97YEOtbcrCb
Flc48P0UH2GZIMKBFkTJHeTJ0ESFsi/uWkdMPQc5xAa8gXLKoLhtIIu3uk0XNF+RUAZgC88qONQ4
xlAKW1Eex/9MI14haE3gZYIsPuKMMKlsdlEVS3N8bQ6Z3egOEE3mZQ+TK8/wUxQi5ca2TrENLpUK
iKSSpHkOt4c/1yDXBGnu6ofplguSnv5727AMrDjOKCiK7UPWEUNhT4dIo/P3gkuTuuqiN86q0mhm
xAgcvNo+qps1bPTJBYwzBRrKxYW0OMtH+2onAZbkKI7cJJQvTejwwVJiy4353y9kDf3Lo8QSiNL5
oFGg5cfMKrit3lVrNNYLiXJbKJzisck8UuxSUAcbnspVZyujO2DJyMy/yYYC42hFoBVjm0QC+u37
oDJ2mn8/QpNMEt+xpFpHeKnJ4tdcVYTgpfmVCJ+q4ccOo7YarwxkRs5grtyLEDD7ItQ2W6TV3EHU
N7fA44bPZB2aEiW+WXURPDaX2L83fU5plqa3pxb+7IWGne52xb1WX7nNH9HTuP2sFR18Smu0YUu9
V1ehQAaJZeSxRagRkJvRucnD8ibIpIf+pp7An7dPqf5erpkmve5AhIVpNM0jCSgoXXCgt1n9n0j+
ZCkxacWXnI/Yykjoyz/rSDj7IheCmS74MCLi/ELywunujGRyLe7R1GUGyfiN1rJmwIoGufgQZcXW
Xktl5SMnBhl6NQha5g9b5ZnluARDnzgUxyP5fbolxYIc+5E4/tgBeAz91N3PxEgHyBv/hsp6cmV1
IJ0EOl0H+tx5pGVenNZnmJztwzAlyJs7Jurtk3+dKpvd/sKShqf/zvjKnwBY87OOEGcSTe4LNxR4
2lZj+INfLRL/WzKPXYpsIiMQM0HSyFn055K/cH11WHo5QBIXVv6D+bAEYnfXN0ACVKpFafdQs4LG
EBA9hWs64XTEekdVwXm4iWpuWDZvD5JfLtgx7oYRe9vIU/Jo+oRjeDIXrvEkpKRkMdQOOx5lCB6/
aPO5GGS0igXSLDDll+nTkuQs3jCDw2ggMRB/KiDJok33cH3nGap4jOcMHeDUUg90jbZeuOQNvjRs
EjiXYDneOrlqH5dhJh81XQfeK4iol60olj5QutW0QhNdxPKRfCFeUoNOKgf4q/Gi6Q779kI3NuK1
QfZ4VmgefOHhvl47AmlqNUhNKqlryo11R7jNr5+EHS1ouraWEZwCSmbDFCjX96JK2jhC2sN0TFjv
hxDIGlUTnoDGA78vsDv2PfBg0Q3W3hyJxSFaRG/6ZZWrDVd2lpyqf/B6V/d3zPwDppe7PI3UW0eH
AmrSP/kKV29OYNfeSyBIiKhR+2DODP2SDT7J+YkvgDLS6RMfEbqMLLns855kz+uB5bJL5S7ry2Bo
7WMXjgJ122aGt7v6lmkaMitPUku37WRs0jGJAWcTqavHy/z0hwap7TMiRAeRdIjpWBhk/Ay5IXib
+Mbgm845X6YpcmIfb67gTwTGD1O+e6JKmowaTQ1+HrEG/cj51vVEDwp055h085GQtzQYnuCIprIY
pC+siI1d57KenBpy0d1UtM5Pos8Ej3g+uP0aL9n6BdxHz93O8AlenWneLz2HxvQuTak6mlMtbOBa
ypGvaN73EHIt0r95yicl3aaxl4BzE+84UoEWy+8Ya1PaIJI4XU76u4uBFvRgDFHnUGuQFlu3W6u7
V39XYbmwQG/I+dwvzUgtCtvBoE0AFc28Q1wwluDJFckOG0OQtKePElFFbobmp4lxRzXd0VJEVhMf
m51ZSalIVOGp4WcNt4c7UNJzTgsuHOxn8KTRAWwUg3EO8/pJ/n/WUUWREQ6gL5ObaSxg7d0C2uPk
xP2tLFx7K+ydQ7vt1aHCjJj/ilZWc+7CdJBr3KPK5cIE/6Go6SKpjCfLG6DeAP3DTkYf8CsWORbo
c5qgoApY9jYDvwHllYOD5sLmPMnnzFrB6NvRrr/KoFDEDCFmPaFUtyzXDzEWCYP70Mv6jOf8HoN0
1IcCa+YzoGJegW6j/tYJc7wRHBOBeTb4XokzTMg2oQpKILi0wOYkONyAZ9hsjeBAjZLUL8BljL/z
6ZmYudzlBk2fvQR3/PE+PfhESRBTu7plXIBPczeHnaKJASRfVb3krzpoCkxPc2TUhBvwrvVGEBIX
a5F1wmDkvA7IqWe1+zoAyPlHq7UjloOJ2ajsLVi9PaYuTo6aZH5sbAyueFidPYFqT/4GNxSf8c9n
VbNKyg3oKSGzg0eurWm+qt7SrhZDFC5XOqz/6r9OoljbN64xYA1A3yqbfYlngXS4CnZAH/FAVoNA
O0KH/QuWs05OQl9TqFyQyDA496oZMaU6AObJSo32AZ77Qizp1c6B2XLSyfRS2kbhN+1ffaz4/+ml
CDvvJDBaCYvTMmSyjggVM4PKNJoahWmZhSbgYPqEi0qa0PhfAQbh7qGr/AAnTtSqi4jDf61kZ9bp
jEWDk6EE1SqeGQ44qFPCFzbz6ZkfXkLvf5bJ7Sd4p0DGzs2vCge/FBe1WFTtIGYafdMJGMQMF7YS
e/zh76H00Czchm9to40AznX2HPwn+qFMqQ4G5QaxVAywEe24efhOrfP1XL0PGXBMVg37WPr/9qlo
h3pNmh6L3Q+23SEMTb9T9ZbkLg2n9Pnn9lO6KdFlVUtR01y/n0kWS1wu95DixD7+x4iqst+AEONv
cmT/Ki6EQqsnGE9b3q6Yr+xVyS8j7RyEfw/TsiSv7p79DX9lrJrZivxbutnQ1rkhVshy3c8VAPxW
XVDpYmMrCkU5cnRgtKPAEwstN/DTay66IZvE8soCVuFXxuBQNMZNq/G9haFMFN/kiJvYIytxNa+n
fRrZlxbS7Mljrdo5oXFzvOSPLgyHvL2+QOC5Lc5vUys0/Gv9PTXoApP2lDQ0WwdleUVM3JQgfmux
W7pNDMCcqeCWp+LElIMYmGTZNZPnpnTdrbw+aou3IC6wLmCNOZb/0idxsaXYqvQFKk7O4647YSsC
JvYSrDcApiBGjJlVEplJyWUGJr70Phr5TsaCUYexhbca5bLBnN09rKOOEk8uN5tp558HDmxdZydA
8GAOUyNemw8hfpbmE1nCKaBXk8BQc8GqbnDJxGxCdk2P1uKCRKdJzRJ7eP2jX6xnCm94CT546KDJ
WlPV697DzDfutVP1MKPQ+5MF12ub+AuhzyQqwLD5mEp+5A8GW6p5incmwsOFD1D36WgbYEZkYgrW
9+unSLvpueukJJpqKjkNs/BXKNUJTJ0kdxMdAs9CEGO1ZJ5Xr7D2s/73KgzDUw7xG5A7N5hreTW5
nq9QLEwQ+knOvWxPkjHRFbRHYm1s8c5uG4qqpJjdtMuBAnG7IVpyKDOVeN8i7gOEZpXkaRoQufjM
Xm8Sf7dTp7ggRQjknP99oeLDsASlIIAXnlk7kp/o53/ykM0e28gK2dHXgTUKmrGT7vPxfUDrzJJO
ktMyra1ZsmIOdAXbstuKWz2Qq4rOiIUXshoiuZCT7pC1D6zL+j41Ip+Mh3mzZOxiETs5IZ8Xx0Ck
n/zlE3tlr+Tzw3A17PjDGZvtzNM6nNLhaWuzQCcp1QiEULv4nzIsSre92ds3EEFu8zxkeC6DQwOk
zX1F/VVD3rqvsilUOTRtykDyIhbkKl3lBTcGG8GuLs0aMPK2j1DjzMDYDFhrYDGILE5+g8ybv5C7
dXeDuohUIEi2RCauTTVfmtdL5Dxv+5bqRakeeZZb9SnKxQOTfudrq0o0jlRM9CRRhIciWkS3Psk4
4CGZZlOYIjkPT9Tpz/7G5P2DGYgtxqgi4nmXr6DSmDWVjmDtOC0V/g04+REDlnTkkQfZazVHKO7z
osb7pyvg58twbG1vSAWRWqlxebwgDpqDqZKwt97nrxBpn44qMQEqsKHWg5ZKeECUgpHTUf0A9pkE
JGje4eUqoq7PsifvNxDy31kVaE8GvFKXhm/+lxJvrx6Krt4eagzsdakgS6hagJshhuFlNDjxP5P3
2Wtw96UjgHzUnKYnOiTpKJqPcjg1LV57q/yNhHooosClF+Q2OskDEw4bdWZqFp208B5kx9ahLOzf
BQ0p9wQc/hEnIZf6HN8MMz8qfO3Cp8UNhS7QJIJpGI8I8uGdnv6LfIbJyAlCuYV06hDag+adjplc
wYtsL9kGCDdU6CCB4lRSFqldML5IlzDPm7h4VN5X4xvTnMnYbwD+y7r8NRtt7VUI5DwFb410jEBk
Almm87IkZk1OpgE7pzb3OhIKcHaHIutmrzEhaaKW7Zurkzll+sumtYMKv/g4PYc/kUVf0/FSE2Jc
wUivUEqa9UF7FK0ip6wbiwjIShZGkbPBp+Cq+SkJlnmjG1fHOHEx3Em4vUhmlhZuIp05n5RoayTo
gRgHEzljqtByrS0QJwwfee3o56oWjE9GCup+HBK1hIxXfoO2U5PI8NpOKdis5aeD9r8mjN0IjMMp
sVPwbvl2P7nVLZzNtEDLO4QdwsWRTDOPfJ5LRklFZegrU0g7mjW0Suj3EpDyqM21d0cAf988FzEH
6luRZ1rr7MleR4pibWLW7aX+PQGv/WvbMz/I/Uo0EIM1SQdFXGS/Dz8B+PS6PHZvJIVH8Q2AMxeS
Tsrcpu5iQKaIKaTol6bNPKt5Avxhb6ewN3wKEUdu56OTYv/y1txbbpJHK4Do7KI4Z3VxqMq5CvDM
eKU9fnICfZJUf5zfs9M9aCp/miifqWbwqGFLSajVrUM31AkLaWT5Xud8B5TViB8WLUfCSEEt6QfY
ogVSPBLCSZt1jO8EkQ+5a89uvoJcR6MHyaIFAmgesJwWi6zBWjheOIWD4X5qDWaTA8YlT+Z35/rb
r0iHuUdqymHHqAeDQkncTLy1y/pGM2iovBUn/ovMmwuatdw9KbcitfJ19b4kK7TZD6xVc8Mi341f
uXQ+akK55hU2X3vtsQqDSau49U9zN8oLc9S0z1tkRNv0ER+YlRJMzSWTo1DCUhnxUE8mlD+dpqA4
vZ6SJNh7WGL3eK/vdIgjTbGIOuGi0cwvp8LRI9MgD33/WFs0JCl/xed+RwEHZIo33VxCnvHyTeHv
/a9pKm96oBEhUk/KAK4bTjvI55/NOhWgvrRkK6c4rf3mdvq6TNE7WsVzI9xXYBLEj5yMuGUxN/wR
k7MPCpGx/fDn+NuHQyB3gB6Gf0KsvaseFIyxin/0BjZpR0qyuTxg4gzG1/p1wMI1FZETr8pkIHg7
JTCC6/kkBMXcG3/4Bye0PR0YxFNt2ApfXEgRhQyn+sTqh6hOVlTtu5M+qD3eeWPM3ygJHmFW8wZA
T4zNKYbtnX/pMaH0rIa6jSPdicRjh2lIOeSb4Ea26BnvbuGLXToG6yw/DMdjBTaND3eMrjJMpOAa
mnTrM3LHxKF8QhapPznr4P3EQONV2lDW5j21CuQ920ncQYzfgGBHxpp5GktoNOi0+a8L7HQMc0TU
RU9dYNEWcxSMkOaJHRpUkUw34kUqrCsjJu/Snt7fhjmN1xsFYWgjNkmbNwr10/qkiYqslTDpQQr1
thc01vWT/jkeFeweH8EGMwGSzrLhq029Fay4OqwzOWep+Q0GPcTV9km31/+hrdxsskUKf0rrrwTj
Zu0RAmFLnmn01wDQnIGaHLPYc3a2E7Q5X9qmUm95xQ5XwetYtpsmPVun5Npa+3ZUkHlUv9Vo4ODc
qKYB6lG+R+iMw87dWonJ52XEJqGSp5i01/s4INGMtES1PJM+LSCytIRA04iLF3aW049Fq9c8bSF/
Dum+iFEzURmJWFN7Ozetwpsv1y/yNIuyYZL4pl+DHz9QmcNyxzzEysaYSxqmcCWcOBr5i7qlfyOe
3u6zlfOHLQ71eYbQLEHdYjojaiJsIGwpNpVdMLokVE9qf1w4qKOlYFQhg+8mr1joc7FqN9BIvW21
7UJknLnCSwmPUNEuutXEBucIS7w4e0m1kwjOwTwmTJjOweZPwhUyNgSIeIURv1varGXkxixO02qi
phXJq4tql4uRJE/ZH+vlQU4eEGdqbImzbeQC1veeCcu82kiDri/f7kHumDio/CPwLAvt10hg6hby
qSRzIw4Hr2/dIFyIGb0UfXeCaggENgN0Qj8c5jucmX9uAacl7SrqCbBmrmUk+afZJzAhnyzlMsRb
VSNW5/I7Vq0zMbMv7S7LqrY0TTWE6xaynnLdgblwJhcWtGKFy9C1+4XhFScY7cziQKc7hfIEvSRb
LWboVUHapeEdiC8i5IAfLyJdhfdPThOUoBEQkizDAjtT/85xKSOOvjiwgKgM2WWvvaUBvOX/cZr7
qEi453K78BPXycGTCwwAv0V86v4ujZra0e0u2gsY5WzHG5tDkV52bf9DVe4mSMDFM2c62mEGc6q4
UZtxh30ijoTh4vrvrtzKDGtrQ5cXZ+2f2HVDAm1zzdb0kEHIKmPpXCFX4DZt+ROF5fXqa0+JE68u
cQg/yxIejCPAHNecodOaQIU+b7M/AYwbvWo1gHxzIUoBSR2Amikvm1BbR35xJEBU3ExAsdxWnivT
rsOTMhfn73X4kP8oqDkg3sNRbmOl5IfDxz1EtgQu6wfWS7xgbxpZRkHJxm+cuDc6DB1iCJEOCLec
CU5DeilSwwJLJd0/5RB1jTfpRPAGMbRH5/Jl7pRCueI/dEIgqjbp4kk29Acth0fukfZraerGlrj2
yO3lpJqdGJY6knfhrXRZ6VnZ9Bcs2RVeWBTH5o9z7NZrOIEflN5K5YqTAx5w43kY7NnPudLBrfwx
EUF3k0a1nbvMmaYbGBy+FQ8eqgg85O/SQhFd/oTkAvFuAHTRq+DVv/fMJ/A0Ik9J2WH/Occd1RUh
jiTt/MfJoZmgkag+zk85Cj9eW8ZMsUADxDxefKsqrnxKMN4ru/Vw8/aJsKBKvVBMp3v0odFCnYRd
Wec/fu9Q+hGKc87o5UKwNm465WMgGZRI3FQi7DQ0eQNjKiZTFKXNJ5e8G+ItTUr6kmJ5B2KJQzXf
fxH4asxFo/TsJ+WuvR1U08SzDrKTYqmAs7SDeMs2EM8MXn/ic0VPubKKk0i9dzeKV73mwy0+x410
Cj/fxOUx2hbN1pJ1riMnWtVvz2uB3AgN8+3vWhWt3y7Kde1L+Dy0oRK/68CUu1hyS24GkniVsrmK
rYB7fiUaVy5Ro8nLOU24v6ZXHQC5Z2/jSNYcdkCWTw3EsLTABlbjFxkQLRm4HqEMxTCegwTKokeL
jJEeJ9jLuDpOntvIjYHvg5LQ91TgwLk9brZJAe2f1sOfobjVNSw5noRbJJBmJbqyucCU12UsTes+
asGaqPjNBgLDERLheXK5dQnjd/64wZKoe6NY3A/mcpCh+Bx0tHPXU7pDsPK8LtBBqmZS1FXV70Nf
fDzgW3SvKBdakvUFvl4Noo+zEhHUduQK0Z82R7L7gA89YwNop77dpfOfKGgdnXVmmRUMXd4Lj/Mt
9VF8gAXOBJH7O0vOg764qbGyMAhsZL43N81aTt6E0+pS359T6CkiSxT+sf02V8dqvgw+MkvTNyd8
8kllU31skgN+yCPsP2ZRHJ3qmur3xXcm21t5BgtoUCCX7DHrlWSlnLH5e5Z5IFHFYT8ukTby2r8Y
8xwnDsjdXMwKu9kGZvzEx/0Tj2coFnjalIlLT9ALIgLJ8cNARYQiua0tYCtQXMJ7E+j+FO+sY3Ak
58Xs4AZWf2xtkk3qcmX2IqRjrtIceOrg4ZK4rL2yQmBt9NGT3yOlXuVoRASkGSesp6hmuYVdglc3
poyCdmkpXe1iD90TKqmedqmZKNYI13LAG2SP4AjaBtiKFFesm13ouQIEQAB9YsBRGrGU9t5OdDa2
vWgS5x3jq+PVTYN288D2WZjmc759L7NcxEXz+loyUzbeqhQUNw6G5mYNr/TKo9NJa7GCYXIkomlF
2m7fDnOPU6jjcOHlWdJL+Lxwewz9Is8nnHzBekCcOK+4mkZrOFLXAIbM38AJriKQdOfdtImpD8eH
05gIYc/6huRYsf0RBJvKI9HXLm1P4V1mGHgdy9CkVI6P8IIuSLHKWRVKJI0kgUFIH8l0QJTQEjse
CiWgasHpS5izy2UbUwytNoEufwVR4gYKnmpklAV9k+rtJe3raNhj3BA3gyRBq3RGwTxUvRu/4nuw
KaWlG3teTS3CnaMzZd3N88EQ6Bcw/48A173PdAmFe+VjnS7wc9iZbPrqZ3aF74+2tBtFxX49tu3N
V+37DA9soBV9WQbzHC7Hus0HOoD1lLaIVoLhF92AZWnnzFWZbibnz1Bn4/eWHygmKqq86NDB2mNJ
pjiiUNvW35w4U3MQW7OPsQ6lCK7TcSp/8dJNiyism0QFHga0EMo+e8ulBv3zb/GMQbNgLdU3W3Mm
oCxShB3LHQhRxGziGz+/m45jUCXmnrzdzqvnZxUNn4qUpF4QfK7yZiLldzZuV1OoxYpHYDh0YqDZ
G/w43uV1AMm8sVj+RG7NPnfr74+1DYohNizh3kgQT0fQySZ8575Zy0z7tyNfKzdjyUzlWhmaIILs
VNJ+zcOqeAWupgE3gTsEY6RzXOlfnQtOyhZXJwlvQQEZzr8L1ZmOX/PpxpEcaW+ISWWRRNrGe41w
3YFCPFs9y0llM75Y+9Slpydn+d8A3pk2kMyO1mQLasFtbaXHTkQvGhi4mkK+2hqrDJJiz+cL/q7V
ZYPlTb1KWBSRbzHqjGYtEh+apmXLnvGTPy9XwLjEF4LTNom6zl2eTLY3a8EIFiPsebfPSouJp+Rp
fZcc2q50Gixgg2Z/Qo9XXfA1iUIQl0ZaEN76eL7a5MTQI8NzM50Gu/8NwO5ydNajNTSs4FrsOBhI
913RtzJN5T9wbJoLZ6rfBE/PzCqYZktvuT/eKAlz8JN1LvuQygTJAGklN6CUBPdS/LSkdY0AjZ6x
WCbaH9lcPcj1iLCr4ZoX6+pICAEsTPN3J2DbnN6xy7kvOHXPejcLoWPQwl+sjzhaoLwgyiLgP7om
dNeOIJHv2J5PO3viNMw/0Bb/wgptfFJXNWrF/BrVdpSbJRdx0UBtDsLt4AuYczpbGY5W7EZ4wTus
CkY0nbL8sQZmqio8pCobBxSlIc+EkppCCseevRvb4Bo2lcf7/gATfx68QZdubUgw1+EaY3Iu078V
/gldRSXPyj/fcor7YLbtZ3ZEjz1Ax6RSfklTJw/wCmUSjbJnf8B8oW/BKNALviOpxYBMq4qGTXRn
SrOvzeL4jFAloKUXwkvzRzHbPDdHGvSL1E1pumn6UixvmIrzReDs3QxsgyZigygrMm81NwLhJj/P
+xjx/B9Mf96DmbDggSJaaz7VhANoj0iWVYy/ta8ycMQTTrS6xg8pQGa0ygRfnxKDaOE7+pcAhNxQ
eid8XOyh8ZGeUT6F9H/vvuD9lXVEOPDzj88qqiuoy5AuETIINz31YQK+u8bCnQShaXkD7H73J/ZY
voGJ+vsb8TgH9ni9tncUZthGLAmfAeiDttan3uiotLq5/uZ2zYnbdho1gkjxr3o1CWjMEfeJiqAM
mNmE17JDHxVXqaCjaNGuoMc5Rtgd9LXdral+ifzOjD/93Sspn8Macjt7/e42CEGwQh2CnbYljLbt
5gnlE/uqPU6UCzXanbt8yKZM29SwVssWoQnaa2041VylShuX2Ge93aBDiv3efhADJYyc30vS6Jhf
7hLf9IEuwMG5Xz6A4UFiZSXnQ1M8G7s0FOvbm7EzKds3dDpRicj9X6puQYoFi4S7kKtlXUVjncYe
l17i+NZ2bgpF3WJS0qbyoc5LIgj5q2+C66R+NKJ9KQWKrYFUf4uqwWtU5uJH+QNk/Si7/YvAo2Hq
jP8FyBEG7IT+vQwSdA0HHoNg7HEBoAcA5/Wbfl+nNCSN/IwSXPQM8qGABp4Sd2XoI57qtnpDtCzB
1KIWro8d5ITlc+RAESY2LNBujOBKqagEZFEAfuGrQJCA+8V0x7G86qZbBVTp0paHnUnw8w5dWqLJ
PQVeR9loTWARkTbF97PePQ5HsT6h032rYlZWUBCPI8wlXcHDGhpTV5uaVJynZbxIj7vwqrrlUzCC
nXs1+m2EEYNVW1kdWMVyHNuDmjO+MoNtHUVKUqyPede9ye3z2VP43N+KUcBoghL8wwHr3cZUqApI
tpFwrr4P94zJ8PhHH6gNx5T29FRsKiLVjalao9eMihPSLt7zuGDKTiKimpD7V3f2gYRXBY2i7YUl
kryoxiz/B+kteByYsH5ijh8eDbmtMLR6kKzjEFXqYmeNy/y/VsgHMHkpYxCCwDw0x+NYF2QmB1MH
wrg4BiKnog7ZqSPgOYb4h0P8nB9O5IvNMjoIApoi5VqzIYEnv5nujRqSxUeR+7kZqUc3DOxQEX/w
ou3p+5cofJ5RH3uHr/CUsjtLtyvSOoEuiiCP6Es/ETrj8Pn4ScmnfJhlS75RjAgvOZbQ9YlmAaVJ
s2npzCa4DYEMzZ7NUQwX9sriYkBvFbkZQwjIjP124Mw6BZBIZSTOzwG3Ckp8YoQQ6chW9/3+LDPV
PLqIK5j2GK+yqmmlOr2KM29v3pHq0LJx+2N6lAvrS0c12wEpfBPzeJgXcKJsNTtUp7HJVt1cyad3
swDyU09Fw/7YQeHHaz60iA8DdfdZvVndzaN66MyaTm+i44vsd7UF0J+R1oIpiHMoux7CZy902Z8Y
xhqtaKKJr1Evg1cRlBnfcEqwMeRIkrRa79XclABpPOjj/X+AsnRLO+jFyqBEoUdXELgZWs5Ga6y+
yoRkv/EMp0J5NsA7JqqU97Yg0DNQWazqMHaj5vydaqTRQazb/5zOs3+kqJkuI8241fZCdEsRvVDd
29E0a4NDEOmH6BVJm4n/VRmkzgf+jJOoKkMDnVIjRviVSz8PX0n41HcurCyCl8vHsPTv2VOfKEUO
Z3fqZJ78cKTzK04tWM024UbeyoJ3F4c0BZZFeVw1vyA8JjPJVFDp1g22xJ6bYOVHs38TRLrsNSVF
vbNZUbWQiLyGQleNWU53U0JI0e0czm2meWfw2ZRVsZaPdQ/87bic7F8NAF2gJy5d9aGjri+QOUNV
JxQxE5fKTTchA2ydQ4JOOF0reJCjMp6rGTZ7RqTpQkTbihI8HlJlXJb77R1Ijj+lTvJ8W2aLnoF1
2cz5oaDV0dVXjAT9DnMgJHhWJhZprG89rU4Ir4ZDww9DcIX3OhTEt+0XpFcp5y/FkG0+k8JJ4rJ2
DMMHJg6h4syUVSmf7SoRSDiHk/kbhvQr9jDtdt9IrAQ7eoQCjmNoXhgPlJDgk7C744lKfXcu3B2C
/3NmjevbQUVBjuRV1AZ3mdV7UPpoohB0ZhBrTKGsLMQmwfkwwqvshV94YC+mlSiSjwgUxgkekHwA
z2UTter5Fe2fYEIkwPdPmcigbTvG8JQThCK0NIyG1+tQjyeLWWL7R0Q0R6VEYHXhriP+ic7QNAMG
rroOGcc0tQ8L8QbqIeCZay41kVbZj+qQ3jl2U5/G8SVgtUQ0ItbkJ2lGEAEemdztz+iDJ/+v4l6y
2baZLZMTYx3evqhpxnIdB+HBRHW12+xrL/+wpvuPW5u9pBI/PWSU5PAJ28aigh3jchTL/Yx5nEoO
Sz9jhPpFwKb3MYoevgUNHtFx8PYwGmOgDI4xLjtIfFMrRuUZ8//yxS/TIJYSz6WgM83Ob4PJEb1G
BrWnkxpMFC09XypV+e48rsZKLMI6R8djtkKDguzP4ayQL3G6yzBVVvMeJ4yImLmc+XRohsIVf9qz
mgIbwIAPaCKAqr8pSNfjFZPSstxzDWRWLQIbOePOR6BRtXun3vGglpXfGf7iYeDunnePifKZLPK/
olqSL2DEdDUgYpyRE6Ze8Pi6PiDo9Kxg36C2XYpkhpL/nj6LYtDsJMF2VQ0gOQojcbd0xIGvOi/O
bA8Kpd3EMx17UYxbaZkJ2knjvD2NgQeK09vL39AiVnEKpFtoqUFESyATsMjEwAwDJ+C0KJUpZ17F
MjnimdRah9qauWAIuUl5dg/GFDZpwsLnlTBK/bTQ4efZAxAlGvblxlVSTnkHVNgbat0zkHOyDr/X
Y5sOgAVZrDyZGwT2Vt/stDFTsPCN3Yuz6bV2iZMEPK7eUaJz/HVbVdLPNEeEHwpg5/Uy5s9XO8Ta
nUJ8X18K8AHXSfC6P+wwzIbyPvGZmorQE9S2olQo6id8+zSLQ255aYVjkIiWlbO5qF2czeZEsbiu
+aj/fHX9zz5Y0G6a5+EBgWIP/F08BdVScjgCRPrarnq3zQUZTOa6zPLS0MCiPq501s4Byhe0Znzq
LwBGPp+k4TUksrZVrzDLZb6zsl9lUaDpFmLErhsozx3pfcEthyEh0/5i0LARCoyG/XCfwQcLfUG0
aGhmUXCrZRd8dQA47etuYrnlSMREqngAexj7Eh+mRkaqnDiT7dd80s4MnujQ2IqYiwPcYLhul27Z
e4jPHZy65BvDX0336/btGuS3gqJcglP3VwRrJyW0aIAw8DAerUSPtUTLHtjU0k3hcA/nLQrOYeJX
TEwLfGCdTtYLcYTrwxTnInwNAKd/90hWlImYrjS3uaHIIFEKF4L3XzvGBboj34Fg2C8PyM1dgk8y
VF/7L0FF8vKiMEhl4j4KkbUoiO+zNnCjMXz/tqTjw1TzADCOdNrgUS782mLexZHG1v/oQbq7sd5t
Atdrlkgu6WfOP6N7UYgLRta9jHd5JKopyasacDZhywyLBUJNi377AYMS19ySA9xv76IhxshAE2lP
x0sSuhfLm9aR9GcNH4rqOrPI92W3adgzCwwdKbyHh8nkD5Ddk//WWadexR9z2YUFIawM1LyAskI6
WuzsKI3Ks04CSK8drPlnjqWih52c7k9rzvKCa44nuBHKnQngIVAUXP/IImSsrf6xlQvVnIYKg3ke
fZMHRXQcjfBKoJ/Ew8Mq6fRunTNJFlVyFM8K9aSv9ZCtIRFubX+1occtCKRAKqvQ8fJInxLBjO9g
NTznUefin/DmX1IT/bxTx+zI8WChR7PactwHiNenKf8DyFALrfnPSUaAfrXRGMLIHgwdSNnbSqLQ
qPGzA6vEMkCBNZM4Z6Regj5cLzNIBUAkqjtGr4AQf2xT9tdqUADvyGd0mxCnhTOYAhayP7tpLGe0
lgLWSf+H8EmzlUS2weKAbNKyu8q67lFDEjk5/xJPPtSq8nZ9k7qq5KwCNPLe+SosGD1yk+ZqpXMR
YIwPze9VRwx4ivKSbyRrrt7j5PxWqD250z5LXRedztjVTPKXe4vkS3FqqlrWefRI/biyw9b97lKg
W5taAwJFoZBvT/dtNxhTQ+zc1yTbUVdx2gNv/kiLPXXZm7PmmKNtyWrMe4h54E0NGkSJo4Wco8uh
9XwSpa1CF+UIGik7HYBmvmCbxS6UPCNlu19VsmIBbuq1HaAOrquL+uP2aNiGQRcdkG4ZOd1vc0Om
eibm725jEwbUpy9S0FZ49LaYt92BU/9nBuuZaPsoJi//qz5nl4+SgTpuDi7tX3xVM1dB6aTW07jv
UKZk8O/3Yvhfqu0EA2TRkDJ41hi+H3OXf5MKCNoY6ydRQLIDDSob3oaEyYCjmUr1lsrGoZ+YAXVq
wY/xLBBwCHRS/oFbcVUZw2Wf2qUa8yokXOX2kWWg7M1klt3o4L17NnaL6LtBAvW5mg4qCj9R2m5K
44DY2jcfoBfBqUDEK1ursWzgzW7DpsQ9wZir1uTEHhL0jw9BbUuNqaJgXa75YJv8EG20NMJu4WRw
fnRb8em1sPyZj6MPP5GPZ4PbppBYQ+RBU9BckTPHpztVGCSIhUZBJVUlBj5AT7gLbTQDub2YSiZT
MHj2TTBXS09p/Cei9eVzlCk8qPMnV0306A2jF7zU41cFUPGaj1rTJlrC4C+yJNSdKX5qsSNHQKkj
0WLtRa5oh2kJUhiNsmMBzIKm8KsL0rwuja9+4THQQodpy0tl0L0yb85DdMi+qnIDTPCdRJ1iZHqy
FQHFmCB5R2S+bWJi2JBp4fkf7h7Weq30S664OUQPPu0Qg3gStTj4EAzxOJD8W1RzRDoW7cle8bXr
AxlE4Tj5xuf+t3iJwrnS2isiIniJhLAKQyI5S/s+Wz6AYNwwDvwOBRtmsa6/1iH0J/FCvO8nohuC
gSk0hws7nEuBkgbE404Y3jbIZvyQGusFAm9EwvUX3CvV1vba48jv1EwR+zkuvJ0AOEFEaasmDwIJ
tUJ5zpIDaTirRcouiOEOqUN2nXfB/K0ZVrX1s6fw0u1a0U9NpmWvBQiKT8QJeNDY9f3rViFX1VEW
X14dCsiNwdI48Lt7Ixq6mVhzs29zRduZvMSU54hv6TU0dBIVwsOlxvCkmnEcR4KrnAOKmaglrsA6
QbFJf/ZaPF8w7BjPKLpbnD9N8lkqX9mRvI8x1OSXek6dz230kmPvPf7/OlaVfhXQDP7QllnXXyHv
0U5ZNDsig/kBoNY5ZJdvZjttuoOpmROm19GjfWh1vGIwp+K2VJ/saCYQtzrCDTy1WjCfBP02vo9C
klVsu7LJR3ZP0S4EgEuW21VBaAF7zN5MKPwux0fa0OziU6l3JRl+jNPW7MYK4eVArFg8REW4tcAw
bbOyrFXdNdMtONAlel4mFW62M9GYcf+j2IJelCQILPC+mDbmhNYpWoOmyU+Idth03SdyD3FLnuta
Y+G1OtmY2pP2FWgy1hF3TJDLm+3FcS4d6cTMAWEiUFtsJn6wI12D3Mgz97DVTv42+46n3XO9FIDm
hAIAhFwBKOCOTGGXM2/8/gb4jm7P3dBrEWcRXt5N2maeGDD32JxJOTzQ9Fi37gU1BrNqyuzBaWdU
pdmgsI6teF3qxQAktBPtJ2VttpzgfxJZU2jEnDYWF+84NA1JTqu72/t61cEne3SPp4OeADWRFzS2
SgsBAAezD3u295il762Aw1dE14LhGdaD6kW2eHaaD1tce00XW9ydem3vcoivME2wfuevKYcv4ZUN
4CioZYobyJo6FZGELebnIeL+/JBuJrEvRwZN7JGf3EFe2R7jw2Zj0jsUp2fyGESduKbQTQlBP19H
y3S/Mis1ZnzxwzglGgCNH1PWspQn+8bkL1vxYI+yVFWduIMCeuO6sAmxzDTTZ8q2N7nvgjHe6FsZ
jUSZp4HnWVanBepf6V5/C3/9uCDTYAlw6A24lBRdW4KAstSI7kwMzId+5NEHyKD7PIGkFES4xwvA
El5mK4kSy3+Z25lDMvuU9SbGksrUHLf/RO1S9hHLr7/lMXtXIggH8QNNU0UuxzVeJJ5mNw6k/1HF
tpMR4vTmDc5y0Pc4zFH1lvgYPAKYaqmok2UpEBfD1Sn4j4xAd1CHtzX7mFEe0WlU0qumzb74DMnd
SqoJM1EAkPT4NjAscCWD9cKOEp7T8WVRAkRl0kXt4vokqLlF3o8FKY+9DdEpilJz0cbeMLDtsX6K
q28ZzMidNSYdQG6k6NFmWjLyk8bkWpBX2yZiXGfv7UV9pz227+jq/b5TZ/Yjce4ksN47aQepqB17
19W6FiPyeXH/0ZMKqW6wMR9ehUx0tn0GKZ+0nits48d41xai7cHFcP9X/osMvkqzwMGZlMKXAukM
RiwaSzdUWwMFmrkIRHmi3NsT642XqQOQ40nCDVR/HeGsqPY3sfmgdNXSHT2vfwIKCeioWw72+6hT
uhybNtg/6JDlqb5d+H86YwXPYj/Oct5gTRf2yu9fzhlsMp34aNJvJt+lDJkrakbfKe4UnAYJMhcd
yjwqciaA3mmBPMBA1+HZcVrrXAuXfim9nw7STEMXLqhknMllYgTw2h5SH7GeBA7vPgVyyMZHum+5
i5hiWFZsbQV+VE0rt1HSDdnkfhK1SCAvcTR+WBec9loTfE8mlQbY57xgz5MzZLVzmhWmU0j0erDP
MyR8hPN+cNdVIAi0DEcw6J0d1ajSZucjXtfT6wzZw25nN/TZ2NAtcwX1IC8yjlypYKeyphaNjoHM
6iiTE10Pwsn6TvLdqyxPeU43chfXDVGGczw7T+rXPPWvzvWBR1NcqhRh95EVZ0/rX/qNPG6Mcgr2
wPDsL01QYmEjU7UyVebucMkW4QiofGWSYp0xLGCHaJNzRKHaQmeoACktZ+ALcoDM0Tii1I8Gg06g
kVEArpP6ZaIDVF5Drut4OXruSGUlSu6DqPCcWcy0xOachO/JHAEIQlZyWtmgK8c5/CrWx0//ME+g
xrXGauzooo/BhyM3CyioBF+8nRbTztFzMaWXg370WW1tqLMQ30eAh7B4WnBnj7XwB8131I+oQXvk
R8e6vyFGzr/sIMzBC46AaeDC4jOes1p5bHVvHavNUpWuhxTdbDi6GVx39U1CRQ/I6bk3qQYJ0B5p
3MtwJaRXOpzjcnVTBRhWwjVpgVabb10PxQNzfsCJNHut5oTtyOTGAMnBoxHlmqVnRrXDuEBYmG7D
/rYcHCdf9MHxI75EeoEuIYQrYcPVajpG3A6Ql4CJOQmK64Z8QjVZqI3n9z4Eg4t6ocj9g29DVWDq
DB8BjWPxaOXl0C2qmERagY5JdJc2L73evlt/eQhiM5V6evCmEc5oN08jmheLQt06e1B9jA1Il0js
F/8klTU+YPHejsL9wdnpAt9FWum85NZ5SqQaJ1JmvgpVxQU2EBR+up2wU9CO8J8pemp7RPgO0MFw
nwuZm6UfyYGYlTB1WPK9WAdVfpNEmUjkJGe50BdPWUK7uI1iDlcbjGzP/agNucG2k35fIvwiY3jl
5norOg93RLJGnp8U66dLY+JeGAsU8XSqR02JF7D8g5yi9JxGldXhtqzNxgvK+dJEtwSkNHLqfIP1
gBipkhwCcQ8i/fmAIA1CxyS0MeMQ1bgCrxPhuARgri8qRcwPNCHs69fgtuP2d37S/R6bH6wd2i+e
eAgd9Aa9bAyk4QfEZoUFhbBNvBeZwUW2oFSD0DEDaZufN97uuDctLHd9Iqf60uhhXovltsNJxwhu
g1OvKFyPMzSh/4+3h16xa54Xh/wN4V9YXCOn5nRHeppPjIDHhz5mv75ATUqKdqhO407tQuzQTyUM
bCITfi25QSYkePY27xozFN0yLRs82JPLlbNNMeifoibThxuM7Ws10wJsxn9B+Ool+4uEsrnSvZ2l
Zc/dAFA41zeKBs1jYTbcyBQWUVwSl3523C46HQcgFld4XENDi7mdGu5rT+Iwd5Ib7rnPKk5ifn8x
ihKL08ILPfeaEuXJ6t3DgIQHfvQwTsC1A3w7wEi/iQnD3JSCFjI+BWJTLqKs60uwptmDlDe+15rw
zsvoDHtxPDF6nGEVUbceBrTy/FkHMV6jXZUu2J6rT9/WhYAAyeSN+JdabpX+IV8K7oO96vb6tnEE
sGc9H2AxMGrI5EInSlQZ4fiqT6DQbHI5DRTKQjjR2BT924z8pKGkQsXNsKfn+Sm3+npgiwg+Kj37
kMqhvRrt0FHJAJAJK10oaPPHemdBp8d0PoWrgfCaBv55Jjzl7gPJ4j8mtDkhBRqaspbc/lkBs329
jxFCExYCeUncg83Is6Em1olf5mdNweo23XovHoF8H9q6rcOUJv4aZdXGmpBpG9caMd9OPVGHTxaS
oxTZj2BbuKqgXw39u2hTvQbxGK6hxX3289QqnfONokqnTbaoC6QMZv0Kck2+JIVojzMW+SxBK20v
8DaD0ZG4EncxGSpBGVCx9yoAlF5IDv7HL+kNK4GD/F4TjsJJzYrxBCaylJAcXoBLIrHWnsHyryql
ndlyRysOhFGjQ3uKz4N3O1ecd6/eSisBwUwT3udUTdaYbXSvMaElFFhQZxKxGJV3rOClE3lWLHfN
QE7+VmBPSCU2fa8KygP6gU2nnYNK7rkgXUDnAVjtuRwQk4JRKRhPkirtZ98lv1C2uPGqkTlum3Jx
lLbnRxKRLWga8ZKPaAPVIyiKhkWAR7BQwvVlPsL80I5U3CnBitfT1MuuvOBKW9jIOxOUqjRDwYIQ
rEweZrQfODFoAFfu0cuS02uG2tZe5usmY6wvAfH9rMYqHzrH1Zfzdzk8U06zjhBUNtn9MIsWaC3b
cAT4bRBdRabu6h9xr59+5zYfz0oCIDPWlwcMaVmd9jHg9cbcdF2ZnjxUA4HdkRsOa1gbADybg6e1
xVscvDzGDvAlA9LTFnIJ35l17Og8Mc+NxUbpzRuT8oRUdrnJLhKdueb4FCZaBsxr6cArNSnlKu20
vo70DIA2Rh73CBNT4rCxte64Tvcf7rSoQhtlqQyl20iLH6PTdP40lrMx7wgEd8pvpNjnQjFnviyY
2VZbZDfayDRCts81p2JpxLRhKKGtIHL0RiY0v0KVFEKCCeDKuutnPl3swXUK1n/x4sr+tnlTFMh0
9n/mYcCclsbGeNTp/0y8oLkiPYfv4X/7oCCejYA5g1sP4tcQ5MxU2X3cCdvWi193P7sFp6XmwBFP
6BARnBkrEnO2ImqyuhvrCZS63zG/zS8LTuXILVAWdtuhbnWaLwCKpwOeJ0Z2swfqbNJihVh6hNDW
g7LCs66gbeL+fvYKhOo31gJVRfdEoceWFA2pfXdy7arAPFe54A61VS6L19ECfhnkBzDjsqmBrEbN
HQQ8AYDejbs0G3pnFEudUo6PwT7mPsrH9XsoroW0u/3Nn4miVBhUC+8QrD0VR7/WgARuFBaIs5a4
DDQI0PzOcgKILYJOCYgfLu1jyuvQDUHVT1hYAkv6Bs6Ze0RhMheFEUr7mTp6WojzgkCnVqErVrab
VXzDZ/s63+rfNl77Zm81PUYgZoS/XijFj4/ouV5eCCVhSNTYD7tJk20f1wX4qv0xTXp9f9htBtl+
2JXxXw6c8FlJekFC1lECZ5ubGpnmo85m7D6S+7dT7N7yIbTpDI8cXRybtv2i8fbHM92qSVvDVPgj
4Tpc569EtxaDy/8LSM95EPfD80xqrTq/gpgTeptvsilsCHPMtQCFFWFhhFXUht2z8HM7TwrVX22n
Ugc1BEMDFvJ/WAy6KYynSUOoAFLYzRVf5F2yRBAsMHg/98MfkUETETt5VMYZvBBJ9Fjq9nLhI3WQ
Yygw4KaZNW+Ul/FXm3Lg+5UiG/WyVit3Lvo3LmKRfWqO3yCDs8m9rvx7/fybiEz2r4fyQtJb6Evg
f0ICD+jvXzz1iUjQimasMGxi7EsbP+8Dwa9rI2eWzlThKQXxYOGUOyLPOtSjGFUrH3Crjlc510a7
CT54AZNGObwb1HMqXVmyl1JKeajVumuejaZjSZJYKPoqz8Nc+VbhZy/CPcay9DYcQm4wyxisPhF7
NMJG5ASFURUIwlMOGZ7NVhAsbRvs6h5IyL5B4cjWeoBeOYDrANGctBInwemhnYNDwnQ5NwTYPcbG
pKxxnaL4oGJogqErY811KnnXcYp06yLdhEx1bzjOzGVfhGNnyoSvTPxH55v/ffh4EV80kSzLLM6b
UD87LVH5Tt/Dpbd2zWJB1P9TWvwaufzxMQzaixhD3duJsuOgSa1yPNPv4of6HgLf67iMxumNinZg
NT3yH1OB3Jiw5qnkg3enC1EyjQiGmy8vQxiVSv10UVZAuGX3cTPegWYgAPay/mNLAtEDDaxSXrN6
zomqlTGZ06rNKAJ5cwed5LOpfd78pPxXb+N5pf3S97aG6j5Js+1hw6od+NEv6WNz60SGTuHPYHUI
VgZytdfxG6gdEVkf7dyr1XgZQT26ijfgx6wINyDckrNHM9VrxzpXCJ4zI2E1il0F9pvrFd1RFbqV
ojciUnQF1vVeEB0vtw5Jn+8++StIQ/X8cr6g9k+eLmRWdNyVe+AnKd9DxmryBZaYrA9pjwW3ONgr
KpSlJrytNSCRITZepXuqnwp2OczCp+7PjxZzWaeNMVefEW0KpQxtSCd4lXUUVXkx+jZ8GuBmbOci
olcFN/IiuCPAvradflz6lHKzbZfrfBZZm+22Pb9QVcLGc+N3Mwq+7i3GC06wiY+/nNZYgUCU8Qt6
7CdCI8ZzUtBVtmT4aaPEu3p5NaaIQD5gwUdLuVnBcjozVieMkXdJcwizzBIwTnekszAHgXlOn2hu
drPmgOCSXVvEhFhMj6VaGz6k75bnkZA1xviWUR/TzEJQPkyvjdYbRoGZEhaCCoXrm8Slgy+LLYc/
vLVHWm8KR767Ifm6reAcCloEa2unI6eN2XT2SF9c5FO5gMpseuPPAjcVeYJcbFnZxCQgGmsq7T0S
1gcEW3otoGDlSrrCAQcPFMEztlc/tbt4MI7pjUtRII2uy46CgeTHxbAya81OFaE2IuHLBhcyXF9N
HFbiQaQ7hAxy/9DndPKTu/zZUxhrFUXNybKVTAI0MK5AdocBGYTtFI+l6Tv4rMDR6pDM3zxW3yLS
2zxOsz2HohQPy4Ap87fJe7nXKQP7/xZo4ZWy0dv4505gsMunNNgtCBT13218mTNT49zY6iAX7Ezw
ZaWTv1NEZIo4FuZoa/cGdw3e8tpnrDgO0FU6PeiAw5+q1wecCP6a+Y0ktEqgL1/4U4hLwYpJgMiO
tMK3zYjE3VqNFHsMcVDW81XTeu+i6OXdmIstTzg3H6knlK3eeKVblvNmlZkZuUG9WmfC92gbh2L7
Cfer5foaJqwaPIJVUYalBHR6Zmy3qZNT/HpEPwcu2BDrsfKlx6+IBj2g9bGFQvKNtR0oDkEb9yDf
yYBRwTSTZc6xoknpHXSocNjyzIKaP0miEohNnCi1jnyDejDny9idhhsuQRKSvzMJj4TcjsYnNyzk
VHC/ulyTBJzTRJojr9IlAr6DbO9euv8C7vdozQlTVW4z9ZSab3YoC00TAWvqLKfGWekJt9HwieVk
WA3Dhw2/uNq9RE8OilAgsm1ALxzrb7kqwHnokiTnh6dwTrwJOK4hPs7U/61Qj59yzUCzwahxsQ+q
xsLzqpeODeB9xKu2gyXW/CUtUG2wbWlXgUwWSq2QVmHsi53dTx5XdaoX7/EWr8ALacuoiO51pq1W
SkeY1AcVthqvmGDI906gqyv7ZAc6egWZ+Bs27t2qgTiQ4FNu56nfOkUhm3rsYFm/DzIABq35bnbJ
NGeuPS5iZ3YDrNMxYubCwBfkSdZM1yAEpZlmzr5w2k0eRiPdQdMbGbG2fHIT6kB7adrkj578SzWW
gRyZb7MylHf1ZbMZTg4FoWEgpvAzFKeJzyvc1boa8KKzaAQyC6lsA6ByCx6rd/v2MmYCnAj9A7ox
lc/vni8G0Xm9/DQ2yEoU1/t3xqEaoZiEoy0cQ4HYl26FLPNFGsqipqBCLdptwCi64Y3JCVllPwmX
6rVdc5G///evRYKgZpG3bKY4SbDLCQo0Oa8lr88A19qSKPG3M4onY0d5o4jH/FjAyOm20llswAK5
sNmG1Yabl4J5BbyFXrjL0disBKoqdewPA9mA41WTEF+PvwiFjntVwsu20WIox4kkgDB0VwM8VYW+
vVZyM6D00kcZzBsmrBkEhVGXf14h/Q8VUKTSvC4fEUrDBFFEXdpWpvctr3KM4YlngHMCi/AeTPvC
ZeMx9neV300ZZoy7qFPd8NpdADBNsgxyNXIgFiT69fR5oFa6geKl8wePFqyw3m9BpB/Ir15GfMc6
N3aXouy3eqdccLzsgSZcVvN4OqnH5Y3f+qhjnZB1o4mn5EcR3zutN4Oi/bng3gWDUJSO9akKvjCW
cPLXzpZsj4nwfxRgaP2Tjaaznejm/efLk1AIERIzdqgng2jheKbjwCWGw/EYSmE4fjoURIeETtqR
cLkCxwhrCypECTJROAqs8LwLh9HRFlYAugjiZsl2w5Z3yLLz81PO27zTmF8yben5nNQwGiT2sKht
BG9PRmARjRwTVyNM2mEKlIxf6hz+q4/8sp2L/29siY5tL+Ap7k4g/VeD7/ROg+MzeegQPByGiYE8
8yfa58dXOpMEcVG3pP1Dd5TAExQrgr/I1f2y87WPEYE+JsoIOG3JhtMS68KoCqt8WVdFSbQB9T85
bvra4CChplIbsUU5sL+EzYIheeSUui1xha723N/LYPWEzRrp1ptUyYjjD9kdiqS58qBSXbSRsna/
0xJbxVRBEiJf2XS4WoI7EiKfMRoBJ4thJM//ChCkGXHN/oKqGQedtJ/D47YqVuLJisVQbgRpJ2yX
8+CaGZWjxrQhH0IAdxYPbsLl7fKuWu93KFFA5lsvjO0JLisN9aE5klKinyC5wVAPb0a61z9pbc6M
VYuWL9ZC5NZkmfMCuMm5+25WJuJE1+mFMI5Pl+nzcIFxnmRnurkHem+l4xVODCgla6RIbD0spQ2W
ccY8l5foiCLOOePXfl1GPs7VfaPRQthb5FsQupe6rukXT0nRwVQ/6+vhzTVd/wr6ciyjvGmOS/PK
t/uhVUnYZXiR3b2V3i1tp0SF0oHYJnqd/ZuefhvMvD1md2Frf8nzQJQRa/MoIIxzvl8GI5sz8K9L
Pz+Kr6urUcTFWb4hQLaZH5g/LWvtYxhdBhqRCjqd7NBCxgDXbA3ZkHs7zLcP68lmmoyX2cYIcM03
NywwbJJx8RhfnhXZMCR40epo1iG4GwisTJG0LV6C55gn+GC2OPLs7UTDhR+a8n6ckIBEh2Ot4eUv
M++x7YH5pHkvvRyzhPbfHJ/xFi1LvpYcqZfrxGa3qQ8hUUgRyAr48BUqf0fcNZjymlxvg1i+3fzO
2HwII5JnqgKvorMPuZWP8J2n4xsUBNZleO7etNA9eQLu9qRSI8ZX7YxAw1LTIBLnrgvs/37gZz7N
ulTW1oUb4lAmYaCSytmDDgzMOvaJTPddCSuk1XNB03t4VGhFft7aWfc/kyW1FaOcCO2EXRjoeEK3
Bmbd2ct4Yd0sm88mLJlKda6GDdAIt9vicuN/ehPwH8+PNvmWR2+5h07Ei51csv9A+tEK5Nn04FCy
9CsJReGctkuWLnbho2D76x8OUPAtnDiyuFm9k1JGw/xDIL0WJ45paUwqS7HejIElbyL4IpeANkF7
nGb8rvO4EOAY/fPolrj0f6Ir7QGlISaJNYbncASLf2jYFX9MIgNmUkcEjvbN5ucu217FEjz5PWIT
XMKwcUWN2L8YPB3y/FFztSp6Y911vI2jqaj0MsAKcFFZI16biyPMSaMQNQs8rHgs+l8YQljTOEH4
39DjLoYxgMKCug8hVKtTb/7m+hPjpYWw/9C12x+imV94m4LVJDx24NfQd/pTwf6g5TdSX9HOeGjj
UBknppdMejGdhw/qY0yzYKzJUH7kx85wmcSy2gOvVnK+7+cgytr3Ld4e4vXcuhPyipTNhBDzBq1r
foCKU+J5V/f2EWa+DoHlDUp7YVyz3AaYruVO3qadprg3zeKUlZQvsQiOYgFn4733odKIOJoYof53
fro9oWMmfaGOEUBJdJ8dAHoaJ2J720pMPrg95SLrKcOuwD58m0H51RFRampPSDPCryKk//Fw6J7u
eCnlzmDIs+UW2Ixau99V0pjaj8z1Cil32uoIfI1C9RFZWVHJS4Pk8yByBlDK1EY0Ry+hUS/ZWPH6
8CtDWITXg81CgWqItfrcWHCHwvafRUgMS2XRMbnwmBgjROLCwXcR2juOxhgY7dZokRs//7ebgWiS
cpVHCmBUeslgkfx8SE8TCJxzyz5HzSiHsvDx+3C/lX7hVp0lXkx/zhDqU+iui5utDYPY8LY3pKSC
+C/CEc9Lar9smqvms/bRpRIQLnLSzOp5FEr8vu7DkXuzFHv4MOVFrHoHL3S5tS4XHb9RiPo+ZVJX
LLdgdA7v/J6W4Cogs01Yij/DjqGy4uSwt1jdvtp0ngHGu8kS3lDOwfde0ryzM5YimC8yHEKgef5w
wHLg8CCNaKs6rT906J8BwI+q2HvkX7UZcJu0Y0PNigAojOU0H9mJWjZEqXqLGbEV/Foe0mZ27lb5
SFDvr5Ca+eoFws3xneqeVgWHOnsJevCGw3pF3FEjXHq7/mQHEcAY63RGeICjPzjgoBp/Inbf+d1j
2UnJdmr6O+8J69sS1imXa42F6l5BJp2ONNuniU86jC9hnlIqz2bRy9gv7+oOhzU93KgeGDcK3GQu
vlzl5a1jOY7x0zpUHiUOGSqvVDiS9xKndEsLdOLnc3CCttTnfzjBDgH4Z73ZwBmLoIVM0x7Sl34t
Ez4mwVU9YXVC/fqJySlo7F60YDeYDCfEiezqil6+KI4lrw7BMPT4jyK6hX8/IlXZwaKwPEMM3lYE
ZYZPD834vieKeqptzG1+mWJg190JtrdYeR1y+gEA7jyRZOzMyvGwFkKwOoFZlo2laNGzJ0/6k+ne
xB4SRQZMfKcfXz/UpvI9fHInpFlbVd0pO1ygQkISHB/fpFHTSMuravAxlIBt5z/dxEpMM3A2EsCY
RKXrkupTf6Erqpo4SgbDBkw+nAKlsOcJIHDxlB1o5xcGd6I/HkjiKZf36cDemP+fle7SfRdoIITU
AWZNsERXeiyonGe0vJZQG5yxqppk1APt3s1k0z4Cv2k0jDgc1O2jw+0DwT3tXk53f4JaXsg+h4iz
ckCfra+91XZrB7ExedcuHfGHoIRwdS2dPE/4zbDV6gleY5YXzGxB1NRbRw71LQls1/X+ChGtnJPt
gRPQFhGipDytFsN4VIKYy+xeszwBH2LTaXuegPjR/gx3bXqjQ8vGtSFo+uK6t5DXMfYDs0wG4mF1
Cgh8P4g+mzpDziMd1kbydnPnWGziZu5Jv5MGO93XjIfLl0q6qH6diNLrFMtj4p4YMaa/y52uyLRk
QIWwzzzaKy2Mdbs5PEa9aDTscNgMfKUApBetLKnK7Lw3NNALmKA1yIHx+veTna5VJpIQtNjuznd3
PLlpdXwYP68vIdGGitkFmew7AsAdzN3+ySoya0gy8WUn/SBPYs7XtKhc5lapqCPz5Cue5o8+74GR
WPThblbt/IDBVTSURQfbChroPBIHYzgeBin+EZ6vwTbKtONjjEOmvjpgM97dR2AqdiGaoTLqbFSJ
2i+2FN/NZ/Kg93VW2eXtwVX4G4xftd/wfQQcgdVqluDrTwZtIid4SolVSwQk/bRY46oMb/jvP0fr
rILHsa0gXwdszKSrA+pYZ5GuAAynu1VdVEewAf054Vv7izabAb1YGwvejRwv3ewS7LGYhOI6Oy4c
LudC1yT4ZCIVExBFKD9uOstnPQiseb8LjIN3Hlvbw9SvnjjWdLK/Gx6IE/Puqzwoz+XaJDCQSmzI
SwwpDrFGvC2RDueew3Pu4yG2SnsI8oL0KsgQZH/wKOTRECGnnBlxJ2J5ZIkGqrkgHCjyVq5+QhT4
ZPVSkqiWcNDVE521XKUpnfW35VT/NGIfXA9swU410okVP0+R4Trfpcd9neRJY95leuheO3z/lluC
4odv5+r9LAe2w06mBwvin++5ybLtXPViSwp+kWt7qQLckf+IB8Tkr9cbJ/kJszR2Idocl62pxkpT
Dr6I2KTebJE3sURmXz8xC/btFuSyw3I3GZKPHxumCcu2OPWJtIlGvZwwGmthPEEeb5iPwJXsLGjr
Z3gUuu5c0JZ83b3nyVIRhCXunpdRXvNdZz8gM3IWv6/0d9MNKyCm5Fo3808gsq0Vkak/D/BIUZqR
wEOglzlYgZoZDRkVunf+OIs66KBdCYFLCT03MhgvZR5+N1P5xO+HOP+yVCwRfcuRRZ8xAg62GghW
rcPxdkr1DaIyabbhFWDGbWHc+sydRhoPCyiOEJ4TersfTVBNgqr5T63jD1uk0YJLo8QMR/PE//aR
Hqg4wootq+4DZQHqqgkX9/t0tMtbqCCH2bo+xk51a72tpoxtjvpxaxALuj72EDwmxxDMSPv3bzrb
33ZD11meVJyMI/ecAwEYN3aNTjKa87ccBt3TBP8zKbJLS7daijqCVXFAj9b8SyAqZj6vCDdgnFCt
NB0c4BH+009ry7dtEChAZHISnJvWgiODD1Jd6fzbXYks/Zw9LY9eY5vhKarLVfP6f/k7czc5nsMG
4KLG0fmmQDAU3tBfF/uF3spcGxHYsWaNb22tznwYGjZ4Hd1l9AV6kI5GfRKRVqda+rb3w7lX/KHT
swINxq8L8AA++ZjoIXwUz0PL00bEYxkpihYQCLRTHQVYYcw9S0U00k6VJeKJXEF4HP+RYoeVHUkb
U/M1yPBKYY1DIB7RFGaxhBpYmVZDrfnvKMaQBwNSFET66xAkmLzEgoGfq4TL31IIqlbHvmEzXWfg
kXQ/CArFLWHQYkotQPp3Yqna6XhEDmoGRr+w3F0wc+CUkm6XzS5Pyl8IOhup30x+l7ag6quV2gaj
j1nGmiT5814V7p0t6t+ZA8MG0mBxx1++dahLM+tNFaOfS1Y+UJsEQaE39pV3qdLf6GrQugxo9UY3
zI1v4WASu8GDMw9SabjHUuco+ekoyt0FoJGb7aKxWkT14RvG+uauQlvFLd8Hn3WZo4wLMDRoHQSP
Gbzb5blse4fNtYna4me8p+n0JEVb8AWEHGD79AB3SsHcYKCkNFENPbkT4s5b5bZwLlSCM1487EMy
DI7cpeixYyqluZJyEBYXngqSijSWmFkujCzZqtTBDWzTfjsQy2SADdPpuMP6YsHXuXsCgxiLfXP3
q6BDw54C2puuqs9Fb3bLvkn0Mvx2pa9VYMFDVP8khpfejOCXY1NoKqXB/R9qKGr+nhDXdQz1JuaY
j+ClDa56F5MFCO9lfHArWqKNxmvFoU+nu07ov2G6TbT009xuu31ZDZ9icwQfvhgn65xULGVgzbwP
lxzqjc+/CqvvOy7TYPb7nj43QTYq6O9oiABiZgLJx2+ItIWIM71d5/tUegTbhqBUaM3LJ91Dh67T
kU7m4FCQJEdMrg4Qo45m6X6Szi/XjeARem59uxHBjzvM8uNmvc+SQMuMri/ZmBl9mqQ28TbganH1
9/hYGt/jz2hHXM/434tE0u3wBkMi+2LiWFysLko3gK4xVwylJIgSQCNMmE9HUSOQumpoa8+5GrRd
QyZvh9JtzElbEAQD2q4ENkRhxW34YUsBSy5d3Seb2UlTB7/yNOvp9ofzKrgARLxFfWS9vcJOHdW9
lhcy9cMAQCqcMXNXR5y8t54Wouk6se9MLn7eFo/T19j3rhWpZOa8VjVzd0C6g4fbCabLhB222qJJ
3XlP3YvVAEWAqEjkYbAB2SPCzGonHZtCYvK+dr++lw282L8rdkyZUtvc9R0KJTG7TqCmZoU81SkU
n2c4Q/6v9kU/36q7VMSXYOkCE8xT8riIdS/baDtfYvMN+Wn2SDuSHLlrDX8WIzqXf/I/3iNGxQ0p
oio8MyqRTT8mR5r8tTwKvZgWuwBC2LpvhRec8C9Vm3jL/XTRjI9oc3T6lHh95y0eqBRurItITljg
UT67IdGLuNglWapy9Z8fIxyImQ0F6u9UGDYu4vi5eA+xp4g/SxtgQQHTg1j8nEkFqElZfdDiR5td
riPhBX0XpyGM7xriGCicAd0DJNsYW4fIyL6zVowXbY6NZ6/TkA6feXjMxgpbGl/z+uKmR4DOCRgY
DIQjnOYNGuk6PBvr+fJLqdOlNaMWFbwjeN8Uf9F+GkB4bp87H1K/SFi37dbu9p9aoXn70LfD4XKC
B0YtAxW9a/iqr43tji1CghKycG0Ulahhc/JUJX1v7+FSaaGVi/ESo7b0J71lxkIF5TT6iqR6AfWk
/zfmH0GoFy/ATQYl5UNsKCTdcMzGtV+XfHJVsDY9U9jWIn4Rv2d3JHFP8vfltW9OBBr0m0pLkbdP
p3NmZJFgRFHwl++owYkjEUi/QG4OI+xfnVFoGpOfBIbwagNucei3kxx/h/TjXijsuC/KBn3iTCEX
YNmbfHhKPFdnVdBxqfmXTMh7ShGVjX9ax3itxPxQPovwoOZpg9IZCSnlMyQJD5DapTDdlqV5VpUa
NVDjlrSqvcLkAQJbWx0chcVo3pD3aeQWsSTYGcqJ4QoSg/o3gxwKfnh6M93BKjtLkvri1I/zdfis
iSyEiNt5bVoEXoMgVzlwkF29E+4QBE8FYEnvXUsAxbWAxyXMRFsb7rVxaChc04+gsY+0VNd4zOgX
11n/86eVFgiJNtOXaadeoxkhhimDpqMnlxhWVAFGseuP/zW0v0I86Dyw+BT7V1XU6LUmL9+Kfgmr
pZqxBP4hsS47O2zESLm/8dGhe7htcXKwwW58UNaCOQajem8s3qZ/q8yYdryiCkmI4Qi/Xm5OHjbz
FVc4lG9Lrz//xBbzOSxqBnnu4pX9dR/B51S6A7eq0pEzAxGST+YchQ1j+hNi7SV04bjzMGAobQ7c
5dRhcAaU3X6c0aOt7ZhBh3g1DboncMT29hpVQaOQmiDEqwXMvLnSrPHU6fAyI7WpKSx6blQv/Rt8
ngnWllCpHhJnv3NBkFd8jzd6Hpg4CPVUVnntWLSEu3K+E1eQphMuYj5EjO/WXQonIzj7oqX36vRj
MBk67vHxhBK0lENV4VPLwKzA1HVX8GFTpdCeSpLcd1+RZS/5Qy5bAccYjak6b/CaSzZgzDnmvN/8
Iy53FboHqzuhueENXwJBGB1+hjpdfqcxRaAyGZLz52PPc37978wUZhHerAI+CsyN6243sw26+rWq
qKU9RVL0kp1xCN98f2wH9T/u79M9iFLz4Ylr/9l58Hij2b8nhvdeSLi75PSgWqHNeEIo831DBrvg
p/qInYY8F0wbVMdCU1p4CK+lhYmh3uXWc7tjp4KGCLDTKcNHHY7/yCi7bHiJJb9MlkqOlJzXttXc
n5wpx+kZW+gK7OaN0MY62PVOeFZwycDtOS+qMAwsG0Z0g9HH/QnQAoH1JgGIaNnqy7sK0BBpvxN+
4DkOaZk9lm12GWzFgBkx5oaL6VFYiAq1MrXTNXViJ1NIrYZY2ynJYb2DcjGsBYGREQYlgYjYjGcP
G6b0j4Sr9e6NHZY09RbVqkLILUuXJXWmZjDLG6EWbsn36m6BlsUQU4rNZHVShV9twetviVuWpeXw
xeiT8be/GzV9snE4PGUbr3rfcwX9ks5oNU6sGPVCy5xWK9PovsUcktXNwcmr+3L4HYTZxUWVzt0E
iYI5luF11pcTFYrbN4AgAtLqjDKpkkARP22ikey5T1ivi0m7jUxu9L2bM/+Gl0CuvQD6+XDz/nFT
bJ/iNqH4bHLU7WzO4sqPXNNxeJIqEFS4Odkb4YZrJvHPQdjS67dC87O1+UerysSzbln1Clwgm8R6
ktVeFbXaon/tfHG1xL+rAVrH+5eMPNvVz9TfnXIfk1LZdYhA2ELVcYnBu0aJ5PTtjJDVkhrD1fNT
OU/y/pEU2KfF+Jy1TQRRtRD5PyChaEZ7WHutdUHoP3mrRUfLU734wNSX87GehaqGWbjv4n8Xg0m0
s5zLZ39qxdiepWBzvM0psJ3JGAJjj5OBVbFKzvS8fTHhhUaic9I/dRxNgTk8iNgjPZH/s8Z1Td+H
/KCfImwUXUg2lNv12nXufIOs2ioPDk/3afsLNXSWM23E6SSs9B2AMI1wrFiD8EnycL5ta5BX7z+T
xNPIjCSt/GnojrN8tNjnaP5MpgApkJ7dEBMuOM+uIzVpxmqG47bWF3o6T7PeruyJ1Oho2tBGocnm
DMzDe+3pwgUI30sfH5f2augY2soxVfh4CyFDU+RKr1hLjdPOKtUeuLnFxhcTnE7i9NrCoYJGDvaG
AV/85ODSVQ8Gmtqe/nQHt+zMT2iXcE7f1NTtU0r8EcRh7CcB8PM3y1Gbk+fRV1NQaaqAt2Dlhz0r
uwBJBKLEntGmvRJqLsF4gCXxPQ/wr9K+JAh1PNpW7l8s4KBi/uE2lDOleNfRJrrKP37TnaNrE6ou
Nxlgdz5GY8kPHQPO+3X//c9Rf//zSdMA1zqZhwNkWiQZGGmsRowJcSFNjaytTloFYmelrn5UucuC
JKdUu8Y7b8wYdigVHoF3J90KZNZ2BlOLJ085uTrbOZTihQqbew89q0UyHjShUNmYuOuX0lYhgFpF
zFsqJLjHkJtcVNC7s3Dhi7eUde9uhewExNvwIYpLdYFE88G9yTCtWoqAs3hFXZygeU3hGgGuJ6RE
1yGhos4IGLYce33Gm4eZnb6xIdojKHh4lxm3FmT/+e6XDAMPEgLHjd9WxhY2Yfwz7l8G7qJ2cENx
XIe5llFoYoNYvxCSML9Wp24J0nsfvaiReF7OjxA+x3PHjPDOEGD8Thlvjvf0UgxeucGwBzcKw5u7
cWd9RthXsHsUXCYBZ2gyVZA3HZmKIAy9MJIP+3vb6IF+zaTeQrx4UsU0DHLN+Rw6tKPCB+g0Ta10
FdBaee/Qih8YdFx2zUktrMidjUqSpgkhpu5LiKll64q4I8kbH3Li8VeHJSsPtWnUpqyHVt3laMnv
xZuRmO14vinmPi/rU23QFMkwogtfuJeb4Uk/FeBa4JrObA+nUNqvFzLR9//FFfeNaeCQm96pHUr1
pMN7f6XNs46zkE9KXNL2RNZnQANSufFhF5j1kfj3nIIFsjVGPQMV8evTKfFqRXZTWnzoYYoHYs4n
KYjQYNIlhFxdOS7xFI5a2TdEsf16IhGdRXHvNdaKwAATnnfobiuAA57UC++X/1oRBfEHjjJTxA0X
9kcodcx1lgs/wGoVplgzeURVMV1ZLPT7WNik/YPQqDhd+gGIZJijPs+15WlyTQfoMrMcZvgVf4SS
oCjIXkRSaZgialpkHbA7s2CWnS/01JlHEUsJg7HlkqAiGv1JqEDN8974nCxfoCCo6Zr4jlJXdZNB
+lSRfPsR2pKe4018wJ/JnH8VWU3kNTL4B1hm7Dq+l3evlPv6SYJwgOB3TA1ZbJOOa0A+vu/PoGRt
PuyrHB5/XZlQf3GKUZLp5K/uifnad5T+BvT/KKnjhB5m3OAPj52oY0X8hmqEgDAREKcIJvNEQLW4
+rxw39bTuWy4F90vpnGt2MITu1zqq1X4K3BS96T8FKG6+5u5Y1ERugB8X+3/9k7YBuIPtu8ycGBu
mC4iK3Vtw6+f+gSX5wrdBxJtJHoV/3D8IFmhS7YsFKN9Ma44k6+17H8SjkW2xzi/2ukicHqotJKK
y/nDjkM3FKCZ2NIld817rE1s7erN94o7Czzpi4ED28sPt0XSQcqQfGyBDUYL5q4DxXDYsNf+xALS
KDrvpiBomqozsaKUygIrBhAm/+Yymnut+XrcbfjTP96y1FLd9LAlNIfnXnLDP/L+MaPxiL3Ypr5H
nLzEHdq28o5REEfvBS/5sZtPM6zkzcAzmDAfI5bKBt/nmH9aSF95A/uUAka9GBiusSf8b1lyUi1a
UD6nW8qM9ZcSDtABhuJMTE0pniYnGjfwc0i9Cz0uxHUa6DMjqBLSDiS0cm1KHl8xg4SWGxB6hdOf
P9KdmDvu1IffDrf2HOg7yfGeOiWRRSH9Z18gPcFnpDu6N8LxkRpfb8gY4dSPD8rKHBXWmNpRv7RQ
H+KB8q+EGxm7VH5b2uNOpcZq2o5KDAb5Q1vqvJtgZv4ElM10+YpnF6Cs3tYaOpXSs+Q6YuQDco3I
h596348+HzdzzYissJYqkRq13h3tGYEG+TXQHYrbMuYvAPsgumDMVO/1E6PvdP4rzkw3yMjNqb1x
5HHEkvMVhYEYSk8kw4NXO/+j46OGmvPUIzqRgC4bQbLy7uo2NVzKrzpKVH5ke3xnsQqJVXfnsgIq
DCELIsdESJxLtYa3fW67jRItedyksnp05MyoxF7QKFRdUAVLus37MCJxeFwBprVTbPCIdSbGYyn/
h/qk0iBRArXeVHCMIXgPPNo8BrUHbIM4RLQElk1Z8/cB4awmB1K3hqgZU9SmdJiSTPwCI4rJ0UFX
mHLmk4rFoEaO11vNkc3fpZzjzCYtF6RbJ97kgT3iFrTWiW95in47/icK1yR05j5eMkk0pygb8Avb
nuM16044KT2t295R7JKaGpgCsZdKydgUKB7Jf/1WysMrEnAMgWBON52kEPhlA4KEf1QHqBjudmw4
qDR6bN/H6XPDF06TFkBenMFWdgFG4Z7KdqywSnBaONV9H59JYkv6XhTIF4v+D/AbyCqoZvzTaZNY
5zZWRQvS152X5qgNEkNJ1SvNrIN61dIyF/OVmbc/DpAQq6NYXNKT+Cm+3vTKiEOGNA/8XoEssIDc
6E+lwUecV0AhU48gR7daN6B0/xl7F7Kx6nI/cTTFMnfzGzrp4afO8pxwPxRCrjny67TSm4okQMqU
FoUaOXYYn/XuEDUbmvyUPYzuAphWEBtYDT38QV0nAOAUuR/ZpCtN00wm+EhHTsBfvDYRixXQH77n
LlOB9p3cO8r6TV3QxwAHAaMkrAzuShZhcmmjKfteMps72f5IMTv0YVcoPDDGmbHyIYkZeJXfnVtR
fmlLTUKTSJ0crBFQ5jpDVFefTNs0ImGHhBPQr8ESGXkuVFaJc2IKLaonK1RwepOlkv2326/5+AeP
ju8tilS1lYdQEkr1WpuUEb7im1x5OVwuSNb7xK7m3ZxQJxXW1w42UwBdTgvMKCpQdQzvmIBuTPSd
BiAG87q+zQGe6HLEX6lneb6MyiZEr0WbMs0KTBAzuiDvfoFqXBDvX40EyHf2Q+dGPaWi2tvhyQ6J
+slf9cjAJML49N61s/MrEgcEpT69aiyI126YSB45M3rxVCX3LEminosCK2e13g81BnT9AZWk3uRL
UEqZADltqhZyEW118VweqUr9vtAdnqx9LNDS0FNvsxe29W89zVRPao2v1l229UGTpLzxjRDF42jJ
XGXsU4nD42zbDpWFPUxtdCPRJdkhagHPc2kEXzSrvXrBgeDi5fqfP13Z7kvf8i7I2ZnTDF17tno8
CX+dzZi6NvmOpvKywRuERMN7x0nvEKR2dfZiCIn6K3LXYjaHXB0ttDWcCfrst+dqhFdveFS+Zo3b
KdldBoBKvq+07m5BTBTeDz8VXilbTrlsFE1gOgqM7QWXHKKyq4U/rNEbVx7vHK2CvauVxznQElxa
j7KtwjorbnU3CnaaxPIUbmBXyOZw/3CaU6Uar2ekZ4VptphU1OFkLbSV7LVDCJG6hQerxa95Dbi7
ncaZJMblk2a42jVwfiQyuFI71yBnXHWCoJxskW3IGGfeuKmXyAcQ7/953AzjZurlxryskFX30Qfh
6FsoeOSPrtqvIQ3/6mMrWU2dfwxxsHrTGExJufOczN1ETYr1HTVu3n1qs99SRHiyQ0tENGCW46Pp
AUovPaVh3ZuNHvQvAWSHEh26Ua37skedt7CEiZmfxwo5l9eSTmu8YfdtakhDgJV0lC965KKrqq06
dzhEsRY44WIr2vLy3NuD5p8DCL439o+UQ1Vy5lkpnOzA6GCmTLADk1pxUYyd9PUzYp/EX6FkVzut
uMALk0C3rT+V05q8IP8tgkuqv3Ky9B/Xu6q71FgQg9gPUAkxz45Duk2dXE1bzbMZxptmHR4+kh+K
W+whyYOevJtnFlPvEsMogc8IwBBm2hrIH9R4UhdsGIzMNXYtegoOLkUVRfmdGqo2IE369jWeYeqz
EANLe6qpHPRAZ0QjC/Kx0HebxKoe5/voSMTHIkRtg+2od766kPXmfLboceAWsolxAkwcZ2teSqV8
On0zslX11aerGQzFKdGZGN8SbCAfOGWIFcAtNKTijkvipG/0khgWOfTh+84lHNKbDjVjNeNQI7gL
ayVXI8+QHSy1Pr6TPk8wEL4kTg57y7XhfbJQhrbV02HBIlBFolcc/m+xwVrP856sV3ap91pVfMim
QaF29f2pwf2+l2ynKb1/U+9ny8jjt1Lz77k4GJs0UU4N0L5WpceOsAOyfDbrYmluKAT5fL21TnFm
TjQngsEdCYhCexdB/Ku3/YDOsaHHWhafq9yZZgajEXDsxQ1lB7bU4UoRWlatb98zNS4P0Mp69jqq
1VAHD9+op/55mhFm0JG0mBUZbu4Nr7U7P631G/0P1jpEkmZXwFObX1DVUizvMDD7tYMdON6GuLlD
RzU+Lz+r+JkyezX5CYwpttxaDVglq8ALrMTQYzgq3IiSEp7uenLDKofG3GDktyibnCTgGKubVCOa
P4qGZz0AIQ7jv5lm8dQoNSkM5chsD06MmkJzldkYKd5XHvGiRGfci2KhSzJhENCd2quYULrgboub
Ifc7yVXTupMxhNi89zWn0M9Xv0BanPNHPjhgRLt9hW9qjuKZf/8mgos4oT3wWK56CcUqKUD7YR7q
hq4S0T4a+qBRpwfQYP7WcIHY2glBnxMEnPla4AYBZhJPPYwcRtKWdBuwg7Vy4tk2DUIpSwsYPpV5
RUHcT4AVV0/G/6Of0lUhiTSBiCJDoQU5CmIyG3xHg/qYRhdjOZpvgXVKH7rs/knEeqWRKf1GsG4Z
Hw5urKaSb16CDWlH6Go0NpqOgKYSUf/r4Z9286+jjgARJ5IWZi/L52gHssJU+Ij/fHA9i1Gakqqj
DNRV2X+V1OGR1/TRcj/r1tUw9b4rpNkL4+X3Blnjk8ha+v8PvQu8fkrQwQSSsQily7rvFYmiH6w8
VYjeFmmrrwe1AYPrphiv+q8wPDyeFV0PH4+sODeA2CeIX01GDdogk1HpPEB12K4JjQx0qCSYsCiU
fsbqF9X4AtMu2flnTUtKZBcTpHEy2SzQjy3WpZ13gl/2Z79JYpKVGubvULtrqT0hSmsXsYXesBT7
w8OX8dLnkTStE9Xgps1GNhs692AJOKPl9GmVmMpMz4sNzBGpFae8ILunJwm8Uo7vqOGS3bEWCMwH
ttF3J1cqcnKD6KYiS04xBnLFz/hBj2vSGtBDZTeGnSIBM9aA/YhX1l/pjEjCGC1qYay5ZOdJ1GYh
6ZaEdJvTOVass4dZ7XpUkXyt8wQNqD/bbvp5OZHNYAA/yctZwkMWyt0TU3hIW7X+p6k2EhOSPhCr
55HeoaRROnEw5PKI4d1u7PuraN46gOKYeSuml2qQpl4nPojWxhf/BqPBnalvdp5ziydap/svmpb7
3V2PATE5SEN30AGYg4td80d57hq7GWSRhfsa5GRQD4yGWwa2KAZJHsjAHx9YAVERD+UB4vSiIrot
F9ylW8zGYWTaqr6fgPK8venoXqNPs/GLZ9leA6p72Mj5KCZTvy05EVhIjGIXXkadlqeXKYzihCuu
XvukNtAZThFtzJBAOmpky/YSBu+Z7W18JS8w1w4vilAXXVq3ZoUm53/YkByXTo1Mey+3MZImMnug
T10ZEcy9wZN/RUoMC529FP/OBeeGKXLgDIxHy9Mhj+bzxEsgl7AqNTWicP4XNV7md8WcmbsDAPeQ
OxvePTN12BhIGu8xEX8eZW3iAODCgRMQwGNt7aHUYJ6ZYF34Ag/PLH/0CLQyV7YgUV62mWrryhaR
0bAEzgT/Ir0CehPHN7oJjzm4Q1D9MC/7ILukEjqufNhj5UpQnRGCt3jMvAZU1DvPMv4SR8IU3jZq
sVhtDPIqmWEmoh5rL8Qtx2CVnlqGLOvVAxHfyDryXDqDwAXQbnd2lFXtlI+vLGOMDSVh07Wyuku1
bOD7j3141NB/6EkJz0HqszOCUTqkVLK0jxGt3iH1toWJC3NAtzG1qIiKKyWACqO3kbjP0HzUUevy
vYM3yOD8fzFfGoxwXilSpfqH/q4QPH8jWXFWR4EvzIf/kj7dJMvibUyxc1lony0/g7MbHC3Qnxqu
45OD23xxJa7RbL0K4a7T2BWNLITQZiTXzrd4b08LNGe1LMw7GF3PQXj/OErWfiK8ULV09oOoN10w
ThP6pHrf79vO9+mG5JCKMMfgK5kJF4PsmEPV06e8PBKw8tUigHXA+7YM1t01dDm0dpGHFB37Ht68
kCEHS4c8x2TB120mZaszBhHkD0DM1nEAZTz/b51IS+2QKpo8Wyn9nvNRXEvtNwWvQyF+tCEHgN1z
WJcoUrXzJvPd5rXKLb8xWqlDLTAq72qO5QXYuUa2/Dz57p/8D4kf6QNZuxMLvZW2+/kKVUaaczLJ
LjUK86Mus4Fb75SWW44UAKde9E7ivAncy2vX/NgULRM5DoXco3v79LtBre260cecoaQrJZNTUlRF
97ewndvyyLzkTKkZ2gOb9leSukxoro4Epr/tl/E6tAiHCufPqt/J9krfHrZg14nCzO6b+owvihl/
BEk55Vm+xmLTBIxq+WOTgcSA/PcPjaLMMq3/NTX7AxiR5P4lIya/+UFxLUK+Yt780qrT2S1vperQ
Tgscx2i91JelA3YYRj5RwGymRM/nvxp/kTt5DUk1WHHirvAunzdBGOw9G0Nw2DyOG/Xx49hRKckm
Oiv9xIVQVKPpqnbn+4vgFYLbuFSazsucoAxKjHj61dkH0KSt+ZsgP1pLX6t3RBu48u4NMXhFrzWa
Qy3dJFPqaFtRcvK8315YxPamVzOzpypzgfiATHqi72yxcI+zx35Jel77mzC5xx9MgTx4DcV0/CBO
H0qFCE0qqO5K4VuDI37UwX2a8UAVN0DNpi29xDBZlx6AjC0DH4p/f8KF4zp05gNnEAsp+QM7ABwH
GJsxlvDKJSIb1gijtXfKnbZJ7t+3ausiluh0j4h5dYtklxWM59mI6+j6CDxxQKXMzPYXXvrOrfMe
Em7obhIt1hc3AYJAYvsS5wBWxSbLc+TLLf54FoOCm9bCFLVzq542kcd+8awlrcU6IFMz/2sdgTAP
O5vGpqWHceeivrTJwN+9LDzbFpVVKj+4RmlGzwKUXlxUyQ60N1beMYJ4jyfL0HLQJf+6JbYY4akx
ViJKQXHSVZsH5xypeEyxAo7IKnFGuHMxAImCjSZvjot8tDXBKxK77EoVxqw6oqTO9+InbuKqQ6qD
G8aJPRDGUZ5RP7QFekGMfBCWiTZAKtFvSywdXXt3YcQOjx/LS86rYhlNYlmsq64UDU/uVAqE7jm3
k+7s6xnWe27gUyddwWYujORtgMixZ5O8K9ArcZOLlsBuOb39uIZYYj/dSC3at6lYt3udSe0fRvmb
pRuXo/mXT/kTmOnxafXfiVL/mWP7eiQwWiVz5yKa8XzTCk8WXQ1GwrR3ZdbwsaeEMq6wha52/tY9
+jtsxzktNTwUNHKueyX64UGnmANmW5oo+SmC+gYm1bUiLzOvZMWotKaf628sHXmWdIlprKX/TdFa
wsN3mFFRWrj/xXoGnjwdsyzusIBR/6wwBYJJVDf+4nH3QK+4WHXMRmPteEID3Ntx0OPRMTsfY733
jDAcKJPhYIYlKUByFnzktDzErJ8zxTyqNlN4BzFeHjb/1JPNftv5IMSRKkVvXyz8VxIon4Q/n5yK
lXanG5aGkcnNjCX9sQw6BgWmyc8QiEMbptsyNkQr65MYyKCgrnKkskbMlOJuZR43rSSS3RZxeJoi
kSN/GqLjVc7eackQg1SvxCttvHhUZoc+rEkBHz0dJwyMHztL7UrKTY+FykRBvaW4a9cR0aKVhBu5
grT2PL7+bYKEVB33rUIhgd0O6KlZT7mVPLGlNF7rhTOjDpO+eiICN90gu8widIeHedqcz9mj7Dkm
Pk4tchH/PWL3r8fHL2kW6o/t0xfvwdFjoA9iHdY8NRw40bV6i3jjqMWBgDiKCm74F1siq/zQ4Are
gDazIjI/EqwE5RKATrMFCePW6e2OO7t6qTIbzWLiKY1koSZt3nGcVlCnQMCjavfRS8nOf5xA7vEG
BzUjnL2hD6HaQnHh7pQ86ExCr3t9WYDRK8YTOH9HZZTct1v8h/CNSq3mWT9v9CUGAUTQN5Yeo3QT
kAq9Yfz41HOOkl5JhuqtE6Iz8Xft5hrpIh+Pp/by4B9GKhh7IC39HHd2QvYCfOtOZeF5sUlnzF3a
DY3SPqxsdjQFyIVNOHbl6vO11ftcUhW/6AiBTl7Cb4PMyk81CZB82PvCubscH1XIrVQXwwfP8dT9
k049YclZOBlburVrsghEHWIj/fqMOfDzO9PHlKtOokZg19T7fprpAGrg5f6V/YYZBNVUqL/IKanp
RYuzt++tN4ISLcHHoVsVGMbpy82ThbUBsn3ajZABXQSoq9YdrdupRHbvr3nIGQ1yt4V3LJnAPlcS
gnBiUcG++TmOdb7AZ60yTexw6/17A59wNrV6vpWWZ4N3vTxOu8Vq/iwdp2oN4Pn9IQqAgB0K/Y/x
2yRs51I47HTOISuTraNQmcTfxc8qleRJXzxP50jDQPqCpXvWydDd4BGgDsqcwFWValN/r8yByLFp
g/Hqg7TZa/350kPk6pgEyZfDUdva1GvmDkb81T6fKoIm1KZLoEeBN0LpdF2HFyLDxBUt46oKsO1M
IzERKD0n3JADHhz0yU/YNFDMsIvaeKMFjmhYPE7Ur5zaLQ0WdjIna7hqGEmegiwTOUxkYOyKYEcp
3Q4SFBhLvX0OURFrRci/PVZsmcOW1TReU7Q53kSGaY2jSeI1025in/FTf4PJgc1XxxdC6qnHalLg
Po4JnIuldgJCZHhbQ31kY2W76drne3XgVVlvQZV1s4hKGlBkPkoa6Rbsmx+2QmY3o/cJFELUSO5s
XVnjmxxW9sNN1y1D8s8Z9qShwBzPonVZjX7ERU78WUcRZ9v9roOE36WyhTfRVu27kSHBD2r9AJbe
+xltbDjAwDp9LtdXvLhYm3mz+/ZQFcvwj7IDlawlwpbyL/KVFXNpOv+5JYPr1dYMvA3EbsCv+9dR
0mzeU8u+CyEaAeTmKWVubirhOE2XB8q4OkBGPyNl4i8NPmDSbhXVPM3yS/niht5/s+K6JK5sCoWd
IM/923VHks4IVGJtY8TXPlbDYWJw+VYKlt4EyVbYH30A0X/HhAdLIerRjdQvzKzCEYmBK2nthQ1Z
GV2xn/EgKQrAv2zmgSMGYz9sWx8X0ofOuMEcz/gb4NGx87riWxRfd/v5Fxk7cXHSnluWjkxp8PuS
YW7DABmdzTmc3Xomn4yd90xzkO+TDyuo5KCNiwCu3+jOv9ewqR6RJl3LpErNYMSFEjH7MzZMsedu
v3HtSpW71Z5kra//WoluYkPSoIu7L6C0HRfFqFELTZx4eosNx+WW+g32hv3yxA5rTkdzXjqQsp/z
ciLxOh8EJsyrNw1MdbcZeKG33/bEufWhtZH18idV9h1RtnEupC0kt2JMg5+qWtMbwRv86VsqALWu
Hw8Mlrp6bPN2+WM4qbWeMaUj9nsRXuG3Krx0OawxHkP8KTR29yw1ZzwUCXrWUJ2+Z4adl+WNLP6e
p1KRCtPl8gyoPyFARia1hsixBGJ0piDlAFzgvDDnBEhXB6DKCyEKjpdZktXWWowqmSF8n+EJmTJD
qXuOxPYTICTfJRCp2neDfv8ieilj9RnKEf/IzKKBW1fv56yJzDCoSfKZila41pyMdF0hWZPoC0sK
sK0DHFww15zW3i7ORclbk7ufIKt1BcgXPHZa9hirtWIN3k4nr8gf2KO8gP85ZbbJpTd0ppX4Bqq4
azKgi2SXw6r2pAWnHM/A+Y0DWEFSsE+nPgDtEhHNhyj8LMlU/Pn3iohkpvRRwRbR50usKRpSwIIV
eQMvAYBI3c4ecntsm8PhT2+eVmU8Ay7tjM9IXp+Ur2CWMFeEzIn+Mw0rnhrPmMi3Mr6dRjimFN0e
7IossSdwECEx+c8m6+Ao7lwxIAx71cyRQYI4WXQ/ttl2tiusUx7jTidF5R6+UFpdsNmBGsb+dRLI
URyDrp/nztN9tcySU6eK269v5cqqRSmKyFGbw/qdzWybzyFW1Y8Z/bBMf1J4bU4EAl+EnuV7AFYg
6vvigvvabOWS16WE2jFzFk9JEyWyu8Ona/sHAR31HCO3A4YUXyffx/nuqlJB9Caoj2T8RDcLniL0
sxBxi5QiLUGHE55BR6YDMIdq0BTc7NUcH1qTrynPuxX4pSh1U+SMiLM61b9iZNhTh7wk1YYhSPAZ
f0sxtOH5Nu8gqX84c+bKCW3l0bmu35aknZ19/QzypTT3HKrACB6ab9kIB08BTTkrYkIIQFN+o1n/
x9ttB3whLv1pSttIlZQ0bI3kCOjYEQEks9uQ79qOfHDrnXrS+yLLCIj2fKtcKVP58UdRFZan/E+Z
+tURZI79aoodHKlLB/4dSx5GmroYPJyVNG//rVO05EJqq8/gfar+dKWnMgMeaUqpC1b8zU0eQj7w
2yuSJqktVN5nKB5k61lyFLYinYNRo+vVe3oZ/4YT+fDJywZ9dZlPNdzQ5UVGXLPDLn744Z+Hnpcl
cXecpoPHZtRq0ty0oIs+LrpveHX2ZDUQvHvt+NrEtSTGcXEeRLryhf/ZXGB6a5NcUuJ287zBJz7Q
gzKN8T5JTu4YQ5CDt0pZ0dw/mKoZRT/XM4Lklu3SkoBo3OkGtCh9Vbb3ipF9ogM8DHU1Gm57hyTm
H+5dWZh3G4mrgeHtUc3jndalQLXC5fyCV4+cPMXUFoTcHuJR4Lm8IQe56JUHDk+3LpRM84llgYw7
aIF9J1mlcqZ10xP6fehmosL1QA/UVIbHINbkNjl/4JYl5ARwLPoZA2CFes4PcQabPf5eyackwLcY
0PMt6y9wvtIsnNLxf29rMnbNp7i74Alb3o0/vS1TFVSxVmt4uUK4fr58s4LTWrvycy8iegcJ92fN
FXplWXexmksohkTMWvYPHZFru20DNzH8u6jjfj+JZNgEMU/M1FENAJwhvD0tIHhaEqYNg3wcnBzH
3pxLkdX9KmfS3uDGbCe760QAlHUh23MUWhJ0IlSOYteqjHOYmkmnyVm0AxPdpR6lqm2aBr1yt8PJ
05uUig4pwSjfM/CN8T27FzKG365mFRcJlt4efAIfguSonVQo3bl5O8dHqQwE+bY3POe8yHUvDEVx
OK7EwKXUjk7ENamUoJ8ls6PaXqTEm0BDUBSkNYgwGWQIiaKUln7P0l+prTgX4l7vqtv8kcMmUJED
863kxWTueD9JB4KWe4HT6X3WU0R837i6EDjtu/OWYXDPF1mVdsf+918vOpVX6kejfYc1972D0uoH
UzpYQTtz1D9tD4xVQK7ram/BVcHuE9oi+05STMVXr21e0jost0bJIM61yjlFRqOEXUjpmK+7Yyug
BzRDDiej0LMYrWwHKaWAZM9LDk5iFNahQhOfOHiLEW5IpBHh/TQi3Wczsl4qKLJ9qjKHU9H5Kwtw
KVzpVNdqAjVJDKBYcSbDvUPMEmUtsKNbPhK26wrAyQyezr3Q1j/7iq10Ji/zCnoxsqKRmL/AKE/e
Q08avo2wnWlulnPcUfe2ze1QA5IGp9ABfshGOiAGk/tflPiARYp9txNQUkAmVIJ7ARmB3PR8E0/N
uqUwpykpqAnoWD4+oW7uZHqxabmHnX8Jjsz+MLhlQLBzLL8Sk6I8eGwllRB11z8rKsakMGwuWLMb
1lh4V3KSbVltFPPjJXHElvQAEspCd9xXt7gIvRYzWHpor7OvM1Ba20JbRUuRQdVridlGELQVuN8M
6MYtc+iJXzzYBiXc33986WY8OJ1/H8brXOFsjExabyAFXT+Zx4Rd+F2M28s6qA7vTWAPQr3ut4yT
YiQ879Ldky74It6aGP7Xoz3Wh6ETfaSbJ0zl4vUYZpI9TH8tL0HentxxKbaA9U9CXCNx+s82Ctvs
PBXL8ritIxDWtKHPsq+Sezh5RAYnQIn4LRsFHr9Gmz9XeQyyL3LT2MEaKWg/X2/uOow08wutHWy2
bm6YQjXnZPDRb1HAKf500kk+zYozkYVn1X+FiAO16eOwiNMaCagqFHLITV9eMVoNHr/5CX1dgRN3
zmA6odhUQJqBaLRWU/Py4dTM76B7SS4Q17c6bfOFBueVrphUhdi69Zz+UuCtsMpmhImKRoMqavCa
nfHHTCcKqNI9nXfo6eBTXS98LdKxDJILJHvy1RYHIpWf7cE/iet9wjOJSYvx5FZL3Kd7Lin8Esb4
5He3HOqG0TA43SGGw9sZK2FYhYodPWQ8Se9vlJ68XiUYWm1UATbli9LhblEiqmc+xeUq/u8gEoc8
7yqndcEs3+/JlW0Kw9pEeVvoVHL0d3L+vELeBTd5SPbCP+c4ERy5cZNDYOc5TY/KtglJJxt7qEfr
A951PBcjhlhsDkYOl20vAHwu/+pbQHOfiBrU254izvUKuZvRsD7W9xWvNqEw8gIFXORyUjNUz2ES
BdoR70qshUsJcB0wbQR6SDzt9E3e0ZH61Rpv4F1h2QXs4Xtta8cwpbBYwgPWOR8s2X2hPirb9HKU
Txh8rKKDxuqiJxbo1iMg4ROCTsCvD8nbBfBEaohWFFlmulSCy7CG7wAq/dAtQGBXHuBrH9GpMm0b
izM01+bLY+fwScPfqiGeAk9rS9FyJ0D4b7b3ljg0lH5Rt48HJDrqOlKiYm4wapSDXSVvv/qHXOtR
zqHxoD1P4PEoJd+xQUqliERoc7Hrr6pyH542AYm/amdp0/aPQ3FrFIbhFfQsADWZPP8kMqUVCXQu
VfVciDd6W7FmT2eS0rctgBdunH4w8ek4aa0f+4dInAl/0etFALWNTB3nszhKIGwsCwvVhPx8/pYv
JzOvjUwaCJIc4pTJR6DOU5LMYIA/iSyIOTVNBYgzaQXlL7ZtO3JTSTgyqaYTPnn+s6Olvp6oi6cD
KIqVxfBMB5MQBWlFnRbSWlE/QhsPRjx5EutCl1J5pwqE511GkD2cmvloWDH8Fo0ZbGC41D6Qa+ci
xoOgCpNqhtml5ZrbQu5w/235m5EkeNdca1c98vOhY30z6Oyg7FnhYNbfta7xNfnDvPNCAZp0NtQO
3c08oyPiQN9CLYYV2kPToUNWf+APhSpp/MXRuEwBH9YpayRmSB/+VdkEiDRwKfSZoXc9hKsqLMaz
na+iT6piJ7LAyL3oxO91tnLakvBWAqKLjbSOWfHXLGWmrDkAgI9aAZJvdgGpIACu6YrVrcdjpJTK
TYbuDMxGRyFOTBj5wxqIMyQcENXZkCm/w+xtsywbDkU5bD4EAnnGaII5ulejUdiqlN7Y13iaMCE/
nPObs2c4Jvq5jdZNJRwZKh7MHwlND7zAAnmtF0nS9Pf1kdPwQStHKxmS0Mq8Nv7Osib7q0qGc8DN
uWVy6QMLxx00S2L5Rxvc3s9WX/RJK0ecKxLH4Sh7OLlnW+NmbvFYj/B4BiO6GwWqPbq5j9PruhtK
qz79p68F/LLZC+ksXidS8rqmEUvOPd0TGCM/MzAdnMX9zIeFVV38oS4VlacnmI41P1Pv5BzdggY2
L2rhVuKAnx4ARSiDAt2fjRWWVeu5FZw5lmJeHJ3F4wGt7PA2UNKoUUMuivwjEL5HrGHUBGt9zdST
ZU9uOVCzsrbjbqpqMGhypWQo9kza28ZDHQ2CS1MMUP13VSaVlXHRNXR182e1SyMhbTJObLA5VCnS
6qlfSO5CPrdMRaZlGyZzI4JaBotrjlgOoOU1v71RoceQ3jwNaeQYI8kRfgxWFHLOIloqBFzNLKlO
DJUw0o94GQGfUNyoMgRxg+GWXdGpGq9Nv0123EVVfvFxUAvg8u8e0Is8NNv5tk3nqEssNmmGBKlE
yzwNbC+0tWx7D6vdSyB8qhJz6whgPaRWNH72fdKQzH/ZKjei5PMRT5L0j0iiKWAm2CrqOhYgNa7r
6GfHUE9WAYc+L7KNt0Thw2Vor9hVTHCv3hfTdheR9AfPuM1T3RJoDmty1a7bwqcN7NS1wTfM1HuL
rzB3XvTL0onE+xvqPABGyPeSO8i/HmF8G/xJExJ7KV/4BTqEa5/vZ86R0eOSPDxnMrqXJIMJVB9k
s9atvex9lOh79UgUhKSzo08t5QeZhvPHIagkAUSeG6JEl2cgpXfh8Knbl78UyFdJWjzR4/wA8OnT
3SMu8PFWs9a9RZw0n8A2rhEvW4T2+AsIFR0wcEhQkakSaid1a/u5oaHZHQ7frIf2vGTbaft9P2hq
dUOgTCnCafaPzk25UJJiU+XZ1OiGPnnvdMgCFqVMZfAXdwUGLSM/oQ+3Ru4/zHnZnyyjk2gGwL6B
X26QvL2TSod48FzVpEYgaNnnSc93eMqqb80l0Y+xCLyyeyF5QLWGDPm9VciQa4Qc+Le/ANY8J+7w
2sZfF9bevGrMqT9yNVdhPd9u721TOAYy7Exo530nuridxRI5PF3ccUlLz6PwvWli3+ER/tl8nmcE
YOECngfUh1H46VO0Srl3pWYL0gma7Ls6GvgtJtTE6hXh2z9EofiLbMpsR/xV/gdXEPCGl7FoPmII
VQ3uUNw1N/t9AUzm3HgQQh7g5itT9mlovr3aopFJX9d+QDAU04uK/GRH71eb6Yt0E9WSHG1yRgyr
A9IfZLbJ7Q/iLELTIYWMKJnQiz/W+ZyDknfSjKdQ5qrVofJ5KUWbDx5hoXMOzYwtTaqO15Eu05Ns
Wrc/3XLvwd3JGXVg6l3OnV2MOUcBUIcGxQ1ED0THEmQ6Dc0qPQ6Uz91irWcnNpH4IyWBy8eMqXVN
tlaRzCNTMHBeThsE3Bvdtnkpt7D1HW0v+M5Ndm4v9Ry3pvjCKkUxsGqfPcIF0T56uySLUPNY3lFq
0Qd7k0jVu+50JumUgIaMI7JvLfyvCQsjZSnzLDN+snoipsY7h8WVz2V8ixDm3bEUfAhi54gdkvMA
8IinvycMPYhAwzZDI+2QPTqUFCW8btz2vDRqZ+x7Ys8qnlCiv32LK4WDET0RqT0GVJ5u1/boE0yX
wQP9b6ooy+NHpd/n/6g9rR24LM8gDB2IRXLAPgoNu/jFd1JGUJxr5LlhbkMfQoqzNUKtvKjsy9wN
XTmQsumonlxZx5KDWh8PXlH0FGF24qm2ikI3uDHWPDlY8GdX9KA9Ri3fOl25s1lwWGLTnvAFiBQ2
G1k8hq8G8h7gwb6zrIp6qMhpS2mwGhatZd4npRzFxJm87MTPQRWN1OcXpzWO5jmGPHgKiI+J4Kyc
JeO04Y8z0uRWcy97JhuXgw8pQY6QFafyLwAiNhoIIihbjxioWr3+pInFYVIk6kuuAFz8cdJrX1Up
lNKKZEkrOL7dpcFXC8WeQoobmcBPX7zLmbfdH8bTmf0i9DDtdy9wI6ilD+igIvEN34e9Vw8zHVkD
jNwN4waivXtNHZ93JGExdr7Y1D+Sp7bo9b5R/QvBwq9VdGHcedkvVpSsx+bd7O7NbE18HRD4uQNU
u3VRQbtQLgyOhOkC7rBC7FvXOQ9KKE6aloloxTyk9++zZ705PQfdmBoRsghriUqy66NAREUCY4OA
61a4HSa/kktg5Lsb63bKAKQTjtydtvdssk0lEND7Ftg4oQbTHp57E8uk6UuXlig0mJExpK3YwksD
lC1MuiGqRyZnfZIKv+r25spMnuZinRUmsthuTJuZuJ/Q/L6/CyafwDfe928ZamFLDNPoGUZy+VGy
vRhqgI/1YA6vtXUZ4heSdtjHxxXtz3KriFl0/YMrdNYCZR7iWx/ivZDcFBRFNN7k8tawgPHHiQDq
P/W3ubvi+I63tVCwGV8pjSCfJ9A/DVnKLk3487rP+/6FY9Bwx6mMQesNbYznq/lSCcTTm8ZfeYy2
OJDdX3kZ+FjgJwuQQf8EIRv+B9KTNZaTzMO1rExOpbEk3FNmBddZm0PGRS5j9O4cOmr0FWYX59NJ
4exAvF5GMD03bXKBTDN4ZBMKp5UxPe3Yad5fAfAWSbfoWP8VRpfSQenKG3EtIMLhYmvinbIUVjYv
2xt1aqg+/ZEDNPEeNo5Z2WcYTXkeu0BApBJLfMd+utc/IOjQq+02mJVT/5jxNDuqy++Dzqn0Nt9d
iFDQ2oogrLgoBGwp0hZ8xmXfnw8wgjPcepDmMPQ6wgsOaOq8GEnhe59eF5e3/QpWATIPGKvXwe2l
APLynh4KpVH1SiQikovrS1BUWfa2NbTN8mtjfA2DimsfhEJdhbINl+kXGz6n4GtH+WlZRyD7FIOm
ioTleQW/ZFiqZ0tAOQGxjclQF5csmAGROOknIyJgdAfZLYxNQk5sEtbgidn9JS/cGv569OJFu03Q
jtxoeGsTrZKJVVM0c+0Qa+N7x6kzZCBMRatocEmQ1mwbRIG1+pfZ/eh3eu9DhabqTJ3Jp6anmlAF
xYsoBmblyL6G23auvzN2HZLQ4L9fwpkb/sDwvQZg4G5iOPVYgpHEt6/5IhRRvA3HJyD0IrUhXsfp
6qxGo5tU91OZAPB55gqZZYn0O+siIx43ZCGsp5rAGzrRjD409skg0TZTY+2FT8Ed/xU00ugD4J53
Pay8z3zzS6l55mdqWH5PckOV/aFP8KhHb8vuSXNMMUk2BfQdRD7ps0DestsYjCJee3jAaSfTZ3wK
O+NSM0qQ0OhX3jY6fESWQYNnpPRCX5FoEYCT4LJad+0ou4dTEdf2sb5fBygZLK9a22CbHx8O9KAM
0K88TbvjFt7bblXiiYABnIFYsMRH/gySF4L8R1swELwDmHEntvXMevAZr1bPU8aoFz28FhSS5swG
yjpLkd5TFbAnyLYKayg0mfYwLzbKa2F6lSZK0MxCbw1/n8cTNbAL5mDaDc7xLNGYmhOdvr/TQHH5
XC3Y21OHx5OFd5b6YNWXlApAyskDGks5Q4t62yewprz1rB7F3e2M/U5VVxdrmUmXIpcfj4DnPeKh
6vezG4zl6OXQ4DkhPsBkj0gF/indYiLAt5S8iZKDIflcUJ5QXihH5HB5xMma8DAo4hUJuNPwGEVj
8Kpez/oVmfzJrYPD9tUw6zDlWCFCc/BBqtAjNU6EXxQr5VXcZg5VDKDsG1Du3R7ds8OpoXphc1d/
WNCZKLRUICCkDnUyYsR+ZwL/F+s3CVNsDgowvoMZouTH+8Q/cLr2g76x3ZbiDtmE8OmfWdkDaWOY
JfXxpjxv8UjSOPdYdb172dNHTTTTQruzxUuqC3ygqdB+YzdYMmE/wnRj6BRaYp0fn/0P5Ew+l3Zb
HQpbXWBtlOOERcYNzrDo8EnqCwcXPc3gK5Z7MilLXln7LF/YqcKbI0xgV1oH3kymjr84+pwfXNXA
9k6UkfARi5Ix60CyYsUUYUUOn1PqXapyOMAmGMhz4vTzyP4He0Lh9rWjYPkTmD/ijOHFi+E+k+Xa
rGyu3N0EjcgOo+UYttfO620inoxRRDY9G5qTADtSuRvazQKMr8/kjlfUredExT6An4Lw6dHkca1Y
S1YdygQZTAUQX3qREvi9bnttC94+cmkTk2xj2nlYA6hoDZdSJfOHVCgBxdaaxpHkOMACehScnZkr
AFAYwjxc82P4dHYbreL2+Kqz+8viuv8VvXoi+exL1SO4okX3mBkhuTHq0EWnRwZP46ewy6eBYmVz
yjoXwalAViob7hzDMWft0s/3pM3fkPn4G9ZymjKgz2T9jsCCwu6zCgXNLZvmbj7w4hFRsecHuVOS
9iGyLaZ/z5qZ7pXSEoIKvEk3vtEgM3/nhKCK1BYx3Jbqv1cT9gfuydDyyGjktayDoQRGO490Wf56
VTbkwseAFWfd4efUpesakHwIXWMoqqLfZpnc8/QJ45vSPqxH1tDtyC21hLXUqmzZXP3Qjj4E5F3N
Ln8g9MF1RPfEnQsPuOSyjKWqAbzXQdwSqLpXyTfnzJpfVjwlTtZNfW/6211yBV4HjhzEPcbZTV6K
DckNH3QoFrbMwcVDVOuVMeK/1giDEzIREHHNlZMCbAAAQgphCVYxxEV9JR0zhdgC3IUAnMf4PvXd
Ibbl5YUJQ9MEVQ5F0e3TpUclv5MwaRI6PYDvWBluAa21uZYM2cB7SuXkCquJ4IKpL6RZgxxjckgE
Av+ozksFyBKWBaMDdt3ue0l/OYVt2ju0cOXS5Xz5/+R/mD71yZ110IXQXos385yjmTygKHQmECy0
9FRJyiBtXMqgE+QYKAPVy65AercnjWZH9bi5ui/dxiL+CQxD6DrOVV9WuMprY7yz/M05u/YsYdOz
V7eRbgJT9etGMN5WO+zSIEigKIp+Y6fK03zL6Zedr+M0K1nTwt4iBfz6PQYWAXM2EH66gsT8ixGX
T7po+eo/vA5uNJ7ACrn9niVKLJaiEEyv70RcN5o9dH5KiJ8wAxIuHl6BIPHNqjnsC2uGKETvFbWt
IBZaDr1hoE1BF4H5ivc/EnXfbAcf7F0lMOHly9zqijI3pVBn9HSC6g23je2p4w/RMzU/RW5C0MVK
TLQOUYsJlE3Kw+/cCGvqN8DIGp1NOJ4dBnR+BJH40KsvJfk7wyZREno8bHoHcXDqH06sTtxcv69R
gC/LGxEh5IAThW6EvP3sz6TG2BBEjE2MXCbGOJxK8MG/NjAaMh1/onWYtZyZn6wgDqWL0WTOKhXG
gkxztFccmmn+5nqDTGftc3JaUwxr8Ov4LVLkcx81ZCTdtFFRoMeXLFlP+JjhjWHUMnTlQHUjKhEr
Wiu2jm7MF+OOHLalUHiUG+96lloUN160542AUxdCraXWi8B4qOX0OlmNxtBEcs7tRmUvp4XexlWT
UvPiGwzC9j5Ff+0KtGbxgfYuh0Y5h4HlvCHlfftjQ0UPR7j/f4yzltFRp7VGX7A+ndYBJRY8dTnQ
X/0YoqBr8wVHmpU+nkz4bfTq1IGlKabU/zqpn24qoDpo+4GwRl0DkAYFtcvFufcjYJp1Dmz2l+5p
69H/evvatTc9E+LF/w9TSLquCJWTiA1OH2YSGCBtnRtwGHyXUTkq67HYYOuH79YzIUGXK8jihvsb
v8kHb8EE4SXiGwqTRoxpQy/BwEbRFY0RR4f7NxjT47J5MUBIBZthKs7H86ka2niyFJODEeAeg18z
YeDtyfWRIOmUDaJjC8LMyYGZWjZUNKFl4lPH5GpgZ+BhmfjpXYJMz8spQ2nDTgP0S9szRfQ5ajc9
Lvghm7NdZHmg7BiT7KXksjG0AFNCbCxfmqhf9T6lcwDWXdgXhfxkFA35mNO8RFHZwxRNvpYZ8+F7
ez6SzYTVZ/iOfvq09nVHOXrvSEqLNgV4lOWgAHOL2g4YVVPAmkndxeMIkshJvnI8kwr/yUwXf3yh
BAMjA1xnKTj+pAlsbSo9WiCYZOyOFwC+CWJvkSbZVyVAVLytYmGLq2LhyJFQzsHJx1XNu5LiUcIX
H09wiJPTMROdBXagH9KKldqUCM0ku7JXNbJK+GGICwvvxmWnMrYJRup+vO1FCtSPt98QQnhzk0zf
qMw4Rb2j2mN2Y+ZxFriiW9Yv/9CSK2QDbU1KjwPNKJVFIUjtfYme5tZeYOOnNUkQtzXpDpty69/C
or/FMDDPQ/AIBC0+3TJwzotEeB+whNH1spIvSwNarkV5see4qjj55eLHZEgDGnVL/xZ0P+3Oib/I
27+noIDHTZHdg4xW2Lkwr08MsQgueM+cdz8FxSC1s83vmg1AAF3BcUiglOSIrTe1MizQMShsjcXy
YPz15Q4qIyc/rwxPR96yn5jDoFASvJ5DuoZPlF0xAejbT7XkS/nedGmglFyVTntI7kVCxctYMXQR
ktn0sOwVRXgcEuGY/07lHRRk8/dXfQEjiNeBMa9udRIT8dqD9ey7k9t0hQFSc3hzrMnptFOMcuCS
QYUKM21QsdwQp3NdVzA6TGnd9r7lDqdpmEKceiqg2M8jjFVeFc7qMPmkFTMOB0/yy94xwipgVw67
9NRsWPIZCjyLXOc5ODsymh3ZV7FgwPqw5aDHUty6sJvHoOe9TkwfwqB6vzBLkDS+eW8y/U3r8/ZP
jhG54Au6+A9okttbUtEEqCat5S/0UZYGkNSq/OQ3U11kY+T/X26dOEdpaCpxE6nXOnpqL/tOqJSx
OkuAaXNUAdBR0t6F16DXSlViViklmxUz/suuGGCSPSdnJcrXaDvAhSr/XefdKqhz764LFAGI95Lr
s4uaMMZQiGbt7OskT514Bt15wd9JurWW8XeTRW9OnwK7mLHoDQ9VWOcIhxKmUknlq4XZxrk45B0Y
UiXoXTNtRnY35DKr84BzNMBeqEcN8CpH+y8gEUsN2wCAdLgg/f11SDWZFMZtyuv8Axr0iOpQ8eD8
+dBPBemxX4oDV6vKutNcE4s9vQqW7vL29miPMTd4xg3iAgK7dDaRBHYnV8o8eVakGgua6cwwdzBy
gpbGsYUCiyNpalevvAsGvmh2HrrKdVohOkJ8htucj2NVIzkoi0wHySHZRoksXCxW3XKN9JJMKgQk
xHzzln2nuuTsLSArcRIgJv8yDTARN0RGEFa4UpPab8E4MyDnZT9bc5TbLJKq4sjvznRRN5heacZ/
FZbl3uw8yPUwJBdiUhBKQSFj1DzLYiuaunFcqCciE4td2I1otCsu+btpvJyhvmEjNZyr2T6GvBZQ
ViWV2X4BtqSXhhGr5hBTNzi6HI/nMLEh5dlJ0oQwEIO1pk9N4zl0iaYRkm7i9EekVJ2tn9yLZ9pf
DF4Zr5VwC9HxFxzQjxzS+KXdVMsDxqSwksENVos0Me9O0q6dPQ0LYVpwZ+RxehruuCbZy5zq6Su3
JKobM2SGsh0wmweHJjSeojO2zNoRjy/ss3ZaMiLyPjQ9HrWePuRYfajJawRTBK7bZhHovWdMBTZ9
7zakQ8LZ50UrC+RCCqmLBTgtbtpSE7gO7K1P7VzRBFraWeP6XIFW2H2odtBBx1Z7R4W8xrzB/UbK
dvQ55qntPqNanUy9PqDZAKOOoztSVrokOD58KFSYyRh28IzjUozGwdwISwDrVb//xDIajgEawQnj
2CzGwh7sUFFeZ9W0hswIPn0jL0zxc05oMDn0eil0zcO66bX2SXbag7b3TZmjqXZIiNJz2dWxggC/
nshVy67lz23TGRHotK9fZ6a2wT4lICeX3IkfDjnWU5vOBYJTYRuRECvIEiO6pwXQhmiw+MMqAmS0
Gj3ohjt+0VG7l5DjWrTwaix7i6jisj1qybRgIq695gqw91LNbKDeszdmDWvCbIbk5WRlD557uch/
QNezza7y59kRj7FWeRy2cXI3Nsot2No13dcNrrXq9N9vRgR5vg4FQWzzUtazRK+8HomG68Gi+Dha
X2jqD9yXHvxypCJZZ3HL6y7OrsVJ53UOvZ3zWNgJWr1DNQT/o+5y+E0a7rJ3H1vU4Z9ENxsJAzHB
lRY/yDBeC1Hr9gx8KVnNXsgiw7GmfsdFCus/pDq0/CUdjDSUeKYUXiooh9tvfomigwaB7KjrYf9O
OquolA+V96K+kWpvHV0Q9NQtPtBvZJU198Dlu1toPnRuRk50ZO2eQS6SeXNuahmPCr9ZJxMvujAs
tSM/lyEKFyq5y6mntdOPehRTuD4bOuoA3RW8tB6WbRFuQi+3pj5uA7TMC60DgUo++E12Ra5miDtR
LljTXvb2S23U7ahO6amwqnWLuFvrH11Tz+HFpYMOawggh9a56Ajeo5AooilRkCW2hJbQn3tNZq8u
iTSFliwu4sjlS+9Kt6+3pxS3agiDKwt4lWhjMkyQhF/ta0e7bMyW3UriHzK8ndMxDBs2u4sEY1JS
8kVBo6Xu9ctyPkqvYdzIhxKq8R8Af/WXMcsbLz2gFTMPV9vMhbP6VCFdWfGqMYNG8hC4T97sOkxO
JUGTlMcCO4YFQknsTIVD75YXrhc5okSkunfL9uTG+7Cj4BwCf4xkufzHnZ3M0X85bmyUK3kASgK5
t4N5XHbCOCQkdfwkSWiVagdHb/N7/2tAwYmCZnD5cmgXsMWMRoEkzvdnl0MHiI5M88PXS3KEXGPO
duHj34zSsOCzTuWJfUA0NcfDdM1B3ZkjkR8EEdJa87WCqJz/VaLz0ZU/xwAPdh2Id9NgVXj7JuGZ
XjG/34AWkHjGoN+MJqu5k1iagy6HkmC27PEq4DpWJhQRwh5uiA59WrVMARg2GFN15fe+IwPCYOFS
TREZ32b0h/H+cmfYUd9Oj30AsQ4y1Kc5fkKISZP7cioOXaXoYm6K4GOlTGY+Ko1l/Cc1uU3ixefx
M/U9O62iulYbaNgBiMFTsdpw87VkZ9b3QZTEItnLL9GbMdpL48zFeuZPRNUoLikluhKi1FebyGze
znHTsTEm/J/9hLxKx5yJ9CfLcbqYjSwApAPrwRdcpawJseFoDTxcTNBi48OENOVSyH1k5KpuVPUa
JwQj2RaNeZJIuXyUHcGPOqAgVWeovDBVLbD3onKeRfCIjFvNHhwzRHgOW73GBIHM9IlCenbGAE9x
4EiaKaccGMo+qgeHoscLvAO32RNjJXyN8Be7DWqqznVIGC2xM9vWMFq/vPoLaYtORBCC6F24IblC
y745Hf3d217pay2So+OOKHaO04khGrzHFUvAIJiCL2ykwCu6mZbyOYjiLyBe5pL+NvVqehGszAiV
7qulbUJDmssrzf/AurBQ/gDNN+eKqcT5nsRJQi5TRN5nwwW2Pj2odhFooqvoRL2qF+LVmcvCiDsT
WZpdy8PU31/Dc1VGeZH3iJD1u5yVBpBSIeahpD6p1oHFbUw5o0ZKcMAf9WY/iuyItdBiF5n3i1ue
eYKYGgAoeQmpg1q5Jxkf2bCGVzL+P4vqp5/BtFZfCmwCXbFdi7YWggTnEJfZ6fvy5m1n39nBsZMG
lA7OOhQ7kDot9J6F3PUx8MaMmrhyNcmoiLcIF6itlVk4Qw9iew27ogbPsmZpl3M7nnm7dF2IHVYC
bEtfLSOpNIC03uAkLORGSvRKUKL5PCQiAnyT195yCmvpfuwlBLwd7MdSjudH4U/1DPWUONVDTPN8
//Km0La6NpXYjcK0upXf1z6LklZqX93QlIqGUQPUJwu3JsZAWUWcuNOkM2uJE5hOd/tOU82mEYtu
cs+SQYgqZ5VnG/XYr68C/2UkMS369oJMwD0tumlvWGFMV09sQqXyLsbocVsAu8acN55C0U/nyJmu
MMipW6Gr0nAuYeMs8bzuJau7nLyaALdqKnrecwsVftspriYSYvbIiN79t24bPkBevFLz0y1x1W7A
wQ+FP2vNwKDyY4Dg+ByrPQEJcWsiiWZHFY0mxd15jv/c3zx+jj4VSzsUOS9xJbHRhAir+CsnQ1QH
/fGznED7ynNPngywlBtZdsbIv4/fiG+i8wuAAhPPoBEVNqMs4+a4r21Zxs7uGfXV0/o7xUcWustN
q2SKyq92KQoS1GSC7w0R6Q+jjdGetqS7Bqh6ryYVoLUzh/KRhjV+gra/nKq7u3FEfVsQrS3icJjb
rJSpCWFxBDg31YjUu+mOoIVqyVfsNE5+V7ruuDEW+l7Mwc2Qk8de1evkG3duV9aJrILY+JR6VY6F
pKK9IUv83zawefRgX8ZOOUe4hEC7W6/91AezshLOtOBIaKmNxXyp1VvRGmq6uMmfumAnWMiHEGW7
Y89Y3hg4FGmFLLAkRm1OxVRlf2atjStkfz5XempAw+fR17USP8VlPrZTE/i/nk6mNEl26+MKa7xS
THCqGVixAI6A+CC4pArKfvg12pxQ8i2RpjpUntzq48kTTwzGRb66BDx+QY7xy6Hcv3Zg5LgpNoPd
z8jKXYT9t1m87rRzxTsipQQ/MpBO4zpgQf4qqXW7nztYDqWnC+tgt7hoyd58o9fpEgiysLmv86qL
6jdKw3F82dwCTvGujFdzoa6xN3hRaQ+ntmS14lWuqZcdUKLeubveNTDICmA+Q+Ao3jsWMh9QpR2V
sZcPbtXkaa8bUEzYAnzHmj2kqy6QoGxQHfOqEEusS0mY1qs+MvvRaKU6u1BrEAbtSZnPO/zNa4yN
ZpYixUrdKf10uJ7y0drL2I7hpHjSH5ayihrA7mVJR8BS6w93mjy/p9TWhxBa873BJf+a93zMW0YA
OPiF0N4MrwYgfjpxtDec0/fIIdK461BRrJzzbOFxOJwSJ33rQoHlGh8xpPzqjGHh3jvOGEb31r7N
QnkdBOrCsT2H2cXufgA1+UTP1LHEXA+aAN1WNfJXw7S6VGdYjusAXHXsBLwVMDt3IR765O5ZuNJT
ovGBYF5ln8BuwoxiuKvGnWZZSb8b0tjwV0fE77vXFv0X4U6MSPhOrkkAmmfRjk5PJg5qpXr7eJpv
VRQxbBgkclzdgcLRl76hrpC+6V+u7ILFpYkDSokpDX8izWUvuxP8JMb/qFx1rGIGP6eWBUZCAbek
uDRrf3WiqYcuZsFBfQubwaQ96n+ajWVnmtvw4K8i33709k3YcQFHqalQ7uf7ediNdusIZW39Ld17
8HC2qQVok/YHyOpxStVq576JAmXNpCd1OOX/0pXLw/MdEsnXpIvDbKoH9T0Wpcsum3dC7kHYU8gf
b0LrgVDjfQqeC/D9Tg3DJnlcf3GIR0dSt0cy1NS89im+VVNci4ml26iQ3vHFBd5VpUJvubPGKhpq
QR4ZzzVLDvLwHtiidmJV6dAbdUHnDnzqsUwqkCS9O+k0x7sFs4SAgXnX2mnXLLnJHJcMZiu4Pr6z
2mvF1DgsZaXMrKZn+dR8uUqZASgt4UppZSHM1Bptwi2rsXN+Y2pbfbtEci5dRlci8tqh/RhqxLvU
meGPg7o0TQ1nAaF6w5OZ3cFUs08QwPPAJSMlBkH1IzyF9fi1GAz1oEkgOZt4HoRNtmF3o1K3g4M9
95AoIL6OJJfzN/xLvLoMBhO5xNhXLvZR1KIksGyPeGHWKwBFMxtlHiuTw8MBB4D0cQXVtu+kYi/d
JEdCQu82IB9Zers+4hlZyA0gzYdDDjWBMWCMxjlUbzJPKkXcS1FWsg9FXgS2XRzUllyv7l3zm/f5
TsTtOlxOlU20Xg+DwkaTSUvBYyHMT9x0eOSk8ORv2a1ncId7WcTa1TYUjseJN8tW6vp9S1v7HeZU
dOfoUQWxlLklGHg6C63R+8NFMCZBDm2Fm1aD/MA6BUvZ9TvJqfywAkb7lssO645bA0zjc7mKsvd5
4ALurLYcu0SaPvlMwiRn3acUYUV63jWDqKLBBWlIfr7fRv5Ru0jwtbWCS0zNfO/ksLyFRzUeT922
XdNsv9GgXBGWhyo4PuNMmCLBzmIP442rNglzpJrfFf06TUkTGI96BbrpduaLK1UwzMabKNHGFz5D
TvTNHxj9PaEJf8xRVSGM3ngJtewZL62qAqYdJCuqXCZWxSTFGC4RcxyVBwQoY7qiwYVvAU/KmuFM
rfDJ6Bczz9sO4pDGvqEgJOHVUG0X1n9iNr19DhnYiVGVfWQDB+gyjUHuEIaSkI6ravLYcciFYAij
r7Ra56XpV1mXTUp1Bk/Bjr9fbtFwRRr/tk6fMxQxeyYHgjZVxGIUGQOGUGqtGjk31NM/1BB4cIQn
NcS5+xojpSyQU5eb/cVEM3GVMeTyMYqmMPTC/uYmpro49XiuoVgB8A8izXM8q0sKeXBFF9wxkDIT
2q2hgFbBIpMmuDmqiCVxDxzqAp0VICf5XI2dLMYPNFIz73DrSVrUGegz+t6qZuUJqpppFFJQScpS
Y76f87CpYzVA4loEv5PxSH5i+OVmpIR534DiUo+QYPfvjAuzXussQktAnP5ha/oO7YreIQqB19UM
LBJdhbyoE1Y1kRDCtDs+FldTajq20JWwgK+Po1aWVfKFw87fgwzeV4KenV4hvZg41KajiQvw10o0
XkEVY/84aKDZ8cWwTgL/zOTL8uy3QHXLnU6K9LQYPltJUDNJ2oClb15O1uX3DcBO1xiL5/G2t6/d
Nh85Pxn5hnsoHDt70zHmTwnAJyFR8NXvvbhMIwdLUoGQXBl+Y0MID8XfWjutmVuUOvNw7sT2V1Mp
FuJoH3UZcBElzOpKTcoUF3KACNY75vvQ0hYXFps3ZkAgQLY9o2/kg1tSv789v4hZJOZlGJGnII8X
/XeDqDKVDP+ISzW5VtOdKRgwmi7whC5m9Yhzr9hh8f0ZH2z5a9LlSNsfashiyQEyT/207zhGmHSD
nDCGRcjKt8MiOuNEKZi3nKl5/lS7XIMbWHAXG+Mhnq80MKb0r3kl0vmf0K1LpJxxrRdEdte5kZb9
vibcSoSEsWrOp75WRdrEpqAHz1FeqQGbBRUrDgiaJp9tIACzIlIN6ZBtJsOJcsyPEpgm7zW2J5PI
H+fTaolCQnYnboxwWlMc1R8FCn3hEtOnl/zxQyQAfn4y5mTADIlg+LKNEI0wuLRk9oBNAKKhNdMq
XnUMzbOxB2r7rxoUbtjcDFH8j04Kw0x4yTjBP4W0E1VAFEmBpcpoMyteOChugD8tgs4Fs7n2Rz4P
TiOj1h7Cpejz5nOhGtnzQ3LgyEhnQIS4fz1Jj7PmyhREdOMu5vZtz0MKdBuMXBpx0/Cf2otSh6eq
uFYia4aW8M9bWy6WYouiQsKFATekxkTFyvF0lvfV2mZyyUxSUbl5PaTUD6lHGTiG7tOAqHKg7NRS
WrxGFH4jSempgOteUr1kPktwQL7u5TBy5n7Ey40wdo8R43x84ONk1wcuFftw7R+tXDVV608PMma1
F5xGS2GRPSd1ETMjxhpVSh/WF+89n7ITNwNveST3CsO/nemcuMIVuIPsfuLr999HAK3CnYScsXxs
Bg1QRYKFBW280VSm7Z282GaEk7V/TyhMNeUm3/AZAFTlmaAS1hyZtdS8V46HE7IlIWO+0rXDwF8m
IJrQXbupZ4ulq+ypM3awinUweqHd2yS/lCfATz5p8OSdfSWo3yZfn9ABQ2EsE9JrYrscMdGd5ZPU
T+UYJZUp8GAzUXSJizchza7CP34pKb/rJ4VHrnldg4yWJpY6BSKg2lafnQ1MO6yx2ovoPlIGJgxy
3X2vDAnn+OkfMCR1AZi1x8jfpjn3HFzqrnZsKG7ioHr06M7NoRckZ6mxczMGxnNawai+1I7jWulJ
/B5iH456FrBeVlRpdZmbMvvozfg93fm40WtF5xGgjnq6x9Oe/3zKlfNH2fhxqujwylMYrmROCXyN
m6lHiOOS+7eHrDvpp6p6jXDWfU8tkOuOPBHzT/iE0HIuO33ai1Et5+gEYzK8Se3Kg5TKxS4F0+vn
9p5K+wJBy3GoUKFsicS/MLH1Hpzf0J65F8b1dDrP2PM+vlNxVZjTE/dCetSEi8Qu6Sq318Fi1Lo9
fYgB4n36ToHSHZKgLEUgx1ZzndMorAYrVJ/etOwU4MsChz6NIm1hPYrSR8U/9JF8w82olUu/QkTK
kWDSIemTTzWdWDH15AMPrZyxJlw13n8mA9aNuQ092BOtequt1W5IcK69elwhFGZGgPgvhO8/Pkye
F3vGb9ZsN7OH3dXSSdKId6PyH/Ltc8WIVPClrf+OFM2K0o+zUc9FegfKNeT/JfbYT5/y3LYLbksx
e/lgLe+aHEqUeEh1fVQ2enCI61Ix8hGzen8+RBcaX3Hw9RyEpyH/OkaMUQxkjoY39rZI3KSChzV0
ze2E/NilyS9Ih2PY4go7FiOCKmAHSHq+tLmOwOcegTTMPdwJFRw6X44dNNbOXCJmXbcluVu8NTZh
X3CVfJa2llj5m9cjD2RsKxvgMcdSo8nropTseEPHP2XsBU2xvT6wE2y2WzFHcfKXqAK53Z/TTQIy
++0tRiPjrn8fBmEmmhBi0oakKp5ltqKJXUgJvQdMLsQPFZAVXBs4tlY1BFwSNIkOGpobXpIVAjc1
NjtfpmUxx80AgO9h7UMknjYg1GhNXyQPEDw55bqVCdQEZPeWNXi/NFnKUBfKsGDgt2nrOK6DyVzy
DP4VQOOo9lPX45n40y44y5PvAk9REvEB4AI2pGAF88x6O3iYaGiWoKo+sg9IfdeoByWwhJ2s0ObU
ZHo6dZ3RHpn+nYsL9WPOG4coT8CeURHiOvhFeifPvyL1v9YOKmZMwdDx7w62kXaq5D1jCNTrJLbY
aesTFGiijYaKwUkFw/rAuSDrB+whVfOo55MeTXVR85D7BMlqFJu9KHrTUk19INM2xUs5dX2ahyHC
tbaBvdraN1t/6LQPvxrHr2bs18S9F2/Ip5JaEov1qaABg+73lLi9eC1eUojZKCm0n6kjOpW0FMbg
VBN2JFUW1i7zIqhDraA1O1O+zoBxAlztU5+FpYLoeosWlplAWMEvERZDIM8ol5uTBqdcxSyf98eV
OrTPiWLHilksMl+4YUBPamZut1RdGE3ekPiVTMPnwB4F9wNUl2XR3oMXqtOvE5bBNXrg/kHl3SAa
6lfPRDDW2yTnegHJbDop5hlGyrVw1PD3CsLk2Dij83SyEXiquseEI2w9HJk6E6iHlhTHWOpg6AGd
CiWjSnRAKhMzksZ1FIdFo9190l8mYj/nc8Ge9eRPuaLfvHLiaC8i065MacaW3CpSDHOrRk0oTEo4
RoflyjrOohMcl6Mj1Fr2xAwLsg5p7uOs7BnCferh8TtmKNux5MOhv4r6kCThFdAMq6WgdYH/4s3h
ZDaUcJDyCR23T6lob6XrzbB/umLDTqfC2OvtOmFUysVEIuxnoNWikz6G01XL1mFvbJwwoEZJuCDH
Qlol+i16wi88IBmsgUxTdb2hAO2zAeLLqzkCKbrgBTvDUhe3aI6e0LrZ/MB2bjUwugWKmQD5zDgu
92mfyzs/SAwBTgrFkZ/bDBOBq3x3ARh08yE3Xcx1JUwHhRCX2U/dTosYsy+LyVvxg5g4jCTSJBeo
AW16E6A8ry7WZgfZSr0SEv6Qm6DM+oX+PS461HTFSNcMxve9r5yzsgTyoRE6iQYwa/O6e4gz9SM2
H+I7ZkjuCaspZ0X6Y82Eetl3RIfXXoYaP9NrIae/8VnXdTlnQQxYuMsDgmNjhWhiNpUBY+ZMLMpT
ISSpuJRlW1TYZ27QiSAS++JWOJaLRIxMGdgZ5/D9loqk17VQM/SwFXHtUJ0IWAM3ZpDadqEuikeh
1s5tu0W1KR1fiAA8IpK/jABmrqWp3ACcK1ipiGYg1ErrryDqIq+tEOQC85EMgLPN/B5Ig4KPCIAO
4zZxdEhVUtfY2jf5qhCobOiqgSqSkTwlLXcmjGBEmFfGhzlFyZnpLjMQWj0t6W1ohJUulTkSBTJX
xp7vfIQOfqVuPj0YvHHVhvnPneRo8ZomkWDIcYd24gTuOd13mNzFuJ+gzivAj75XzxW2ddCR1QkW
FbRHvIvxSnl0dZbcpRSV5souPfk8BD9Rjku0xgYVoMeW/CDjCh0uhSzENWdDs5WSz3yPbZTJAXUY
vX8kLBSSU2swzkcFcXvDpNJpm0uRpO6z5orb9FLfxlUAhtG1LaqxHNkklyis9h9qqahvwKgWay4g
qjG/JgmqZ3K7jdmcrcumnYmvXDizO56NTotfcZ6AY22S1PC6naYcygdZ2PQItkqi6DS0cPA60P+r
c1JGdCfPngYfJoHu5qWgtP5Wv+cAffCb2SLB6abAxrSBaZMzRGxDfz4xVVJck2H3Hi1M1nXDulKj
mCsCcWXQiY3ISKlQr9L5ERYhtxasv+ctdjpKTbOToreacra220D/8l4jN51G1gbJc3SkgyuzMrmS
GqBT1NUDy45YWhRV+YZ5ukQn8bI0238P2FAuTEPL4D0N9Nv/XHXiYxBog+bDwR1POWKRRCADobL6
i+8nqJEPK3EqBO462jeG8nqN5cafX9St0qqwqGRFTMCmZHzysP24AewahOH9tZUSPpyNBzxpIEw/
bQjYL9dsT0KzYFGuvow9UHJjHlJ5/JyVpM1kBKQZGgRPU7GxbvELde/M63spFqnQURlp4YoMAObv
MXohFZ33nAmD9NXHauZigNqfbegrPPDEzJllnJaWYo5sF77TqGrVFRSmPWmimZ1p7y114PF5/V+H
zI1LUp1fN+ybBrAfYgXfdDt3k6RdjYAKFTLn9fsAjIpSACWxY8wxcgewjEPCX7ikC13gSUrkA5DQ
NlLRSzIzIId0FKB55cQRgk4Svd4091jYyq0NZQgc4+4iyqRuO+tKqtWVhXOH1iNHJpjC/CUU6wwK
lZVeUYUbNKgVwm3t5pjG6+S79n7c/2p6mITBb7Bl60DjFd+a4i65JAJW+pWN2y+lzLZdYhItviiq
Sgana9gXQJW/Ot5VMeb5BPY3sB/zYtUq6BR1aHaDX4k6ANWPEoMq01rymJHtkmKqYW2Ybzz+5W52
tvakqNVt4JqqzXBs43NR2WlILxX481nDwUOUTqERNJkgPBfmd6lKfDy3aXNCQ6ivrnihRBEX0y/q
Z09oR2jHRgvM2X9XxMJzO3uFK3vigewMv329n+Toi0PC322MUtM6BecyuOUL924INOh+I+8ujB/W
cOFDuOpmhG2hkRbi4IPIoio+qcK9/QpwZvePWwX/82dkxQcSSXvycDzmZo/xPQ3IK2Pgq8vm48VK
KVq4nfYYN7wkGd7LTpY22J4WJuedy/q9bzTVp3yQtSBNigX3lqMZeqh8EOUvcy4moSaNGCT9VMGD
egneeuU/Of5CfmTEtiJBdfK54C+UAa/Z5CEHJYlnJt44MScsNCJhJqSOtxc5DqEnTbpEmBLw7DXr
fFCg5D1mFAvkPRJmLyBnKW/9AVmWnmMk3436TGys5FP1+HQ7TbYJkBvE5hUtYrP0KD+E/oPUcrU0
gRygb6AtEWSmNCNPjzGNp9lM8zVJ56MSugNnGZUPciPo+3Pza0a7iKtqBpak1QAWsrdub8wnKYvn
JmkY/TIwX4XCHAh5UaKiw/qJyudNZuao3eba5BK8G9rIemN2GKhvlpz4Gs7Gd+jlk3Vz8uowxifz
fiF5kwFh+Nj4cC5wpTk6dTajK7btWEo4/Jr3D2jxtZsMnVSTD15594DlSWQ2MpmGTcy3d0IlEI1W
D58rv93V8/k+6VouqEF6X1vAnhI+colNMRRzSt2vusFw/q8bCrZ7oT6VJyJDVwzNMb55FEVkjtLH
Hyfe+dFyGXfcoznwRyC6TpRn0SoGdYvgfNtVbopgMcsalm4TaaEtVfZaF1Ey2k8oufedazQxu+WF
U/hGUiI0PQYjafBRbC7YvFblFJylSj6u7dQ7aP6Lv0Ac1YqjIdU7bCFXuCW9LDth5KMUSOtmZyxQ
oFpOIehdC2Sz9TzBEZkqhNucHdhD1afnzKBWwEMPCEcJ15aOxhTygHAPXx9QwrFFm8O4pZVgVSpz
hnNaL/X0oubTwgZywY/ZAEHlPGBidI75P2IcHvfL2lrIcJNCcFjV4pFP7OdTbk7dkppEZGCrFS8j
nFnhBbXEn5/qu7+u0FSrBPeAjyICG8O3YNaecBMZZ1BExQKrn6yUsXkcM62c2DHTcsz9exUFWzCa
07f0HWppzMQTM8ewSDOzyyBPC+MQKVbXmVGFdRwNExqtKl9tlyxy/FRZ6qa2WqBTxhgeSqN30tKJ
Kyu81c36JCjzGlUUusAs17/cat9WXyfRT4Qrxs2fAYundPiLWHEJyqYCBZ0fYuA8EJUQVWIFsnxS
zDnmGHpFRaNpArxYlWwdEKVsQQfVNRhAWNsjpclikoAtaDnu2drAcSQmOF/mB1yts8ra00GdKwrk
u+VdsZO/0VrKBneR4794jFeeQHdgCXIPq0fvWz6Japf9aTf1OkMlLsNQuLhAQ+Zg6J69rJQaJ/C9
ZnVaETuVqou2H/nvk+b4gwVbbYL7JxxJl4UzvyaDlm9FNgvT62GTHw7Hg6v80ubAO8R8Z4TuJN22
s4pYlGTdoQf17SsrnQTr8MYm/8WZLDu16Gxc7NEOx5W0iHp5foecfFAxBG9bnF+1/7zxuWHpZTL8
KFmCxFDJ5q6czSwyHZHqEsAjAVQa1kMTxQRxqXd1Ra/KUNGgW5ZFevAWMR2lBFEUU+DVMDhsIcfd
WBVnMVnPnO1uzC6LEhjojUKDeqb7CvPOkHeira+tSvWJTJlyPoXtzeWNysXYSvHJL+NRdG+fxy8Z
dF7iVeCBlYJ7DZaqKwK6lh9mRWvrd/NMAyfuTdtfmHZGL6g6ef6HfzrRhQG5q+UiLvXzQM89scD8
oV8Uo3rMTFTGQaleBOEy5kEyqsPxa/d5Z3UTxN91ZeIxSdml3jcuYpwsL8gIDfiH6uQMy9wtS/o5
mDMtIU446bgMwVqMdBL5YEO8xV66/80subqOpKEEqJAcCd28J/AFFtWBTKsQE23viWjSDSbU3v63
wd1+zzTu/yVp4/xn7xgAFoVt/GxHfpB7xZD5r5Udac5vTkQja1Q6ZCevGJr9NgwQ73iBVhagliPL
knJKLZULIhArZJqq7RTUlMty8jzEZGKZ73uWsnb7hlX7GVZZjYw1DPOJKIFFC64+9UbTMc71O5qH
k3VcxBQEiW34eMsewS1qpbcgG4HnxsXPCPM4oMvCXWpJlVD0TpkRg12z7zfjCABMP27tsXA7O4rc
+Xp2wdnc/cvsa7yL0DKIJ3opt84VPiBYLP8F1cG52kxFBXS83z9MaPy6dwkJXc6CBl4ZOu9kuQOq
9g30NwwjwPndAJVKIEg+UhyCVln6t6hbW7Yt71z30tyARgJ2wBZEKS9OvZ17DE6NyX4yxYpQRYkG
+Tjj1ATAjWga8y/F9H/+ywfZYXuMLSzxHRsLxaTZVS8lPOIC3qdsss/7IcoqRd8E/325ovQ7BHGQ
LM5sQHCpMXl134bo67UAuwY+MLX1Bz7dg81mk678N7JyH5zLGxYnv11vlHeNpSpvi5jUJlL6IC4A
3Co6YFH3B6izd/nlbyj18ApChili0xO4lfmGE91ssMJnszk2qXWIjUFVw3OTalolkPX+gkvS9Dhu
nO8Vc0E461QepwWU9KYMgRS2USUISKUiIu+/HUkRYNJJZbhbGy/Qk3x3Ti4584oLkYurL/3/sWIr
Vvu7cYBvOj/tlcDiZeXS1Aj7PwYTRVs8Lt2/fGx80HWx1dLLpcoZSPmthwVu6S/czythZA/yPZk3
uApa82kxUFw+Zv/DT4OYwPU59XdzsokxMMYGqMrfMSoRW8I2gL/ICIvd+ri62e2V1b26llsLTfyR
dL3MMGR2FsYlFrYPdKBe/2UHBv7to59XitPmT5bwkrcTiTnCOcX2t3mzy1Uhyq/dwixAyPANPcON
Rkh2h3Os42wufkPkbbTUcUxoiZzHC9mX6dCqNYVmaXmrQGFqSYdgOf7NNShegg8w1bh2pMQVtwmB
a5wsquoRZH7zbkEtCs614fqKTZZ0UK0mA1BjEK2KsylcIbUf2OgKDxNj8ARXpIGXIDQnMpcqIZPW
JmfECXgaaufhK+dckTUUGhLadYtSM/L4oKsIhUytuyVDPbyrx8TewkmUaSHqJjzdADcp5jyU8UqG
RAWUDma7r28RYRnEwx5F/uL0E7xyVt37pWibNUvFV+OKhl7aLElh+ckOLI+mUknkVvbAwM6zHE39
lTUycdkQR2TeMBNdaP++nAjP13LcHTO7F/sfxqQ7UFUybSRpPreAAZZx2Tc5ioHhRrEIf5I+o2u1
vmnm+zph2gqgo1/nO29qjhrPZL+SAqBPZCtV2+lQIY+72eHse3RZoPd4kcf12l4XgyuiRb4/Qef9
indsWNd+/MJXp9aNIt9IQAWcaz0yaL9dZSmN8AE9evZeZvAlhE/i78bUnK/SPmJHokGF8wJvrDXD
S/YBhpZBbadsP80HJzlV7PjTFATf/9w55q5D4qO7lMJYF/DG4/jq70tghxpO3rUdanpXwurfyImn
Ao8qnaMBwvdqvIEeebfYnepC96v7sW5KfJcCRQ/icHbx6LKRV6XG7FEPf7C3EDu4/JDUU8MXmemZ
DQLTrgql1QoWZc5Ywwy2qbt8xArIk3sRC0SQWtd6nk+guAPUOpjdlkbjQ7K+7c/Z85c4iMwltV6u
JS1kqKh2KDLS/1RMXJxLJ6XVSnQcRTaAl0ea81hYTwCnZiPvwMN/IkIXiLtaL+dI4bCK87GNs0ps
pURNb3V5QCgtsfv477agBXA/UR+KrW/pRjW9pdI3yQunqWDYfQIJKkiDrg8wvogVyvc6fQfhFGkw
TBmBNrzrWa1SUA9GgJ6UDpgoznfmZg/1Zy4rILhuIcnGkC+6Ymk8nflzQwyszX7VbulaKGTH4DfL
w0hJHPP+Db4wuHMQZkpXk79Fvt++IvZmj5jlBx/lD1RGmiisgty2odkt/PpTGhhD6rep6MVu5Bi2
LRpWpkFU8AL+JeOeI9+UIiEXi/q2/JvnBdZtIbXc6/UQlcbDbzL39A8x8XlLWv+w+/qg+OskzP42
qqx0yoge3NXZh5rbIYtT+U/Oq2z7FsWIV3Ze+wfLdEEK1H7U3mZdA7jJpzocJ2fxUs9PREkiOjR8
1mlZzUYp12/dupSefG43rCa09G6SunEQlCM04d6k2uSfSGo25nOt9sikpfycOoA0D8rTzHaclfKf
hOd9HDghZ8Poe4KBl6v0lHoydTTybisQmzLQ30QIYnixhRFYVK3/XweXCp0E+DIe8mV+5t6IMqKl
J7fSaJXJOSGPcsBpRl7gdKj+9SgfTljdr06oLsAjnuK3H92jvZ3Ob+HAw2oaMqsaKsd1fvXA0c4V
su/tyTZscS/8TKBXFRQonEqvqz0+ax/8u9hx46sOGiSfkvRPfGyVzKtmYC3w1pVYo+aau0djww6b
3pCIH7eB640HPJUTFvUjLyCh5OeOU3M79jz3T0hFiHlNWD7YB7LIy3/o+pW1Cme+rJV6LkTJ7rTj
8m+2SfvKxU38SqBLk7ETtw3NN38rZDKCU2OhDKPYf8Be1EHNyAWA5KgAcBM2k9T0zsmpDurvAO+/
SmURWPGMDngNjcHvjO6y53P2AS7z0AO0VVN44TPzpNKGY/9FEbYcrxWAQFnog+JMTDiQYt49lrh2
9wjvu3skAgtZQzq9xkzmbStHE8TtcxUL5/JWdzoA/WN2Kuana8ZEe+adSIl/Z8GMIoY3mxCzeuWt
Ndwt1Z0vz9EWcea0X8BBS0G1AXps7r6d04/3fhIgcs5PJH0hUtpBEF1orVVYVyBLYl22vq6U76Vb
LIpi1gxo5fd/OZzjf/EYJ+XbiG21mRRE4CtA3vX2XsYeHKTfzCqLDuGk/3FXwh8hUamPDDOpdQct
SyxMdWyCSaebvfB9vjdMAfKmd7dQjYiyOrb2CpJ4N09aQWz1IM0uIH4u1RnzCYFJ3tg+rv91TBSZ
LHU9wIEXcFhwfWEQ5IhWydAUTnNIaLVb/DT4tsGyZ1LPwaxlS8MdIiPnYPMBrHmtYUiTVGV2sx4w
PiQY9e9KfxeSibJm82cGTNLd4d4yn8JKlmLs0J00R7id4SMPgJ0yXxd9WYGtHRw93Esgokz+Cx69
lDr86CYEajBv5Dy45gYF6Www4ROeNlaSQpgDHEvxbSGhSwfy4pTC+g78VWR9xhM9OmqyFVLdDgBM
uQ5iwrKmYd2uExd+EDvFO80+KPZ5udfrnaV+CrKq2gnkXknZ688PnUSE9md0YtAsMe3V4gwfNBpE
XH9zR/mtzJEcZrQ7cLTNz8cyRBfzgyCF4cm5M8rSggGTKsFKUiWCst52URY7gbThwrvOs6cb7I8n
Zg3q+WxeNQiSg2Tj/TNmGSxx4ZbGJX+WKwMeYsZmdmryWYVO2tlLCcA+YX0rFAiJ72AQQd4Z6w8Z
axe/6oUxHWLVN8IsjZ5QKwsucGLNsulbm/JYqX1liyMzqF1XXhz7e4yD8S5SESqYprc09btqos+d
vwLqohOe/TXzjZ6ecNNDNqpmi9LHuYl3nX+2YSXqwEgtGDAu0MvCh6Duwm1m2urfbUG2QNZ2DaJo
woqR6aHgSsuUTqPj8gwpfSJxGAe9dQwzjZuos6e/UdBjXc64t9UuHhTFEZJS4ZQ7dg0J2KeC8GcD
SAXX19703N/q9pJ0/nrISnamWJRE8jFbGUOEzP4DD/B8glW4/Suh977dARVA6WdBAV1kRQB85cFK
2eE9BB783OIwuH0K7SCLiWbKL9fWaPDpYllH3MALzXDM4lYzKE/+Z/0TRliuD5PASNeUzNQ2hhsu
n73DGuBoPqGBXGFUAMmYMTEqTeGV7oLBJScWBOX/llgYVSBklLXHxI/CYSwktRU7Y4/KvRGo5OSF
GeRr4FC1i/wKNwDomTQcwAcHYYn13nsYVn6n5szkmKOqZ8/uiW+Uyxz2VIvhlMoQUa3nP0ns3qfa
2f+clzJ7O3B2X1zuCmWcJIRYbLIMTbnf+57M5lee1HqgBPtTyxi4Oq2pfIMrpXnv5Ce8jwnxZstr
5sqQmaZ8iccCL9+Bhc2aN4aVCZYfbWbyA8hFhqNBGoJUTRQ9cX8uSVEOscHvEZvH3QcE/JVynROC
49J3FrVGwadc1xwJYvHJhmqm1rOzs7KU/ifMqcPk/o3zIb3NQ9YUB6gOaJ7TkRTYYHRkEN5od3t0
310TsWAr+jBUvcO/lodMRPj3iAm9gy1NEnowrjrW2G2ap7nlD/YaxQtkTRH8RyGFXQd0kkHM6N2y
jdH3gPmkNtbZz0LnLD0OnqXhzZZlMCdoSOoFX86PfOlwPHc+JT7y6JNAPrfJA+VJms61EIhrvFTk
81i5jEA2Fn6HEXVcBxZOVedFtf1xjCFLGlDHvwM/JUMvw4L8+/c/J7mbPEzIAjQt2i03orzvKXdN
Fw+ElHGdIU4tExmYC1jdwfGsxmJ75GdsozGZUYt77kuUFqeZN/OJeFaikpsRHKQEpR/CZ/IaHPIA
zP0v5tDB7RReez4Uk5eu/1vvcWm7RwD/h5vf8xB/7AwIPNGo6hY4M+Q3fFYe7qsgk83hS1apY6ua
IhMcs4iTShV3GKqn3Z+NQVpLRHGH8lyiAg+RNzoFAgyBmsNsnHmjcEnjmdz7394ZS/0B4E2n4cMf
Xe6pVlvgMP1jS2cjHWNCBHSup1XpK1vTdowku0YN2bMvJOYsX60koQ4pV35DSIB8JHTkEBNC2TPN
Ud9tcWfLcnI5jLQ4HtOG1p6VI48G6RtBERI5m5eE4cv7AaJzEUi3TICwhMtPF0r1D85us5oHUEAu
Fw5V+vR5eg+JRyAZvKaFNUsRBBfIs7JFwmwvxUvpkrX6b1c6dtcFrsDQ4r7L8HlXTLD2lwGT/BYQ
NgArKpd9zPNOadF/sdGzPjGmy6Z3A/2Q0RGJD4vs6C8HDzu6zGtDLyz7STDWjqV2tUTrlSfbnJL4
g3MdhLB9MuZyRb+hqyrVHyw/svgdIhwxcb4ruAk93nDpOAC3ZIBEixn7NJdkoxA+uKAoZOkXUKFc
oJvKAPVShjDzAkE7hjqDMWR31uvjr/QJgJ65b6ReYs90cdFgzrTj8DEGTbIEIF8pNIQfWsIFD400
hBZE1iZcgTcmjuENwD3EIgWEWixq0oORj/U1SIXN5xxRJpnBc4SLexMPfLFA1Uvk+dwi41RNDy8S
Qsj67HrmJ/Vzql2pWfi91KMOuLs+NQdx8Igh230uREf6SOrAU/0l9AJlFf7mMaT2V28wFg5E16QU
RZTn4OySosMhsWfyUFHWSDPTo+V8j4vYYDdzigs9VIM02Tn50imVd0EtJXxtkFTTqXTM/X3thZvd
+t0gt+LJRt/AFaiU6qNQrgBTCGbqsws6C14Yg/+UfFY3zuf03kXzN5R+noVdv18MOZ9qZ4z+DNgI
a3eXzzqVFloKh2ZG6ohERvpBZDni4N/cdhqwCgzSSmykc5ZsA8KaedvzD869Nk9xKjgd6cUT68IQ
yioFpCV4t53/PYAoZ4wJPHvhREUAJH0nc8htCs3Z2cmmS34BBQQZNLRpCXjKaXMLmtlaym89hlb4
Kb/QppQ+p6bbGUJJatgbsP6t/YiVKP6iRK/1dRrSNWXBMKULdWOh2LKmQXSPQ6c40bC83LLTHV2A
YHKgXfBEk3yYZDfvd4Hj1JW2bZqcc6tJ1/Q4CfpV/HLHYBRYxAvwWwnsEluLRkMZsCodVkSHMkbw
8XFa0MUUK8R44gRxRZgQExMpb2VHYCk2WW9LlsAnRmhDaXyRcQl62WxE1/W1EPRtpuN/CGHpL7UW
2Sxcy8A6Yqa82rqVOB7YE9zE5bjNiEHDg6JgWz5UnNzOJLMliGAxd6OHZbrkBCwVqeKGQnXMo1cz
4kagSZj08EnjdOCymkXv+RThXANvk61LciZMKGA+uwHK/6l/wXfpOnYwzjjUdqR1X4zlY3xA7Dpe
UpF/20vjqdoS3H8sr2priHyRypz3jvPJxAFw6HM1XYa3bbzrAVBnOV7tMxNK3b2bOky2itTtr5id
KU/DapPU19T2T1QhmDFXzLtfiW/iiP+BkzFwaRLmzjai/EFMDRLMjNd6tppeU/SfvHxi0LQPq86X
ejW6L1R7jEP9b++Lp17nSqEb7+Tj4OpKX2VJnhu6DCgAhcaQ3f1HsSUBbEUNvJ8mm4Rj2OATR+Ev
2nZt7X6qtIBbxiJrGyVVl+3tx1K0WMEalV+n/e8H++SAYdjD2YpXNrPDId0X15wMCsWljOBJ9Y0q
wXsDaCCjpRgvG1zFU46EhQU/LOvVoBcQC/ylI/p5I2v65msYDR8cBEbv2gZ4oE0fvIwUM8CjpnjR
hUDfRx++XhQRX0dDR8OrXFTur3dkJqE3/jh5ct/lVaJDv1SRLhNkz68OChSnrvUMqsNx3uthQAE3
lvLBXVMpPI2kWPEGm3oOAQDmLIXahewmqflaUFhZF/llBfR/2BiARg+z7qCI0LfbfSxIe3RuYtDU
fciNKsoW9cHdo6SdLQ1eMqqyblkpYL2bU4EZWj37mQfNjg/QElfVwK1URpKzuEV4n8lHP/a2WbDW
10PvOwskJx+///ZrTyGBBH2nScAf9a4l8xFx5Wlley5QnD2Gbz1VV5t3TkfmBYS3I8JtpKOrRoVf
Ds+GAi65O3iOuaHmlu6ZSM4R0sPQWeHiaea3kTHrRhgxFodGsDx5swV8EJtdEJ59dpLHcuoFXRHr
dU+GyzGmhmcUwS7My86/mCzUVlNxzkbpOPwGbOGtZGpfmZsTDrx8PsyMxJj7Cd7T572+exJiUDjS
ztOrixxc+Tg/FNzZFJUg1TGM07eduChcs4NFl3mXqRmrzIaCbvdrapvNmHYnYqJzrdy5574cYvJz
Tl8DYvBWxD31C7KaKDL7PRRraeZaT4hP3boxMmDYXm83CIiyCTVK03DiURns6Nb7MUnOedHNK+I+
RWyy0HxTqCwT6qCWHwxfuHSyolXQdhpYw5BxZNtr439PuRV1JHmnlG6cTdtQKre07BSZw574JgFU
2CfPiq1ykSUE3+EeubN999o5QXfe3CBppaBteVCiIqROCqI4kzEPdU8bpzTjMKU/OrQu5LxCehQ6
ZwWWwJpGN8Q+/EEclh2dY4oPQ1JnFG2Hg2kA/ZdVdpIqACItvfZNllEG/WXgfD+ZXaxpxAzqAzBR
RjG6ZYt4MQxwo/jayzAVvqdR88cNbj+vzS6PllqgVfbELVk1VPzepUibu8hqX2JXcv/ybUR5Nzfu
oWNUh4PQCh7ggUDptZQ7/fRxnZ9B1paRxcAylzwI+QGsUd60Jq67LdV3A1BfzN2CFmB8kH3CepNM
83SPg6kG3aRr+DRWA9b4e5lYMyb379voC+CL3c+bWeqIWozM6Ei7tVy+ZkUKawWr3nvgfmnImcFj
vVbR5oz+IOzhfydx2j9BdK42Ny6tqcvPb9tf8cKSMl+sQ7TlZ+hZ7PjCa47JHJg1cv1DnHMh8dpv
28NHMEF148b52zB53nz2bxc3qd4qGmdI0WjIJwaW+9UqPEiJBIW3U5ijcbMdiqQE0mYw1OQTldES
/g5G+oYmUocwsfqX20gBwb/xTBB0UQXiOTMw4ej0eVN13pWCSZqkA75bwSn6WtN6hN8x6KWF7IQ5
+RuMteQElplulEyN1ZW6qzQSKmT7rQ+MVzd6Yih4VnEpB9mWaiItZZMjMuu+QDGjedPrsUOYDp63
d2XR7GNPeSE+ImcATLyjG+YqR/s+PLljWmGDs+Qkf5TCkn0ceD3/r5uIg/B+piZ4f4yXbStdF0dL
F6znQXGowE5EqU/A7KRP+vGKSwkFpnnveMrZTkdsXCq3ytKyI78HgnAo751zkomOVx/sJiV5LE/s
HeFcfu7pNgrLGiMqaBO88rSKouri0KzXgdcoZqpyN9gyJl0FoLRQlHmpcGbeiMCM7dbqQ8KHcCPu
4KxhvmiiAMCMLm1HjZB5rIC/RarRa/B0v5tW7qAJ1MWUb1i5T/+elTXeVjRkiZofrzhLNCJR63Gi
jxWv2D0pHnJIs9IlQWmFL1qx4VOWCJDfDSYRjdALN8SE7mpK30J83LCnlLnsEIG8eg3VO36M11+N
DnUBkaBUZHsjGx0g64p6vdz5rtv//Z2MSqp6KISbvJjusiFC29458xu6BbkX5SToPmDI4wWsAkbW
WZxJyAolYAYQ75vQGFe+XDLicd8olPAS7xkkppizfChjFABvXdYB9lcFtqQyrZecU4btbJbPoqub
/XR+Sm9G8+08PaL2PtwV1kGPFJyDiryv0sR+cXuHItPnpgNnXcxy9/IP5nMyMCy1n3PsqAtYjTnh
8pqS3UuoYNTXE3dAkWkzjrvsPIekGu9tUQGSf+NMeuibV6/2wOsf0RkMKPiFRRuBudYH6TWqlbRG
zqZJ96cKeFfBiKBJ6AqxxvfQbg4JtZgEwUQ3uk9AtY+2nyHKAHt81lWCldnni83Vvu+NUBamPdXz
LMX/e9nXQlXzhxSWQmP/76awQ/OS88rZZnyahnDjMv14URSt/tQxIRMMyvvV7eWfkXkFhDxh9g0b
nwt5mTEReSjqtuPM4TaXwbmGN4mnM2NVGOWq9QVVlIDqtb5sp312mw/+yXkMxFWJqBiOqxORYpYQ
SR4WKvc/hilr9roVQyD5Bbn8XA/gIys4Hjf43i0AryuAHf21gzYp08CkMH1/VabxsCVqjnPGCpwV
rBJ//6fB9r81EOpNWHFuWOFj3y8ePQb24MAYPhTMEUK7lYD7t/qMzrhVKbOlKVdyI7sU1T8FDtJk
gR1PvGSVaJWGI2lC/SmjiuJhGdjHjt4tDJk7crc+z4fRENHt3xzghSYtm+lFCHdzRLc0S8BtDUzo
OHS/F3j1r77lOT90cjxyOh5oqHT4pq7Pq11pkIC0lPpqEZ7tqqPlbhyYjC+wwL98wnWt7eEnp5Hy
uDww3wLObp0ZufHAYS+5FLpmwTTCsb6LqBj9eTkgv/fWmGMSFGZJLPcaD2R01hw75tpPpOJkkLnG
XfyRlMAgPOYh+USiggkOFuQR6PzeVJhNFbFNYZ3BkNvmDhO/0FsPAm+ksu53uiNt9fwkJ3r1gGrX
2Nsb9JbDF+8e+uFmGhfGRerXJMklFBL5XIgwUhZDfoJzwhw/pDtH+JYqS9Aa4oHCdtEx3U+Knf/k
8vg677eL1Mof6y1kspXCusXFFc0HthZHP3TQn6puF9d7vzarR826IckcOMCuZmrAD6CzovHnXJ7o
dd5VlhFp7bYCSH3jzsdl1SYZHvaQJcwuDMNqLn8bYuKhbYNqfQZqye/z5/Erlu3UpdU3nf03IGlK
9r6uNB2WZ5QdhdyibbcqQI8G5Ubrw4APwvXA9nPNvvtjebgFGlP/EeDCyF1z2tPKWnQannw6BUbx
QIBO0WFPwe7pR8kgP2stWkL/AbZdJIzlOdFivxv7GvLhJNUNN+R5I52WsUcf2AjCyxEgaSvYhTg7
huBoZRPycriO8waQ+6IQdzJZj803ZuT5JshXbeMGVMir6SsORj4e+IS4LQznVjiHfVHYH3GeEpzX
Cybd0kkeSKaDWWjix8lyOUZ8ZLy+TjK0s/j69kK8QoagfIgyNrH3IeUm2KLiKdpa3qlPP0IiIObn
DHm7SxiDa5l9B9OkrvcNZz1PtmniHipMoc+OlIxx4Fi8w2WBDiMGOyP8apj4SH+XbQvP/iMiBKhs
KUJLY7F5I4DUzQt9xgBe5mDcbz9M0hfOuBEyfG5gz5QO2Iy8VgYbDCvkUSPly7S5uWupVcEXqWyz
zIZ/1v1BiuZoaM79+IWe53opF5WS4Uz3ij+sPTdxP04ZNtz4OHxBqzcHEceFvnYVlzd7BHXloL/W
tgZyqbihXqmj1zBXrzeFgzUBaKXmBSLLBdhTob9D2QtakJ4MQ2ZtgBaqa46jku3OM9mFh+zWSpEK
fi2/AT+d06s9Boi1+9tg3vBBaBihEyRHw6PIdjzlH9SRBJHhA4gXih5NNUSJ1CP6ISYrNyV0J3ms
KPfEXUkylkyssaGKKyub5hY2Ft07h2qWJhOr9MaRybyxBViMY7tsHbF4CsmBQWtlPD/wnxaP+VdV
qSN+uANkQz5RACg67Ys0re2GP+DS2XoTYoGA/f/b/vvf74GaKdOwTGBYSJ1hX/rVrgu+c+/EkkqO
y5joemhWkYiUrZCjs5dtEI5A/mefUw3ioyZAygu3Fgx79xGBOe/nY9pkJ4vLptISnbQ5VhlgJOkr
b+c8/MRpF0Ky2xf8vroWngHJejPnS0rFl8e8afu0u+8HtJMnsHque0PZ+UO9jkey4ZM1LxxzqPKO
dRwsPiXQilDiUv07vzf59+MR9dnR6v4omHsh8UlO4xpPqvcCyjdEii70/Snu9zbrSWY/IBSg3VF2
i7+KMddZSfKrykumVjlRQRtVqnvU5QTMYEg8tUkPs/v7vrBWkXGw2+U7RhCQtHhioihvL31agVbj
HOztY36wDM6GMz1JhD/fZ3y6jMxFW80mHbCb1dLaMcJqBobF6oW9aquGt+zOZPhjeX91CcQaPJMW
RjzVUhdXkPWlya6QLtX5VlIJTR7LOS77ce/1K9aRY8VGiIvSEiXBr7e+HR9RmgR8VU1W9lF6PyDl
9SKv8Z31DWSwCfEDoUNJSpJD1f0TA+E6jqhVUmvBFuamDbm/cYKCFRASwLvmei4K9ssRCV/mhhsI
WeOv27djhyL6XfAyj2loU2ftelZne4iJqZZ2+dkM11/qokPCQnmg4T+nfabVK9o6VA1veOiEyxU7
T5j++DPSucssXhH8n9wnuWpt9TEV6cVg0aKeDd/yIeWyMoHNf982IWgrK+GiYbmYf8YTK/Qmzegi
3EJxUAbhF6A25gSC00x7CoyB2QDljR6PbnRpF/tXBjpFwtxZTFimKtwgR9+eOv3+eYG/n4q3Y+fb
rxEHeJ+tOGwReIrDE3OsK6fn5Jm8IuEvv/y7AuZKrp948goSV6OWasCC67brPmNeIbUJrA2Kgt/Q
46a6J+h77CWJAWOcPY3/L7hPKIp3s5T4HJIJzkng5Ue3n3ScrDCiORJR7sNyzMWr++zi4SQz3Djc
XbClJzlPxRxYuu6U6p9OnnSrKyKt178OTuZnHn73ThFiCFeblMi/wDu2r8ZofPYrj4tTBdOQhP2z
8aYGkLw5nzSj3oSsgeJ6GHBhafqstFY5YqpRiacv4/3mzM5Qdw2Vhj3G8IcOyOTQYJQdRoMz71B0
anWPJJnu6ba+AVKSvo2D1zIqHa4ehx1B8SPoeoXQtT5Elf3rJO0Dh03hE9yXT4HmqCwTNjamqk/0
ZWRNbdV8q+5GJv7YbqQQMzi/l9C2cJgS+Ex18pF/TydL1HyUO6hvPLtHSdp3lh79OFgxfGJV9Pzh
xzA3QqC3o633RcWBCEpDISq5NegiNcN/Y9gUyY0tzYM3wz9jcVIGnkUuua4/I9UU4UQ6RDmNTpHC
RkItPl3uSGOTz57sd4/trM2XCCW5GN/iBeKSqN4I2hLpscVsehMZIPo8bqmNqUYOvALGS5b51wlo
HX0RRZFI0SYb/NJ2m390F/v8oFvHz7Jrz2x9U+wRxFP1EHaO06cyz7LH/uJ9pUsZ8uBshqCe2iPi
Y4ICkoEy2czzZLO/fDkrFxTvBnSKIe4fCgyeNRyYB0w0xIg6PdHMboR2oNps6UxtY4ndHljT2tS7
Gr/crwXWQX2Qihu0EPegJ/dhp7N/aogMax21jRxHu4Bknh8O5tODg/uoEFsaguXMTLtBMRtaBZSm
S4HDZdNsPKQ525Iu+Vgavpt49VqSTyPl2l4WhIt1+onBNqbTIcsvqFILryxwcwTxEDL3gcM4pvDS
CopWuBim+5keYtcvdrQjfCkjX6DC6cndU90glsOWx5XKBQwI0BduAjFrIDqWDThs7j6ebCbke570
vLNn1wvDUFzgrIp0WN/MneBhKIk/RE0j5tMx6Jsm38GtICinEogeH/d0V9Cmv8iJP9ZdrTcBHFBM
s+WbmqiKgrMcYvCK/HKhk2hnU7D9glwKzNS4DpV74SzUIjavqXSQzlH89CMV+s6/CX75s6WExFU5
843EW9Uu1Mu/vxGBi8MpTSfWAUV/MuFigmMEb1FcnWSv3qd3E0P9BcNAXFMFVe5MhvrgRm3mTF66
tIgALiWE5BqH2S2h6dgtNzh8hczLeYOY0emGDEqoB9roCIqg0MJ5/6tibp4J+IqFElPe7khH0OdR
JwLk9xhmJLzxqNrZ3jGZU07uBJXdVJl6YF0DU81b0gBvYLenLYBCpJvuEiUged1aPL2CHlT7WApt
9pFH+ChpKneOEdT1LJIiQvwoSGnKKbCFvjPV8xSaUp0HPv0cPcIZMlepp032rDZQOgF6om2xxTQi
xjy8mkv8eHnP7SZYMovDf4EzEzRQ9oe9+NlINCQnjvn9vnRxkdACIBxHqUkZ2uDoSaHC6yOPcygv
ieSJDVRT4mtItjgsrt+fNjkRWKm9tzLEO3BY/JMF80V5eNSAQbf5uGNpBvnafEGyfADWna8bmsOC
2++rDsIXfwFXtGD+q+CfBMDCIK2mpkNjxmf4xAh6U5noauVOuzdHfoWWk0IkpS76p0/APB3Sv9Tw
p65JCRx37aJh0g8m5hjdIz635txTt2nvgYJfbKwWyk5sU1rO4icx8K65cmFviUXoBCZLChhVceks
xBW+DearB2xcJOraA30oNTvVarWMTg0m8ikHzKm0jM9NVI5iKqoa2/1cwIuswaVcXKCQb97bLcE9
6mI7UM7xIb1AGcYDWpHccInV0WRjMJI1Yj3cYgVygMfc9iFCIFV2TRAul0fONA32C5B/3sl40+Oq
7A6Z+AcNhENalOYzLRTy/0DW6x9zWIHA7X3HnrNFLVl+ieRM71pJESYDF/O7tL+pdJ27mownZm9N
E/hQM+cQ89CIP9YJXjJmsmbC2SN2PBXAT5ubVJjfBToh1q0SR45x3YK1o9CxDysONBqPNngaigTL
2m1RRfnO+8tBW+FJ6cYB6khnYVIn8SEj3Ac6EF7XWKyQA/VrBRJg4H0cn4MArA4cVP86UzdkrKoF
tteCY7ATaBkgVYhCHi0tLznucooR49lvV8FOibOuKJeO7pwCI5bKUlhgdlG7tzvhcCyd1PSD4Uyk
xxfagdHaJmL3t/sDEf6QMa8gYopeQFC3nUl/hHhOFSXf+5IEkWf77E0KQsHvBtfnyHi82bmvgAm3
EzjoooYoEFSFhDw6aDCcOMx2FVwPPSToVBQxSoZlpx9tKX+THWvS+noT6dPW+mUymOrpMF3wvohN
l3MFvN583PXEg0xjiBMUA9vmtGrYx9FycP3V9ous5FKMNZW1V1CKvaTW9Z6TPHi9JKlspA0BJ1Mq
OAqnwIxkBL0Ti+Kf/ZHlQWVgNf1EIy6qbhCV1HBKCqG+xEUlTPcJkQ4yBi8SNWGooxV6FSaXXMAJ
fee/EAwVYc9YK0sHBqISmHtFEmW2Cdaf75a1CoBuc59rcEEHuuN5D44aNgZ8cA1zK6PyxT/u4+sp
FVP+ieO/NZhS2HUhI2+8XBPgkrueKwyTmuhrVUHwXa4DIYIXqpL15R0KrLuFv0EF064xkpIQeFBQ
2hhU7gCkc9GlQa1v4Z9hPVz0mm15XaFMgCa5saVDDmBfz2996OWfqL/P6zp9BsvzJB3ZSSkdpm3h
K8BKcfwQS8Bb+vaEFAkdwH6HQKaNyFlm92A1/2UZnWu2w41OgXaQNL258iMrXS7nYLRutViFjQLw
/9zW3fxtl+Ea9oj5Ip67t/rbpPC6zCgKrHlTzNKQFE4cJxQtq7qLDf0ackka4/NEhJTi/in6fuMs
XXx9l90kjoHYvifiIxx9+Bb2eydVS9sXYhAtOqY+VonPtYGQWuZ1+AF5VTgU9pn+ArW0AkUbAFKu
xq3ZedjktN46He9OnD9drTzweXy8IBfbiXzTXTIh1EpNPOpHVllIIZLAerP9vNYJ2Bpuh9WSFCQC
9dmPqZJ+JBCbjJ5V3stDj7AJZNOwrJrkh6L2xszQIxRK/3PFBJBwSifMxbYfLVsuOgIqWBf3jsFK
xGSBOWbeuuxhb67FxUyzd0hgUyU37WgZkrZV9vE4/CmGOdx/JDGeUyNAbyghAy/WBuN2k/bt+Biz
clIm53bPYYR0YShaOItp1g9jG6t/TqcoU6ZAeZT/Wyz8W435TTEhaA8QqcDG9K6NiShDHbVcfs0g
LNT1J+7or7gqBDuYKXo+JfJRvHYAs8bW7AEdt5vHtsiESnsH09+8ccVmWTsCUHPTZzIG90Bc2tAB
PT++i4y9akAhXYI4tmhv93ufhn1NFNRO6D/sVoRRoEKcb1hEr0UxL62DbkbqaAhBR1XQSd2tt9Cd
AgUSN2bMy/r1Y47P813tHtDGbapfc6T+OtdB2sKnreNdYTsw8kHBUMJ9M2MsrgJkzqT0p9doFzd0
7XqWN0RuLwrak9jy09DFMYzhCgPeNT9ByApj1qGwd4/0aX3ovTGVgeWurCFlc9QUeRe5e2rYBpt/
fWNUqMJ5Qhp2erd2KQWApl2jcJwubVRLLfduoPNoF5H8IH0QZZT2WqHS9Q74eWT463FvQkb8GcKe
lsEM0VpBME1PaP6Z9iLHkqYuA3hxthMiaL3F7Ooa86RvSfGQPXOGAKVWz6uS4KshMZOznrLi7czf
XlStP5n448fo1D+U8mWA/1QE8frm1afQNUEjBsK8mrm+MRjJ/qEFFnWTZHcY3eD9xn2oHaIaJlyj
cMXRjgWyRVpOTZNajZxOK8wr9ZvKi579O01ljKzSm/oTqZrH1KL2m4lSwg88iaNdaCfN/XWnikxP
1xrmbeBWmE2+maEnUt124FGQLEkd6jE8Rk9Y8TUV36cxsL+zxlaWhe+f6uKXNH9GRyb1mGW6/49G
2mf/BeeMrTX+ugAhnlsgc3IGKzr4X278bLILp7V5xG2Xp01rB4QHOpLJ3lx7affLqYC8g91izrO1
EW4AeT8Hb7Swq1gG5+kg+nBuC3dnz5SqJg0Da2bvysVaGFlU2S3RqFrJW7HCW/r0pi1GkW27ggh0
K6seaqk2nEHbe32OO6/GeHMaEdFdPL2br71tZ5v/mMxvmnYiHGSIQIkFsbn/c6MY8Xsu9s6IplZd
IgZ8y8jRrx4FKTnvQ1wDo7/5ncFIzNfxOva23gmS4bDmkvwYCrTvb9MEssIYHCCFER49d6aC4Zxk
2XewirLL7qkB33/IJZoOCEUUC0n7/k3Z1/7M3IwNej2S3CEeEWlpS+mVuQoKRyti0DZd9ugdwyWC
ruVNU+RYKYq/8aBKFzRwZypTCv/vlYApSTn/N2Cje4KqahHGnTuROUexXoFjB0b2nPmsZF3faq6D
iz4dQUHby/8PldIlq+5syWrDn+ULo73ORfjlPgtr0ljzVGJ4fzVBsIPmJwvmkKSNwwylBNVaFVac
u7itPLRCH0SascpLkf4Bxpq/Q7rsFnBrbo6VEyt+F7e3QwgsaOKGrTzn36IaUSvknGoePf4b9/fA
ZdRcOYBoCn0YjAKl185WabmUtfCDlBzwYHzw/wBWZ7q8q56kT9pWCKGuQNKA8V0HoSKmXmGAmBLE
80FbpMNyoVn+pUQZZQBk0NIgpQnbVFMk08jMubIZrzWc+d27Axgrm0W83GurR9Db530rm6TPztS2
SAK4RQtDOeo3GyidBPNEC4JkjRAPHwjI2u2nbkyV3bQWNBeU5bViYQeJ5fOvhcKHyxYE03MMbN26
9sdcCDx1jZjN88htsRjBGYpSHBZTBkzGp879+h2+ahpcLIncnoqsqlPSlJ0VI+zyohsnhrDbL5qv
SLFmbCTKew7m9Sa54HAipDG/O5P//qY7QwocYmya5LA8HHrzLdQgGG10gnMcFP7VU5RR6aY4rWhC
c2nNv7DlV8OcbcNMRkOkzTAp9eyeXVRPnpM1DUiJXeI6pFaAyKEwiDrO4nl1KBtEDNVYav92U1KG
Vv1A7H6+0ZlxSA8Ype+jvWpvb2Yzf4rg9ZaZ0JGG0K0NrkNNxpC35L1G5XVGJDtINzqzVRV6F6Ii
Up0lOZ8GwpcPVBMxPe0k10Avh1dqTG78nDzMfc4DWNQk8izRsCzTDSPNnnqLxhUySA8T8uk2zwi5
BZ17bx69OfML8RzQ3VoVQ+WesmD4yGpn4mFp6+wjaWURRshx+jA4HwQ8knhWmBTYqXB61NwdWc39
1roIBt5GKKqeCc/xDpSy84GCKOsjQxxBJTXrPM3+B9QYz8kK68D7rrOySSBQlb7ZyMpWe08WJ4jj
5QlhKygmEW9rTqO+s6ompiGP4ihYT3qEDN2rb8INhoRegpcD9h3Q0NIYNCq0JcsJGo0wGE5VRg7n
pNtUiE+WMUa+AfO71IraViU+33ZWyaYJxLqVec5mEoWsB4uT7mZGe1rS8vHYy4d3kGMgXHn7c0LQ
FllBJ8UObB7adov5lfkB9RhTWM7NZ3SEqDrxuVKwyGzRLUkxCmMRTYLMqtARU4Nt8CetAuE8ba+j
FrK1Y3/2PbHEUJm2x1ng8nA5kiQwpWy5AZOnYqveUYxoIOfM5o2qZZ3bnVoCAZ22pU+GxMlTZhRd
ZGiZGYRVwmJg7ELZsYkOf4T74EUtV/Q6wUc/eAoiCzvNJU5XhECCFmhNGNgTPpOyKja51a+FgETI
yGLvc5gvG8S/oTIUvk2O3yb5iL71FO2dBEix78pW7VucWNvn8g6QPY+TKJDIKkHwju28YcKmnwsB
7M8nOtTX2LHumQLvNoTFjYCuwuB6Qs0V41dOayBCI+TcfxwkFTlwV7HFPt7Z1E+2CoTSLPpxgHa/
PXgK7+d62hT5PG/HKuaLx/qcz+qw6Lp515LjT3zabbIKaMEeM7skGeYmHHGmC7Qy8j01Y8saOUDg
ZtAlSkE6Eu3hDuQHPBY4CP2uW2le20fuDkwMC1sxf/Xug7p+piTBdl8ZRX8fDCJG9NPs7rN4ys0B
ZeUWJrgHTUBTfrIGTd1CpfpWPzTVeO5m/9uwnyD8otrsS9ue2Palgc9dBAbZgUZT8iC9RDrNs5vo
hGdu8h7G/JMowb48AQxfrpze/8yYH65IwQfqLUKGRJn/Ek8uhQ7M6SXEaYbjeF8ufTVBzZSK9x3J
xmI67uDThTB57aeI74xEEVRplqPrePQuYdjveUfAO8uuSNyIJNK/wsuyJtHZv5zeQi/M25yT6Lue
U8NYFpegE5F3/e17FYqwoGREHtLeIltEXL20XS6WtTuWnzyEUF+SzpRZb5Xjf1iM+7GcLhh9lY/i
gjpDHDsHCxI7tzXu0j1zu8Tj67NiQpeB8/SkeRecVJAnNXsxzDEp5nlXNJ2FF+jz2xZGNLAuu4Gl
LdDsgQ62fmMKwvsf3ni5GArhq0bnqkw9nIOB+BmepyVkc2Ih5lRUVQzFh8g2d/8kFWTCxJwG7NJw
vqikri5pLmYk8kUxRzmp+WNIWSfIvgC5aYi5RS3FUjCcDUw6HMKKan2AO4MmjcY0P23aKPMzon0G
kxflqR81AWyQhCIq3zkqspjPoA/qdgGZO31hYq8ra/KPZr6ZcZ3k5kQqG51rKUuwwV5NmVgLBn3L
Um0U+xOx1Jcu5cPSerdCiUYuu8EaVhg//p2y6bijWWwHH9vScsiCG9+ezlYd+fjCgfBFLfMSitvh
B8Lh8hIowxdzLuFdjgs8IUajge3aXxmsVkcScDddffSdVBgSkZS9zPQOeTfXdRu9qZfF+ewlvV9G
Zyy4yJ4r1pe/YIjArJJ+W0QRUSk0eNeWGxRev/oIEpjlqvFRUFPpqCD2CGKGhkA0++DW1DLbCJ4F
Jb7d4adcVDlqEzEuFe36rezhz2vt2pS2vJlREwMi0O9aYW2RtQgPsuOUFl+sUOUrI1+JKAv6IsQP
2iKM1ABNtlO/qXTKOx4/wO+BbLj4q5vDU24GNISW7lawFdlvYgSaN41ieimu3jUpB+pUCom3qtv4
ntqm7kf7TomZqtYeC13EWIKSzzLzE2n7s+GXTzGlP+EP4e7jk20DAcxhO59QOx19gx4AzxJs3sNI
zbuTpbZr2x/22VeW70/G5AxdxEAWs6hbDl66lwjUhQ+pVE2hjY1mOlVVw4qEHwkxounSLkLeRBxs
jmZcVfLyeiyVnZa6dtmoMikaka7fbXLMZlSPYYk7cWrd2FQJSU4GKjaXnYaQEbJCXnnQIF3uz7hW
1F/qwt1NDpeGqPLcZzwHFpIvmBcWKjJhLo7mBhf4IX0G+49rkqaPxhXIIXhKYnNYvm54Mzpn4yB3
DWCDx5/hbBhnYDWIN7alQhbo7F5p2RtN/SVH+ty+NGM1CWGKpYBdmMHrYt0RUvQyrLtejRbKXlPf
Y25w7vD1yZFQ0gZOwHLLM1BrI0NkoXRxzlL0CpxUepAo/3MBZO4LhmawlwV1XeehEsQ2/tpiQWvb
fRUQ/43nhCDO+FIcho5jQuhpIj2rdgUZ1PgUFgk/ePbkUfMjCbPEDIjCYps0Mw5ERxueCi3YdjQl
clBBvhIIz+586xg4QMx5XH+hXg8DhtKtgFXFGnz5Zpgsgpzd9bUbF6Do3FSkjoEcJoUIrvrzN8Rg
VDJHIupBq61wqnVeNaKcT4TSQTgyF8Ounbd5F46pZIvLXDXcXge1J6149n9ZCZIxi3RpqyCeDiHw
8dn/waYgFJNHEXi94GwG0y2oNS/durwCiLze16nyCkqv+WISy5Bhkd95AVSdJdQXIArOY2dgFaJ0
PP4Ii1j+m8XerPsDw+N96x/fQJVUhbn+jyI7yTqVapcDaoRamNvdbcZN5TfMezuLT5GmPXCRJfnj
DWUjplyLXYwEbQWGIxF4bTYGe7vrTsdNe4odG8ybTspKW+DLwiITWVMdEnw1afktq93MKTjeWFQY
f95hDJ/gu7YqnBRaZn/lZan1OOMMYfu+VEZcz/7aWEB03+qROcNyW1wo+BVJYuXPjmI11qaorh0Z
qmKaS7ZNCth1qqHuWDUHUTHZCxSE6qGHgrYpEB+fifxL+1WfZh827FYtT0VV/wyWa7ODFbL8NipZ
mMXwndLluJjMVlJvLCMibqkSBBkWOw2iHu4B5X55RpwsBuoTF05pYjTRUHSplpJyiZQ5I3meF6Uo
48fxBtsR8WsZIqbWN18gvk22FRy2KAOXskJC25gztuAsJ+I5MRnHVefXX92N26YJZJNJlqSTvKs6
OEvv+hP5zI55d2XHj/95EqeZGJwzUqRUfi8eKxvDK3WxGJysuorAVY7lizVS5/FjUCaUf4nUjl11
LVcmXuSe1+FK3FIgar10Kb719DCwdJ5BVHLXPo3HLwudVkFKBj4F0niWC/UtP7kE9nw5PouoRWjD
tP5rNCJn/Apyb13QuEQZhjiK1zq1jmiSNRUTViU3VKoWpkKmJkxdrsvbn+AQApLxaa7e7Hc+llUc
7hAmCMHu3EVBCKOCSL6/ic3B8vcfhGw3ORkbAhc4kSswJaMVCF41tfiFMzBp7I/c/jDcYbjD4Uzs
AxMBhOmWHmgVJYAUjsPInYPBvEQeFmNfg1zzyjrJkbwXl+jEXb9evU7UvnG+0gQQn0VQUq+ce39F
k6BlfzOnVxQVRhoiObho8kkxbIk4DMgPHLZdwixq9WA7rSEqF5YZ3lsu2BF6Gl1clbZcKratHv9P
T20+enp419HldkJflNn9wJVJeyrfpbL5tmvhY3XpAxlwMwZ/vz3/qDia1FsvoSPDqYOF7DaKrRrq
dBL6wuN9KApjJ6eKdq83ooMxZiYXJHzSrYLrqgDROr0VNnzEpLdpREA5JRkPqFsmXdyMG48ERKAM
AZmK+NZTNytyhnCvpDRkJ5yxTpgZXriQmXAqiJJfPmyMUDpKKTaif9mYLlCcj7tuHuFPlhVB+t0X
gZREEzXG6G7goHr3yjKA0jCAgFFG9xejs99zWbbzx9a2uJtUQSZTH9ZPtvgWkryiDtE09QnQWxr/
r0sSMqo12Lqf4rlqK4IbTz5qv1/Ap6/8/oHOAV5lXWMBVhNE7csWqKWRNk9oeC8eC+0yIaJAGdK4
V/36CuSL4hbs3JPMx08MYyuYYAoX2+4fuZcQXXjiqKmBNEQboaMdsOzSF523rGhxOfUYe7n1hj+H
y9V7PxfJuI1+4e1V+60gg7HFFunA79pBKUu97AjeTwGfXqe+vT6UQMOB1h57DKfSoKE+iScDQb1I
HoYU4MpY8ca1tHpyo+JSewYOSFPrmMe4bbT1uTeQ0bmGS0m32JKcux/yMUUezNEuiHdj5x/Nw388
oSt2f3z6j+wsus+trhxzCTSZsC+bXqdvD7ZjumzoPpMJVhHJyrleRzi5xKCj92b2aTbiiAKK/BHg
989UeoMrohI2/PWdyF7gUpxZyJfb2Bl9724v2+Q4ycrAK+KDlnSdj3yn66/4tDMW7uWPOFR0KyVn
1FASJeudtuXQ8w9mTCcHxWneLkmaOmdl+XKCO9WeP/PKFHhodC/e+RQ8+DO5Lj/jRtmxnQlHela2
TjR8rJg2sqYMb3kgpwmyYsi1yzpp1KM1Zy1ZnOfW5CkNUw8pJekjW8b3lPndeRyU3jx1slJ49Mrj
bqRGDiVeGg+DgP73JrXZ0b/7k9xbBvamoVDaFTk70kpgFevYZ0+1/qv4Nbc0c8sYoEVxcBFCQdmD
q/E3QRlfKOJf8hEgjflZx9rqUs4D7+zgqJKuCzxYDNAx4NOmI5y0fhLI5NOA4x2RojXOWdvH3fT/
ERQPSVSKTZQIKe9tTZcAI4fl05qTkgXNneyqBcYlVi8kbGZvgHvrEAjGDqqO9leAzEHcYeuTeoCS
uqaXf3+6etl2RmdJ1lXwzdQojnzS0jRLAvGXRMdfa2gYdYqVtmKHMibCFN/8DRAjD9+il5GEP2Qi
L5J7+3xVrVvq77OMpPybtkxhRF1lGR5jowLhZDQnYOFAU2PXtPH5eUUmwdsU4NJkJPSnDTyBxQCW
3i4OMylgyZa2MJhjXSZynttuzBQEf62Sx7/pEnDDGlv5/Rrp3ISMNeUeO4mk4Q06SFxpU1Jdr8V3
WR7fqBqm6GdKJBgsyRgNzgkDY8ajXkXO+ktoxWDhupo+D/l/T26OxMy2CN9lU+ee80zxBi41KQWk
kmyiA+zlDcR68eWGcKcByQYL17mLSQm5sYx5uKGgFsx1z5JfKZVPtMDTI9tBiK1h/kBVg8jvRyju
6dHjcuaKLxA9usRy+Q0D5i6OC4QfjkAHA5En9g/HI433SlDcTpyJqh5Wb8yPdtHUT83eOBzPg3hU
+QjaQi2q6dXRhE7fS7mFSPat3Y01qxA7fgIfztfJbCH4IIgffIJY9W4Umhj+gnsYaqFLmqFwli5Y
gDp/0lLFGu88GedpOsn4iNXdZZfo8bjY1NVbbzpe3pXkqfRR7B6o7I1ZFnxrZAkrFHfAZvnPX2KI
b/yvRXLLl1uHopqrxA/cTW1y8Pjrthrr3rhwDQgLpmy3kAQwbIpCtowvny8rk43kb4M1KGrRYpuv
PHulQwF/SyCAF2MHmuzDZaCS6uybJ8RU/YXQSoQYiiyCfUFWGInzuqVTVCOuUOkDa1BEWTWf36P7
hdx2Kt6bggsYdCexGLZwp3o3t9OPBJ4eCaVhfEKrKEclre+XCFU1aTYcZ7vLkZIwvwZpUg7xUo/s
IZvxNktb0fqSUJRTezvjY+C5XdWEsoWxv+xndcsIN1FBP51sUUXSPgQrhbDMgPsqgtzQg7hIZrfd
zsM+AslZ6k67leXIvKm3EmERkxMZdkjsGxkUXbeQ/6X1bvIika4Ih3hsNsq/Saif1uPEtn/V0HQi
M7oN2by6E1lAxrLpg+hgWa2B6vSMO2VO7Sx18arduToOZ/HawutsDY91gtBN0nXoM9bA5qAXmEj1
7lCag5RM77+/idfRANQBfZBxHqWFh/3jW9+lAtqbAtrEf8+IPfVKWIUgE+gPJddxEIIUR+XcYWba
fxD1jiNRfyCA9R6awAirBXpEnZOu6LAoMeyyKpGSNGqe4u18aWl5tjj8U4kJHPA00JqrkkskEg7Y
vmDQvr1UXdWpd6YmmBV/VeFQa/NnUw4vhOZLdXL5sKWLihNiY48g3AV+pSH3sr0viXFbA4obZtZ8
4gixDpo4mXk8dwYeDKXnhYeuayJtGjzhuH6EpW4cKeBlD98UraZTlSwnAVxI3/v8sNGIPRkpRFlq
LZhtSzkkBeUw8y4aZ6zC/dUgEYd11Je6jAWW+z6BgdilrRy2weeee3N9OqG/rSBENZkxCPlB85L8
S9DZNA89TnfRvfcG8xGcpiDvfu/3phOO1baMX9/niDxoJjG3hTHqJw8ChNzSLSvVQQy0w4onH+i4
thzZyYr9fm92S2Luhxq08UrH8tPl7uzxuHY47TAxzO3+V0UaNVRHpVshVC9UtNTvYaMHCrcdwoNT
gn6GBnhMReNxpVgmX7NKhB5ndqOdmlT5r99W1CZCYfB7CNjGTwVje9bbHbpB+unGfdNdfqt7i/qM
foQB6znQKKjvh27wIAHSFqer3u/GqrSr3IpeDUiA56LeusrwO+aBeTMq68ty6Q4IILojnlnzxQi2
itEwuMtpcKxsKXEc3QbPFy8N7LO/HYLBRaG5ibSe0Ol7JHiC0qjP55IajVJXqw/OjS0akN6Aqjue
iM3kX2yhzT30Bc+AvVPk2GeTT2LE4cJMRXFpfALCg7uFyjgG+zSFicR2r8sXUFkh3LYa1waco4CJ
2q9xvBfUa0rYCwdfeIrQsNLc2cupsMwTljyc1Yfi+TiI1r5yU+mqxJ3TCsbQR+KwHL+rVKGGcEjZ
zpgvwHKmukhTs+j+ZD3ok0yAtJ14SpXIk/qEecsddt57uBbTXzTrAI44XUflo/gLTmoavkQ7eCku
3tKm04Om8897uPBUOOcT6kxKqLp4A+AB97lniilyRUJ7NECWtinLkSkqm7KPxq14qQWHiWxNvtUJ
D2rKUSQwmxApBv5DfIUs6Ff/Tww/sFmHB/k7vNcUFGXv8/6UTQwKRlT8O6nbRBnK7W/qA+VYLcNy
KwxpcaPItbKyUickUkOkF/lRfiio/+q7+Kkbqy9oSvusf4RQByYL3djRZteChvCgw0hQSic3iEM8
CM50mY+g2yF7tcszxMSR9QM+MR0cwI86LGXS6jAzFd2NPQVIXgJ8rKXitKs9ZZTX216D9OhQ5B4f
hkOwlrLFlbZOflOxMqRY2T6WopHdvMXMl6WBSw7IzP6sqZWxy2+g9oeDUYncqN9j/6LfIU12X9wl
c7vkv/fPAnqzIbJa/O4bielMEEVON+v2kfKaSIEHugFXB4BSh+nmCOOUGwd5WaB3t1wp82d86BGa
BFyb0O0Kl2UJBHkqrg/JeFbXvi/LKFlYiumUY0uAFB/TjYci564I9svfaug8CNKJh9er4nlSg6E7
oZxpsvr0b983/25/K/MJGLa/c/f3FjIbR3OBewuxvdT2S+t7cMlnOV/aCFMQh/qyodsSMxgM/wj9
650aK+/gxa2gjIf3apjHSJVuuucfvk/wQL8EH4RbBeTZXGT77gZKC7NzPdHUjPB3LiUzrvJUX7Ta
UimPStPeR91j1eIx/lh4K3xcwBTuSvbaIBz3gpaWvOjxrNmzwz6XU7NLPOntYCf8nsBcrjKSHniS
dVrdXLlFGG8NdspaalYwg6g9AJU1cwYQ5zyvMERMQ7YdSpI1mmBXoJK9vLQ7QMGIu5GJVn82p8c5
mBESNT9ki1OG2vJkx51UiocU7VoRnGy+ZJQ4EiaTRiL2Ka2FSa9Y6JTzjdSmjdIAEDxrsRzy9gQi
3pFoKXGoQdw43/PjD9RNSfq+NDEuba2FOL6P9Ddw82wviBRok/P3dsJr2SH2XdfP50TcSs/kHdRz
mAkY+zBpKNI0RJNDU1AV5o2/l9bZDutZ9X0pEgb5EGebR9eF28/GhjvhyKfeWjA3lHDdSkXbtptY
M7qYiOAXZ4ud/HoeP2Pqpf5PcXiuXyLvMQU4FSJPfmSqvyKwlbpG9qajBQd7opWN8K9p63ovcRhx
8FwIE1lgYzWB4JokkPPA5U7GN1lmM1h2W85QNtRJwbkqEj5D8xbP+/+kjqlputvOqOCHAUZ9bRZh
oxNWgE5ZzTtIBx9BsUN6AzprZ4UMklJlX2w9EgJFrSBc/2QriC1yrZUTXHfEeY2nULSfRFjwMGxe
AGkHJQK79jQG/C6fvmNp42lNrMDEhKKT56tIqnaD72eyLL3Bsgryg1F9li3CZmOuILqvy0CjZ/n4
it+gotuXUKioaIG82nDr9tC45EItR89h0e27MAXK59AXKWNgI5jQjxmE2JtPiJdUspQnfQ89PG41
HaxGtZn11ZB00SfNRBEwKiO+pK5iyX9b62ERLgf1LwfzoTx253Z/n62CbUIyaehTcWOZSwvQ0FSo
h4//ZCXo/D6HyAC6p/eXoCBjzQggNk9gSZ/WTw09wzfTTXr8R2i6vzesY9Nk9kHXGHqROyp+mgkc
9owmme3xIBPJm7j/a0SDGoiid4oVsJko9GHf2sBqrzIJvg1D3D4MjRVhAwo5pzPU6CSFl/kVrmMK
FgisbWZVKpNWc6grS5wUR69C0nnt6jWKzD0edRkvErrD5m49ekaQc5p9gItJO9jARx6ZZxZB5PGx
5ykgEWCV7A216fwOSWnq6Cqs1Jca7JC2HNzbCzPugNgCKgJDAu9KrnfWVpuXz944UeEER5OouJnN
oqkDwc9AKIDVKtzX+454kOhrOyqIyzovrJ8bpfCyDgHxWIqsaSHou7JNTG6ISV1UPWrzc64sKdH1
TP9TovA336/u7sekjOVaKzA5nDmOt75E2Z4dmprgfcFxOYXSCsjpBIQwUA++luInYmeE5q6ywdAV
KaWNJYS4hXJwmHlvOAUKY8wQFJN7IaXPWnPVBMse6WWd39smlhNcfr5rcOlzlTS0p3g+FEh4tkgw
iJqO1XON/ApO8pkpw3p0oAF9pTUm4+s+3BCiNgSb6LZcXcthWzlsON7R5NNOeFUaD/Y6zYYCkBIm
a4L3pges+2V9wXBvxMTGybywMTGnd3AWfYNDqYEq0VPfK26twbXd9ag1ebXkAFgQf/TPT8h9gm0H
QSXNgIAfQWV85RaLiq7cpeLKfL+UUye+04lH705IZo1z9/XW1/gKqZ2E+mFArqjqlQA4ABIJHhm7
ed57kwShXuCMy6xZmAd/J1/pY1cTcJqWXapwhrsoLflUix0eRVQH8WD4rGX8hICgoUPSCg5Ap+ei
Vf1dhYxH/rODKTEgKAcSFKzIUOLJF+HA+BRxPaJEudLfFOdWLY1GhJhvD0XW1KJF7QaAmimboeN3
G6C8qpYtZa+bVM6JgZL/bvktbb9VTJQYm4zaJ2QfkrJms39C4XzA5gF6+rap2daizMV4kGTsY6yW
HvC0XtrSGDXc6j6a28sndSWgpMoj6viKsGeAW9hoxHuVuyBvef4V4NfCP+xtWZoUj24Ds6XebzKd
YcMmdd/w/vk6x6Cs7unSaJwpFxY++PR3vWtihZ3hyo6jtXYJHeQj/MungamrV76FQx6dxMOl9e6i
zNxNA6y1mkeMsy8qEv7Wb5ePHfpoccLokvlngknPI4pY7NFmmw6okW9aXnYx0qkTMayfKgkY0+lh
z8kF5FTGI5zbnjOrtRGC4vu64ZbFYq25vBy6A/r8BOYZRkyQesDU6UPa5t7lE2+fneSm58aD8at2
25NAdyIHeaaDJ5bOHNBw6bJgeWqgWV7F034ZUz4MRwu1+slE5NQWNBCfhdqZDG4IYIAlwW0pOMXn
ICTXxIln3gPhKzkVqs7jDHhzA4pBTeY4tbkKUCBBIcJCDkdJIdyJum/2CDio3mGAxxVw2dd1aw8M
3PUGdnthYtC6u082HZAlvq3uIvFl0p4itvGO8VEev3vmXCvTOThVRcgN7LcBe6AarBJKum+Keluf
IvzfLzx9p+oy6nEpA/730LOh7/PoHcCW0qnLoiuaNf6+YLJxYPX0Z+BV+ssDglVZAOlCtwKqP0Bv
ZLA4H+4dx8JfkcCeH2uoeOg+prS0swB/lBjyHQD8VhNCB0WaNUcj18o2nCkPv5+HXQRMKHuTyYwG
wTPiw3WPsc5O9kwdfINm6FB7G4+ttw4ui5YZJxKmT5Fv+zVi0qBvuYTG1Mlzj0KlxuFe5NMKKaKl
adc9TBfmWYHDXM28ZgWcc42Pmk1FA3itO4LRHFgjuazul82638VI1ZfsY3/PhljaRFZk86IH3UFB
wL2Y/RWz0pOvd3ovHAH2yLn4I8VAMVZLmlR6srXLmO5UkHeM8EuZZXgugPLCJ64qUY3j+n310yp9
XnX6LsSTjtUVg69ivTzIcHtJdTRI8eRstPNra0cPw2T+q54NzWvryLOzh1nw4gA1QpmtF1Z7ptYB
moripHxyppO7XjWx5QUQwi2h/yXh+Jb6aReoOGiMAUPoax+PolElZe/yQmM2G3x+KrXpRY/xtJP0
tjFpjfU2jH1sYmd/4gPY23dFGxgLZN0vn7QzJxfmf/iJPzl+Gh2DvUvRoKMmvxLJewMJtpvKzgkX
TRX8sVUBd+EQNbLfGLmuCfC9/ATdjQ3rcl/WishX7V24AZ12BohlyMBUw4GCLo9+qaAvo+bw39zj
YrN7YjI7gBDqxlmrw3/I6pe3+he0mSdm2IfFUwRHNZ9EyGHtZC1K7TqhdfdjFG8Wt3P/HHKhlQJx
U0BUFmKn63DdqkbHTBJLNDhNmGlse4P39SWgpvClPxJygDAuVhACWtiCP0hf0YnKz+60I/T5cxOf
iiBKuHiINKliaC6qtdqIpyolcW6cjTKHq6r6STjMSw0cSv7V229eirL/UIqAn8Leo0mokuI/k9pF
bW2OP7JNWs9P0hn+ECq3ilme3T2D4RM5s7eOUPrT02/iyYjIOhEu41kVJTL3P+B+8n80UrEnorMd
V2dkg4fDZfaeD4v1i13Sjfq5pNFoJSvEd3XNKe5P0DJVskW/8ZKI7Xu9KhkhQrqqB9JNZ1zFgybn
FIrJqnSykrEsQSRmtEKhvEIuEtShK5O4sIc74wZdljXyODMQ8z7HZ7R0rb5rRi4pezZQoUveAyuj
q1sXz/BqUsGLA9VLQTAHzirWYg1Hcppu53DT+9nh9Sk7ArN09v4gEWxkRhPopbb72mkujWq6ups7
s96PGWghowMapCf9csb4S4BdkC7TPA/3oALK0DrF1PGGPUTdYzz2sTVL/trdFCi9BDIAHBwG4qja
YCiMAGlTBsdrJMtMCTG3zEP6s9sG7mnVcB8n0xfUtyb0/XTg9s/83WUF0rwNhRMQJB8ONojEnbOi
tizVUctN/4s+Adb0eoRniqgh9PaQ5Oa96758ZkVD7KBnWMJjMo7e1y38y3MMJUsTIFRbArU1eKL7
x2i3JwoyAv2w+A2JlTFxN0SmyOaQ9p3EQ1uP2MH6NtwgQtRSR7Rw70THFO2TnWFFFkTHA5GndRTU
zsbqIV3sIdJiqdz/rpkwEsD6E26eKpwQUhYSXy8WDD3dxMlnZbfHkZ029T1e6lzKpvxqjONEuFyn
y8JSElPyUo4LK0BJFQTFw4PcXuVQ5p8tSAFyIHw+jzsnTGUXYYEkEZcJL3az8vYlVmvM/Iyqlcey
oPFIBrw7E9hKpD6Jo5Vd91gM4vmtevHF81FX8KAkkYqXM3SYdayZ64XwUhuSPTpHEoCHItV4SmaD
mRuIrQ8JOEI+cm2yst9r6sy94fM5Eoxb8kN1BwnMy6GMZOnuWj3BzfK8X4rBDgRL92G/QHHdrtKM
INDij6IVDnpNYEcMjQKY/XoQnrvO2Jp2ocyIC71CDsQL4KZw2ruYwtR9KEZZu8eRKe7jSYQ6CAW8
dySfVeVHbnzC70O4Lc4rD9FzghEF7Ri3yP/v2OTXroVuKpYIUPRrjWZq8BQEumya8vP2JasGwuRv
Da/TU9IXUAIT6v2sbtc9hn88KhrVcqkZt7I8MxIXIe9uXtKhW/0SYVJjiDvwsyeaKQJnvmJUC1rG
1TgDgwcoDlUlCfrqwjNCyJ6xWym+AZGYTuK/3Rsx/2WurCp8TF6x/p71tlXWqwLBrNZbwRyaHKY3
cNUIVDq+CZ+Ue3tTjeioEIxdkK2zsMeNdwAVnQ+NxenKow/vQ6Xn8RRUG1AHJTFm5z8mtj3Hsjs3
5IUiFODOgk6r+6IA8WwF331mKNTsbqgOXCqOMzR47NROa4Q0h6WU/JyQRVfVpvtQJrdq/kQbiZDJ
f++dmm5uOPU22OWrtbm4mz4r91u/SblLNYUMdvyO1FjeKPKfwgzCSXv3EFuAIY/OG1aLU3VEw2EY
Lchg1kgO/worRVJifu0CW5GQoLi2C9+3ZwbpjXhP+pa8SA2hXZ5k8vJ+5Xm0KUoE4EadcvbiWzPQ
nMEmlFAGlj2GkFoQWUgy+Aai18csurvxKVvqBF9IPShE2e6uXO1Yamheqrf3BKKutolKijp4ikUi
pMO+NcVC0193tQ7g72JAOLYOUr0boOf2ezJdsaqGFcUj13+zRoTfA3fqtI5+/9NrI0z1oOyohdKZ
aeBj+VhWGpNVdCuCRMo4rmX7Hk0NTWa6FP58qwlQW5LD7RrtEQpHh8G3Vwk7eMm+eoIJMbhjngDc
2EKx6r9kE7k3Gl3rTDzX7YPAb0ecXp2Essb99sN3HayruYn4mfDM23/C09rbNInlhUmyhNx4hJyW
YzcgHkV7jQOYaDNbdWzK/EAxDxrSIpnzzMaTUofYAiajhLNn4g+9UJRqoAh9lG7MkDUOK4Zm7s0o
xkRFaDl8DXR+/P82KlhBQnW6uY78uNnaJ7y8dGaAzbbAbrLUdZrbW7+6bm3ivnEZ8v2J9+b3cX5B
XIqgT/DMo16bGToqi7/c0wqXj1D4y/4wM0r6V812JH9qwr9o1L8LWErDlqvDfNqkjeyKJgMzymvc
eeXj+pfH3b+Pw94Jw6j7HdPrMDRMSDxXuBeRlcikoZIFdk1BzOnxSyoWFPFDDWYjoCqfJxMgAJ2i
Zh+zFEV6Bpl5gJzJ1226+pmiqwpwDDRg+NxRgI4eL8QJBj56tCpssFRG1nS+oS4RaE1umFq9pXVH
2RDyCQQ6Mj7s4TH9h5vHiDF70xP3Y/4AhxDF1c01SyEvS6pC7PnKxd826A1yytiMgS6h5LERQsFj
YqCjX1xc4nphfQavF82Iqi7WPOowow0dwy+Varh3aoQPFGMNJDDRLpEwUAaDT1GCq8s901XdNmsb
MhgeCA8R6kt4LGxRTqj6zURe+bmrJcCSKrqzDiLn8tFjke70oTaCoU62fEal9UvOJcLX8tP4NPqN
bzedTGcpJr++DEISmg5RUNKbsjJjMur6auJG+bYQlHkQVFMHLlMeTQPklKfp2GbNKdNdxWbGrP8U
ku29xhJKTxDIRiICj0zkBQKrEuVT+rb3u14TEDAFzPO1ddLVRuzoTihRe8v4fT0IwJwCgs6hHqss
HiMEG3H5BF6UII+X/bkTVCfd1hSr5NIivLKQlRFJyrGAlduIRawfgH+LCMQ9wq7zbQh4Yno0Ke1p
hpnwqJR/HFKTaedTtxniSL2eipBZwYsmBMY4+ua8swRasJ/Kuw5uwjOT0piQioofAhD272qFFfWE
YOAh6WRuTT9dhjM48vbk7/F61+B6CdVIQgSsb6/0G5b5dSTGlITA/a1XclZybDDSLwLshkFwmKTb
nIm++PzMFlze6CRm9p0pY+BTvUuMlQh3fUlKkuyd2JBgHaVOvcXdTZYOwStCRwoBshRnz+xGrGvk
a0Oa53O6RPXz3sPP12v1/kzLCT0g7MmP8r20cm3F/raEMFvPNlk9HttGFQhSa/oSC74iA6jx3y0h
jXhvndPHmIYkAW6J2sTdLFs5fObTsqjSLkyQgNVvA2E/8MJWIh7I51JiQcxf8pglj9Dbtn/bWUEw
+bswbx2f3nI9AlfSna2b65RvLq965sEfqGDt8dn07zmG0sb1bBsytIghYWPVTSal+t3bd87QKmg6
mLn8VacOIJa/tl0Fu5sDIJ0tXMRxVXhJ4WCO+MJm5KFzISxVll1SeD0Tb9I2wfs3iWY4pk1QolhE
/JI5FGSO/yTndk4oIE7p+5gb47yu067wZzT/2pyypWH3XN2i3iAtFBzkIZDn2gZTm+mWdzeZ2EwM
q+8t3OtYU14vcInilDO+wjgcZj/WvFRt3TsAG4l2JF2aOMJnCW6FT1LxCOXJKTydWqQGZCXUgWfi
WTLrxUImvOt/QGY2LMyrMHVwStAOaWgPUQrQCRjMy3gYNBOB48KmJMcWdEKkH1jUgoRvS/P4Y9Dc
zPiKO3KTDx5FRuJm3iQ6ez754AtJYbXiLXoHhOlsBjeMWJoDOmxHn4MxXGY8tsSsmf3JN6vAeGPA
v5/cGiblVYBFyCcbz/CsuTmGaCZRoveLA4j+OUeT4Im5Dquxkewn4pamdcWOSmFdk7gvUNdgvv7B
aCypcm/YeNeVAG7X3JzHUEWf+fb2emjtjifu3I6X0aeJFDjqXbNtT1kbuzsNevuJzRgleFuxGaJJ
83Leh/va3g3F0+sUgLxphCZVcj4M2KFsm8L0ZKazdHH0lk9o66v5p0VmjGcIrneD+LKM6vap8Zlm
0BjnBLZQ9cJZzJuedEFZOYGbs3TPopdTK+lSHr1FpOCL+JTe8AMNFjyQBXE/G7yzF3Eyn5keA2Hv
43tk/qsbyIGofnjn7++MUzsj59fnzvJ6aCeO4TNnuRcUz5XXEpbmEg1wsuw82B5yJZrVz4BHO+NB
F+dpXRvhwx/z+Uc7D9pHFPSCT5AV1j07hRlh05IpNHSeEs6Aflydb09TYWtfBKd9/xuQemJcUDha
TlwC3vCPO1EE5ecy1mWtV93W5eJQJpDnclxWbHMLiEZT/heNp4kh+94Mhbjyi5whzRvrq3rsJ0Z2
0EHg7wIJpoxDW67asA4mvCRgm6o2XE7x25JwThr9OlagSJpc5961w4Q0FHuGxpdTMDoqXA+oMEo3
Sxgw9NHgjbhuixRIFUzQlyW8OVBTVjcMI++3ISZRBm5eQ63Bvh/nmi1+LByYWNqiD1vVUEVt0r20
QvPeUZEq4ukNfES5wBZceaJwxHUgEtrOtKBrPh+uvzvNgyIycG/n6mbIBaNB2d4llRtrckYYX85M
tpD+thMhMuCxEzKuG82dnQ9MZ3Ok+oV/sPfzmP2C5I3UkNpcsMAdd/w8njsmP1WHNd5hd4Lf8GCu
PFmxkEu+9ugUw6Eyv/IYI1vnJO/ZO3NDy5utautEUgcvgFve/MEE4XVg64p06+WpORU8hfaQJzLq
puQmCsDzyF7hf+W4l3TsZdKtHIm53Dknqsb3TFTaxGc9SrCZTvU3Ezrwthh0gXfrXTmdlTBi1xQq
11jWjdnUeb5B5AXkHQlA7DMiv9qK00eSiyoGwCdpC+G6GBhLd9PYzcFRG+SA3+/PPUBIbUWNrJy/
s6L4oOQk38XVpTJcIjRqcvUvK6Etc9XRDR1M8bu6FZdZOGWePliFjoh1w00zu9A+0x1vhyiaC0tl
+DA/ln9D+95ZwVopMvJ8/Mx9vc+ZyGLaTe/X9fJPYY59Zvo1uWwqtmsMYGGTHHPxncjg+CIuXtZl
e4oHz2p0KPgOpTJB8/jHVYDJjehzvknxv5w1HmiH0pMzQuevWzo1NJZYbOso1jdaRb6EA0xozhYp
oPy/e2jEcoVJV6ZjpwSKIySyW+mvSpwWzDiKKiCltG7fHj8pJ6uxUNJObVCQGtnGhLv7lCwOhqO2
grDCEeesbO3I9GZ/TNFRC2V8L4IJhNKLW5ty7mC+/ZYxzVA5Rj/S15LvYZhXOG8wZAKqCsHkOZbZ
wMbHK5jjst6SqrbtB94BTTWxlMRIlNfhZNLy6uLxFypMfweZMBRKh9svSxjO6aFi0LP8LGrFu7jb
wDDxmWB7aJXT8HNjaaLBp1YF+jY5E5X9ATBzW1Dawjw8AWbRg90fOvNx3+UHWth81HEt/+FbrOPl
0BqPqFXnKh3pGgRMlIYJcP+Fbbhko0xz8DWYMghrHaWVkJo+7YvKNsn5uqq0MMwWWqdwzDxzUfgk
UWdWT6XDGL9XT1U8aKic8sWm2snKGkAy5QunkBGCM5j3kgcGBO0ZOLGJYDNbSCt/fpp+z+o5QUEF
uYnlHgIXlyXqb9DfbH3vIdD+/km8K5xm07OSkA2BxYcsJbR9lTxmcf352RE1FkMvoRt+uNAYh/I8
+kBBCENv3dNWH8tQ5EHsxkhcWMDOBVuKrf0Z8npOZdlYGfuZDrbn+L/qSD3VSLekjq94UhSUFAaF
kc2r2LAhpu1Avo5GYiJ/bccQngV8sSvpMkhAE+7xQL87IRsuvo4C/wut0E51ApbYVTmPAJ4Au+QR
/BPPYnIkoYj2AsIdm6pxldb/KyIwRhqjy49tzXhETK1l8W695HPiRmUfdTw4cLTIy4mnIO12mQmo
pJ9j6BBXUf90ms0dvw/gTcISIGoEC1Tag22/DTaDoNGeJ2GrBKYF6vFJ/rR5LDfd83XqrPQXGnlh
8AA2lcYt+1kt8UpxCwwQ955kctuq+L5EtcZwT+Kwf3mO5RuwZNx9yXOJluTLfRWUhKMccf5coQKv
cm0t37zP/6/Z54TFaeNlxK+rz8LgxzB3550JECYSpNAoumGeLEkZnzMKyCFMCfWbwdwCR6LwxQyl
jUVo57KL7kpLJUB1yBsRcnJnAj9g4SLTtIxdTB8jyKksnRfW7Y8Wd2LrL0+kCxbCOxf3fZTq5Siy
CL1UdZSc/L6oNttP4TMNbZ3yffjRpE0QfmmiAieqRsN6d9JpeexL6qfjj23bFsVYpev1jn6ZwpOh
JP0Rbqu1uHbq2yAnd+T8NH7x8k8uGNele3nHx19MwIynkSPXbBTewdArPIT5Tk14sJ/fdF3ESOXs
Ym2Uo/jZng48qiP/v0mpjr32klYdizYG2zsdQ7dLIR1461HCDKN1lnXhw7sGKZn3LQv+8RrKbbUn
rhJ+oD3KO6KEHt1V/ETY+Pst7m39paOHIZikld+hYO6U+Blxa0l7ouFWTUPJonh7doRNJJM5DDNo
RaGjXsAsk6dHDZiGGoR7RWqqGbK4ejCyQo0EatF5EV0tO2zQ/B+IcGs9eL4T7czM0Td4z1wDLIIp
N1zRRmxNedtjUzflNVLufHzQuFZPoZIECQwsxwfWAux/Fl8G877HhzI9ATrUntNX+S4s1Q1Kzwel
CCShBqBTwO6Fyt+qStBhbwGg4ow8RQ1CgNKJrlHokCoGiJ1MaxTXVolHsES5Kw6EqXFpqMty+1tf
PSNe47s2yTFQYORZUfp3fiUfUn1yDsRA9DrQTINfY6YnDO81MZ7tBqYGXYp7dESVbPLv+CTHm42u
pW+e/ZBSPDWQzNXLSng6vTkYRIf+Pky46InboAMxEMQrxL3dNtksfc6peceeM2iXNtkxT96b9S/s
qcX+jxyi8/8RmW07VNgu+UpORhG486o3sJpYgutuSVzbxLHPdU912mhpAk2PCaULoA0rR1JSbs2Z
T1t73hU393KePLozrSb757HhYbnIRTwAbulpwOFurblYr6XlptsP5KDieiZQYUpDisbygitz/HZQ
AIFSjaAcjJmPSqleZDFSXlXnvjbJwK1FDxUA/pVMLCsg7Nlg4R3izgCTz2ID+ejHhyWiS4lZL6q4
C2A+/Nu0LoC69/zXNFPIru0UwmUm0uW+4mSpdJmAqWNNg8YPa8ye1Rz/hwPK3TVX27dZusfa/69Y
6YGG7Na7t1DGJ5zq/DXG6ruPoRjXFEwxVw551LWRdGp2qgWFcyOiHrMlRbGMn1hvr1ehkkl+y/6O
GAwUpFL3VWgokvwM6bAyPkaLf1dOCnMKTBXqIQ4u75iBk5lLGl49VJCxA156qov6NitfVBXcPyrW
iOLdZpAJUFKngDI023mvWwvWZcVhtbx69nYJr1/edavDXFljfOXBDg4LYQs+ykUZB85wp77twjhm
n/nge+MSzN5dI+M9LREZ4YRtjY9F8sAXbncEHhC5S8vWCgxcVJ+8/72mhnvcAKAi1bahpIkXLeD/
pbevgTKpnqkumOgbJ0ZHc/Ib9eIi5wXa8ny3fq3XRdLS3pVXB6LZdKjS1LiqdEvDShTdUb/onkhk
aCNt6N0sNVnMI+zlyXZDc812evKjCAO7z9R84vKN97RhGR18u//IkKsRwbWr2bXe497aEUfViOOZ
BBOBTg4LZZphripOmZYB7iedGdhkRAqr/lk5QgWK+Mom5ZmoOgBwRsO0P2MUmEaGR9k756vcZhen
BDmEhDZbbBqoKQI414s6Pr4zJigUslNpauI+3u5dIyI1fkwLy9wNNTBtj7ELBpNogoumjpxilnk5
LBZd0iFOEua0fyAA/rkqSe85F4wL5tTybDyo20v2YSV9eluN8DYv4wSP6XMbmF0u/hku6rEtvPHB
rMnax9LXQGwSLflL4KNSTXEWNjOYS7m6ooODZejZu0LfwPWUsnUGsJ/tQNcyALwN4tbw+W0lM6sb
NWw801uRx3wFOhl6gYlz1xtDMTWfN7Mh0JAdp0tpz8WrFOw6OWuIb9uv+hNTqHbKyGhjAr19kFI9
nh0kN6u5ivuHThqB91sXhwZRY8zxhyjY8tadJo7+gQEsTuYCrrqZpHrL7Ink2D/takfQ/hYgmNJ9
lHJgk4kP9PoxrcKdzbNMbzTMuHE4kNTM/btiDYdmuP3ji4EQ3/z92zM5R+6udK3cvi1fjSwfLhae
sIkBw3AMsGuzLpaUAuMwWkQ9ryuyl96DSzEuPlz7PgMx4uxDTTU/ySlff2W9KyeJkugdspi0IWV2
kOAJnviZVrpEqHgSH18o6JJ91vUvDeuLaWOJciDT3z89UHjBLSPD8Givc1AfzOKCZjgRrHl2kGhh
tChREVH4bMnCK6jKFzuNLzmBVhZkg9vaivp59G4VuhlFRrGRvdPwgtwmCq/v4qq0OT13Ba4R7W+l
1ET3GlLYbcrGY3pDRwU0gxWhkE1Z7xidw/Hnmx1wsDh8+lF4jvLcPyYFRbUzNggeIsyI9F2M4ssm
D2zDQx7qSvG3au63t4TSuNWh5BQhfPVkPn6l+jvA//BUkFrPxsXj+St/tCjmzp14QvOPVuT5nMIa
OxDWmzQQiFF55Y8i+dbESKdg5q0LXmMorSlNszN57Jsy2kecj99IjZs85PKGGPmBv0iUGcBKEInX
K37zJI06WeFN6Q3W/rLD1/5ivIBqpdERyjE+18wVT1/1oDuIg+a+XFwHdbNU2sC/wpQ4afTPZVeE
VHA1Kk6HPxxX/qZMnZhyOXANwSOBfrHKq0G0n+c3a0bMcdu6vN9mQU3cf2mNScpoH/HX5Y+fviOm
3MfSz2vqmNHMPU2q2GfEE0+PsXNla+HFXTmzgg2QEl9QA/PUzoppP2+w1r+CYY3pnxLDP/exrFuz
UcMAWyo6zWeqAuT6uZDQnMn1LfSBDQHvPVNa7S3BypfCeaTTgVGM+RYtmpIb0hctTxUkONyP+8rq
I5vVjHaTlq+do3zM56/VQ1Oh/XvgyZHxsGZFwfjvoaGh/lGhH7jxuo4ds74eDOYD4f+9N7fMg/gW
Cb+j15+P919/dKhyITgJosJ7uz1d017piaK1LYZn8KlFHJfxO157bFI6enMzKYc0wsjWb/vUEe6s
MM5/GCNwGQhMB/Jhx2W4UufmMHqNHVTSRCeiVnY9MLQckGD75FbjEiKD89YmqXKDjG7lkKYEM/o0
doVvyY0yh/bM8nsWeVifzrSpdDl4yZifJK+XRr/L/zDLzlPJaGdF3sCPd9I9mtVxl/AQ0ESwfE4g
DW7aujklddyGeuSRBn84jRMdD5ymgt0XN+UHgrrb2tELcYhqLoBFKrG++S+F4xT0lVZoNrbOJ4zB
9kw7eoD0CeBVJT1fJZqOK2xT4midxyyDHRicMu/uA5WHnBgf4ns+K1zcwS+sr7+90WIT+kAGs73Z
Cal7Ijkw56Q4cAbmXaZtXUxyksr0Xq1Vtd+Ih0Q6HNSgRAOaxqWCU/YIg9NqPXzKr4+fIHcpsKw2
5N5Ce9NCUPPK1hj6NMsDLKCaE1qB7QIO3/SS4Two6wlbX+IEdVC0vaLBwPUacKavlxtH6daUf+bO
IrPC+dcIqALFX9QamAMstBDG4JayhIWJuMJ5vgQ+kA+dO5LEL0RyqPmydra9mmwgxKILZ/JbLQ+n
JCmXiS6KdR/X+exEEZAzpde52djcXUS4q5rXGEVN0kLDWECCVjcbgCu4gcYu73sH/SzAmuwVe3bH
a7tNG2MrKgqfEwnUAhNyhzUyNrZMXu1oaAe+xm/229KcSizZ3+A+yvknonvVtazLld6lhJDyOkQt
nQgPZFOASF7VS2dZ1B9u3Pjmy8YYazazrCIvjbSVYSVsuEPPVOEBJsJbtbRqXROIuTVG2/nOMR7j
SV5/eWXDFJqdPKFgMU90QrgUy1wY9mF6Q0bHambbUbJsg8fV6AbjtQW5M7/dEPsME0lKL0QPZUCs
Gx/MlvMDnTFQhHQCW2o2dpI9qsdE54PD2CJpA8XjC1daUBI+01vPkU3XQ5h3TcmWwMWviIdRz5Q3
VDjm+fYJT7oOOTy9dxvcpsDF3EmHyukTJiB5TygovotKXfRdSP9AmPi3N5EkOVqkFEyqVZhTL1u8
9y+tg5Kjsg25e3rF9duaa8wOxlBWcK2BKFrpcIzfwaQ2aqY2WomaTyXGtinCHY80mvhGaYlem8Sw
2wKjEEfeMoYhXCzLQwdszUQ1kyNOd1hjujVQbeVVSsMEUAmcalGlKdk9elzfeULtSWyMTcDFOzB9
+MFd42kcTKrXrrX2mJyRvSPc2nMEIDqW8CUNPBgInjT1il9AifCG0I1AELnXCQcUHuN1cBVOYj9A
PuOinXl9VRaShdzjRzwCK+5J1MluUkcXU44qdqDbMRkEMldaaLuMhqmi3ZzqimmPVGwkOAxWOp/2
4h4zvQlQ6e4cbHej5b78b6tl6DvIvS4JO0cp0kqyb4UOn36QUYtIPOQ+JeUZrJyn+VKxRlEMQKcc
r1t7ADJbOV/LLV63TpZUZg5uzUodBu4hHTt6oEsCJfcmLoNpUNp8N9LJxmPX/Y/bVns1G90kQ60V
84UTRMiqbfVkbF/9bSEouE0u2RImzfuTP1rgW4GZ1t7klRTTT1SI/jWzpqZSsEhTQfeD8e52g4Ty
q0hxcUFnD4sNIWxZE3ZumXlQYGvwXnt46M2FiX8ltZ7VonkSXWKSYLvNvtoUaQ86HPjLQxgDw6Os
OhToJHoWDJvvUNq6kDJLTwxuFGQtSwFDqnaBvUPbyJeBHgGEsl3iqQ0o3+6tx2DMngQSdtZtauEI
s3EpsDFP3mlI26QmFrlQdAdqy/B/ZjTjd/9Pk6/cw88X0ppoCYB4IbVkd8zBSS1Rnkh2hoplKqN9
cPwfPSQ+j7yI6PhSVCtCqI6crglyGt3gBCG8xFzCYtvqnllcBIqjJSYyxHbIW4IqyURxi2mpZXcA
8dnDX27vqnxttVcKyeDtVaj8tCzDlgq5+lRYj/xBOgMbU3dXcJqbrvtY05HZl1A9XJfydQly3Tq2
iFw07p7Q+ZRjZdxWDVG/TZkHkJBToja40VhyxgbJaFQvloPr8+5TgGWPJKJDC7tcYS67aoRkPOeM
1YUHAli+aiSMEt0s6c96ib+cbW2Xvoi+RANEUDamiRCkf4rpCYvKRFWgHtVPLjyRfbFPlTqGdXp5
hy0sRk4j9h8CkXVcv+dWPgKMbk2oEKQJBEHAsvFPN4xW7mYoPcD11igMmlaw7mIZ9LLMXfnJ0pLg
jH9SFshP4PAd4aUgGIhGnO77sgKyhzzNc0wv2WU0G8zEKJBDnBS+k7WO2CHE0BiTuDUYpNxTTtrF
s+n5vzGxC5WMYx3XRAYKdzGBjz9x14IITVsWKl8eqAm7cDqsAND8R45BXxktzdAlxq0wvNef6y3K
8R8iB+Yl1M/pEioExkcCtUN1oY6WknXURXJiAFlwSTmDj0m7JvilczgDFMK8bibhQvD4UMC4t/2V
+WbBrjP191Ejola1b7NYasLZCVYJcLhMpdREQESM9fn6i1XXaPddM9ZA/OvFUinV9RVBl0iCrcO5
Ocp2piwFLePZRyFjmyeNTwjk+oA+FPsI9rKkBHo6dbRB1hj9rgJ+2/hTmmuFQKf7URkHffPrX27I
oWzdADKZMkO3AYzo3dLGSZ/kAOV1o6jlLdSwCe6f6eVZKf1Z+uAzDa6K6fqEfZwwQBxVwt13/A85
PbrwwuVQBWtsJgtLS++Jo6nBggePfymUIpb4v/fSdnBeB7uuK5gEpFY/2r1c/pixH4tGACHxNRrz
t7u+gRcEymlZLRzzK2gqMFh3aI7r4/WiNy0eRlD2APGEiB5C339OvGJIWTgR/NxxK9+ToSReyUxi
rEjhnegzUjau4ufgB1chxb/CBpLL5EgKfbhFrbBqnXCFp6mBhNQjiO45YEjdAq7CqjqFAdbQhDAz
vgy35ouUnUCfZXmSegCFbKgsYTb2zLMJai1/cjg5KnthIJqYpCWOn6oBkGtpho9ibTYoohG4mvyJ
RqoRJIqE/FRrCZZl0PLl+QYcpt2zTgsmVsFYvv5UUN5YESlxYJYSFhWDQwHS5j2pbnscWr41utub
KJfBgaVVE+jVFQBgfZ6TzWbxZfJaH0aUEwOkU1wLlMImPzXPtfG/6nIYAEFuv0S7VdUGSb06Ccvp
xJGDD81UYG2rNqYI/UD9eAsUpWF0UcTswceSLdIV+BfNnPC3ZRsR/t6HOkF5lDuQD2Z8bL7OwTuH
OzLqfEqm/sM07dwmDgtvlW9mBf3Y03M64geAanrDMYlHRHrhFBExps/2RYGPQLXHOAf1czCLsKT5
T9EjCENXZGAbgutGk8yXoRXUZruIxusSJpSk2rD8BG50en8G5FqT22IMeuBNbXx6KMlN8g9BXwJP
ppPpitm77TkUVChxjCyhpZIInI2FdO8xyRGs9tUz9g8Mztd+LeE57J6A8jcY5qmhLEdXdDkPSuN0
CGWWIIxGmpujJaDSege5XLYZCGxbRoe7m1xtOFVSayPwfxdloeO4sFCiywCYOzOZYj95F3rewGfw
YXqDjSiXu2qWbJCniKQeKFlT7AmOSL22mUPwJC2ExxzEne8187NN9XHv4h1ZFMSZFWScpWntk6jT
jNd5L6Soh6CjBe7MSOIjJzlqugpZItTiFWqVtsjPf2urHO3nUpH4rvGrqV7ypkW8Si5YJnCq6l9/
IjAdY66H469d9E3MQOSunsn72wTuwtO9cA+u0mYErfq1HN8hmaN2tfr/WF5gGFIkt1OBX0HCpQWf
6v3sZjjrTPJG96MV0xOsw0XGECwhI2IjG4S20tG16I2rkKNFJ5WvHK9vdd7xQW8ikf3yEcWVHYIP
NIW/1NKir04WjXkblS+jmSpRXuYnS1RyZ2DUWmO3Q8dFZx1ru22ba/QpYUXMzBcLJq8fS1w4xvqd
fflaX2F+jG/HXB20p2kaql48wdaSoX7WdvzlrAs+Ukc6/VSC//PRYRdJY+Se4FTqhNdQGGCi+V1d
adIeDIjFA08zKfvCdFElSmXMTAHUsvaQ6kPvc5DVeF1KI0PWEQXxXW0PSijFnENkGxP/Ai0fRKn+
s80rmQekHjFTimaU8w9rUDaMn9jLtop9xHITAA2kCEpLXXJ6/RLUVs2LSJq0SiYko0dlYJ4wQLCH
HsoOf+0YcjYCQ1UpM4ainxL33VyjXPwPXK7cmU1itjNxMWqJZCdRk85xIv3eQ8jvmOwhEPRQTCq5
EaW+SsUlpkD9bW43g9c9vUmCGQTH4puwDfpX6S8mBW9u0V64GGtVV/gqOXpz/ujQF4N9L9a1h9/p
ZuAYjIpgwQquTJMhhN/Vfi5ijDymsrog6TWGsBiUuAzZPbGl82KvAE9ojL1TOloxkUUxr4z7+reH
/T5k9R2G87s6kBOyoWrFNgBq8qpEuhmRwRIG3bXLJOlPeCz++0gISLT21tG930VBfZ4Yn0NRu+W+
jS3KeDXsD75uPiigy0tdyG/DFANxb70mvKIAqPPOSvtd4EnePS5r3ufBji1qbL19nhsWHLKrEffm
ZvoOxKxe+0LywLAcXY4URpj9Kac1104t8fRGaZovOatwx6969ijpnLoy2dUms9j1d/p9KM38F3FK
hWOOYfYWVqAaSJ99rgLpoOrE/tgD/YMZ7os2CJi2bw4dr5CfxBSbcMiYLLDrwhNfA4FeAFztYzBk
+k/RPAutoHjMdh/4MKCxav5tAFTEzljzzhl3UHQuW+16X53BeBa16rud5gypP7ryNpAinHgHTRly
sLCbyPyy6s0AqoAnXLhqBH3szWjfVfb27pGBrsTuCFnSoZ/NqrCFuOI/fzYQXg8+yB42FB2EZJ2l
cKOjJiDJpXPmTWPHjGn/br6uJKSIdmhy8pePWAdUTYItlGfzexVP4Z+YT+m/5I8UDNeTOeSTXL3l
4qiiOfF+YaHz2Pox/uUPPPYORaD776uF+9Z1gz2PV+r0qcp+OHNotA4jxuRzstGQRvCjvPTZLV6t
QKa49x9OiJCV4IjMBRHFYg0ggYv/pFpaaHZNrPznWKQ7bA370JdkMbVQvISu7JwtqwRjF7AvOm0g
XH5PCL2cuRaMFiLYlz+9EywZNTKTddhGu1VFe6pYQLoLOo2oSPgrUd0sASBgIEP9+rSWmMkI2C8d
x+xkjKdba9Ci61TH0VZ3bBaa0NqJIi+zkhVLuJAbmzov52hv0l6znn8gdsw4dQJ/nAWo6q5Rc8EI
H2tct3u+GEHkv96+C9JpevXXsggBmanF0xhoUEkH1C0FePMeqSEO9c8c4FeBCG2v+VEzsPTqZpLd
AMzDKFTJgAyJ/tLrN37rZyMftz/biklf6sn7mp/NoqLuAQT5wAe2nU33c1x1OcRC7eu4RSht3lOm
ZMGZ7SoP0qtUw6phxHwh61tN+EThCqbN0ytFsRk1QALEdwkS5oFCECR5SO+Ti+N+e5B+UPIOm/dI
dATq3nEbvvVjm66o7bh/ZP2NjkjrUEnL0KG68YJomm1edYMOHAhDvCVHozIgd786CCwmBmnoIvDL
G1uq4ISPdarx7CpHcuSk0jW387GmgbhKu81ETyeGjHWuHgqKhumA4g1Q4y0Ea2b8MzlftT3oVrnG
xph7Wzp9B9URzLGCW+j6XOErORnxZJaVpaF+s13/Flf0Vxix3036k25tvo23s91hvaZ91+Lzg1Cg
OTCLL/Ptcw6z527H1hrotMFzQ25iLLPR8HZ99vNYB2z48nSpRX/i+hnJUs/c+rNBgJ2jHc+dDGfq
LgJF+IfNEG4b+v617DOMklatDlpkjwkzUsDSpPvVG6aa4cA9MiV3rnOWVi8hseMK4V2Kh4zehXYP
MahqP22a6arDt1UUJL1ZuchyZXRq5Mp2h6h3aH8e55zQxYaTvi/E4w85IObsUiekNnKpWAiG0CAn
P34Ux/SyXvg+atEpwIMDoV5jxSmGxDGbNWQNvCZY8GtjGZnXBF9fExUNKvesFPF+ypEa+Iu6SsBw
3t+A8ViT/THsq1vO83NUC/JKin6OawIKWKnzBVJOqbLa9xSXZhIDInQSsUSqTALnc/l5efwBHq0w
0ro+bd5Cn5ZDwhnr45Lucbo9PVaIrlLBuR5uMjzswMGv3gP4VarwZYF9zH1TL3OKl1tjg1+4Z+Hg
KY7BlcWDoZQNI+kOVnJAQY8dh/o9JaxjxO0s0bDVJKarRmxUV/e7QPYOGzCyKGrsT9jrfFtDPqsW
LsSA7E5fHSvwGvgviCU/yDALWZP18P3OnjEZgPX7YERcpHZJqHhcfcyR2cyjey8SJeUvuFYtzS6H
Sx9g6eg5vYO2/1tuOFKwmbYWZ07rIuL8Pj2Up7DLDup1aDDZg6mHF459JY07kE+mQmK18ENcpbJX
yuL5uY+nmJNK6TMI3q3V6Oh2j9rEYng2aFETdgptM4ngyEKJkz0ztx24XXeVSONgV0n3BF8nOfXa
fMH9oM05Fz/5XfANWBYPN2CYdurBD1K+G5rBMjo9uaSvA6c3AZv+6L5HVfL86OnkLqGn/I/j8mC0
0F8CMUXzMjFrXW7ny2s4y4DfTrQTMZk9SlyAdX6ONrmjGU8t4fI9XN4hjwy5jAaw0gpBQdFnzlyW
clBaLKAyzwWnckQC2RAkFgKrV2XPv2ub2oIG4nzt+D51KE1WcPUiXbyAUFQefAk7WzihKH1fFuc/
lqOEQMhMzCGSpit9UXFXPDip12x39okRpGCiBfb/CijQVqmqEDU1Zrt8okS4uXb/9Zisg72TojcY
XLQ4WdAmaxjcIsReTUd5/lh8bpfWrgSc0LHxLAcct3AFbcJNIjTg35cH2aLfIUS/hOyCiq9pKos8
qOADI2IQQg2vnBnDwpu3QkMrcVE7d6zsrjIrx5lJ3DfY8WHkfSDUQKqiNZ2bZjQbK4jFVHrKjCVr
2vizJ+bmOCoXgIlKFlu+hRsmjWqzF0SZ+VgAUIYkwqr4Ygy/hYEFLHvQHPsLQ5LgOR1DOqkK7kBl
pr5WOWsiIE7Wb9x3jU+kN4az+Xw2KstHCk0PQVgB7p4p1QkhzpCd2dbVjXYo+4F0Xg8/tC/W+pNi
rrDQq3Mp/zpJF8WIeDNXysUmHEIM5m3qgfFDcW6ohoW3jnzsLeVkU4whpzvMTMnCOrEzHIE8rk+m
y3KCgShJhuNytpk10igyCe7vImshSP/JstZoJVhzYYZidn93aT9td9F5Cb0twwoaX7Ph8eogZmIG
yDeHhl0MTWAa4q62Q93gUvtKRvw2h/xGpieeinKkKj61uS4fWqvTsuKaLfdwT/50R5oRY5TlGkPO
upSXAkOfomtVu02Wx2b/b7zMNn3Nv2AWdTPIUBsLPL0VhCa+ycrImNaKdvHFj9hUFeTge+vbeTOz
APIVcI+x1dfFLNX4lm1N992hiCpOCogK9hLoNjzlH1mgnvnwc5pxuIAaZHi8HcU98lAXjuy81FB1
ZNg35nQhaVGrgV/OZmrTExb+lnWDpzMWHlYLnnJm4nIms7eYK/b3P2gCD9xVS06efRGqWQeR0zmd
Tvq/GV/oIjNx8ovR/XcNEOtODw0MD6A8GaI98bfNyRcDPPnB37y/YlQUTOLdnyPxzO6NT3XnlM1I
GKVct3R1ihjD938SJXA/osoWKPW6bYSqIykTS7okeZ/V+oxBvsaCezAYvXDw9gUIrOiU0BmhRTlO
EkHJ1rbq2IQbjsBFClLuWvUOKzbLVXBsQXlZ1S67l0U8y8u+gorKOLSQpzCzolthza2LsuNrr54N
buUgJAz7DD+pUAGZQqr8jBzK30WXAfuZv6F3o28z/wvzh4FGPCcMyI4rjW/35ZLy5bw60vhKEXIb
zrikiSKGdX+97evIUEHaAKOqHI1TXc+gZ/3R6HS3n853hJN5THJAvd7m37o6U0WtD2zCH1tott63
tdRRMZ2SVZbQX0b2dwxt/m1UjMJUTqWOa++6UxqpyPz6yM1z7lNVu1f4kSg8Fy9589R+wlzWs1vF
An7FKAh0OQVjOTrnVGDNc6JgGGjG61T5c9eu2zdT8EmY7boQXpyQ+3gcqeYjT1jM3Ye/1sGjO/2i
mGeapUouIDRGukYbqAx8cnAIGiQUqmCZvNv4+BRdwWeeecJ8zhCfSwEjBgvV48Vg5iTjfuPjohDY
4yApJ0H8NYykbmEKT8jm5Pq80j4xeBCsJhrvvLVuG98ccuWfa/It+2FiHh4zTkb1spxxG5xwfDBr
lFAPi+Voh6JCBv72+S0xo1vMu9reZ71ip1rdkl3W8ymyo4tRziWCTzTFcdVJAoOMoZoJE9VZXJHD
Fe5Zl5nl/3QrsOqmlqXkcakPaPKYBqEs/QWk8PwpbVkN4U4zRkCu8GeT9lTgLpx5+uTT4p+xh/9V
7utL/MMM1QuFi6BFraBF7AgLN9H5aZGEIdHk36lZHjNu+3GHDOnH51oKk3C/VmAF+sbQH/des/Oz
yCzaIwJknIl3+kZKYN+JB8Ii7V1rOtwCe332Mpg96MDEZG+N2SW8n8AIC5ZlhCyrO3wZm6JT8K9S
SjA7XeJFD66IEBhGljrx21IuYgv0AcW7VHBX5vcZy4UIGfW1JjboT40XTev9XSaAcRxGZrHtYqvL
As2d5CK1k1y89pf0sStr0D+Q9FZU3sURUFPiJmTQRb+UuYGyc2H3r5xf02ByEc5yiQb0UYXJ8f+g
OktscegY6R6dMK+rPp012qMA7yUUTydVqmmR9CZt9y/OshSGji893bDfHuNO3SjTPG1Eh76zDNFU
g46RjOmbD1kRNF8FZZWeg+i5Fusah9P6m9DnDsF/ZoX63wZzPaPkKIbHq4OX/1YtT4Db70a+SOyf
myw0kFFnbRe255orDGlCn9NFzFscsaq+YI5jmXsA2x9hLKr0WTRVtLndRIDlmZLwvKDOZav/c+EH
Rk0N5lwtFqAEe5cIJUZTnfaVisiM1wNjv5d/lzIoi0nMy5MLSkgugTpY4Ow0Ji9yPkSjfkIVe6kQ
fByX7k/AVnw13fwdF9/a8+EE1T9u+8b2Kc9xBqGrt7Kdkdhz4SIaqhAtyd++OpuF6HPYgL0NoLSQ
jMEWy5V2sryiJdVgylGgGDL5eleCUJ+7AypJsD/X0IljHLsnkTKkjrJn9DqEhTEG4j1HCt3lgfZD
5EST3fCEh7UJvxvMMA6egE4Ut+YcU2XllJzchuCRQSC9nW3GRRrPktyz9921LLM23dhJIIpV+Z+w
m3Osd40+8c95ArR0qQSDRgm3cfs0XsWXXfFP548x8CI0CJjzlQVOdM1lHfbD2imhTKYcBIYqxj95
wSTkoObPNDvuQE6BMo1TRgLLj0SlINL71PGMmY9Qnu5Gn+/g4RHQdiwdf87AvW4GvoV/++VCBUTU
qAhXtMuP8ZmvtbLEXxArMlDLw7pSa4Wbmzmc6vxgcVfujh5/7TKmaRxlnbOZcg+7UYYx4jrqrgVH
aOiSr1M8bZwGrEVE8masVnbxKxaP8G6662eUsvVMn3Sph6KHcuxF+gmvR1+jjXXnBLsHdyn7ZmRU
R2d9YpLZmhaVUQ1UvK8X8jo4Hu5xpiKaZUqsAOZz2ojrrUP5jhe6AByfo69ya0qSheOubwoTXRqU
DqUufHarOH/y9JO64hXqjbLdeOMPz00ifQ2wLLkMqr9jARcyWGRVij/i+/MULweIKye+FYPAyssw
DSM7LsUX56aazJGh7yfqtb01FQyU67SaRVsQFVwtObAWQ40+aeYw9BC/bsHYgIMbyuqdt69wUa6M
bjyu3eYD6DdRc1CA3L5y9EkYqaKEYE1eQPxcs4HYUIuRhwxFgzecp4q9rHp14hl2EC+U99tBGpPC
MfvkaojzQFJVlU6sacN9JzFP5IENyhHatfVKo5raIYA4sNFrbrpvlbJdkZmqzqcV4B0vRUHELAtB
/h7Eq+/VsSZtU+f/kr1ldO2EasSfKK4EDFda2gi0qH1NfyuUgCqCb191ryIzD1Xg1M3kmGhbbTxj
lGNjmkO9p6npqOvTtJKXaGx+skxUjklEtQKHGoGHOC93FsECidmoB9JWlj/QfFxGRZ8yZ/jFbxIy
VXGv3bET43IsBkqrYv+Zv6LLJp9/aXcQGPg97wW/wAEkFK5ojLab0w0wh9hlCSsnUcd+nhnk2Scr
RFcfENvLncesHe5rDxdTYbf7u8NVTbGG00YnvRnnI3Otzqa6bvNcostoMRAmSwQLhQ9DfzHQtHJ5
6GQJHAiDCFbJFeTA4RCv2j9WFQBRXvewouqUFgXCVRYK6O9s/7cOCV768cT6wrkxBZFOwMvW3ilF
dXvM4GkcB38kV5WYWkIwEjwbqnKb9HkfkJUuoXrsEBllCv/8tn1zEIH2ax9RuT0Kd0N+dAyp8xbw
hujsrSnnO+ZSlqFrDPuiEHeWaZIMPGjDOJxNFZ5HxclEhOFX1ogSjAW8TAsclZWnSgVxHPun2Mcg
+I5VJdOdndkuqkKwfGpFcMsMu2MVe55IyLtlg6fn3rBf6Lzt7qZ2XB04gwyxDOv0/D4fgpanMD6p
jgGISsQcqMEc2TILGyqLnMWK0B2jTKBe2UbguZnY3CLekNBsrfiQbZxdLEoBiT+7NyJIISNgv9nI
Mxso7u8wxP6na09IswSh9ljHqo/JOd09784cibIXlSd8cqayCK25djZdlMA5uPlxuKzwD/5lYBHh
rjD7oRc2WmZfR+qi1sxQMIEVEoMKYswnG78bCUypkPdQbg6j5K1JpNLa05OU/eFUBGF+yuN9iI2N
Bpu2nkfFHr49kV2bJVkr9bAgPlSGpIARZJacEwheCFFTio5gN0Maaxdg6XEmI1mj1BtPvJh+QkYC
9xwQF1J6MDi7ESrtz998M3fEuY9k57ZeYvHsNdwIFf+273C3TjbJZ3Ju07jZz1/sbcpnCIe06of/
28Pbmvsq+CZQQ9tzGTSmcgyWp686gIME1DpZwtC6+4hgjdZAgWE9O26r8Loa63YEuG0t0biS4Bwl
A2U0kNQKRjZT53WBPsnVapke7+8IkeLRlYM1U5H+wf6XrYWlMJkV3gCyatasVaywhgiu8WxRazXF
k7pXk1SkQvP0ErlB3kbW1ppLm9xLx70cKkkjc37aGQc9PhcuznxXRx0cI//sFbu8N3UZ/G3k7+Lf
f5++38HJy1SAZajEeuuG+hgs4tjJJziBtBGrlCG2VZMior8kUe3Rn06AZIfTT8jg5Sksl4uUvIW/
DsJZgKvlw4F7fE7tMIhJYBW3WemiFkNsE8QGNJbUuW8weUv+zmojzSjhyQZkcn867ZCJzRBcHNLk
0ydTJvuZK/nxmY5RQlIje87+W7EiMrK+G545U0n0yrgG+FLnuJETA+S7gNBx3T2D5jVr0qAcXMz/
If6YR5Aom+lcPOR+LQNtOGUDxSeIxMBHTYbz7izWSTdxcscEYU6MziiGK1T0qPuaswwn9/fjS4YX
Hy3gcT7hPFiFW/mJtcoH6bzJId6kXpyZJfXVPWsqwM6p/OXw6SbVUvGvpckyW0ZN7tDo9/Ipvibw
C3/euC7qUyqAizBgVwAZhm7EfcOMTK0QRJRD/ktKvYji0qsALG6fyl0XZxKdzEixG5M8qdPXuHUq
wc/Sm0QkqiIzE8eFswY8v458tLd3nT31Q+qsITVbzMH4afsePSyXb1K++ApT9puSmXgCojmO7gek
fLB12RMeQampZkdO7422lj+asPwQpqSW0BrgFQfQxISzVWbujY5SeayRTNrxqvpAIC7Kv080ProD
Cd/R0bar5VV3rGS0JfJ2W5BSIC/B4l5yHk3T3eAbQ2DUgZXRG7St9+77ngaqZlg/7A/xDk0hgfb0
6p+ZvWUEt243Q7pVVjokcrz8TwnC46i30ggW3USNO3eifL09r8pcHbf2MTww9GJCDtWnbfaZXohi
dg7ywKC0XrwfTXP6pBK5U9b8mE5N0ONWWI1GlCFGbxfZaaRd4BFhoKLqN6gNHuzei1ZdpmUpDJw/
iZHlbZaBDbpt5jEQuF3Bwhq+KVLZ/RNlu8sOiwLJkQ8tuYgPOxBjH36V0oxAsFqvboCwx95vDNUO
ZdUDQWYz3/7X5lRZyH3v6BOW7FCbF+5zV6IVsoppfuC3RRkelJllcNGxdY/pQYXAAOwim/+6KZUj
DRgkvSs3U+4n/o6Bwb0Gabrg0XKJrNbwiwaK4BU6l5Yxh53eQijXjsorHoCsYH6tMNDJCaB/mUIN
7ysIwwMv2SVwzZexYOzS0iaffdL/JxQgbH/SCsimtK1aKeq8FkDsIx9Pxb67HiAzHli73nhWVe8B
ZxedK/mM3rOfPZhQfIeK38A/OaUOfmgN7MDKfWYS+GVyT+QuGczVL/+7swHET1vwSdhqBSuwAdZD
flsV4P9MmQbqPP18CGL1qH1nP3yta4782h39EZEPiVTMxBZlvitaukwy/6ExJ3GhZi+fNsbNuIwb
Fj1gWxHWMnbIPWgPjez4kmWyqYwoUpSlWjim6HcBtukcVmIrp0VYRWdlmeb52KfUMdLQNBSBpjz8
aXJrRkUxJwcYWdjKq1Pi/dTQdRo4yysZuA9T57rrKpDhh1OYF15L2FBuRX9fXB6uVmghOyBGDIyu
6Wd50P3BMS3yrbzw9/jfT+opshl7g2uaXTWz9i5XRUC9hL3wZhsw1e0A64rBR8kOQ1ZcQ2JRY8gF
6fPTDBzVpalKx1Y6Nm/S+eVCjwn7nUyefeiUhRYTHnAR0lqzr6D79QKWp4iZYEXpzqPuR/sW2rsd
K6bocnzejSjiBGYouh1NzjmQvmVhJe3M97OXJdH972c7iqdvdposHJMEDjxgewh2+1bMvRNYOH7y
ohNblme/olUI3/GyC9A1Hx7K8J3Ht7d7QVBBbuRjAQjBTO2ExpQIgA0PcuSWGevycnfJi1BSi1FE
bqA4g8ltHAIrcnQgjyPV0T2VimusPWj195svB5dEDICdlfwMbH5zEEDoJ9CmAxyLX4H74XT8Jef+
pnrBU7CRFeim4TNWttWXB4eGZKcKnxSWxaG+gMo4qad0O60SSjnyvFUxYWc/6ok89LXOVUM9LItA
tO00DeKvfZAQkBfaIcjdLHATs3J1R+n1ieJWjlMP2ol7/0FMXboVnkBdPCN/0ng3JotmznVucSAZ
zH60wFp+eBeIwCyz46ZxNO2uRCmS9y+hj7BmIfr/QAW+a9V4quulaGhT/QwYrBumdD+RBIPi5UHq
IRokmecmwjrSTi63fxtPxUvotBouOVaRL/pB56NIIo1G62FMTSwXtkmTgLF5O+JrCnEywR2z/Unn
KhwmXInT03+w0ja/zwYHl1sh13rvXZBUo43np40lkq/vn5MaEKLoUqGKOor1Q9IiVBPv6uk4RiNR
ZilRGWgL6EpC0ABqLpqFwp/41tsaiU72sGev4MtPGH5/6DqhzQBIS3XZgTcRzwRblo4LjRGwbSIR
D5PXVGwnQRWJN1hZvurQIpF/SRAWhbzMaz8oEIGMy3LwZSxqLxdDbU/IICYKSrD0H2rmYba3+mGj
LCC5kSozR/1HVOcRmMDUh4d8C0mGKtHjYDiNQeeDgJBs/UD1G76HFh2fqFZWFeEIK2SQ3YZQPcHR
KZqUZPWDX60GI8RuhN8MdSc64uujpmxu5s3f+uL/gb1rjHp/+XiCOJQOR6FnrxCuOPBT4JxS9cxd
KIw6+f6ceDi4mD4EIx+yryv+gnRYH1mSQqJZhUJQWd7MSzfHTcKw/KETjdso5CYhOkMF9aJIHtTX
Dn6EAF6LdetezKCOT486C5gzwM/jDmlDCO0QnH4v2CQJ6FipANktjsd/Q5vP+fT4Ay0xe5kMk+8b
zGJTgg0Uoq7l848hXZvm5NzIn5z6HwDnXW99m+7jfJgnfLrXei9JqKoSwX9uh+/Uu+yem/YIj3P6
kVd9E8BzPZ41KR+siQiJUEb65CjLAlusKH2GLhc6KkbJ4rZElhWXgk2F+aA7ku0CL5KCWL8zPdjv
/G/yIKTeSreMtCfpAPSIQi4kSRSPecTYKq6NLR9HK0kittJhmpJ/7x6KgV//MT7Rb3r4R0qEcUKX
eRt16LjbhFHBtwfU0EHXl7WPzfsIuOLXHAmG87IlyJgugPvkI7HkeJP1apf3Tgvgt0vtlYYCvnzr
xSeSrJE5qKSqZ8YwXPm6dp9PTZhwQq8CaORDuw+0/AynAwncJBvO0E+nLCmJ/WIO8qBDnk6s2WxH
C5qUkQL+NiV8yADQVp3LaLgFfA2IP53lfohMgHYBzH35YbuLySNKGdqFVluTCfuJghmEiR6BWwJx
izga2vhJ/dEvimyTllMWqD7n64puCcRPBpyVYBKZjsknUfOsGWyO5P40exI8+HgXhPvRS722r9IB
4KMDtU/HdyJqcP5PwgLcNTuMSVWm3emSQzUqlj6Xz0S2AtcshwdnkTP3WgJFRvvrNIF1hYwATB3+
HGMpUCNJTWfVZgpoNM9FggsmgVBPuAzL/medaJEukwjlhn96jnbJQexene4u2ua/xSVtqjit5Ljl
jkG91FUQpA0gh0UOmicmGgSHovYFUFlZrMTfIZ3wTWzA0Vyw757ieJ2dlGnAghGWxOP3tDvsn8gq
BnPUPVqToMcbie9vPpI5ceCcJ+Vycl0sK+/T1mLQLMjXNZ+VJj4EwopnjfviFaBFuqODCrp1qPYx
aMhKfPjhmF7Xdfy3EmnmgVJf+y9MAVweVAsDi+lUxX89TjZ3VZyCky7DiHxLrBF2YnG4sZRFlYTk
wisi7lA1EiKqgojdwNCBkgjN1SA14ehpV7CBPiw4lKsOIK2VyE0RCzrMLrDxGVrLrVjJxrtDsulP
yGGRArmbCQJz13YvSTWj4FsWTEHY9ed/w5J8yIaxjAlne2WwL56OU0cjrzy78UiF4fOlaBWID/mZ
nvhWbJPaUXoFXelI7yDoDw4cDBrayIWQDWSaGCXFVi0kcghpzuUb66RlrZrAZXFGazQ5McG2vjNc
sqih3p43xPBonpMVO/f4DP+iniWeJ+PZvZC0EKTrFHpb/p4mdLghtM2CcGqycTmoE64RCOCOaNWX
sZfJL7JtLaGD8gRcAR2xgIfY7fJoPcuh35W92ClUhu//5EycHcNAP1d7U3yXkLDAdhRTUrdXnutt
9pfzB1ZBAi4rMuT63JFz55vG0napuyb7rMm0kVs+6/vXGRBz6FnUMkhdkfyUvOFphVof0C+fysQa
NCQ3iny0MP7vFTtg5XDQjE+DIdS7MZWkRaBmOCZW3ppjs87FclPrCvDNxyFsG3mHbD3bhQFzjkw9
8URvWNE/du2NKMqhLk/wtuPfEr7FHI2x4D0EFMxAVoHA7D6l2I1+jWseV64hzFWAr24BR+1R6Tr1
96bLuV0N/BtZDkhXaOlp6E3lius5wNzbhmvFJx7hEHYzJ3zOouUPDl7IjWjyy5AvKBM4i4wtv9V4
uSlJrUDl0F9w4U0dipYyEA3Nxa3iw4HxWh8lbnIW6RPoaIpVOvceV76hbEuOjq+4opinw9HswIqj
3mRj9km+8hHtrgISFKQE/Mac0hhNvgkfIq011e5Mxt7q5YHKitgbHgnSdRQm8RwBJdBLW7bqulyK
E5EWSVgob2ex22mFnZ8IsAYXhH6kC1DM66SjvEFjrgjqybvfGq8NcG/OR4BfpxFmSd3XaPTirKRk
iJgr7GOPi0SI8JXjcdPPkiLCrD94dJ79pXT5NfkgVECJ7yZ44R2enHK27Bsuw8mVFPLLverDk2oP
vELp0SWmMVSyJrmSv2daBqUuSG4MRG6o6DaQvuJ6LkQCsW9BwpKIt8xlzOdmz4Maa4kvNlzZ36qG
hU7zv0F5CC82klh7Xfn87OKQUq5WioXxxhqAq+CFGti+fv1KvM5cg4K1nGkirxn9Q8KJEdTfdOWN
ti0cFnDPKIKUWDMLOqh8Jmr9O0X9HQbXnB7M4p1MISXZmmmViPiGYK0K3gIYexLsBUTTypR5jxs2
87LFKhgIXNSXMqR2DjKYMemhjHiR9feTfXt5fWRL1dqTRuXtb7HC8Qm87XnXNDV8CkhyzgHDMQbC
4WAQHXjzGVKUofwvZZDELE2QuKbo8bU4LslnEG2DB2d26r9KjLXtPdFNC01SbHZkBEB6hzSmLoKo
/fOP4NqFmG65zzrwJpxdKMJTgqa8brNP/f6R16xkYzFuqzdlGFvDNb+jDePhkvKIlOmXiJdtFaOo
mblavuKPw32OzH1neuBuUyMIIXhJ4dUKAKjziVZuWs/QiCD/nv9YnJ15B/xWtdOZApJQOlEVkhKr
lEIMILPzp6+qFdekYxKjKys7GKs/exEsr8Tkp6dDIT/uy782KFZNo/F0pQ8ezrBHoCV/mGWvGCqb
uCVAbjwSKDAHf8/jaqyQOHulSP5RReFjYpg+e2vcE4hhLxYetR5yERsxK5KM+lcw77ux1J9rdluZ
9Yhb9q3JWup4ZcXiKXF6NGIP7PyAoBTknFr0KiHzLM1xPVIQzTrZSsu9WLS3ZTiKRlhPol+w+/ip
yQEP6GoOXSEXt4jP3Yy0OR7wQ3DlzWr71uxrY5zpJ3xfgWZSRP7deP81J01cKwYX97J6WB3adHrR
QcYoPtQgXqrSHoNlIGfm6RBb8bCuQv0ym5IKDL6VGWOrwqfySqIGwm6RvhX3W60/3Fzfpn/FlCbC
oW33jZ0gZIHUWmsAUdEYMVssyIlJuyaw6PMblNvqAgzfvgvXq9NFFqWkvHJvftT+o+/+dfDuX39w
7wzAptjzTDzlzuFWChUFJtTnqf7ORDGpuou5GQ6UdBrw0nnZ7WAxHnbvzANMrMeQGWA74C+QBO8Q
2cN6ZA8y4R4xI7SEoEhBKKJtKok912F3mFd1s2yM+sddX2nGMfKMgxnolgGOZOD475MPP118lAz1
DSCxRNglodJvq6rYp7ugjBBhU62diB2ECVe5R+hHo1fW29xQtov4hX1c/beVtYujHD+jZKjdzJcE
kJzlsjyztWnYVWkyP0JwUobxWrnD3sj2aG3Iv6s5pWJGZgf4EJzOz8d+suUHgqUftLblyPQm8Oxa
LGhn9FyaKWpVQecRcwSI8Ei3XEvA0BbIwBoUgZsDA87inbgsdptiJHzVSl57cC2882jdh6A6Tv6/
uwyk/06dMxAeN0lx9auIVJJYeZQdEn0fRsWO8/kKZt1HlxSDq8/R+RuE6QJDYWBPUGUGu83h/l7F
z6NKYG62SI4U1UNJVS6GQe2CmGHDXt4drMEJMbUksqPQYgyR34A9YWd7uvUja7ie5O+8PhS1USsD
fq3Jw82/ZxbOIz5fgBDs1n13H2apD9F3IWHGLJeh9Xlt0dsPZLL0hUaPt+ci8OWTmFZoxHu4NIjj
/0gYvfsOK/Z3UxUd85SdSofZ3X0Ld+STOtYvzwrIMW9kGZOJj3APmrENxxCNVsEZ1IgXaN1SeVU4
7ZhcKXKque8W1DR7taBq6gwWO4UfjMNVimCnP75pP423FjDSIXRQ3Eol8OCXIyARrZCzf+0tg/9S
cJ/2mQjOfHzA9auTH4IBz590D6VmFkl7KoIXOuGrcqbyi2hdE+sRkuCSDJBpqsDzVbVbdlgeM0+9
X0dVv6wY1Ns1oCRcOn0L7vjxnFB6vJndNf+2kUPArBe3cWv7bfjdwmiATDFwH192LobAoYj8nKsl
Rc1jc8zocGYQIroOnY5dK8l4Vhya3AzcXGXA0YfEyIRtIESmPapqu80mxxAtAnsoahdTIiBXxX7Y
BFFPoI/uMQZy6AHRh76zDPCW1EDPB0HeZ4gYGatVKDswuxfwQuc30Ugxf2VG0s1TVIJkSJU+KVen
XRtTyHN+M3UsbjLuLmTqktiKlNwS7dpCvU5PzhmcMAikNwgLcyklXLU2UmJeYkNFDtmiyAQwKEnA
ZEbYmpfqf2MU4zK089pBSOLrMEQNt0GgWxmNihkGqELHK7wrVw3h51Idd1cZIr8Imk1NYphWAZaW
x1qLpS9M4LjOn6KdZkTw1jOUv4eYzF8ZkumPAW9ftCyYlpDWiaPpjsAYT93jKsBaNEwPicelRwQ6
unnyzyYPwVjUgsLSWKLJDswALlwc3rNPI5vk0j/lR5X/9PUThBZJZuIdh3ag3R1Hrhr3uQegxgW4
Sn1pVkPMmBYtNiP1jiAJcCOvjXbSkFaBStchHyd9prPvVUAM3pPHaTLkIaTKVsCgTnRU6zOkDZAr
SCbKh5lcv9TRSQ/j9hCUfhRPBp3HKu53I32GSCmRDzPu8kQC50vzy6zjZSobIJeIW6ImBepbIs0K
jpWriwmvg99Dq6MMqYaNXf6zoDccWpaqvzAoPxZeBVp5NRjDTOKxrDBUb3tFJxsJ6cSTQnfcwYjk
8qSs+3pxrdDrxHRDyDyiCOnzmelfM0HMbtnAo8UDXy9eF+1E4cjg0Ni8xM3EpRnAilqEWSOlK887
PxH08atOgfTbeojNWqKCaXbFO+cjo+ogYvl7QTxwIrKa3/locRFq00/0iByBVzi92HZTmt5Lhr8T
0jdJG609LKVMnEi4MnaTQ0nmh0LAwynp6owL7Rtcj1lYCSJIuoisqtW0fwFzo7cwGm32BHWxwKs+
3RlIVI7pnKHlz/6hEciVnGFqjhXrn1/BJpVvEl3ZlafNqBW6vF58Sq7CXrhbzOea1i4X0OgVU9FR
BN40p0KiwBBi4vPffDhzlGeG5ZTqHzimLgezAYSbpOkacB+0HFOEIqmcO/DwhKmAROqa2jaoO/dM
U1SeSWQxHUx9q/e6GaeZ3fXi7k1k/RYd5Vn7T3UuoXgqhOZYyOuzeu896Q8bmRpfiCnNhgLZyil2
t0FURNwYW6phW7nK5L79vsIVkZ8uJMFSt3wxEz/hAT2pUW6dEoyorptvixpzPdikEP1cEyjROMhO
Q6pXVdarh4Bi2LiXIriS5wRX6Is8jJSIMjIccRkm2lq73AWNSphxhUmNFvC+tT3U9KcfBcUSpCdT
rveLwmlLIxgUZvGVf1VLS46XbSrdVLWTFO1jEvSvLdRHbb/Rq8QY2c2W94ogPs1NDTEBI6OWPBDh
5gfmXChSqi1ag1OJEvJn7WPGg5sTp49liouKPjHdr0pnZ1mOqd3E0S3M6vcUonf3oTQeumt7YoLZ
IZpmVhnFE389rBDvZzdMTfJK2E94q1DHDSLJPvjvCiK6t9UPgFY2j18wazlbR6JILPUSNM0iqs2n
r95wN8dpUyjh529b/dv4NcF9Eq2/Md7XiYIbybm1CYMkdF5TEloCscFiVgSqQDyYTl0aJwwnYh+H
LYTPoh3tqjRj4PvaMVSX1fvJubpkiCUYnA/kOa3zDYd+/q2dJg+Do/jooBwKYuJk/3bsHq5+B1XH
I3pu0tI5YkNJpMsPc4P30A2yDumnNbj7Ks/G4H1zZhITE3CKsZ7rdPczMmiRF0aglrrGW/Kyk+Z5
WJLV7Hm99qB8l1PuuchS0yMsKUKHnGMv/PCRO9ik4uawFAtRaJD/ovSxKQKBWAk8zSjFG6WJyn8V
tkY/PKjj5TJagp6j8oaeA4h2okBl5arSK05pw8+l7yJGbyhP7vxWy2h5m7LcIeXfGrpI9pHWYOA9
8hMV+1LCulx+5HV5JJ5YXuWKiUNcUJuyYnQdD6YeCdXPVZcr4uHWcUA4G/PXW6uM2wvXW1GUa/ut
KbAHgdA4IgSl5ro7q9qzf/KAIoBjm5ZhYfRKGbRQEW3v8lxrziFXE2QnSRnxSD6XeOzqockXbRTy
Z7Tz4qr0LlI1i11dVC4296VGlbEm7bn001GxL6IaL65xS374BdtHrGWvzBc4OxiEp6IPIEP+33iJ
RLP0rnwG/hr9wE4oZY6UARJAI+1FGXuUCLroRtS5kglFANnIuj8VZyx1jlo/ZNN/p/TAPPESGiVo
eCZxa8Dzja7TyaCixY7FBucTVN3XSiQ20KbT4+2wLkLHsm2WElqHYiexpS0sBBQoJ3i5nFplNeG5
dqKSE6iF//48X8Cy4lUTPG2G0p5Qumrzq1y8g93ztNLsgpO21tH49CPvhHW0YmCq3Om5RO1fQaJ0
E1XqwRQiZU0IBrk6QEw5l3Bt6f19hnfQ4Nvo4URQ8F/+OsZXfxr8IBihqgtBHw3s2zqDAN5ql+eV
+D8cyHoABAtZ+QxpudzlA48ZPQXucvR9dRv5jb17RjerNO2yww+BJyc7UUEKGMGfu2vc09Be0zFw
gOGyCbs3gwiPgDbqS3DCOrlyh2TSxM4L0r+0pzhVMUV5g4BY7+P9HBm4qE9OTVhC7eLIFfRHWZKM
3OJtyLjIeZHh52L+JKB3JgEEpA4n8dmuA1GxAEMAs2saDp2DHJB/6Y/3oVS9QtbQqjHkJNT/ZfWs
rUMT+8Nx9lc8LMiM3o7alR1knrrsMEZfSL8qlQ6qvJ9nWY2PwVioAD3HxIFTdw4OSpf4B3+4lHeP
tRtJGbvuv7O/F6S4gKoKeRqizroA7+uxsvMx4lq/7s7+tJRIPV2cVnLu6jYksmuRHd0mwtanR/fU
DvIzzI0S4P1zSBu12Nwl8fQny2liTo1yNHP3i+0Wef2kzu/IW3HokdcxR3rXMeEdsA7RAph8WMQY
ga2qZwmQCkkYhLPHTmkk78zXXViYFedUeIIf5xwlkfBJ+7KkgHAmfKsLhQEfIhFUoR60gydJ6jQZ
b9awZP1LbR+6rSIF1d/SAvgB6lNfLf6rU+8qLx8rrU45BAhc/VSf3rYIsCeIixPQ8Bt+9pp4EXGL
c0gaDpXJyIaBA7q+IIjToAJqWaTWivNOz0/15Hy8aF56FNqqkROP+2TS0Ek1zO5O/pkUCZlhzAHn
jjdW042tpLS1ge8mE1qETqh/Uprg2mZ9mi0r56ELm8QSWXzd4BMj91QSQS8dc6xRUdR3g3KlBs7G
AjkQQXWZOH60hOTgqjBUk3A4RpMhCbssyY34pKfRmmJYlSuuPJFSe1jzNRvdmg/l29QPO3zYQpzw
JsHDKExpdmttqt105olH8ss/JGGD3iwoaKThNXAQlOwv7Qkt04JJ0XL/1ClhKrXo1Yr/qgeNNgIg
o+uZ8Lq8MXbdcQQ9IG2jWXy+o3WEHddSvhBpXLRy1bXOr/nEHHHkgQhPvMOm4abngYdEa/+rLWSN
ET7VXznIPXQIkzqfvpuUgCvXGxRXaTMlu4JfW/xVkrq+ROhCTJaOEmHY3BBI3sT1jRL2cGL1aO83
Oaijw/oLTeLpepHiP4C7pSrP658w3hIoLHbV3NGS7Y/9IoBM6kBbAd4bx76cTcwyD4GInjkJq/Dn
ozYfYzvv9AotOBGeH4nkC02ObiOq0MWYs7c2y/0JQDswtBTKx0jNXm7+OZOLdp5wLf/MI7CX8UBa
G+m05WkKhr3nIXQ23T1KJnsBbgP5rYXoavDHZOecUj9G/7fVa07MP9oTzt6BfKexnv6qfrGPKaM9
govj4s0O7qoPCZ81Xyvs4+dlUXAidMLcMdrgrq+7N5FuMMP/IxrAXDHRY3hIEeUVDMDrHCQomiv+
VGkn/314B6Ah58xw9d6RZNUGqFt3+D1RMOcVwWIU6k04HP2RMd2RN6fY2gROn1HTcMBsrW9eUdfa
v7pmRDvAJ1LB3BkEtIplQiG5SE1zHwyn4R1VZZ9nVumTX3BWXzFlKoqBOeWtgL70MvBq00xrEORr
hMjRE96O48PaSsT127DXjEvfAfLBJhyQieavQPoLNJwed1g9R1g4hbccwPeTAoDEnTiOa+7ciyJM
8xemijbIYhov7815dxZEZldshmg/bOJ0pihilr/0W1zRT6X33kA/5bHgS/P1nruC27E7MLBQ7JMV
CbC0RV3Ar5BbySxZ9uLRfI1ic8z+p1T/qwrRu+tym+aOqjt8md8qhsqbKdV0Ngy9KsabripuTMuI
piD77Z2FIG12sNiZqFL9raonOrqjKK9GMao1y1LK5U7EEchGYzzHdVmptHOXProEBnhssKNdNhtR
hE5ILTPtocELtWZNNyfHKjLzp133ba1mLoOK9rdRijEmdLx6+x1lrdvb7+b1vAV38Th/23Hbp+N9
idTmb9tA2tzhR+vP2zihHKup1gUzc16OdwVHCVhp70e93tLehkePof+Q8xJNEf09JwMPQV65gEFM
2xOfMl/0DKl20oYv1+bCAvSxBazx26Qys3gRrgX2ehhlMW0FhqJ58A3i0G/EuqYSyjNtuEI887Wo
PMLRvch4IXWDM6ajJy1UhozV1dadADNwSZyZaM36Eftxzjqn1oE6JPi88tL54AtiFhpGy4n53Ok8
uUflzXuG8OxQexmCx2I65zyN16CPY43ezC7bJ4I4iS+z5Y31vPeKdP4aPmwTQAvck4bsNNI1Dw+9
xxxjqALlRBJ1Bi8zdojaKmi66Q+TpEklR5E3EWXDRjohc9inZnu7UC0pryPs8xHPo19xSOvROX7M
H0sfZ/ZCzd6I9SqmV+sXpU1bLuI/WVNDtLgbzY6XpurgdkL2NPdFBKVDgNH2NzH1dm3iVqsId7vt
1u9eTlUX3pgNDQxWUrvVSjN7GgHORincPaoVpFJV+UKQvSiniP/VtiJk8/Pldv25hJeawcuqtbJU
I4dbSf6YFkjob2a/x/2mUbWfdt2beGtXvoEqrhIQ6La0urUCfz5kYML6Y2dZd7DZTuGse2mqn5wp
yFCpVXNOWutEfxzZWvqeJbf4isqpiBgfc1GlQEAThEqHrtX+SIBVMYPqjnHGGA/A2NciHMGOgGKH
PJHA2dzS+MUnej+BdUxLjG6STplN4ruEoWcw4eZo0keIETVCwcXRGuuUoh5lVAGadXgx+2exXtIi
D18XVRsmJaWEhCwiFLBAyumNdIuWQgDSoQRiU+HnwbetVv8e881b3Uxxlji3jFulpjf1TUwSJs/O
hsFdQyTkO/Grw0vXsH05YHU/ZyosiIg+xPwjpRV4R5SQRwwdKiZjxJkE3KdlQk2FW5TSiBA61p4b
4GRZl0E0/P2Jk9Kw1W2PyUMdGtIdW6coqK0XGeA25/PZUI01wQq1/reZuaCC3uPNr/p/UB0iGVTx
QsCSAXnOs+WMTPMJwq03b9kFuRAIUL3Fm52u/efY1FvBNA3rohooqRi1OqL1jtzq45h/UYLLohMW
ojRuKZNNsBL9S66yzDmQCwhubRGcFmrDUeTCUh4C7QokzrQKAEm/TPy3NtP35T00fN+Fx/buKlKm
p4/epX2JjhGoQWbh/WUNK01nwAgAUyPL2mj0KtxJdYuTYR35drFknjyr1F6v+nQO7aanPHK4jjaa
/mfvIYREfjlHEZwaoxGaJnrV3tBJouVwep/EhiJLXHMbdBvIRN9wJGilemFIqe6e5g4Y5wP3zrcT
LxttqZo0+JjBLv5Rn6kyEAMrM1bQ7S9MqKRwk3Nzt1ZF649NjIF5PthFVlqxCNLJgmyP7a3PgXGJ
5yc/hY27jPLfMTb4C1vwewDg2sNYCN7myGG3nTCVTnWLOkjnka2wgOUUaVwzFgm+jJuxYzTeO4Vn
mLniwbNLxs/21qCVo8blA9R/R6cJ4Kqrx/FGgd8Qz1QfjYeFh66D3vhw7ROL0/81KpWfOwi8+q9F
vkEDO2LaIK9llAT/nSs4yI5pP8QV6zoKsbSTCAvGxVkchWYimhhKT4MQyraF7TTC5Yhwjt4xGqsY
MDpHw3PpdxGcXgENOPVIDHT5mpWv7LcpQ6G80GNBXnDibQNHN0nTuIUiSIuUKRm1M4dv5CaRpldo
4KpjIAdulyGPN+mwTARRq5YMBLV/QAdj54iuJENkK+ic6epaqHZ+FWB3zoRgWlZ7bLgg7jvNUagG
J7iA1CaL5zn7fhgAq1dyDVOnt3iUkkAhIfhHobYF32y9lshkLsnHmVtXbv6+7FcTw2BJQYxHg3en
XCmRSJnvzXnjkhs8NQk0vDf8kwQ8/RxbUVpRLbJIwJEc2Jc8tomNnuRGUJcNF/geDH/8w7NVrUdu
dtuB/4JTi9hr4WG43S+dHDygb5Yd7QEGrJBl+sjSsMG2FmZ3QzcytP5m6JR/ypTYE8WkSIDjCkO1
vGHK3lNwt3qyZAuAzYyXOWBLQAWq3Yr7DXr/YWyoGZ4UQCc3CMIou9fgYHTnpSlpiC1A3eykCP3r
btIJ9S9dfG7bI0eTKoU9oKOTUu1OPECjP+MTCnyZxoiwTm+lEsowSppY7nq/0K9fgCVCJSdkJwnm
oyo4O8HG6TFqKDKegjlkr1kvlboi/eMiVhuiNuoFKhiXZf+qGPkbxePseqPA6xkV5QN0tSAY9syn
KsqJfk14cXW9YtCHXztfzueEhZyYFSOP4B1EAKcczFuRBDm0lNSZl1Vz3dNwyZYw6E5GyH73W8dz
oyZnJIkwQNNTQ4f+ir5RaD505w6V8LmSZ8L0tfmj/2E3cIWB8239K07lmlsGDyqDLeMocrPJE/2y
JMd6YEyPX2Kkl/Y6tOVNw3oLmvGirmSWKJas3bag2VwWsYA+rLyI5WGaCDHYXdq2JUH4BTGW2nRi
6Jy5zYJNgPgsy8Xk0mEEDToei+WCXU5X2bC6zPbadLgZj7rBQFBSO2ZQQmTDeXjZUzYdU4MeZAU9
9nuDnPsxuudarwFY2GysTR65bSsAPedcxkFx1+ZfvAA1Ak9CjxZ029ltdzziotD0xoC2tU9JifUI
syjK9YnrpLxy/t9Dvkzm/5j32XC9imWcIYcXh3X/fBOBIG1m0zwSRdtmgT76lMKxuZnZ1xTX32gJ
xSAQQTbseF+jRv/l3Q9sjCet5ljpJWwl5l/Pf9ErrtiHY5TRhb59kFyYczSgO9lKovq/uAdLwvKM
Hq+OFxMzcKWa8FLWbdGY7ZM63fVNAr2y8rv19wQJYfzMQ/sEeGDrazqLE2bm05KtHoKWoCULtMzp
i+G0A+7Dnn1xU9wcmpW5iZwjOZGRhGQtwv2buTp6mTTJNvp/3QK1JChSfpaupfTyEvHmSIUKSMgP
XQJZtgqI5zMYvc+PnJmTgdWiWMzUnZeJJ0MFCwsiR28ArU2kIGsh0Ji8TxoACHpMSMLfS2lfVN5X
HW9XNUB4qs/xaCRs5TRhcQRYji9/lui6nQwdrFnzz4vtinESdjoM9sGAy23TSUcnVNg1VBaW1Tdf
tpdRZwGcaaVnPt+CnS0noeZlOBNV1cuu1yS7AM46Qasd1Jh2oSfDe7oYCmqvTxV6EZSFl2ULtlnc
gRVskBR+suJZX/UMi9KLcsUdJg6AMn/H6CDVC1A9B7cofnjZWKdRzX/8xacmbzCDM9sBkp0bbgvP
I3iPk4IC7aLz2U9mdSsEct+ZCcUhSCwUPpHDOZc6jssgi7q2UltVOvpgcZxzlbq5vMthtZg4EEvy
CwcaMcAjQr6s//i0RGCWDwakg5kD7xE/2glzpGaNgyMTj7CFvN6qCRlbsKIY3PrmYcAncYtgJo+R
Uucj1JZqtfZ4hSUbSTjH/xTrC6vsI7EBClTa0b+XSMxrGoKoN3Tzg5zT0cA/vWiPfcEIGIEPN3S/
yFQDKuRHyRtOskkVmyuKw6y7KHo+CsjQ9QaxZYUxTrImxtgrRoA8Ex0dRx//k+Hb9XwB5STWnjAg
2x2r91uJ5B4KaMV/vGyrMH4S62F/yVzh7LW1enrZLnjRBbz4iqcSyLAMHWFmP/I2G1/BhkGERnOB
SbTASmCvfrvFjlCrVyKFARxd0aqnOVtCrpwY7lvJydLPqmkp3d1YuKUL08MGo9Cp4huU0bSKfRzE
w0xqMLQBOsEZ3tPGNsJ1tRPRXkAlH0xnkl4YBOvdWckXJ44GLdm93YRVan4WavAtwKybQDZSTYSJ
fht4wjvW+zrTmAk83lO3Jp6uU2E6CA67FsIyvnuEZg6+fjNzaMAi2vkr9HkireFc48xMG4ak88rZ
GAUdWPPRV1dMEno/tYYo4eXp58rnwuybtE5tOHRes2aq2iLzYpQ4+G+1siLEsIc/pT/qYGZ39vja
Fw29YOayqdj5jauWZhv/u7Pr3xI/5KuydJYlWuDZRoflRlkaXkCQG9KYjht0b7XpRV02TmwoA7fr
1aniP81DCmD2hNCM56ZcirBghtyQHCEpD51ZxvxFUF8KBMRQVrQ3phoc1qP3+btboNWE2Ta5XyF8
wDSDWpfUfhwhl4+PQ//ioURlsmpbdGjqvOCt2SXd9PFO/D5KVtQ8QO06GmKu6poE4cdsUny2ZAUj
6VFxFwfSYacV5rEawCswBDFllA+c176a0xrXCdEqAUD+hyOuI2B0kaFMeJqkj6Q2EuMWnfyhOX1o
KefV3wY4eXZTPzEEziloM8SmwE37dtJqZR+aZUB3b+w0OAE/JauNvKI9PaQGZlID9Ubz4/LYtbE9
H0LodDO0GmVXAqrjzIVZOvVN11YXnvT1WLmBYetr/eSW97a4kWa4bGfh/ya3frjtIvoa6ESARcxQ
4rAk1PKtPdsBlmXP7YWnXV2pf3qTDNMc/BG47QGyMdT8v5DBb0mtxkeMm2orj98K+AeJXYDXGB3Q
QcrfAWnAnPQGXqTy8TFRZkvwfgOKqTW4HLHm3AGm3NAo7FHVg18+givnqd6X+p0Bu0PaQlwi4lPG
SK5fh5/jhpCk6hhACGwUFJwIdHuh3nF0RBN+76X16gqVcpN6ydi1ZcQfyHggGPyJnUz0atGOvL7d
NT9Wf2I4/fm6l04D3V37XTRscX/ixVLynClLk6eVrGNRAjUFl5d1KjENLNYOgSHiuA2siXjj8mGh
M/sBFNfb5RdJYGHPj7s/2fXhuy2+70XmrHzXjYgsZu6sTkl5JYa1CsbE79+I11PcQVf6e8Z4gkHC
qmWQNs0R9j1yU8UbdUgZVBn7z6puu8IxoDj2GFbPmGIMzqqwIZLnJ+CLlYfkCcqx10r6duo1UAGp
3ch+tgVorIG+WYn7H/T2+KmT3HcYRUBuBhoRPEOvwoALSyBvCXWerfRkH1R4uS2PsGpG1HunP/hG
Ehj+ylEYZcQI6CT/T7/siUcX1UAnnUMkpNWGPG+h9MkmipT8pSw92p4VDAIfYQu9ooSrKvwy76Jo
781E79UCMXPyhu8uIWepPpNERAKwqJdElRb1sIS6PuvErSdG7qymYOblAxC/4TTVZB4uu+0DpAJR
Gy2vcEGZqM5+jbSp5gbwDAtXuUqRCMlTMWNbxjVMDge1UNDj5lIg7WwaJWnt82ZT7A0S5BYzltO3
ALq1S01ZXsUhCy58Le4S68mjr3YeWYW9HjgR7xzuPWAevRrlShOtYUA1tJPSLGSLWbzHd5/o4bl4
lAOOXW4SBKoT9H4feuM1wTtAtEdz1PE9shimZS53Hxc1enJSDMUch3zvYCxJqzu19jLhKQmAE7mk
hKiyaeQIlIlU3Y+OW0JutHdwxSLgcXJKlgpvtChQyBo/jwj/e5MqMTT+dY0x3sQ+MbxR0Ku3mzy1
4zFe0xbHEyeWjYoa7a+fMTx0vCew4ntxX3cvPrEEkqHZdo5wFLC8H3Bhu0jS5pPpo/7VUhxd+Ltw
0w2+vyMPz8ifZb2taBqOa0eWCt9N6px8yeuwrV1GMua+ME3JhLRLbLcx2ORhDkxV61UpysnH8Jg2
YyLYLu7/LWt5n+C10JK28E2FDKCTlMHe147l8JCoWyZa9UQtkOKHW9hVyhHJze2ZjQa9/sBWF7YI
zz1Oh6tedA+lKYqmNgIpi0xIVYSYrgQjYNpaKsO7ZtUVE531S+RZ7U+UH3jT5CXkjYTF1HpLcyp6
irUXVp2Fv/4Ruf33Udn+FaVOMFKnVdC2Iut27Gxu/qqSSKEyPaLyAtir/6JjVQ5R3YJo5J/7d5R6
NP5ZlsC9cpy1UXgIiKDkifaQMmS7BJzg/LXYfjVJUrfCf6UAPugcG6PI1HmN/1iQUUgoWxlZN+03
UxYOgFjFrQSCeaiqLlq1qPQoNresXSWMWyfXUnSG6YSbmBrVwqewXwLiiXXbsuoczj6XF7KasErq
8/u1FHxiwFKpe8Ep5Hli2fBdSbQZEfTyP7ZrHS5SjAlXxz93cxVe5FbR98O5Q17iBZ/749ry5Ay2
dLEE6c5p+rl6KjbStClsqyK9snrQOg2oz7SqQ2n768Ed3UvdUggGb7wLU+9BzRSR5pJeC0BpfksQ
Tp4HFEGy83t+F2wD/F3X1lxMrsyaO2Mplk6eUMrcQurk034y144Mj4bkTeLWnOC9sa7EU9Gc1CeW
UGdEFbn75et7B72Wss97cy/q9tHHwIrXxZjULrVenMqbW7BlfrvADjwjVc0qmsWpyxUB+vx9y0YD
Zb41piYcg09qQsLrHCnEEo+0bKnBn4ZjDbJtkcIpKI/qqGowpcrgz7F3E48VNcf9Yz/BIUs9Vtrz
dLnF69O9IP9xsffD/ExNyBpX6Ik3uSmc+4WgKYKMJ9+RYp3OdvOeMucSNRhHHcmFdwVYI+tXylS7
ttfbiF2NG9LpiwIsI+l461Qt7gtO+Fu91oc27FDARxPDZJVBXBqNSSFKJYyA6jqb85JuN3cU/rSb
Q+pKWQJhGNRhvs1/QHizhWX/UzGh6cXcIigHWQf4OGinmp7Za04lRA3Mke3ygop00rTP5nucKGGo
bvbS6P/4HH1CgyRhJ3loQfehjENfY3MKeH4795V56giGifImOh6soo6kzDRohnTrOhs94ENh/10a
9VLS1ICsk3se+NsqPmqJ//vXXNLqGoMl0ZrknNb7NAzZiBrl2UVbZSj9HFZhN/s6gr0zqcpy20QA
Cvy+IKw/Rkb5bO7mBl0knPUYONNoT/RwoeNTUWJs3Upe3SMQaNBf8m/SdqsftztH8pzfRXruMviv
zEgs113eDys53Eb00klB7PhTZzwGhE7p9SpCJD+YebfHT53uS7mTDtreeA47g3Nm2Y/5/RWPZCvs
JOtH8R4C6jJ6Ie+jUToIlxwv6vDu609+G9j7ISFymtnP5E+utN4JgN29FcgrpFIUZ0NuDhR/N+8H
8VZXpXRJJkjWaRcSf++ahoef0CepBZhSo2HizCmPKtsYVsGO7u/X09D4Y+yJTcYeHK78TtrB/OtZ
RMBKIQlRwcjGJHREqGxwT0XK5eLemsfdIY8Z6uouFFgma42Veuycw2GjR+qLRTcydZlVjta6katN
55gu/FQFHTYPq6DpVzH+PmB6ZDY2EU3MkRe5n4gCsApSHTwdztGHW9TdtY/wOlVkTOSQr+DIj9ZO
ccbvErx8v5ljN6D7KAypvDCir5ywiA52KAStoRV6SosolIIYrtZofiDWK708+w964kh7Tep8pVIh
U3vOOyfZ09JppM5737o6iUDVW0q6fXkf6nObslKn9bKKdtewYq1hpj/AfQEIaxVTBsO5cqb8bZ5i
Zn3BVEBwu8rAuLfqVLTcEl3UmflZFrlhiB7Wq4lkytwQJF70q02biH276gXesloUdRaOV9fWGmC3
TdKTp10kL6QFYc0imvsONPAmnRoyEmYKU+BuhKJTSL+bFhMuBwt0kti6Dho7dkxDh7vhBFas26mG
NNH3HhDgxJm+pVvT6bU0FA2yh14PUaaoKVK/EKYV8de0YC0HpTeIdnYjJDB2qXk9/uO4V9z8lNgM
x8+aK7JeqCoLDmigzGrMqcZQ+cFYO5KQ9piP+5NObLTSIKtjX1HkfTzq6EZgC3s0C90MBoaQ3yUk
UCTzPbRyPlOHppuKt7lu3Z3PR0MT9dYwdjy3/9AHehp4GSTWcIroa1RU3YhH03CBvN8dOBgPqKOD
AbC6OMcvwkcF3JyEJ1l/yTz/UwjHZw7T0G3eRuKu597gTuWoNvFNlV+W0DFlSdOA3FHm5RYzgwVr
S9Z8yF9GEk/8y9+FYswvKD/sorSy55UHzjcW3jY5XEebNX3xlL9DU2iTEmAvtaEJHpLX0JllJR/R
DjHSZWhCASQj3gIDc4Iaj6bXI4UVoH9FEpZTIBjBIV0O2Wr1g8FZWOQA1YSh0hLqdMrssKhmiMLH
rW0W5Txy4qI3BEwdGhuPpmdeIOXN3AEuNKRxmyf6Ck+xfqbOIGnMy41qjWsLvZBr1vmxIn3+ndE/
V16D6SurovsMQP/2VmcFdbO1d/ErrdQJ9RRi5WSbNlgx5HuQW90wjF8PmvXPkNG5ahy4Lx5OsvZ6
GcFCkX4uUbuTHeU/kFK7kgXm43/EWSoiZv7QSuvlceK/GlD/Z7t8ni075kxAhUBy00p3wAeNtuth
Rhy6Kp4lChT+pN/lMlGwLbqq0lmmr1h7l/i3wGS56+TS5lmHpN2zgaw63vHbf4F+vri0/e8SbwxJ
sJf1ORq8Q5gGlU+++T+u2K+C4ele2XKG1Dt5taVkF0UCHdp5WgXg5WvOSmcVNZjVhOlkkXC1SPmr
uytdWx+RRyExWl+AgZ7FrYyDP8Xti8vhFJcKZvOhLQ52FREulLYQVtnqt1apmwW2LkdNiGA44hin
KYrx+eJvjLpz0dh4C7LVqA2EKMclStLuvWiAFUghO3dgiLh1pVAmX8+wb57yLocTmDoVY0FLRwcZ
J6DjsrV4BdvRgHklMOFUHlFZVvu8HO5xqM3B+6lh6W/8dHSMgFgrynL6mv477WaCX9vEFCVi1UcH
qflnCvd0ezc7lJoB3UAQi1dZhBhGdH4G8qc2d69gZxPhl3RDLuOC3RXFoYr5TjVhhi5tNkznI8YJ
CHQ2Pf4x3JBHxwL3oAXmPa9pjY6h/qpr01rAiXydUhPpUzqfythg2IJbruKEmRLgjcI9+LYcxEi9
nIlYq7bFlreOA/bDsXc3xd8h1pLRnDo1JTbjLQA7r4C7K08KIbQNyCRj0eY+J1EmS/LdvUTUYHuz
Bitx9QH3SWBDmvJlCaf5KwDrGc4ic5oqD4r5rZzxSUU4ZqR3J1kxm3vtWkzMDBytw7/TubAiUHag
xVMS5tAgVFgKW8iAOa9StNMEZRS+zAyGvMYdtKakfdDZuLxqVTSGAzSfye80Cy0BfCW7Ok8vr5h5
UuV+ahsKHO9H6aN1WYwI/WWzfMoBafKg+Hjelz/0K2zxXJAQyWuR391WVC9Bgk8nX7eS5fLiGgGh
USM9rET0QPG73/l7HcJQdDfQdoDhuDVWIk3A7HAUdxLmBXjdC3UXhbHAa8fm3Z9PmXPs6EYZPaKq
HdbB/ox/15lxLcQFcoT3z75E8syXOT7lW9AXrn/HodtCfjoprCtF8b8RgEmxfqSSkpKGrwFS+dqh
ihwORVo2djmJcoHbg5oFcQxenjiTco+L3QvqYxh8PV3y9AeXTtgs+ZSGnJ449Sfi+mF+bI8IwbVK
zbclgTfvJdGr+I5L5tw4rBybU2Tfy+BQ+MgG+6AEKMj1j9iWcqbYymqi7GEPunSYc1lR95pISo+f
+QZTJJgVQ01dUA979wozBy1rJVp8XId7k0rpkUDXSvi+s37r52mZHU1WKf60HdykjvY29jBmAoFv
pP+0+5rgJVWkEWMM6ezodFmjw4TxbrgwBcLXpgxhhqxgDFGnMlrMX9VvYa2HgJY4g+mnl0NhLJlb
rAvO8Y8SAnCVY5Essxopueg4a/RMUSqMTjPToZGtWeT9uABE5TbDYqPD+0MRibu858ma+pKavRRv
20PKIA7kdDuQtpyPmF5BOXdGDIXYwu6+uiLDV8kseyTV5DZ3Ewu/1NQbJVB5M6VHzfu0HOF1MWtf
Rv3qhwmOlUrBxdiMySeVHIG25Smu9nYggdzznTceHNXo3j6bMZ416VSLwy2eiQSWyfGW4ovaJ/Bj
O9tG/ctwBEIf/W8OVnE/sR03XVWr6FEfA7nS4RFIzXpQI+MWG/H6kMta2KEAVq2Tf1jE0pOn7Ejg
V9ZzZsMp1fjN42lJSZEGw30yPwNUkUlGOxpKY7me+K8HPeOJpJgwbyZGCkD1pi8A3sHYy559553c
slCV33ZB4zRCUkifE+SkbcLQeeqrMP3aCjcA/lxbFMO/7AIUT4DkyjkLvhYNY/uCgHnUnlMATior
scztZJX3bF+6KGrYKYkfPuIGYYPVjKOtZKhDu/eBdUE/EPk1BSuFirKLp1ILB7lYpW0LjZqv+ilZ
7qbM67VRas/YJPzTOenjtLQYXJIEz4OUhyeE26RuZrdDOGaYZs9R4c2D1LSLwF7cTL0BEjBva/pp
Jh9vlT5vZZyJ5XdtlxRdO3zfZijQYLtPiN1grJptPf2gZFUzS780aqLk/E3YjBHlpgNHZGvLhyZn
z64xgMG9MkIufhw1BcLKX4rp8Jhw39eUWPyKazIivzVobvPR0rqX4cZkU966MAtMAEh3OiyN1sig
SJ2PYCib/dl+YFeRBqzDPkrVXdyayK+LuxIVlVQtIF+qDyxg7KPzVt96DQxoyNONTXuYjsmfbSRX
UVUauN0JZ0dntfKgO86BtR5bjeC4qrqkDL9dCRuBzU5B8Z3g7jsPwQNJPcDVUyyo+XC2b+TFlhR+
x12cKZoQD0jd34a0SML7UdDANZTEyuJ7qG8kxJiL1un5kEdPFa2Wcs1emjwBUGClsFTiuVmM2HjO
plC5v6FPi32OGqrPfrb61SaLqXi/OUXQf707DSTNeAPNgMq0/T8dpVK/eaXc4KsPSS3IyMNcihq5
92/FEE3HdxqEw2jrCSPZBeVltziePOvzp4U4BnTE5OiN2TYuzrGDDEvFBbc+WgBgNWpOLelQQIY6
VS71psqdmtNIEyShNq6KW+Rq4VqnlJOZ96jC8/OSO8XVpMS2Wf8IaLoQ6uNrS6sZATbrxo3dQqI9
YSbnrVDPmuUWWgjdvOzLoDSDvzF56QCvUfphAndtaSPl0QW5Owdyz0NU19YlyvI+ax4QSd37Iukx
gZdz06C67ok5SqrV7o/DXN982p/Lvf3iNxge9wMzs7UqwkHOFlkR5hgJJS1gtxKis0EJE7P4ihUL
nrxtOv6IF5CSMe+Q5CpNrFe0nbKvdnSN/mATMikU2xFMCMPZ4L43pWDEkdD5aEIn8weui0UxdBNV
P1Nsd7A2z/oDIbmCfcQqIX7MaAhluoR1T8121Uy86NxfFn5B5298zf8Ygwg5eOz7hPB+pAKh8tVt
JpDtay1O+RazT24uDO0DFGRgg3am25RZ7jEWioLRl+OiaFOXH1oSXsceFZ6nejCKJ3uqB/6vfIUf
80rn+Cew/DuU/vHNXAv3DnjnZG4L3zrr2FTBWttExnAw3rUQE6M1vnPd28nSKvHKZW6sMgMfN+e3
96rsr1KU0M7yegknqCS+TFWV0hNfumlNa3hdaQiRpjTK2fEmmqOFeHggH6GdRuJi0s+709QPLta4
qPKgzo8axBB5KqP+ElRQYpiqtqz0ZT7gO1XKzA/nqCAyW7L0MpEcj/fgE46UDmlde9JHx9OwbZHJ
6jo48DgHDtkhYrk/Hew1ibUu2U8GHmOLETB6Y/lwl3Ww3lApWitdekreOvGZ6Q4RTXwYAvKY6WEJ
eq4vWxUVf9LNM0L6ZTzfQCLEWTUaeIVLQr/sP3gJzoI3+oZ+gA3nTKobLKQ8VlX8/rqvgKDA07oQ
S9knqhlaF2n88DDoTI3lxh3T3de/Dec1o5H9O0Wg/wNQtOhRKA3R95SZlCumMV5KkY7FqnhN6YX6
h9iGeXxpAzsNes6CckxkCdV0CMknbWnkxzAPgVbdg96wos+Km2jLT1ri3KATttpaQoN7gQ6NloyA
jzT+W2n+qUcl2KLxJLPLd1HzOJQ7ViPUn5fA12bCgVT4LhqyZbFRltrcJ6PzJeM0GBl0bmudX3B7
QBaGCG2fdJByg8hugOZSUTjUPW4i25qfg66SPBV3DQ2ck4zBDGzXIbs1I4Ehwffy5lcDC2XvpIVW
XgCZI21idOUexxkzqA/qz5FPEz0kw5VrWFefCGlEreM/V2Etqd/C08/UWZNWOSn0dbkvVONoqmi2
cfjoXkesHUUl1hr2ArnWXWg+AS90xbqP1lcFHYvpJjMY5KOoaVNZQOBiUcMeQ072RhJaZL86THrC
tpvguB8s+lJS8MtEm8S8F5+uP/oHUDY0p0CvamTNyP+wxzh0OdA/AM3fMyOgkIyKF2cEfdFM+S+M
3CduEWs8iWg2YE6lFb0IzvK6Za8jmzmY1XPqNa9XSZhuOlA3HkvP+zWiH6eg7oAMsUsZLXOvVqlw
slzQ9YiRaNSQi9RGJoeakVcLjSA1x5fU1FwE8AJVnFvHGVNyc/AJ5mkq9Xms9hRC5EYQ4dU/DO85
ss0mtOamEq27NWckUdUvZfHOgmV5W++7OyyetGnmt6nY6KfGHex6Yz5AYbmcKEaUFoX2H//pvckj
aGqyFIv0uCUsWMQPrwjcnPKtPz0ft/V1AfSvjPNBn0mbx+MudS8XjTK2W5lCyfrzc+d5kBYkccks
OoylpykGYJbrArdLWMBCiT32wGpOgKqVI0xznxkXpwBYnY1e7cGQQ0664ScQHIkNreW6A067na1q
5/mxlC8gBI19/QVmq0hpbQS/vmW/YOPPlNqj5G3V8A5weMDC08hIJ92O3IwMmbBiDS9An3HG8qY7
1NWqLrxFLPvbDaF+Ou46HtAw9IivHoeoxMNaM3b7cbCV3rkXuV2QRO5Wivy9ppV6oZ5y8HvgzKkd
VkQeWMAq7uGpMR8d5WqvvAsFHXa2mhz3bdZl5RYg6vLKQNUSN7AAzEnV86zupMTXlcQuLQJnLSRe
mLg2tt4/fZ6kBiUUyeFLPB3fKMjxfoiDUjxFekTBhTHYKvH4AWNlGx4d95AkbnkCYfrIcYgfJEZ+
werzDDI0tpxIzjTQdMyXjD+jXOZysPtjMNXsqOG9eOshV79lvmNpxaXYr3q0Tp2+WQqWPJh6pVul
8IRCnJVYv7SDk5eeBNQoGrAmuKcvTXeD76B/qshxlmGncZaDsx0XW8MzaZqP9PE7WZL2qXvMO5h1
ByrNo4pwBLio1v/j3QxYpZI++TodMZX0MlF8vPooPxQgvAW/fI2wd730wwN6oCkbkSYdtmHQMMjD
HzGU/SWnRcAalPMDP+4S9kBL9nf6VeO9JOel5eGfC/m1mml2hTMHHFXeH5ZqJFh6X4OewRe1TJa0
2oLeDX3UPzPpUpqu1js2Xh3VmyT8/79shxnunuqQj5KfL+tuZ1s7+p97Zg/Ij66ePQFtyPVrVG1J
L5I8ayZ1YyBdUidFYdv7uZqlFcGKJ5aGuNoXHa0jdQwKStoGjAORzcMHxn+Awgt20788kzJia/8S
Qyhnaq2MiG7QnyluC30NuRfyvmKXn5O747TDfxjww+bubN7jq/9OWTNsD9uzNzhEySvJoGxTM41I
ikjzbrV9QYoImgrmNrnKsPARmmAQ/vpCjdsuykjfEffdurySDsKfAyYEO4ihzzylEtHXQdNL9/pA
SklxIElH3tWhy/E+U7AbXb2sS4+tAAH16Q1PDUFRdN5Q1gMMJW98fSpJE6PgT2Q1Up/+voYV1Wg9
8xmbdPWZ7a44T23QZhwj5mraW7LqvriTv92g96jntMeIDqkPDEc5fwEcnSolxUeN1KbSq3P521N2
QlSU5paPT6ekZpCOW4Lr5et/nw3U6Yyr4vp/QqY3fJnUUrlBvdnqYczjEKxFULvdEuXW5P31zn1B
fSqryO0zm8xxQj443ewis0sxKbDBs4UBm5VEzYnprVDI51fz7EN5VZxJlJofvq7sctkrKa+ytg1h
/8pkI/O+HT0OJIHF5ue1PUU2G7L2bRfv6rb7/8qTCJOpci1KxDCLSSqGAJAXNtweN2YLZ6OQfm3b
1G1ITlWfce577ps9DtKcs5N7kLvrl2nyNmNdsofMwEztfo3jVEcSl9uCEkY0ATzG4HFyEwT+l7Xv
MxL+mPQl2/ewqNilf5gw6ejWVJPg3VRLfJoc5oGKYChsf1+4FlwQfP2rXswQBV2uxqJXZXFZQ9jd
PYUhURMAsmonE9dlFKp5hkixYyqb5uhNUzm4+lDLRT22UgFBoWgSZv3c1ZjUfRHaJtVDU5d6fquZ
RI4AmesDkDFblt6fGpQwziR0wvJQu47wOfQ0FZmUvgEw1H8ZcEXxIp6fy/ouqXLkpcr/GXFsV5L/
uKuH9xWmOOmL3adrYKtKnEDA/jVoUQWTUYdgubzkPgzrtOc09zBzFTEp9sAfaKbhJ36K1haOglf2
Q4B2olvgQQaT5Wdm2HgBtInWftZY9NRcovjtxmrnyovDpySh0ZRAcqP34NqPS83AItA0mDK+tFz6
FyKpDwI4UaLiTNK8prH8zLIPdiAhLy/022nP/p8HIjhX+stA/Glkxrl+x1UpTrmw1+4XZviSYCZE
1B9gq0mgVY86CNH+n7npoPuAs+FFfI0Z6reMJkD14L+I9XGFW05TwBSuL2wG0t5n25Ouuc3V1jED
yzFzlIn4puYhRALwf3sm2B3Zeb1mEZX1n1oODuXP/o0aTNFsiH3lKU6VrAqHZCmxWFiDHWQ5FsNU
0P/OlpzNBMpSzUNpdnzdlJv6Pk1COqRnaveYOz4eBZxSvUKngi8AT47Qm/6yFginGFYMPSyw3FEr
qijL5aPSy7SqQmCSmXifALtavmXl+cqTVdsT8LXApFtfildn+wrmRarOjBJrch9DTuqecVQDvPya
e8w35nb0pTcVE9EVNMZoSfw+n+wHlovIGl4AXAAQPbNJ32lA9tKdcs3ZEYxjmlFyxXToAn3qejuL
Te/j4hQHm4p4fqCzRgoWljS73BGKlh/t8DgMMWx3OjeyAMAyhEzNnh4k8/MPlocKgLpTxzCgKJ0f
iNN6SeT25yEx9KE9Z5fsocOj+rqG9BCTanFatQldbLYfWvmAnETl6Noi7Rsc0lf/GLUvx7dc5CLv
qwLCTbedxkZ5gT1zlelMdDu4/lXPc2fuWPPEDmbZvbtYA2ywwQ9zjjfBiIn7xcPhOcK2fOgNDjVN
WIOEIPNSd6VjOu7m/HOTv5f7xTh50Ioo1cs2OU0xD9RSURtQIx3McTt8Phmvm0YjPxQ3baKtrREW
gkYKW4tPexXV9GJ4fPaWvkUUM8QpkG/FxnlB1VRjoH2DDEhzV/t+/TQzIh/D99hG1pfc4AXKIwV9
WmM1GHY1bozJN4ByltJP2833/OjtgCNboVR6cfD2ZLTiwb0nA3MdhTLiuLyoG96l7+3wz5LQGlUR
NWvH7iVaqMk50rmlaMbjHZiH/u+MnZVPong9eIWWGdff2BFBEVWER6ihckTReDB5Vy9A1WIVn009
m7b3nL3uXpn97tBrMm+SvwP4Qof813sjje/TKuNe8FIESjCeOWSYcfnYtwjaRZIiHE8UZNRL+4js
gMWlV8JtaFpqh0S8c3Og0JLsQNvOVTcSEx07sYzj8XT9Ebm6e+K44RRa3Ey47/DEjHtk+tCAzLn3
xNqqnkDKdTUiiLRRtu5oj+NpqtXCUG/ve4F0L5SBflKUUO6BIfmPJZrZMZzNTJxzSBeGMo7MfbUX
mVjgJf5fAljLU3HmScQ0IVGcJguh97vJSYmP2RbvF+AlZXZyiIUmXV0wp5ndIHs3s1DaZqiM0+Tk
hZzaTbk2BmFMQ2JuPKSPauUmcReI2f1kb3DvPwwyCpvaW06iA03dKEQfSjh6QpXYpI+LF6AkU2Bs
s9BOqaaNHEvdE2HNs5q//t39F+f/SJelxlwqgjhx62CO5WoCRDzQ9vL9/mxSrSx5j2AgC/QLdnLv
fSTS6M8bep2vGRkqjJiNkDQyXPHGK8faxkbpPuNhHreb9clLGxjAx+RkRB662XAcH3zEplJZ4cW4
GLkckBWMMYuUTDjcr3JmaIBqxh+fcuGyUAWw9Nlyawv4ZtaKwbN5jbcH2cr1ZqZPFOpMY+4QafQ+
+61m8JCUBstImiI6i4l1OpksgWvObnMxVgh7PgkS+04M3LysvCS/rXJ5stw8Dyk1azFQ0gSAstjz
Gzj7ywwaGarY/Q/1YD7Q24xeYpRhvS7pB7SEu4KU33rXCw2cBGyJghY15IBFFNbUV+3ZH8SWlGFi
pqcjSBXIf8Gttjbc8nmZcUTxmN/eOxGWecCGzmbfLkHyl6Y0KIYS1XOAMEw5db7kz6wMaq1u+vJ9
Mf0pYthAhsAvuy/4ADiYYxacqbKnXtVih1BNVC6FNc8O80dTrZRpzwhlOm7OiQeobNDLJqV0d6b0
r5KL4jj2DO9e2pSNwbwep5IpmzRY4yaLUOoJtskvh/FVYrz31UzmDHeXLJN5zKQ0MA+kZf+bBkgw
IqpBk2z/6PnoRSlyOJBYNGvSA4Q25D1Kbl45vE98vDetVhOlkGO2YJer6xTMocWA9XsPXRWfTXA8
pB3NXDJpQkhqCnyWVPhUWw6L1OpYC76f+dnS7lEORAhN17qfqPcARRTemk9r2r7qlV4BxkYrDbn7
EzZJhp4OGCtsMoNqOcoOtS69chXuCFeJNLBmRxN+M7FyCWgF21S0sF5XdUi20uZT/FFS0mnOjISD
YHemeVBeXQhp8+RAuaapYA4bdawkyos3LuYnNimRKlSGFMWJMsQpphnOzQKu9GeTBuWURAT+3zdz
LzqF9F1ZyjpIgZRRLSRvUtZpb6u2oLuSkK/HILskHqMEb/Lhc8LeeXk5qTpxv8LOEILl1wsckT7Q
lsZ9cfqQg5uKCSITFQWkIoktdivbv90ZgUgCjk/+aSqt1eXY1BOZPXjN/f6a/MRAJfGNOP63Jahy
oOskA1DHhwEICu+JbCtKliNCbkMDbo/cHNC5+bvftqBZzq9Ks47Vp7ud2wq5R2DA+7eal/Ui/dyX
jqqd7fFoSkNYBMl6ndLDX0XZ3LHdKFXKy91sFQw6XMat6T5F5MnPGGU7boU6vdwji31YtXMaPQ9L
RYoh9oDUlhfmBlr09cNSy9T5AnoQRVyIWmG8PbTWytLg7aL+/7QXIXTXe5hBAvTcnca2OriJtjb+
ZOpuqRN5mKVYn3H5iN6wH+81vqRPp+78BLOkr2Wc29NgsaXcTR1wh/zJqUUjADkYRbq5S9h2u+gM
O6p9NI6G6BOE5EGtJDhnGAjYEivxkxqBUFczTkt+p3pnXQVj61xMlwWcb3Beel7Js9GcBCmtVBbe
TS6HMklqn1FYOwmbxzkGabEO+Op2Q9SiYttmOU+aa74VyrE40zCVZxQcI/UhRRXd7oodMGbQBj1o
WNFWVvCT/5gJi3dYYQpSE3MP6mWCrNcszsVwSQEACREYpKKBwCpkz6ohm2Y8aD+mVIRKe7W9BrEe
7Tkk2TAQQnJmAvecRnOCXlWZb4O5LsOCD5ilwkngfpf5cLhivHDluJ/A7rrVcyu151+OiRlge5Or
IJdk64TQYOR75BMMY8wF+mXMXPf7fRaolYse15gb5pDdteeRnYX0hr/Vu5oLSSybPMul22n1hHM9
NQuLPxE0hi/FgfNSbezHrXdgpbOBJQC86z+1073OuCWELM56i2mHS9rGFadmguy9X2ItThrVRLuo
1eixe9echmFX7C10wIloaHpSZHtLVgNE+BgehWVRcszBWRUhzEBvEP7Ccy2seemkSPqz6Ce/lxkT
rAL39r6i9hJf8XKXR0bq25w9iqU80tF0jbUIrped/oHGWGkh32a1tEzU2QzpXZDUkuKvKnU29sM2
gv3qxzCXs8ID+PQ6nYPPQuVO5CjxVL6+ytsxTAJKd1uyR2OQGzl0mL92HYTc/n6ZVnkLgq0ZcJPG
A2bRyGToNEwKwEeGTZI0EHqTfiKJmMk40ZJr/MG8EbgsliOQlGaheHcJbhHOkCskJ0M8ETF7+eAM
xJnG5DJ02oxPm9IgDbdvziADHLbnUEzgDw/m/MOm9O0V8O50769+7HcMEF21fpmGeMgMVJEZj+bV
/+VAWJM2ljJqnRMdHpjFMOXHngwt1k1XQQ95TnpDG5vbkuAig8ByiCWZthUO3PzuLBQOV/p5qFiy
vKDvLL2WWMy5rxC5+9YQDmwtuanzojoX1OaigQLTVAWUcoaIn00dc4q9uIOrinTlxwiKIGhnluua
Zgvg2mTgmSFIE+BSCED7TDiA8NWYbhopmuKYVaJHEGASrs5TPqe3yuCHK3k34vlGIfFzUw+mD1BX
oxPfjvPM3SBUeECUqQQPibfxKsdXcO6hZpzHIQK1M3NYYycoyAhGWWpQOVVSZjtvDlbnAcwW51CC
yPeB7TXhWjBb1fWhRm4eCXS1fVLdMGsj5je5j44QrakCTOgsVwYmAzQK0JFkJ89GdiLIgXqiXEG8
HX4cExO+8x5J6TWcC41ggEU/AFHVbnqHBnEkasWvHdbdTPQ+xwVEo9MPBoCRHhq8yIL9voi9zAu4
39x1EKOIIpVMGSdr3W83EOHpX06C85fYCIme3H/UxA07Mh7HnggTYl4qilEJc2xJJkssyCxdR1FE
eKv8ut6ItSgKqWHAVhK4cPZs5/wo6PtLeLGHI/Bv5kbwGfJiPeSQCPj5UPKSAl2coIdGwunUTcXU
Zxn5/iX4piQT2DluPXFofmu1P3cbdHzB4ZlZPqrJ6kdphcutUd+KHXBoWQEJS+025bgdvdUPMAb3
COOwYYY+uIHLTNZYPGczG1GESxwaa53p86rClbgMBiLEXC6/zYfdWphJoYG9h6xu5H1GdTRMMnRa
brJi357LWUiFR31pTcwSniuUKOSAC7/VdwQLN8NvsGLp0FAj6/dm4daO2eDE/TJoXKOPxb0O4bOE
TcfVBjYoRI71qjQryHq5kLokjzSkoEHSB4YjDscW/lNpb38/Cdhm7btavsGtKlT2SIl3J7TvEt5y
u3THoqTzJtcyJmsdgF+M2Pl09OuqrPCwhrfrrs9YPEpWDZGHcQu8A6eBAzdL109zd+ulmsdivb2n
f/U5qTAtywMVt+822X8R+/MW6ffs65U8TsgR0WalYYh2pbrWWu2U4ZwDoLHB+u2x4K7mPdhuv4nP
lUnWayCaRcePgFzOfnM9xKBzJpOUqCiypX52Wd6xbJNxUd/A59bub5yZrwjU5jhf4DHuJTFC6BgY
nf2n4FmaoVbyNxmT3iyXT7vEP0/hSivic+eIcK+eHEDHUSRJxqMC8OUk7CATTNlZGC74DC8BUV42
JWjBrwIAqXVrWcF1JV9jskrzrYesLG6Gkqd49EncxRPR1hkhxuX+lzSoeHIMPKUmdryPuaHMaRL0
SO6nUUx13f8VDj7w7yHv62nkaEtLdMyx/H/JBF500YXUUHdF2l7MxTJ1Uxg83Niz9vW3t1k+GCfL
Krq340mOsl7j4WWAc1o1y6H3fW6rkO76TBteo0IAUepn20yfAV6jgtzQ2SB9j+HKhR5kezspQqD8
C6xpZXQH/GC+HdHuU+wNZFCAlaRHsUjN2hJT3taBDCAA98fXlHnl4nWi1pZlacewT9ZcErQfN2da
+d0t40Jd0AvfQoVA4BgAQS0Ri9UvgK/IapB+nWWkA8oSBSc4TrNt/gazRsW92GgmTSP/NkrPnO+I
LZcIif6YrGlqNjnyEcq7ZG9/c4rc+YbqmHnTXvQ+O10KWN8yBxxNG2ZJV3QOzp+9TxI6jMdwwBaE
1hnY2tUrOHPE2yQOZ6/PRptGk9RzswCpMCVOU0BiNxIybF5OXackvIjOSun8Eeouym+bLoZ33b5g
fqOYNbugBAg01AHd53yJcLBn0PC7CC8utZ//gj4hNt731qmWUavRO03RhcYfzaxrEcNj3fNOy6ex
a2i7TKFq8wTtfZOOT1AX7V1kkZPBp/l/3hYkLUdB9T/Qnf12LSWg1u0x42j7wst4/7tDVeH44l1v
d28mgBAWqTAx7oHpSRC3uhJfjp/fPeVmWXmcKMr6B0advpzNT8lBY54LJP/yjmmBTr5f9NB27S8C
uDhnZsXSTioQ6+Wf3d7sAh+oI3QFM0L/vr8ntaLof1VggSxm0eKaK5Gsn8XpKDkkcwtWGi2Qja6G
z57Numur3S50keeS0OkxmRKuWZowct4/phlIAu8X3eSuDa++p1KaMqlcsII/dCTL2G93tDpMDQmw
HR/8r3ZJ4uUi/s7kKRvq4UVu3GPcxXw78FvOj6oRhkeNRc7rfcR1/cjpNkR2fzN08/XuYB7RtcEl
bWDvuSDIXmD7zjqPcbnXk4OCnjIBbSRLXzWMUjcAP7XqsEtnGbc+NmmFvFkKoZuBwLyjbStW3ib9
jZg0+lJTQXX8C5WPVjtCrtwFCEzU/1poPQw06HnquWW2vzaj2vvexieAKLGsMvok1n3j3/JqbEsu
ntqfBQqm97EVNjvQgYBQfql0bajlm3kGctaRsmYQv/hQRuB4jRAHkaeqPVZzUsMUBVePk+wrrCFV
7Sr8ELmr0WSmhSeRVYwNwjN9/TkRJ2zkzi9KYedWNo0/UpjdX3Nwzt/Xp+sdebtY9Lr27xZ8tO96
JICNa99v/Z1brjblhxUHbpkQcD5GaGURXgSb3ntj88NtMBb8Nysyj91pHsXE690OjhKQ55HvYb72
O/rurPjNt3r5wuUUOIhB5LFuxOgGCxJJTIG/Q8zZYw0m6s7t63ZUhH3A8MvZaOC4iYXtIb44cD5B
JYly6RSRf4iT4I+J/bWaK7KBUrK+qTt2edEPelNTTt5Pc/WtHv79PajbCMOhDO1Ol7WdEHzUva1w
QM6Qtj0vB0Uzv90sae5atwR7LbLuWJQNTn4Qv+3HEN7cRwM8eDspf5WQGlYBLOKaWlx4t9VAJG2t
QxpBbynRrMGdnK4+foFzRSEVO1/6X0JVXGyWdGY4oajosUN4XZ5k+8Spn/6tb7ZODYibtGLIkqnb
KrBYCkzq3c0GV9R9TNQE1BnfqXBOxYWDAYRnCxu0xeR2yDgN0A24c3i7YGTQAILReuos3089udba
h4qNnD6bbf0UpvuwYUd/YCYyCpvNFEJWRzR1JQxr21SqJuMPNNWV5e9nGmHCQJ9LZcnM9mqd/PBH
EuOCyQvmqYtzdhmj+mnjnNsEa/H9R8dExaeFW8Nsa5sVRdAcmAltnBNPIBwtothISw7JkkLa7lq1
4/0Z7PKeRtzOekGnU3c4vZkfBXuQHqRw8jR/wxw2fL+nU3XGV7Gj+2c+qiYNs9H6FlJOCdh3ekiL
K8/ByULe49sfteX+Vp5TMutc4fMmT1QiuKiMtSnU/rkFdcam+IbM41mC/KDSZUvhzYtbT0M6Hrmh
ACOEqwgfZt4arCCN4dKCnXGPUjZOnYLV6Yo05tbMvUTYptAJ+/XJ+iKjZb2ZnRb4v+Zx/rPl0ZyW
vNrq+r2qwEKWwryZdMu3Jhg6C9uSlsYeF0XsB30NErba5uOWyYZi3D4CSRHxAa1D0F5F8qxA59UP
2yuinU8h0uO5wUl80MBjFfHrB9NiRQURGFQgbdUrl9ZixtvueBN+HnQZU+3NiphnGKCfnJ7uFIjZ
Kr2OFXRKVY5rGhpTApwAiF9zy6ORQVtiQZvf59MewFeEaWUkilTGT7s7S/cUuR2Kd59GUMpwBD7X
AcKjN7xJRvKCIC/yAL4D5eSKByVAOUtT9vUg5oEm0fP5WwW0WByo3zZuSokzauH5VTWSvdO22CDq
UmWYI4hIpdD3FWWotVI+koTc5kzUhALMatHztOs92KcQdWDpopp6PGmzaQwRcjr4/L1jXMhXZndH
bL3yYg8Q9cq1D/VTWgB9FdV1Dw74uJACq9EvjmbGqav15Vp6fnUEXlO9xbOW8xm+7nBJvRl2W9JL
6fLwrKI+/jgbaNgdUWqvx4pJnxiuxgC7ZJofnaK5SqOJjn4XZxemzRqLMDI8qkFCwOucDfu+aepG
DU9un29aUGEQnVUCKz8fdOUVL8+Pj3myKjuJw+JWBlORFN6/L3JPN6PocPOXJKXiBcFvPW69BbxG
PXma829rs78Fx2ZYfs8atqh9cs1yRdTM4poNRWRrQbUecYe8bH+vOwfsXVqUe6pEyWWiIDpbnFE9
G0swg7UK3hgtYHmV5EDa0sU9eyBrpVmqutpJi3Qc5obi/p6xBjgqkPndHNtxT5Q2dulXjkCuorv0
Ztckd6vcxcCsIKpv0eNAQX0l+A2khxoa4bTUzU5TwmmWrf497alhKuI3+swhywvmn8xht0HJUfzt
TWfhtlPB63yYqx+XfVgBm7pROhVSKRGiqIl5RSQhb7nSMHFWGrljF7nOoUAnG8XkuK9L8uqT7TDe
kIjmt2XIDo4CGmQgBHyHYNjVzGKYUCkYqOwBtSu0DeAnZ6kFSjUIQSaNv1QuaVn6vKwghwMMVvjr
oZa+aYacZUcG/Aqlb/V5eOnM2EChuS/NiBsehuQLxVtIEOyISd5mYC+OB34Hs6GFe3FUK9q20jXn
ErwwJSB/8UsZwBG1vcYQLHVYPfKbEsBLR8SOxv5LeGZAMXxwBv4zb0xbo1AQ75Y9KfsaX86P+a0c
I10U0GR03WZrcoimXhML4uTbvul2qmvf2yD/jUN7VfTfYwA5PeL6S9Qs5b+cZluIVdE7tdI4aH7x
4K+h3f0+J2PDDRbneWKPdzlDgZMMz7qALupyvlpUBJqOn8Z8Cvx4KldJ7wVHtua/HciAM+Aow9I1
dyPGlkGOmE8PaFjejZDh9PYEnLP7pSCSw88DuEtlzNWMCJrpmt1FcExbLZF6S5Qj3pzYkQq+99iK
wwOSHwx2oiIkQ4YZcMdlHmYfqH9IyWfYn4W+V2mA0gYrSbokgp4enwQezJgQvtGQ6Umb2GO7Vem+
04AnXEbJ55as1B5Xe3BfBIS9QghbcNAxzl7QDPRXmT7wC8WLjvt9xbfd69vmGgEsvD2wqnRT/dDG
YjSX7Thm0ZRSx8MWPdWy8zqUtcmz5MX2SJJLMyapExiatkELC3bhf3BY9PFR2jmEZkKMj4VmjmKT
paMwyZdtSs07p3bTw0g+GOieDoZZnDPacVMNw35Ix4+rFHzurJjGXOvGGtHvrnXINxcr+virvO5Y
gsNgA+cvYYJ44ueQdSVfVyztBPNykrJrtONjKlO7R0q+p6nsDi/pMJDD2mO5BBGKn1H0HvSQfyt1
sHguP5CLUUsmZ71teWx8ImPYqAp+jVB27VPW2s79W4Md1jAtVdXt/Il2x5/2lEX6uDoDXbO9k7ur
91wZPkG4ow73AlDghli6C1IRnUuPrqx1R0BtKI6q6ZZ4GIIQBrRxL7ImYYK2PEV//jd4h5G3Z0ZJ
iM3uVFT5sicxYYxJp8XmQim82+Fpk4iTZosLJIGon5+egrgmV9YubrSyQPXSGjo4eQfe1Q/APEFe
dOv6oMrH4HVgpSrkcIOVIaWxd6cdTzI44P+ynGHqn0P03YkJB96BfrPecshQj9sL/tyudzDLUGQx
rd1o/smL6iv+BUv3I+wEBMT8eIOCxSGm3Z5rUxSoL3PRvX/oM+XZuNuhtYRzxgJPn2RzhYH0s/6I
keul4ypuaAn5+b7V9UkRR7m26W1jlUO7rnkM351tBwe2i0yGvzBn++2EYtbH4zEe32CNxdUtg45p
BegQMzRa2hB7pkHVpwQol+jnW2zuDzvspdmkwg55Vyw8yqSWgd9mtDGSJWcpOXMexuLtxns0UkTl
CvcgtQgVVMZqP2+WGsehqKghmyaiEk1wfkVYG2WmhGkvj/dSi2kdDh6WmE/no4WRaw3osNDysfbh
ahRbi0ABquhDik+ooqpnu1lEk8MSz3LTo3zyZ1X4z2D2QqJ6YSLWArI6oyvWx6WanG0UbcTuVaPv
GSeA5+BrUkqP8bwbr/cVVxpteo0pPCJ+DFkThIO+twt4D+zK+UhsvgP3aA0UIAwBMfEk4CnfeGTW
9T4I4G/SjwU/hN5WmIQFbUcVdKMhtqsPA7fwrALffer5xOpwx4w3+dE/zH1Oq2c9aiwumnhtoSms
kbN/8OI58usG6W9dOpjkh9cEKyN9jZlmiOIHsmMCPN22tPrl576HQ690EmTuEIBwV0xp/zFUyQmC
j8OKUT9wXqNfT5lwyuqynLEXGWFcWV+lZhWTazxGgPCypoWy4eEi8qlO+mu44fC5igmX3LFifgOe
MREOEQVL98c++gwjlhMMqnjkIdWhRe9e9mx+CHBVvmmQdXd20lFIj2mcwr+KWHqFrCRrofxvdzEO
Sa5n+gYzufekxNncIRtuMBgY4ZmBS6I9MlOHSw0Oqfbwa12Dec1RQaYSKw3UOgp2rHQwlKwMrXvZ
Ja1v7jLnCSKQq9oBQVgvV7/wheuo8lxzsIqtfJWGRup+zb7HTyvf2mHj0WULlNzf2A9+JB/Kl3Ai
cOlzSx2K4Q0LxOoqNUv3TRucTuZGAD5VHQP3Vi4Oks3uMGrmh67sZjkubnvogm4EC+dGY1zaO4Um
1a2sXs0N89bMpT2Yl7/ZMpH6pn4uqnWv1Bu4/sqfdzEoIcpowOYQx9w387OG8eGzPuZuUwlaMsR6
r3GzlYvZpujuIQwBNWtVmZwKlTY/djB7BcpmIhFiVwIsmZorB4Bb1IXC1uWRjZmCTJ+tRtIgaYPK
SJVSZOOvqiDH4Q0CMFOIQF+GYLntyGoD1tCx+CqjU4JCEFSnJKfwSAiF7ANkG/MmA6/qJ7ZAvqrZ
Ull9NSxtbESWKZmWgZsZhDZ7TuXjaPzezi0MGK9yk/i+gmZjEYMT1pgjLjvqr/ote7nBhgbjEAAM
UIONCNZTiCdVXa0ntzrBk8Jn/du35HrqhqaAS6LkK7TFgYUJTD9siB4+vh0RWmTluBmpsmf+Q9w7
7ZVz0qbPpYq9d7WMlzdD1/Ym1tMKhg4y+pfppr/36QxzDW17l24w9PEVtAydoJN6IIIec9/VD4qp
xWDVL7kOkOM2RFKun4TzjPgeXHipRMxySGRqE9Zaf4hPQQpx7UAw+ye79XWUviEn3kej5aVwxliI
dogWBRpF/PvbDVeqQ6swfsX6CU1iNB2io7bc5kqNe+zZVEOkUgW3gZLPaViKj2JLmegJXVy3Akmw
08zhorF6r2E0eKwhG7SIBn1+HPvxoo9UIFu7J/+igevJl8MQ8RabQZMdbUy6I31rqlcVRdTdV1zU
ki4ukYf9GXruuYG45hm2bzD85dSbdTNIhoec3tyaDggfn/8R80AwM8uQv1W3Huj2OPjrKvNywet2
+HETebMS8Savn977RNoLnQEZ/xTcNxL+3ERZnjNppqIRNMmY3jKMtmRCIENqC8mBuWsuYo3U/gHR
BiP9vGIDceNZK+yJKJ6+J9YPkUkfXqGrR5KqXkBU0+rH5MY09lJwcxX9kEYgHJe7DOhpGgAvu+iw
PWNSa+y9OBh1vZ34ncxwh6jfZWhBGC0X17cM8Op6+G1OgPlx8999+hOaldCFYI4hM13GyVNnv9yT
+8rUukl9W/7MtPpMY5Cu7iyBv6O4wyYGeXPvDaceVeO8tQfrU5BCD1iUcyQuXewU1uLd1T7ve3Cx
5sGfCbkHZOnnjtU9zch9g2eFrFIE0hVGypVh7xCZ+Y4ScMBvFmlpmyKGb6bZ9xQ1waxJVq80z2pN
mj2II0SbdV8aHVDWUoLM9HuvMJ0LN1AW1b9nF3gkogLv1j+3TVvUjJhUslQIU93io3dDfcMobPLm
arDs3v8giKdRnlLJeMvUBh8xKZXHK3C4o37aoxPF5vk5z6NwnMNd0NpUCEH2cxxgjhxegvX0vLUs
E+exHrgKLS27yZ0ISKGS1NnV9/+sCKq9dU66isGAsNr9aybNwJA6w7zajxEazOQCizWpoL/5XaaM
WuiDtedUyfvybQQ/InHVrJYS4pATeKrKnDY7yUrD/R0khJ/kDogWw7lXJ4cLDjPfz6eTd1/wt44m
JcodM8b7or+NtCj64BZ73Zc0nDjdW85su6N0s+WBoliaXGmREZaYL16MvfSRiWOzRKIZUoxSGV1F
YiUyMiJPA7FBgizyu8wmlfEsWrmQfcmiFUHar/VclF4kOEPnSuxXy1Cge4jfJqb1Uvo6umJITaGn
ke1Sq74KqsTONSYN0RaOG6BxRBPV6jKUDdkPfx9Yz9TzsxryRzStjQs7TmdgA+XqCI27xfcsxyIA
ycUiK/QUpBPZMSDVIfTsaU7eJspWAVsprtuOQnjl4Z3D026i6qHWXkJPFrau4mbEzlcZrLUusB9L
JdqolU8+Htj7L9KjWsbkd1tWMpV6KVdFHYs5P9nCFiTKsYbUzRWbeQ6V9O3p9FWsa5ffhK5tgu4R
JjEnqzK99szncgKP0wC9hKarMIgrDIY+kRT58MqtJZQJ6wk5FTIi+SROHZ70W7Zu+Y3cG/rE18xW
xk8WVQfi7YS8qoiQgx5msFCRJKhHej6LtTcj3qyvaCx4pxbzqWcrKOhwN6U9IttAv0yurYGX/8v4
Hm7kpeFxnx9bjhlMV8sfozdNWrNA1ZULGqRSsap9M+YmoSAdCX563D+yYMVrPezFe9/WNnBplGaE
8yoDAZvHtgvECjQsllNO+7tVXX+YezYXM00oPlfKNy4njC/Y7DdgGcidCMpSEVvfmoJhbE5D/pg3
qR2Xf2vfG6UvgrVmfrEAnC+EUDjEplCYfAB7OIBJ54at+zlxvBTq+fbRQvm5iWeIWfEjB/FoQPdZ
xFW8B2CeVxYkVViZ7jg1FqsV5Zak3VUBlgp7V3Q34wykC6inE9dLVMJA/b7euLqs9cPtVie7cmKr
9hVdS597doM85EL0pD2xsd5rD4vDqQmMAXh+HsiacSQTm7cJtGx98YI/ebtJ2koo+KsTkblxT0PK
/UxJUmURwvAHmb5ZTrPdL3iaUiOQeTJL8yTwtWnaTKX2i6OSIo9+/OeEy6Tc5lcmpTyjMm3WiNDd
BXjkvhs786yMMtOUrrbSiht1saYt38pOpF7CgIislLZPM5lRj3WH7iBrzQD0mt8sKn/SuKxS/6U1
CBFRaaF0gP+mfvxNKMrrhDH2ryPKXI3pQgbHTDwGoFfSLRYHV+32TE5AScSU8ouNBnp32tioL6NM
bonDwlXB6NBi7lxAVuePLvpSJMxAvKSlnmAKt3q3xpqA7YwRwt/m8nnat5y68VPz5oM2d9FddBSj
75k2xtK1smbZEVLzcjYtP/U/XbeMlrM+Fuwlorn3HGy2N7VswMpJ9WSR2F1M7tt4flLuq6jJMMxE
tawMLLeq1lVIZaWg+Wrx5PV0/X88I2rqfjPu0MEC4xDsnOron3mJuEBZ31FvAO8YgjEYxAhYUIDJ
YBvEYVEU/ig3Pnt6dRhC3JkDPo0z/R9LqllByQ+qlWgob19VTOjO/GvyKqJTz8t8k08rVs2s6NWA
TMtIALSuLhVF5Jbgcgsad8L559ANq6TzfaQFuY5pi+GjaG7/kKXM1/z5dvM9ucsjLT+tk6pWpldN
Jx2AaXrJpHsRNPyi53G+73hapheq6E8kJ4Tw96iyHiPdz5Z5OPgc3oHOCH7DuO7smO8ljPCwpj6I
UeGvInZsoskDsEVoa/ifWqJVdU9h56hNlziq0pFUFPvWIPoJCwAv15GOsSt59ALXdJWJZ8G7a19Q
60emZm5KcQ4S0H5uQomoXYBWnzejc0erKZLSYY75wVIdU6CQGm7tE9r6TzGmhDeOQO/rdxoqbW2o
OVl2EpDKtVk7DXPIX4UlX0kRW8hFgLaz5Oz4R3MfwcO5nsZMeO/tTYu78TeRHSVGVnZ0mI3ZJWTY
HUaoHBpemGECGf/vbN1ATG8rVV7NqLynngyW//to0xYSWpTEK+2KRrm6/wnG0ScfeN9Wm2wmN/0n
uqY9Eo15/JswgfQtIsCnSpyCV/nJxfsUIiQ7WgiR15PW63fcZBxXbHdCHZGdGq3gGYzftGH6+uyI
GllcHEUM8UX3x/IXAWLu+w97G1+5k7+9Z0VvPeXGqfGzDRPAjQVakdk4TYKK/ul+YEejux3lAayT
pS63ZXcisl7UuvGobiWqeb3jrqvPYDPzIwJbeD/YHId1FO75SrKcWLIPBOXSkA2hA5DteqtGxVV4
re0k4ateKJ6537RUq2TKB8dSjvjpyG2f+ZolJKqfdmwmaaZ8wt4DZoOHUgnwsBLn/Ws2RmiIDV46
NWbaCb/hXwt7aVfQIufSxfcV8WOOB+N53lWFyLmKN21fvaxtTGxHi7otOBn+16uKPKQFwfpy2AkB
pRfttWFNL52jE55akN9snwhEcvYLYnlOKNdhBk5cGK7EMtphbngqwUmp2SqYHoIDovJ20NtpkhMk
OgSeA8LyEeSVF5CO20azlMcixD4jFH0KRj70m0GhjXkG1YMsRu9TiCZxjad3cYCMovsmX7o9E429
7wMWQWsT0lUtmGIMmWG1/cQBv2MJOVUOXH0201wARRDp/+9k2YTBWI7hL0whBPZ/fqMNN0qPuZB+
fB9ASnfEZ999RZmcYzEPy1ChfCa9Q1UxHQFcowPnRQuHHB5apRC6iHLQACrSL3asmZcGfzaR8HOX
RmO5QQtb22oE+tVZ6QsrMW0vh73nq1ZQaxp5p+90ESmewJg4lqhL6jz9Lua8tnVe3fqxPwH6d5t7
pyab/N2lanj8qGqncxt6Wfqpyrdis1+BRUHRjFP4MC4bVzmG0nLKTJPCGp8rqEqYyQDsXbW1VCkT
sYWMRnBdEKBmLardC1xSJ9QhoDZTqrhQ/HIdJ57lxa4O+1QWDD3bU1G4QTZlNYn/+H1Ai/g4ryZd
h2qFvOm6H0kuPL+Wgb6J+hcN+HYRfNOEKhhorwwJcSq7I76CDg2qqo3UAbgdV8oOp1Xxh/NVSSk5
AKf2VwWC11gamOizWHUX6OqLfeagTCZdMZMpbtUYSYtXIAABc4WNym9P4RnpGh0oyd5DVeRORgTJ
cAwvwqUTHfviHjzdGdLVnsCiNcV3Wq3gTEz9/YhY5AiBlV3ijYsA3NXw5qq7MonQxg0ZVs/agkX/
TctEBwvqZR60vtPCaL4Zvh4tEHc9IqK+TqcpuwPKR45uT8cBAmiZeh/5VPkwMO8LKQNYb+Lsa9Fs
aUVJttyZDg/UbpPR15WUUYrMmW6/FyHWcipfDs1loVhGKmkMsUMsmS/Bdcuu4ls8DUEBNUq/ciuP
3IDk5ePBGUxZRjcg/A3I0Tf5niwHpdg1aEzzM0BMkycxv6DbncZac/q39fb4GaJS8F4bmwdS1LUQ
O8pwmuPkO81eP54UQ2E2iXp/S07O3qyR2VWwbZK0/Bf1hVJyd/XJxjz8CItEay2n8b7Zr8C9UyzY
/CCCUDuLBdqVHwXlvRs/S3hWY7Lz9MisdoscCjIAmLLZ+aKhy5I6JZIuL5NqqF1hUmBozWdcBoza
zAo71BJGIrHQkTZB0r/yhjonBv1JOSgUzqZkAbD4ZaL2P+CzqzubDKGqBfR7uYf8Wy3mZF4ARFdK
M08XPytRU+Ytp/tRiHyJy2WrqBnbZIYw0wgvdvDCVNIexp5OQuBSPOfhCJ5AxA6o3PPeX1xJdM+D
QgPjRQ/H+W475aQ+S6rnejvrzSaonFOjnEG8tICDNe2dJb3rYbYcl3RKQtdD4suKafvQO/+T5tnE
2Kv2YGjQyzYdiYnYHLIRIKqbAwSOdRiUtDorCr0L0/0OW+TvL3NEJRnP133bLugR0xQsfFmEYKaK
p+3qzgNQlXd4oCRdbe/JNPxM3HxMbHlqtuOcFiNnTmTWlhaS46lXwcF4HX19qjFrIbE613a4XnI3
BcXJUEKW+mvqkNhtre1tAVDSla8mdZmjDGPwnbjqlsu+ylahnd/KRG9h0FCZhK/HIwrIGbv4wcOU
udqMcYypVi2g476Kb5oSaN6Nk6c7VFXCVDU5O++Lw85zhgD06jXM4Y2tvhEcNchSyOrQXEkD8x+O
03WyqM+YeRyDWbXg4/sTis5f/QXoDdsDMc7tDR6CLUTJm6uMAn/gT36pbdXYYw9FcV2cqmStLRbU
Ln7b+Iq8JkYYd8g31QH3hK6KWWuIRVwutsY0J5LW6RHPoozT4RFTDJ752T9yvlwyJAFavJN+bmnU
j8NTM/8rfrYo7GzzggSCY55YEhEpVEPnnr1lPf8q8lTEm02hvAXvQjeqrWV3l+crsA/YFr82vudD
yqQzw4Cwcoo+Ob9Vib5LPORp5kWg7OH3zrV15Nx6PDranLhGZafim7DsPsbaJblFkogOoyFjzZbC
CRpYEo8y0I5yh4W6IrItAbETJ/jNw8hL92JRe+U4gpsSXfFCOcpfkvyCN8eGyffsJ6vY0SMETky2
3/BXEeGI+FNhRxekAZvGBzVNDctL3tiNYwPmMpS4WvkFnehdLG9SCJXRBBC1Pngjhl9BdLmrVyCb
dq9mACvb+QuyGkNGVF0HOC42uxWbKhN5HnQhD7FLZYlU13LINpSjzHfWI8WLL288PTJq1RIzlHej
wuJdLQa7D6GctnczsOZ28BKwyDiTbS/6pdsix16kJMYnwSGO/77A++D00i/phmupV8FOdUaj9aT8
Vg44PRJjl7bzxZ6+CN9OWW4b9InuQNbNIGpz/Cu0MaxBtks6uizkA/HMk7PdbB3Hdcy4fB4xlAv8
pIGUhh195N7zP6EeADIwbDKX3hHt6E4J18OC/U833iWf/b8TtEBGl6Iyip/YS9kN15NPsyG9NsY4
pRPu/fh4lZA5wCjWjTn5CO2f7zbboCBMP9plmkABdT0oq8o2mvA6GWfgCNX/E4X6D2TswcUbUsJW
ieTeqRl2Q5pAAbfW07TQ9c09dGQBsAsdL8QYoj1GYT5fhwLhZm5jgbMrik/t/Z9ACJTBuvSLHeYd
Kd0Kj9evhLLgq0N417GGsZooXhhGmRiy/wXcfdn5Jqh/h9FGAyDMUwFJFyEQd0xKcQnQCUuaesPr
EAlZK3N4b7VHECAF2kqIbJZRRVaV373zoc1YSi6jIp2NddV7SK4LzghBb1LxvoCExwIYocWUBpi2
PfAfhXpk8upzr/1LeTny9eG1W5dV0Y94llqwX3GA61oTRbUrC56vQUhFxn3nRuQ5wQW15AJGLIrq
HwD2IpYEaRvgbmBhJDlghwGO0fc9TeE6ayz9OH11+rg8Pm16YSneId/MJHbRbStci58xE+9mC8t0
4RqTbd6FsFw8Evwv0xl1/QQdgOmBdatmftMf31ZosxV5N6akQDCVz3OhIc4gyOL+Rb1Bt9LGsgWk
OtLlbRZHsjlxngo91VU9RD2YTo0gPf2hAhTXbk1isHuKQq3jIAu9ParvpN10z74vfAwhohNBLhq4
/IdArFAIvZzJGeqRYpm0+nF2ZEUFKrOwfsejtvY28hhUODaq7SZNNZqb6S6iPVUGKDbAjkHSlPCc
31YhAo+S8lmPz/AgjI21kd4CQpXsTdeIDcMzuMRAT6KYCYi7Rmjaaz1CKqB3Z1KfGDIi6zwqLDoT
Z4mryh7Ld+J3Fv1MYxS8nZ5ShkSeqil8PIcF0lI3thzXZ+/WCjZuF2bcTqk0vJRll2zE93GzMqrk
qHFahq2kKAN9njHxdmfhP9MIdx7UN3PBcpoa7l2zC6cqAUldrVM6Czq2dasq/qpmS1WiVDbzk+CS
/O3+cRz70n2cGwvvYIyBLL3vw5hLdD2VfuVukZaNTyD25m3yGRNi8hQAV9w4UcBwkKbKWkGPMSjA
Bt4mzLMOL+Qw79aJgKbSU2OCjm73IfXg9aJXhQYOAZuBh1Qs0KZTIfYJ66ibqMcxa585LvkIpHWF
hi81txm9qf3FGLTGfOaD35460OQT0/3vfMfApz9aJGcgQTJsBeWJD6Zsv2oOjrPWw6DJFXunU9RN
nmrnhFaiKyOM/zM2tNWNGokfvUx5L5vmWfV13EiR1oW/1NUai0n75bCjOpOP3eFQysWyt5c6HAjb
Y3WSER5L0CLRZZ3+drRfpmQrLNHSkH69FtUmO5fDWO074HVPQv2PpamDw+Lvo9JQORc5rKR83XcC
rc4NCyT/uerKUO1F7Reu9lCXwErFM96ibkIq3H58lTGNdQAekVpvAiDqE3U7rBZbVeUCVYH4+Ywp
H2LHgPPi8v/eyROq0W5jmPBcM5ua/uptPv5w94xB6scIURdNv81Sx2g9sUpl5AOQVk9Mmv7jhBHO
GHOA1mJBWwSiN8u1VbpiZTll9HgIIMkd0rss2N2itYhjCISWgcefzjtf1pUI8YW9PKGIvhaw8sgh
ys7J8gtmnFph0ex/ChVGf1ZWPxkvw5z+xD/pvRkUGFXK3gkQF2rLEPdqDBVY6T7UUCEudfQvApRZ
uOolg7dxhoyM8vTGKELXs/X0AL/tYLUeBK7/XADCoj73GJilMkKirnU50hEsfRPzVMmvPDjQvYp3
Z6BjnrcFoO21PRYdCZjWQg4DPG9WaBbbaU+8fjl3ftsYcjSR/dmD1KI8QAC4EFeePZo88YvESisq
BcC2ANTmMd/D8GfC3jKb8Y1PUNC72mxkvtzQ89KzVJkXXgxLD787RPhbUpxdUXDzltXC/977SLl8
cYLilLF4NebtOslc6kiu0QYczwmo6j7YuGtwNvHo4pn9blaEOlDB70AnziVeKzIdddeSlMJBZ15V
MIX2eR37DXCLhoxhUkA/rE88FDwy4KDVSSBYWI9jYXyVHeT6IKaFHANF0nzjudct+dTSkan2ws0Q
q0nmnV/RHd/aEieo8EXNPAbD34Cz88IsIOsTjmO8p+PMT77lU7s9PSBxFt77Vt75viGtGt2yERJd
ALtFrmeZBdK2wotHfHqrLwLMciQJg2/VufOSVJDWVCnXEhUOhQ5Jk1e+nKYVTxsitpG/+Ls73dIq
Epn6T3i0aZxGa6URoa+llSnnNpDCEutw79FJlRUwFOQPf2NK5DYRxtxx6OkpC9ti64KOI0qqF2cB
1+e7g4H+Ly7bONaLK3Nar2nWVZujzJAtoksmjek3iaYqYzplElii919chjp7kXL5v+Bszv5AkQSj
Yi45rFist8KSVq6uYEvEqlPBYPKt/u3KoHJSepPU55cjI/AxRvcDw7eEjwA2Mj/tAR0oRnrpUO8X
7PWpyjrqrrojSkLVwsERcuxkF38aDUDQ8rP37lSxcFN802VUh/attDMhmXNA0k1nX+0dIBtoNzS/
XgrCYSEG/D/bmO6B3/e4/qGBhLOyOVBSbD7B0aoiZRZOPvnBMpzNI9yBohgv1L94R7D6kFbbqtB4
hcDFZIsyPOavlI+qO6IKKUtz71HYNCzQZvpRZ9jZNU4h0i5YhG0XpLIb37fMGvWomqzfL579nE7S
gpqBUpsgJka43eavWjSNjMaQ5B72STu2Khh9kIEz3gxFeEJHUOoHHxXig+jP4DJeInPzpZ62XGMU
pMOmpFGaAbmhD3wNQbk/kXFuxiLfVGxQPP6HxMc7OccyWobonhvAGMaCyS9RfoLxUCSZ0lbf4qO3
POP1Z/om3Wx+5Jhn7HcJB11bG31A0sgO2bvMz2hpN+YxUQ9Pv1nM5t+Lc7obB4W+MMBDgcnxChk9
METnYEH6lVUyefJ6AFqDG7Rz8JmAgxV/3KQKI7bHuY2cG2Nx1OSvYNlTMKewj3Sgp8fOFxTV0GRu
HDgztue4DLU/xbBVOofYYLIWOqp5yZ8x2M+AMbejCRKytWPTN8EC/SmSrPi51h97WSyuz07Ixqys
Th1PXpZ894IpPJMYuvJx+gnbWuplPWuZi1tKppS+MlqU/4IjJPX12TLZS/vrWtew6cpflQBBphyX
pNmSIiXkuW9uXckQ5qQG6dGFnoJea7r/fCCT7VTUKHoQSJRhArw85DVfmLvHJHPm2AFSWyOhkmfv
I2rGn7HEHVEH9GIcrd3bWmsVDeeu9dW28CXUQXatn/n/NAN1Fz83Cs7XjtU5cA+UC09Wj7n6mviG
LWLKe+aKrIMSs/b1uFcKIW3ALmVOypYN9VmEbmEt3Tg7Q/4Emo7A9e0ayOSYN3PEWGA3k/1SsE4D
WoL7xFqOgzwfsn+pKTSib+8On3w49rKymumhmN+9pCnkhe3JE/3r9utOqR8w+PNKXRrlMQR/ntle
8fQSnhJCF+W0DWl8FUipTm2y90vgBVm7Luw/TklSn39PZJfvhdMrKa63GhT8/KwsKooWndWS9Fmx
j0GXBTaayXJl8mYaZCvrt8eDC+y9E1mQy8OYKdmC9kNy0c071xXvSuE2L5UOOOTTAkpFIvznQBaC
g9rjij5vQnmr1SKgFVHOdLoQ9EnoMIjB1LXKFqsrwlCE3NW8AvCF1LmOuTBMaYZDUXP0lERV93EL
vr0q7pLYRyfoyQKAIwcznFwb3cbQQpdvYK07whmMAjFA3sPby9y5E8nyefpp9glPruGrepl+BAoJ
ZVf0rcP3pB1O/0XJ5OWU51GrxKJ2MKRKzzDsE5wnSeepku0tRXMRC8zGs19ZuBJW5/pT66BSm9fn
ms10aHQCz2ubWkp+mDuD2InvxPOjcuilKxvLwFaDewvUD9edmpBiKYzuZLHgkuUx38S3ktASQJ/9
zX1Qh0H7P49rpP5PVT9h8czS5P2yK7nGGVuhPAu/sMh0+pqSo51sc877bqQ8Mau47yHiNjZFlX2G
4DVfWvg0NMtR46jVUmWGFk5MEv7EVjl7eB4Sx895L715IpygB401rdyWrqQupDWZUI0PymQqpblJ
lBEcyTzdGHXuRpNF7NAwMjHHQrDP+ySU7/17ee5nD4MaNaMNpLIw1gBlUHO3QlyeCgWxb9v11zBD
NV/yGk5ah/YZlhc+zDpq2HQcLXYkzikGvWACShFn52pM39a8gWXr0yFAGtJMOpGDNOAwMxupJ1HJ
c0cGedOo7ZsVbN40d8VYCHAcPK5H1fD0Bh6L62fDAByL2OBtUbgWCF04ryZZWNFwd8bmmenfuStG
mcplTilz0kvhKU6CWo7UqmwtRnhAlhQk9kgcKkTt4A+jHvlRbtY4mRtMEptOTVN15qRRm7ejEQb1
gM5U2Kkz45sL5sA970nODY9dL0hMdJg/Btlg76Ao6wK1sS8nk/Uq2uKqyWmkmVB1W8vexvLhS610
z5CSgAr9SdmG3rT5IChSn1TL1cCUO9JG59amADM4UUUGKO0Ew7Pd4k4McuHNvqiRdMCHhfgvlZBE
R9EK0i0I3APipXUA93lLaw4ucpntFbM546dDT5ImRAaQO8hBH8apu+5rA2jO+OUSTQyjAscARgZA
20vu2oLjPTyrOMREZolH6hNVxxHOuiFjVefv/oVMZS/jqtemk/d7TrTBsGy0L6TGegEsQ08DWLeA
9CZNVSvcmk+AxwwM8VQdT2ONjuRw8oSEU9/ktKS1YBm2h/LjF0lvMCgQCJ+f34ghx2xVKMHnml2w
MLS+y5Gl7BTEYSOfJHcxOR6n7brFJmSLzaNue/nhHuEXq9j6/Ir8nZUpbBDiyXdwqCj4zFEeYnjn
X5ZDi/2wINdgFGMmYwhM7sxGLME6sJ1koNxvZLExGwl5MBS0HnyiyP/NMY32xzzh2GPfu9qu0kEv
Lb3k/tspb5DP9VvSimph3bbcMExqVHec2vXzVN6N+wTPxQWZKjrCm4PBnNICpFe7wAzFM0Bc2cP6
AJ3xg48MpSukYgEkDrDvVdobMj0NXwvKwlceY7XR0zKhMTon/l6lDEioPwDLslhYBNSw74mpTMvy
TOD2c9ZWgps65/QdTP0kqymshC36v0zI6cuvMnQZiHMeWhG9wfADz6thmsPIO09CoE8CNCsYoBC6
8zne4HEBmR08a9BPb4W5zvOQ2MGpsNGcq0ZuD/odTuVK63GX0yNmgo8jb95csV9YNCAFWAzaRRiz
gRGa2/wBB14M/dSpZuNFwzwjHoao+chDRm9VV2dt/QCPMOsSEMgIfuacAnukzhr9Xxk6fzBUdsOj
0jeFAhkAcwiF5RP/ltHsQnq4Kr6WgFE8CnmPHtlZEmnjZSnDBD7EmyJPe4lDd25JyzSCXAaW3t/o
M9/XhO9ZZJLBofeoclHCJwaLoQ/1we9HVVOm4mRFKSv4GpPrSK+1Q9+N0QWI8DmtyJ0a3iddjYeb
+dUXWnM4gEbyoNd1ep1JGKxKlF5elx0PlYq/2oT/ETm+xX9XazenTm8bNWSXA0YhRixSddQi4X1f
YHbkbs6Zm54UDhiMraQAYCfX27FyycxhBS8sY7U6SnPdGN5XFCA1capfgqFbA0Ufhjm0jFvI4YaD
MUczGhQSma+q5JSD+W5BdDhmF1v+o9xIJh0lqq0/RIPAwYyihGVhkTnBYQNE9++dY+x7UiDE3gVn
O4lZzPcdm/l8/rxz/Jp+YAGK9Gds9euXzvLEpNZDUi6TyJ85CnopFa3qMtoFbdboQkmxF7A8BoGf
TuuLjlKJtI+hIl+tpeI/0HA574qW/ljn2MG/1fsMVXreH6kOvspf2Xu0pDD3KlhJ8+bLx9CrhdXu
oTUW1c4RfpKM2ITBkI+deZqUG8i06spT2rzKU9ypNLcGyz24r+siLr4vkNyQkL6EPpeUZWDWscLn
DiAXoMlECp3SJ/ynvcBq71CQuto2QOT9oaLiV468hvZJY6cqwX9vTTcNHLSRspgBb1eoJG0r9OHT
91dVJkRs/Ih7IAFujQ+2qQfy4uaKNWX6jsGYeAhagtx9hBTdiAAVjCPn1NqdJOGKgmgvt+QMwFix
nkWrEZMagGtXlRsv6KBsUcED9e2nOmZiBjA29qZoODf9ajvpuzmKlV1NWM0F1Szxy7LK/0E3ZJQ+
D7Qz4Dmaj/y+L5X0an1Bl/aqobDXbdexQ3v8v8asqpVwa5DgpnQ4qyVXDfrttyQRlW1pZY5UHwPx
yAbN/KTKwLkVyV7UWtse7v8rDZ5TJrM7ssoYEDxz8/Ds6GDUgpYItt+i9WbcQ67AjxF9d8vM0l0w
4mZCpBIFIx0iHQ93QxoZLYoUyfoyPIrwmrzrRFE4Ytwg0EzIysAj6M2t9W2oj4YbcTXMq+xC3Btq
VWGclNwH1JXhRKbKs0ObtcEYlLwGosJBTRqrVvIGuvf2x0d9FXa4XHLjRa+mfCY3ZGL6PSDkp/ZK
q1/pwexaUrpqq/PbBcDCgF2vPIoiU7PoRbTnmt1RAfKmOZx+BWylK2nD8Ji9P6TNsUP+qNR1wAR3
nYU4A/60AYJjSzUf7o1DW67OovRZ83JUoryoadOlYGM62Ni8d0NwqHh0S95RfqwWTICfh4Z33b0g
V/G6dotEBJZeiAglgj2A8FF1BS1SvwyDCbCiZp/FPxdd7G+WE/+6smFrsd7iIp5PqO69bCpfi1zg
PMA5c1zqENvgWcIEd5nIHq3gnkdI7FnLButd9EeNnAAq3/SydCgBB/JOJ3Z/fhmbkvXfZ1TMuCf0
AfeteYAnyAr7h6olEZCoDm7ReCQrJa9QhdQ21KHjV51vlkqofT3J1z27RPc9f4haDHWSjID7lBxb
svjoWeL/wcN4YanSVKyuBAT2EM1zDEQOSCReg0SnVWy7U8FcRNub9iY3bNHmlG1gtFaHCewofraK
ZNXWWrsKCNgvhWqLX5I/C0b1MrGsqBsR6Cbykw567PzYuDDBs8x0X9okKzfuPmMYvRk4ERbfeKRS
iTp/lyfkje6CNKR4HKJ5eCuPEXfclpJPSCk1DPxERiMtDq6jV2blzpjOlHzrSJOdJ/LkypQM7ZmX
4WvpD5LJjVPFZ5ltmFPwgra1v+ASeW3Vl0thk7Mzwr6uOxKA5sC/zKK3xfi8AgBqjaV5Nn2b/4jT
p1I1RWl6CBUIgqNmmTetAHiPa5lh6edJbbOzW8ueGviXiWPrHNaqh6vPvUWg1PnX1hHRLMqkdODP
SUCeBQ+rlKjl5ejUg9qa3aeJn4vCqkknKBNggHZf7QJbadir1/hAKM4c5bc3cAPZtHjLuEeTccbH
HE7/UJW9Xk2jrobIlxnImy6t13fjqGWq8SMY3gaWr9Jhh55GQ3ogH/xNKPfdXffysRyYI4t8F5qH
hhAMV+oCde5T3JYHuM8SB73t8XqWYVmE5KiJ3KBci+A3vTjKFVDmoT8JIwB5Ej/EPE10Jt65h7SL
HO9bIj1qd7YZBhaCvHIOzuoMz4oFda6EJrb63MeJuk9W/4cduu9ADkOXXtzKEOaX3Y5O8j8g47oI
vuojNvO9r7bIBxU+Q9I3q/xg6lzboWU2qQTd+8JIEjSeQCLR3Y8LWyT+nTMUqS4jxH0JLTLhhg2M
9ao1a4xqJ0gIO29UCg6SzjUyMo/9zwyQ7L6801lncbqrYxzbGFU4SRp8G5VoXZNx7zBb9FMru0DZ
UR7Au8YzLIfYFdW193+kiUpHz8r0L3WtR5nVmo6LNtBuxxd+PtfKVX0HdWHCz/F5DCX8Z1ZqHqEL
ZARhCAXOKYUKpd56Ax2PCc7CU4aCrRjolQy2700dICLcyWSrvXZBOXXF8CHhcuAe7E3FTtBnKeMi
kdrKZPazDVyCzioPl7zss7lSI+tDf+V92FghFOq/H/0NM1YU27LsskWcshgtTHFCoaILsN6Ifi+8
kxUNw2ECTDLIv+sHzy2dd/3caz+ykNeauAFGH+mEFK/QoVMYOahZTZrazLKWtwqOFZDSpLx8WDV2
07a8BnKbIrMHm4J+WvSGI+PQAJ/xYyOaE1c6M3X6UEMBIEZiKdwGNzMCeovFaQd35ftWfZdXvSvZ
L9TtbM9lSn6bIVyKqmulL3CQqEJi9WGa8j8bDiszzZpLML0pX+tFd73xKE1qMwn/A/Sd4Sk7qe6y
i5GWi+CoSNKPxVSZHbZxe77Inhf78BO4Ke7et6FHMMuRifAEH7WPPE7DQJn1rl/WgA6OWxHIfbna
F5/BB2aPzR34A0aamGzWKpNzCwT8uvn0xxO5h+8WUfwwydm+GDnmD6/z6MSgKBEZ786s+EIKAE0I
aS9xMJR4ZUmAD52AnBl9XUDf/diFKnS5mOaBbH6TzNol7rRHIwuL5zGrKYyNj2vk8u38CDRBftgs
5OXxy3EFfEHZT8uTu3yX0RlC5eLh4wD2/Dh4BXuZu0wGomkgKcOCgT+LJzJwI4O0bgGEV2a714LZ
WbW0ocfD3ZkEKjRJ2JuKNo4VtqC8LVX0ETnqHB5aCO8ReYHA3uFFrXAL8pZUcdlq7RxUmEcBNB6I
O8Wbo+td2hGjF8K+Osk9urHCsDQN/wB9qwaCh/pHBOpcZksAG6P01Dsh2qTEXxAd43YQGOlhswF/
36bBnQ5RwpXmN7bK7E3WA+x6d8yTbESkzNeVH72zUfcEycJ8zb2C7J0dD3wBuce6nOXg3SMuZPct
BMKOIRs5r5zN6+9DMUdO2vg+/+rWRdKeV2ydjQ8Vp+pYxFef9oYwlKBgypTtAlVVCKp3aZgySt2t
MAzfHp5qpNzC+qpeyHYwijDR2HekcAuzzLFMjw/7Z73QDuRtPyUdYDzaLofTB7PCxT/KkW4WHAKQ
+y2eOgU+bDri7W4oYch/ZlxkWQHtG6e5QDnu+kY52NeFVhyPvNCJ0dkxrAyjVQvnjd/6yxoQa1Aw
SKpHrFHBXjRdrt5CTAiF+1AcC3fm0oSSwCHJ5HXlbKUuprJCx3ddUPhp35Qg5Z3RSm4Oop4T0OtT
tDx0jrP2zmiJS4ulgp7XmJPObLLuT5naC0mooUHWJjOltn+CevW1AudQaJhE3gcNTNQO28hT95++
IGxRSIqKhN31p+7JVDvc7g7pGZuoceEiQ1B0Pns2IOmx+DDQaJOFADL8asc30GWxAdAOKwmBzoRN
jNNwcGZC7khHiXZwV14MTW5nP1DbnYCeFifbaB13fdXhk8+RPmm2CFKZP0vNrVIFF5hL57/fsTxg
tQ652d8ijaOdUd565ja1Zex6OSpkgJKToGlDXd0Kw0sJgMBWVMuV7WeGmTUkbwOj2YGJyPNSk80j
J76GhAKeEjMZATUXXboZLbH3NTJQQVN7jo0TEWJNwqnDYfxFSw2Ms4jiU3udkjO++rfBwy3TAq2D
Jf5OVL1Vv4Bqm36j/B/B5/vh/ZQ0YuZfz+8yXj5CYxtJWk1jIzWoUiCj14r9CCpbT6SL5sm4EBNx
6epl8JV5gk/pyFajLYW7UUT233JDLaj5xbAynBSFcacC9ufJKTiLgrwnHYOouthC4p/IyurQ65gF
Tszyzvig+PBhUPUf3JSJe1l+bNF/rQBPqwdkXaLfoOo7tOlve6LThO5d2M6CzJvb9HJPnpmcoscD
Uhw/P+sIucdHl0Bo4G6igwKZRyZiIXXXIxcOSj4gTTvObI+nEFYF61qY5o4AneIgTsEPy1ff3e/6
/pVafS/tMmIIW7zThT3XXvDBcGGt4usdXQ9tO9hpp8gzQhOWe3h/ePUcLTgitr1gvTi/6m/6JB6O
wWP83n8ngfUDkIbTWNoyHBCdw0hXkvVsv0jdDYcK8tMFCZ8JCmTVYhJQmt6eE7FcWBz+AvWNl1Bw
nUgu0oCK9eDi9qbHWsx3rwQXilcSrZFzSET0Jjt99DW9Ir7P/4TCUlDiTxPR0ot2Su4w+ihBzN0u
2OkuhvlGXcdI8H1LHE/rgtjVO3vZlRmFMXOiXjRoIpMF5rD6HbDc5xW++C43gtVeenUPUWi7zILX
xMpwGiqj6TJmEmXmLywCZuSd+Xvo0a4w+h4p0K0BoENZGFzzN+z2KaXkQ+19GmQotTDvmY9GrXwK
XdieJYDqOJrdLhps9rpIwqH46exoda3cXS6y+Mhtz/qKGdLCYIAq0EjcmpWF0EL+JVUZY0bQd3DX
61r+myBp6UAeckLoI2Z8xHo3URzIM84++FC21mPBq2MsTsU8cAHI+/ogpPzM55NdEknYIXq0lCk7
k/Ru9lTSQSTJ8k6K9YYODfdd+gxxjmFfAh8VkOLl+OeQs/9nrUHKEChKYyd6RXcDTPq/U7S2x0G9
QOssP6Z/GOuxRJQP4ScXrxLDPd5CqtGGsbvS+48D2jYFGyQVD/wrIhNyAmhAxyzqkdVevRpmzWS8
7lsV1boOl5XsQ5rLABkwxTVtdSaAEXes0AHpkjx7a7wDlkmgGQ2Ncxe6Uihc6UiYzCwaoc27ARvr
yQRB0xMjQqgKXhNP/WSgvyufJfgiusR2gWukD6Jl7ZzQwqZ3i7Ta9kFCI1hmuu+ZF9+Jf+55OUht
RSt49qMo9ADfLkRqiB4iSYCVRzBbDtoa/KtkcXZuQDObxRWyMX1xW/KC/hhBwh8OQlxUUXBWLnyZ
bmGbvDs+GD1/9j0gvA2bwnTgnjYF79zH0hb6F/xztVN9ndYqV092NYMsmJk0FgygoL9c8PtRqllA
W9WprtAJ4tsg0EO58KmRaD6FLhfr0dznXrefwYDv/w3gSQ6q2oDt0sdLRU+gbKUsATvXPDpuMH6J
9SeOPab0JuLmij2pfBy1gQrzg7I9QFxMmtwkooD+rQzs0KbqCvNBGWO/neeaOoP2uMPE677qgQ91
a1M5p9zgEi+m1e96IgMeJhLePthSscGE5XWWDk+OxzS1djozBHW4l4xHVJ9nZY9hNm4V3WpM/Hwd
XUf28rPvt57EqMY/YlwgXt7Xh51MHzy+64LhMP5LVpoG+Jf/ER8ySocY1icJUSu4f4xhlGU8eNgN
tgfXIpdsuoR1FWro/cxHOKjNON7Bjn3NNE3dBaKC8fUvsf3ap34tlXd2/Pn5tC5UDHcOcRSeweG/
OEA7hQfAkXaP1kJnoai7foSuFtrvvr4hjshw0+5AVfEaUNxHphQnrCG6x4UdgZsCAcCh4fCYlAsc
vRiywb04NpRjSAzAmNSaPTYd3JnhKQlhOHZ2HB2XFFYMHNkRNeaDimszpgQCmiA6ARexTXEvqs0x
4HK5YXMTeOGI9tw0vX8Wa0q4aYhYN72eRGZHNxBjuSJglIA5f/d0/dYvHMfUUXu1jlrShN/f7WKB
TSKmg9dRvMdBUlX7RH/S3jkz18vndXxNTWjfuvGD9WRGPhGEshYNrKrTT/DZES+aQLaOgnZAdMUj
HiHJNQqesPOBZglqASo4/vy6W23I4qIKmliIdkJldhIeT7xF7iA/+kvhHUl4hCCYZ+Aznszcb/Ek
0Q9JCBHU/DewosQ60IK10SPMM6kTXOF8ki2KCESINYW0oBYSpiMmdkyBrejkfTWNuN+Ya3idjzAK
SNJ9B7eLI+OvVZigE6kkw55Cadd8B2pFx996Cv33Qco9p3nmS1D9F0ujjO1VA54BXqkpt9AjJJwY
Aby9NY9UcNQvcDzqThg8Phkxzk2mVdqWPgks4N6KGtjxC1089d9Hcx5Vr7LC15LFg7HJo7T7UWq2
TZroXqliYh9MhLVrEuyTa94o1QmYMjeW1gNR3Q6j1+qKl1MZPf3UORnnkAXpOo8FN7CuecC0GcJH
8pa7st4sADYVgo3VSpFConXq5FUE6B8dduU7J/qpeN8SlCSDgbaOLy9adE2IKLE/0FPOMrFDQuZ9
O8HhGsFe2YGBi+ADWUfL07LQPVJfD5EGqJHVBnW4J4v1jKYN9uMcoU9yn9t7HeMlQmnkma/sLjPg
7adcLqvioo6o4BPOhIAma3Jsfr+/JRCHb67cXHlbkEKi2r3h2cGkDr1rjrTSjaTbhAv/gn403DL3
kxvpMgypTPRMGeDJ2Mw03MJVv9MWGHL3hgAvELAVAdeyU4ZwCg7QyEfM9Eu7q/BGW59pNLgchCP1
+PIO6j+DEkOQtOR+wt8CGWo/Xn7Cju6KnV7cd+teC7GB6X2JnEpN2Mu2fRHIAXRQB10j4z+X5g42
Q7ip04wfVyJFFnhIji4j5Jw0Vlth5tCwT3L+p3uL8idQQj0rojuNoWE5avTSahpt3wNwiCmP7LCu
FgKqjCnwYXwvAlBTIKPMbA0DsdzBvaITJL3+G51OiB5o89VZwB7dictzZV5Nzb6L34Nrmb5czj8h
sD8OVMyQVnWKQYJ+f5PiUW8SGq1FiSgpL0zPmxP//39y5djlEo79iCq9EsxX7mUp5eRpm2JTYRfe
zRa4GIc9rT3H5p9RGAAbHmybJpEGpfPq71uIUoNY4T5cr8oj+JeFQs3cOkWXoiiXsyv86EuYDVe8
TzjEbB94isLaLRbmUnDLsYlMSFfv5GCAD9X6g35+urVPClQM+pziZMWnpBbJPqcVyoF9LKX53IkS
wn04EirTlTxmrbA3ubA2q8g2uZbuXfDrMVZAutqBPg90Dq22kSDZdMjgukbNfYwC1uwXS8UFtjjj
apQHikOGXjJZ2wYJnOb252PCeabe8XSbezn8nrho5kyZEIfdFWDLzIBkE6ZE3CLeyuk9Aw+jy0D1
Ywm4CHg68A705g9Jx8WH4DFWrp+0tleViR5uDeCKpYyS6dTcLqLCOUtr9tjcZ66ZKDN4vBmHI9+j
8qybdytp2EX3kOZjxz3hzD0A22WeWW9QdCcuuzg9a69VR+vNkxmQnkyaFXeuxZPeA1H3HFsp2DKp
A0ix4ryZXUX5sK09n4CIQo9IGgn8RRy3a7AqqtSJZFxZwJEIA4Kz/+qBMaLQGdvq0HOc4jnclqNb
+tQDtK+3XEnyiyT7IZD8//zYnE1U2g5DOfF5xuUYtzvTvTMXJziXv+qRcI5ppdoP2BGRNsUhs2fJ
k3mwv+aQpuicYPk+MfYD3R+ytxauTryIsmXMNNkqBXkhrXOE0Y0jBCXilJfFOXgROi9nnNcLwgvu
JXNxwvrpNefUVP3x/ysqTOCLa/tD/Q+RcZyH9sIOOqvHva0LRCohpNqJLYCWc/5iFRbZBxB2TpBv
gZFZUNrCIGXQOlEfj7wm/RQ4VOUbcXMiU5LfuHVl9HMT/DVcl3Pbc2b8De/r29Y+XPqYAiVw06QE
StUV4Y8G3MX0MuFLxb9czPSlEhO5CKRqKUA9bu55m5CCb/3kmy88fdK6WlGWTec3AaaQidvhb2WU
AgGMXnV4ZRq7WNssIyreHtk4ojwtV9AHAEYVVyn65YXBB3UEEW0OWWS4kZ5jVd2WJCwheUTbDmJD
b4P07aHC1b8sYJqTupvfhoHf4AISX4ilYiXqIrWzefSQF6YE/YI0t9waXvVl/Fzc1zYNGBjrAlrw
recuxhZ1duqhDrGhcqdTmOC5yYIWSVpXXfrZYIGNJP0rmcb4R7KNcwH2zYLOZivm7dtngvUcbnXq
/gBnU+3Ue4LetBsH79li5abejyI3a156htRaHibp7zTMittAqhUugpXnOFOnwoBliAH/H/6ymZ4u
/77WdcHGO0pqwtcOFJIJnK+Q0iewztuvLo7aL0EMEQDSjMTWu1h67X+z4wVRO1vWczsijJwNPIgZ
jFIbGcZ9StpFhXczxRfrQ4s33xZeZ+zdj0BMkRVFxc/e9m1baM37f5oZf/QpwSLLwNVyqs/6EOcY
E/iBRKdOmhsSnFDCQB6epuGHZfCiftt7vRWnaten2cq+WIz+TRPbWQIiVtUJ3WB2mr2wbFbkEr0d
u/TD/aY6bfB3Hut8QykY1TjkTLThRsjl9lsIMjRfzuZXX/0RzmCcaGsFT8/NudfdB/dHbBvgDzZC
3ehZ/O+mJWozUVbpESXs6rIRu9AHRWiQHb2Cf+i64+GbqMyLcSiwc9ijfcxX+0GCguY5xL+SQaxK
J5u+iBZ2m/coqraaia3LrI8A9HuLSejThw6VEEiARtiGJNoeYHbphADPm8OZ0bSfvZ34+ZiFkmHP
zMUzxylGgMgDHXq4YFanhAcIMznoATKNBoWv/IOjuTvQD0tl449lXY4Mh5Bb6os95JHqOxVeiwZO
Bqg1yMheVmek/WPuTRmleFYU6d7NCI5SWvBHax+q1fvdU/8UrWbmZNa+/NQgOKX6hhvt2uP6EfLr
Mbhyrj6Vjz19ND1S2Uv2U04I+Lq4cDeNp4dQ8V0HMqDIGsUKPp/9I/EveWMWqz4W4wN/1KP+2lvU
/hDQQ/Eprw7JjG5c/SLEz4BQctZUj8Ug8cY1QG3nxsA+kAfjfQTxvMR/Kb2YzhkKWf9ihkcBBnyn
6Xf73y/GGX+v2HdUg6Naz7cZh+umM93M4S8IaJHIC0gw36lvfE0zYf+ZiqyEmfSwk+rD6SWdzcBx
W5P+LIebknBKEWvdATh0iCTCgkQL/cA6XYsBQ7nkhu8z1sTyzJcYR52c0LVuF4kK586ozwbrv6L1
6OBR72F80od2ma9zS3RoQX4aR8eo1bIrzAXCbRIoeR91Ujh6Z4C8wra4OdKvoH//iNeokyXj2/Tc
32jIncrfxjkl37HdlFcJKoBhewm1r46Xt6HRb5El2qL0Cql+oHXC/p7cknX6uAFegvus3yo0Lx/9
3XSqLC7DgMnozYwiyLtALEDCTuF3iKwJUnjdNCdHyJCddYzqeIsegXNVr0ulwfwwiKSzNd63qOeE
vhNkWJubLR3nW8du3ZVAcjjN0oNyqZZXLjeJ4WA59N/VKWdJw3Gqofx193gCDeXHxGGCeXmB5cHC
p9DZrofymmfnb9Jq/W7zdwhRGtWB3w+NHLvFafUIzsh59qqm9j25sIkR3mllUTA9K+MCIopJN/XQ
k9vur+kDtNlTvRNV71S7e/OKUAzx1OZs76scl6OUfCJM4rAzPj8H/k/9FkDtJwrwA4kulkBVqvu5
vNByowKkun2hqiUPMuUEmJANWMVYwx+CspHtWyOy+XqyZjDPc7RcOkKhdvaVDVpVS+ajO48KiEzG
McR7inln9LqNs4oqe0N+j4VutphzG9intFOvgKOfssUYIo5zdOKxHy2pNFUkm8FBFn4iGr99KDsH
12kTPDF14GRIeKY5Xp0hzE5nfH2X8Vo0kVGC+qOyVO6cpQ542Lsa8M/kjTWzArGeLPJbzeVU5hB6
z6q5hVRs4OG3nbJo5P9mjVE0T0Hn04YJazxdDnABsoZd8uOK1SyXJ6ZiLG4sfREReobRrN258oGT
5P00zN1lhk9Gz5HtGejRA3HsxSmjePFRdVS9q9l91KAYjs8k2gT/tFXM32iZNZivl8xeHoml9ZOc
qNJd48I6CDz48KUohteXH1ve4+nH8RT4m4Fb8hXlcZkQ/S8CcL+H+ItRg4HmKg3UvB5CiuXez/D+
xKtnLj8i0O8xorwqNEPZtGhskYOxoOX/2FN/kmKyp/4ESN4ZK9hqc0QGrPYjUckpso5zW0u3pBsD
JfWkBVZIMQPQjsuQ0YTbhGqdWCYDfymxNKDdzRxhBxEYvPE5J9quFmYxUga8V8J7YjyOGjZVP64W
j9DGwVHJo1jiOB6XVkt3mGV1uNg1JXke1Hy/EF3wHolUBmcmgLRB5hzFg40iO/7T65ayOgo3HWIs
+m+dmzDqMGjEg1z/Dn0U+71l8+1CtoOcUAQvFaI6f4qSU/XmUmW+1nIdwE4a5biq4Vp9W9B/LKh0
cs3E9tHrejUDeHWWeDZyZ19Yb3LzL/93fh/FuwAEfuKplL7JipHWs5RqA5xcVfRMPfqV4h5noPyV
eg7V9mmoDxNPfSf9ZVhZPJbLmjIXIbm9Y96uPKfCXDdOtJbD3c4RwfMB58vuOqsBNElDX/KQw8CR
pwYnKDoIa6L4f6YA3AjRn7nSlOjr+xpNyHex/25w2KmDOM3jBhiBfYyDSsVpPrkqeM/P2LGXJui4
tSc5dhQ0ZmxA2Y0fOfhBZWUYdqx7vzrtGmtSBbxdKHQBuwHDBy2TrNfqGubEl5r6EPWXULywxmMM
y0rVImO5oxP43rQ0UTRf5ukhAKVWVCBQmljqukReXnwlfyMBmMucVSsSwKY0vglOIP1oVp5HyELh
ndHHa4QelDUOUDzIdXn3upPvUgRQK9KiFuXI9IWks9x+T+jWMj0p2pO2V8fsfGNTK3ScAkk4O8Cd
MrkDn0IY0uYIxLZExq1OBfRUNXMhno2osXIFpBK3iJZJCbfn9N7wHF+ougAgLtvEa576YVCMjuQt
irV3AJtWm6+lDFYGXsW8pYrMOBJ9UTum8md+h1VOAeGif3RHMC667rt5dqpQVrYQR1GOvXmPVO72
e5QhGA1aTlBORN08nEtiA5q4v2iNJfMb/Rp5t6fyYeweeQDP2c+he6Blde3IrOO9o8fhkvoKLnpF
jLzRTY0YYCoOMWTCAvHlMJw0CpnfUMoLQPYTsp8lhjnkMX5h4Z0AvHsmrd/bH3OQVVgM/9pieCb8
TqREVm7vbudTsszPKVfaSzRMVAC48Kt2soHKShm8j1594Y3eWWbEHl6BIg+VWktn/k/YBh5/Bfkd
aCVMM/QypG4U80YBwQdzMi9Sx755dOjmi95xZ4nzv13+E5EUyBqw7Fp0P5JfJMEzExgHBLqfcO8y
Gl+dl/70S7x7BUuKrkIjDGbhAZnq8uKGhAb93Sn7qtJeRksW57za0lO5wCr2BO3us9RICFU4DmwL
CixOWXFUr++ctYVx8LG72qBoSNDeq/BtGRjX66kLc5C7S8iCQXSo0O4ByaAATcE4vmZ6UjrvZ/PT
amgnZIa33g8ejgiKmU7qrVMpoiEHllMWZBWnxNjSE1Tggtb3UqrIVhtnDsSo7xRJ5y1NLPeSmWhx
VVGrRmUmfQAeq5Xjs9TRKcJWS/CyvkF0c1jUAA2nal1z2Ieqz9w18An2qsNiL+5y6vlXfelnYUzM
vSymKHAT9uZOuPXadH0GjW22BOTldaIntVmY7iCBmuIaJtDefNanLFARy22X5ZMFuZG9xNBe8O6z
C9KLiPghQO/QRmUu+CGFikeSSiBCOa2dCKN8/zQHt269OlDGWtxChwNA6i9uknRfH3qiPQWxfHIa
3KPvS5J5S/pdv+eVS2kgw6ysVjbK0dpPe35Aou5bEl56hRX1Kcvdc3HG+Ua5mnExjLGV/CRTY4zy
SqGeKN6il8zrrb6DnREECB2IpIH7RkzWxDbE3EFK05Er4wTSMRW7x0ZmCKlY3yX5iW1+LoJkj4kb
2gGUSNGrphGKp0Q844AKXUS7p0180eg+t//24XAjvayrGweOuKyAaanq9kOETZIaIf+oB2++K+IB
y9OBS41AcUFXejAKNt+9YQKlVssvxXnOc6a0bfwbI4lWa6WLlT3THLKBAan4sJ5YMD5hh1kfkTn8
gfelMA2gfHp2WAHIXboDX6VnLWBz6f7gFlToQW+UaFWWOKqIiutFqzvTvBi4Xh0EO/8nI9T9j4Vh
UT44D/VyzNtYHewgk4NSgs4KNQ9r4uy+8Ytr2RaqsxOmjGT6VNEkUVVw/pbzXeO3GqtDJa8ZkPHQ
m2oKWgmG1sScDRpIuIxodR73n/6S0yisEeW3/FHyhdY1udGJmilvIPVhmSA4pRhBg4QRRyRBDyDb
CKbwEmrA/1IhbxgNMjutSCnSMbS/0IKwMP7MSKyi8/8ZMNH7LZUkcOub9YUMX3Sy0H6Zk8QM7uiM
f4WSirA40pqYjd0Q+W1Ppz9mjIciKkJdjsmReId/NMfKDO3ngHJ+KgmYmY+kckQ/IQp/3Zet8PTg
NseFKrrayQrpfzcAh60SMjy9YPBe2+1ucuPe8xT77XEERC1ycQbzjU5pjE3Gd4RlfmK5xsZmUmzo
YIDJwFjtvAfHKQntr4U7hSBWVQIJ9O1luUf0nAlBvodrAta4EToeBM3PJR2Ht5NmsGywA7HIrpFF
iOUTr8fxcoJEXDuAYnz/gYB6exm0C9SBgfC9DjB6nMUYoV2XNPuzqo5WeVWhIqK0yoGoY4dXzD+d
ERC6xO7HuabgvbGDs/ubZCe5YJomKm8vTiUG7RQjqWj31ajAUP6XiYXc/CU9lpqJaszCR0crSlyq
2YV7LSMGhmCXX+w8ypD0qHICa/9b05Vb4LRNGdXJt4j/nwDAzofDMlAqlJS3Cu79m7MEqkwXXTCg
pdQC2vV4JTjaPOCGu25yZ10nqICX+7266SJ9Vr8bQ6wDfXIFkXLI9rJGy4XW6UGcvl5eCaUguS1Y
qq0KV9KKLl0GbPO9cXERhoehWYXj8c0SIsDm62OWvGCjos98walstxf2D6LWqxsbpHk/6H0aanmm
Vi1aJDz4+rQSMmw5FuLI2ygq+rBzvTT4xL64yhnkcx3cRp2d4ehRNP0dOyRrpEXnhTI8r66o8FwX
QCxzx0N/eFpOfh2I0Wf+pgXbyqNULo8pIbijWVplWVhHD3KPcW2Ui6pVNsTWMohy3+lfrfqtpPQl
q6i0myk29d3S+NjRISwIgsphk+CgSmZbctJtqOknfKpXbsLU5E1/385vwdXFQidAY6VcnZRayZwb
n9kvvVpwGm71+9cXQfF3/bfEA9LsJ/dd7VHgliVGePyJ8U/SD0DDvK9sS+FYnMZwTycOGr/d1faQ
Dm7Mh+2e/ZQUQQN5k8SoL+nCUJBa9i4pPKJ2C/Ou4A+HAluy6E2BmIkaYXW7otCrrbu2wR+399Vr
QL15VtaporgP1ax9s/Fz731O5amaLzGcQvL6GLLBSLKSzFz3uMlYzxswW3SsUMifQ0tfujC0/xHQ
KveExW25L9MQE7rm1zqipPhBMytN31g2DuHraU26YF1HJr/a8hSy1aY0WuNcIoXmHFaG26C71YZs
sP1sjsGKqVVOaMHZkiVC6dn59g62Y0PsnL0vdEO7cNrj1TeFU5rWV2lSxCcvmsEqHt8LTJ2vuCaj
+aa4wGkKCzzkE23Kft87sLSdODL1vtZwwrfZ8IuqwsHj+PZyLyoSM3O7yZhkuyjPkwrARoLNSUU3
RnEh3eQPPe4P6Yo/1q610KFnGgpDUqZ5SQKZc4bVFIAbNWzNggEwVPAvTptCoaAD0Cf2WTL87WK1
AXPK4XDb2F7Obng+l0Vmfmh+CKu41Is9zuai03vaPLjwUjfyT/7QLY9ovwUe7hVN0mkOQusrKnuv
A/HLC0pxdAlKXKHjq2p/M5wF8rG/x2iqbwaLC6aXMAJ0JepA6t9jg8dHxUylSCvR3kOlz79Y27jI
Dp31mWkJNS4ED77XIF6Zl8o4awti5gMnOduxAH1+tAkxGmHRTfta+Zpnbu/MhrZQj0Sw/qB2Xhk6
WBL9P6Cm/D7GGh/Y2s7CO8rtLlE4xveN2C6ce/ZtUeaozARJlEkqgw5nJXKBjKAoD9O28s9fL5id
dbghtRuznYfSs6oSBs4o8Xm0liHl/TcDwscVousA0bO3SjDfURSjBi8gwCsJO19bmI3HRfA+WWf1
rOhNXhezuPQ1tPg+Br8rXMuGrJzbSL8cXwRAmZojR/N3llJA5zvqkt3EHvSsq0XoWEzijZ10xSdO
ckXoUsezDcXFLbQ+XyqrKLENhUdBGxqG3SnwdL7mJ6DY2K8p7BZYkN0t7qQ89g6RIhPSWxpDjmZH
8WkTIBFdUeKppYO+646c5P1gI+fqB+og3T7pURNRXdiHTLWezuP7Vv99Gq/Wb2lcoY7mevbS5xR8
gt+DQR7LQtB01/seAW3XwiKhOVzUzaCxITYU96FWZF6D/Jf/V1eLu66DAH0pu00+obV0RXF9EuCP
9k/M7WVx3ijzDi7VrqGzoMeRHnTi1hvplLDtaTbtb8OICCG8UFK2sz10JOvkDTqZvyB3EG1RedTL
lTRmzvUO1800oyjivLGxdNVY3Svp/HJjqZR+jgT8kI8dh9e+Y7xQflqfRdr03lDq21j1EEkQVcJn
vw0U+tDFE98j6rwecpUplLZZq6IzqPgmZF/RMTg9T54bTbdUOOk8uKASAarHsNqPOyiCQ3Zhvoys
WfPu8z7MNd58bXHr5KXEy9TJWBrcS6xPjc8B8v+7I1KpARuyiONA3/ptYD9NkFf/IEbJs1dtBh01
wRbz+qH/F06toFGgqBA+keEa/YqemoX9qNrzL0FFC4jsKRojGLY7xH46U+XQPIJe74ZLeq2pk2l4
asLYYGs4+WRoudumtLRdP9DOBgw9lFz6Zp119F3XooRMHmVd0gka9N/hH1BwKIA9sYAC/p6Y2ipE
KSJGgei3RxMyfbZwWjkiKVgIZPneuLSW3ziRiituETxufLEitfyfpyQwhPtZlYrlvLoH7r/+X0V6
++8+khgdeK31rP5Pweu+PGIFnMhf8sFgXn76cXFy2Y7itYhyypU2V+RYBGBVeT+C9xQF5nlE/Mzh
lYWhSO4qqF8O/YIHrn3Qp1Tm57hI3fuDl36w+DNtAr1aPH+zzBKGUcO0HIpiHzwNAHXZf3DZ3+9H
1/kTEnhZIlEESKBIPmRgtl3uAArYpBKSJUlArZNXRCvNxCznH3ZWXWhnkpfgjtRHy04BPGbHuiK6
/VgNqL5HE7cAar2iBEEb3XGf7q/kaZM+/ZVvdwrBoljnPW80n7I8cNwNVN+Of1yyVOcQr00wboRG
gZrAHqgjaTKsCYgycCcd9gwEKQPAUuz32blhb+9M+SpuB/AFrTIyofHRl989cvrD8kjkXjsUBkyU
ZcjSlr1wgC9QHfSyro2N/sdmYjURq7dSrIycdDGQS4dJiyhIoj5fy1fZe8DGPhtDzx9VgaOnrCkF
JBRnrhBPbLQxg+98cSCqvHuAVWVXYolSeDAL03h2AwH0ukAOQGVnT37XVig5+UeSAqwCu7cTFedH
zrtIzbEiGKcW6T+HsQuFvSvcnHVL+xOnq1Sfjkgff9Iil+1Q3H6MBE46Vyk1Xarps7ZbWFK0uSUj
F8rn5SZJYWxyfCUxOc2RGtLB+zeRnQPuoqcjbUAzKJmDYFUW8ik1Wsyefa0x+lVf/tJX+RmqzkF4
Ck32fvcDsz7FEb80Nmqaf2mlORz/S1hY685V5JT8G0srT//0Sch/5lqw6Xmds2KruDA0ZnQcQWZt
0K9vRUHX8YK2V9BQWPphwR5Md6kua2yec9h9ZgqPymZUoTAslBqlSS/v7LvGy/JXjFz6iZiqRcN9
MUiKmanm3neoZckTZCwwvvdD0rYOkG1irZKUeDh4ePF5PoaYw2uYlmxI7hW6qzu4ndc5iQKADA0L
1YwLQYHUpucZwdn+V36S6n8jaxRrAiYm0pAClKcX/6pjOUzvZnuNoZAqDRsz5n/XsCqnYlgC2xlB
NLoH9RHmJFd2D7oKsSF+mBKwhoJnNt0NjZFianNFRjpJ72JIzaBphiAvF9tPDD8f0tdDiyfGyMZJ
Atsr788KuS7Heo1zWs+CGf1lL3MjwxbLwrXBth4stqZwsvGffBUlBilRwytXUmj+KdMg66NqFNnZ
ZAOMQGX1ORkyYxFB005C+Uq+YjsT7iM5XHE1yopiZ+kK8z4r76avYsi1122WoItYa+Q5IW3ZE+aT
FsJUD9kDWn0mIBzbW7PhydZ7UBpgOn6v9dRaWlCoKKA8JQ/19i0m/k28Wek5BOsWLrCuR0uvICqW
qPteOW3NhxMGZNBnqGx1VCxM3Ty0jSRpokLFs4VqhzHgq24vkLpQUzIvn9dVgJCZY6nV1Q+Nl+em
+4YMTjzOTcUsHzn/J58c4RJdGtOgiMzid4Yw68cc9jvGxlppbmc/xdsElb4lTd3vPJTc/2rqYt1/
C+vLzXOdoTHtoql5yv+Youj7v0NxQS6KolydDdPH/sLW4Sw0sBD8ZP7iAj4vRLsStfKdKSY8QZTL
hjY+KYSx6Ed9NYAePfKgLEnx+O+SGEo4aEnWBDU6LlWqGdUa6kzZZMfQx9/TkCFI37Q3V4PW0jZi
HO1LbWTViYQigSejxMKUlIQ4gL5UNYFYFW2b+xc+TcdKbYID8h1Mx66LVIUnVZ95eqjw+DlQt+lG
pVQvvIclrTcuJ/9zfMVdzQ1C8owSsMKZgGGS2C1FQp5cOlcKjGWgK6Pac8ohrcwDTdN/n0ehPCzQ
y6amKqv2EeL20XlunwOLA8MBx8Z2sgNMYNKVJmOcQiVATCumN9nhi3FOwnDxoYMB1BkRRs3NdcqA
LuRQY61sFcNeAbgH94gXQ7+PQnjegW/ev9vuvmEmilVRjA92SPNeMndrbPkQiGcUpTFjXmIn3sBm
ZvckfyYWADfkyWo51GvKnlnSSv+JPjPYDgaTVcyVTZbQdRpZvzJw4Z/emJAoVISRWMoLJTCVgTXO
q+QsDpZvu6l3dLsm9p8tmcPPI/4UyKUcTClGoE/fpmFBU9s+/1WR3kEtHBrs3s6P5VtSnNHx4mLV
xWjd37IL1nFP7DXqncLBpSr1hFvJxaEtf4RhoymyKJQ9d3ql1euIRxrLmrElkQclW2Ck9bQoDO/L
qcsGqKeQAF9sek44cds2TP66Ns54fylrImT9v7aKjo5IVxGoI0Y/xSxZHvUe1ZN9IfUNFy0wQ+iP
0TdoB414ItkqdOYs/5heh2KwyPxN6CEwVHPIHDst0LhKovL7N21fHEP/N5Y+ihzPJtsUiGVXMDMt
+DyY4Rz7kxsKHpK0VThfg3CGq6zu0cULfFaf44mDF1ZnOBNQO/VyDyMWkucdHHtAzrVkChQzSKEz
G/+E/oyBxesYqXakoasLv/jU6nkdhlmoQzEh2PdrVOBaWHLrccDQyI4UX53SCv6biYt4o9N/21xo
fvwta3l/zXjdCRhFlfzbXQA9u6n5PcAIyuWraComrkGVj2s8fO3GMGCIzqo0twJlzzFye0FPVsPa
gdhxSnSIk+8jEO9LRGlWa/mB+4NiF0rWNI1zHTf6Nr3/T2mOJz+ATEblJrkQh/oPSghZ+P774a1z
coUufjt3MMUZ/3sABhIISmiTsmbJiLI3LB6OGfwU8Tb9vadYrpU//3wA5sZNmw2jHQbEwzuIVlgq
zksCBnDip5qDZcylwjQ+hCLAHrsrLrSP0sy54Fra6UNIED+JPmEowV4v0uMkTIIn8NZ1qaXzh/ms
baP09+1ydB1T1+sQwCfdDuZerZPMxe6bo/zk9pxYSsIE/1qfJZ4H/hQcUSK6LN273yJjlEJXm3XE
U8PY3KSEBZFXtAcv/sWIhMguPkO6iJZi/C+s/hgVLRzYq++eEavkEFxnUUAq9HmLGYgGVPDkx2mb
Pinb5YKivlYWrWFN7NHrbK5H8KfdlVw9/+7ly0XXxEJ2bHO6AO4rs+VYlUGGc1IS9M0R1itiFLt9
Yj+RenMLRwvXijxhrG6aDGhTGKy7LboJpqHRWk9Rxi7hVrwSAW0Xbru8gtUQH2zbthHxbvr0Z5B1
zhGWhGpYCI+AmKbegLzQfXauEacYRnR5jLaVl3yFL+rssi9JtPzXNSN5fkls5TNiubc6BppG8lNc
Q49aabDl/zJL1xLnea6aJbGB2buW25Rfu0HoznRJ6urdho1RXm8pbRB/JkAThN866luS1/gyE6xe
xiMQk9AjHF9hvwJaTzAjsrW+MRZZ1cmiWCnc5+xjfdLJ6HTyjbUVMdLPVQoHV/2jnwKt3bD5waaG
8ZyQd+fvrgK9Ay4M0h1PI37geIJ8dM0MFnDMIGsoBUYTRDbcGlrCbyNbgslEYIhIP41iZF/hjUwY
jKCSrl8tZgxsECav7PZT2Jd7p0D+TnsPrRaV6GW9twazDtfz4JqZnwzg+P5rNxj5dXN5Oznu9sxP
+vRRcIWN4Q5vYxvfFwCwJsl77nIORBvSvxaDCoC15MzkCjhEAj2eRJ77PscmJ3Hyo3Qafxb4hT8p
YE7rTadPcaJ8y6uRZhKWWNuru0YwhhYHn6b/4drLHCoEVXQvR9ZjHMlgoYfuPEtvEjgwwyfT+12N
otxOqUvcZ1WETM3zD0Y1Ya8QvRCdU1eZ6D1UJU3lshkukaaeFKzumoFgfCZJM6f/DLj1vzj6BKjY
SBvV+vFOwdXcoWq0CV9tpsVm96J8W6IO2ZU9JCe0jLorL1HqE7x8ouNhEOklrbML56v+IIsnFuZ6
ECCgXegEU4QT2p5p+669Tr9l2YA9VTU05TXWmVqGBSEAxwtlrWrYJY/VQREJ/PAEGf65Sc9HvPS4
4qv2p26Ady5ds/Z1cskGcQ/Dyw0l2Dc37MlSP0kydv5xPT6A1/wJCQqVNS34IRQAcOCZEqZQy9sr
+kKiqolfr7JZZ6OHEM8H91Rz52mxu6BDhHcpayM2DWz99W6bTh5/VzJHaGqVaNjmB0tSv4kPoeT1
T/1I0/XjCEwmoUu58OWLlNcjNcA1WsegUtBwQWSVcG6gnQ5/LKZEv1mNPKnU68zzrunMBEsXzhMX
RgFpG4Res1cx25fKNPICyaA3QTKxgo5bt0dOgB+hp4LV4EQ89b95eQy9ffhQmz9w9+f+0SQYxIKQ
/V5FOQxHkTzEG8AIWgvxOU1bCUhnc6IUgHJxlyVo46X8uV5Xn3ryx7f//6HlN8Rot62t4OYm5muF
225QOJv7fafINW8jvLSG1sRt3FsnqTURgrjd2Oec3+2RoYxQhZoOUuQRzjw4dxSOB5rPtTRvB5OH
nWJnrcG26Fs+zBo2ONFGWcmZ9w+YObkPxaHbtiDY3U0lXBiBHh1hGufJjGnP7chOB5Z0aX+0Et1w
BzKYCB7NNxcazun3vNv1t94WLnz6Wppu6ovRUeyJOANL1f11+R56qD2OTwTdQGLSq2OpzEg+buvj
aoCe7kDjAZxatBQfX062aVEpAgj8bU7XJwhWj4Ecte03UpxgMdvQ8hB2DvzlFaovX9S7RTeSap5w
y/5U6KhdbDGkvXQb8+sqKdueY7iVylkveJcpJodzNoDyFvqVqcprkuS7YYl/B3JV1vSPqc/1zrwM
SJqUaoSm3NqXdyx406/gR3EKyEC2E+fBVEPkh6kShVqvqAQ57M+yZl2skUNwOmz6ZIpe7mYP0bqz
M13pLopcnjOax9MK3vfaEGBs8helLgB8TP7VFacvKX/+/JrMY+QKg2uxzN+iRgQbQ5GsM6Ef1yVw
KGM5Z8HanJX20eN4sKeeYctAZinCzgaibUwodO096zhJ/zyuTxdmu3SE9dOJRorJVr8cG0SDCJeo
pYzWHdQqEAcpQgaT3vnpUWh7Hykz5u9HZHhuHp190MFF9Um2cbBh0dKx7AxvMx/vw5yn6uh+AhrR
Vdh4rzpjvZCilKa2vaGvD7ZnmZ8DyKH8yJZp+bLbeK9aXzsC91/0lYrvvv4LwG+pRZC+9SlRjnoK
ytuW5nW5YjFgayhF8n5jz/tWRxRxvizfA7T2+btEuMOS5ggBQ1apv0H+WLmYc3cHxNhB/TIHpNSo
QaD08fqY0IfMyZ4pflB0mcXS/WYiOBvmv6KJa8apHiCVV6btgJea4ccw+Ru95m6/SrN4rSXVAPwe
YCAkXNRcgezKIvRy4w7eWpE4K2nXbTbB4pdVii4kjIvEg03pVMoQKAtyF5KNjvyap1LYAfcI5E0D
GyEPLAjBWnLS7tjCUDinOdlva0fmcECWeXQdgZRHdQXZa4wWqUOwShCuOVDizwijZtjHqj5rntpm
eS8mglanQRrgJyrUrGRSjBZ+KkSx6EfI7UBoHWCsE7FshCjeYSRT6NHe2FXMJ36hslnN/FVYT/nL
EIhWEU/pVeJu8HXw5CSkFryNHUxbe5KoBmdFUEPRDYhSvFeReaNuTb/sjygmu/RYP0YLupJ/xPED
OGTGjmAfMcOzPyPEvyD8GyWCCgFY0XqhSyaxEUJTGAA/EXAKfz2Qi2LT6v885q+sHGJWSBO9Azqd
gTJJ5JKmlmmhjNajQGQXxbGoeThS/8Qx2Qw4AaN/ZWeKEj/mrUTe7ylHDzZVoLkXlzEe+A1iulP7
XzyXHbl/3uKQkVfR6iXC8gY01dfWYeTHCr43ioBel5KE+RP5Z+KZ4gHLgnQmTtDZZB+ZbSr+msFG
iZvNNZWiM0DN8jBsVeGocnglcJxuf7yvP40U56g2Hmk2hmqEv3pg0FQo0ApZKDm+FpF0+FxUwgRQ
aXNpFAdJaHZ9izgjMH8n/bylyz3l1Zn5R5QZyVi2V53JZVWaG031zbzWg+qP8uaVRejozfRIt5u4
yRBiuCPqI1uhEAXRRnN30SEx+c7nzSNhykdSx3gIbjrFkybHln/sxPvuDKXFH4nYpb/3gn/H69jO
bIXC6xVr+6SRAp+mMQKXA5j3Na9Z9VTBdHnjf8a6gTsE9VScLFWZkEPjonMJZh5TgXGFbHnk1gIb
SNaxCLcqJlqqvMcHkW2qXL7RqMziG1PtHqEfyStUS4+utM9CRxfKdj0fzW813WAAW58d7VPqL1W8
4Jh4YXpdddpCyV63gPhhKMm8/qUA6a0osYYuGhbEiV0cti2QV5A+fAGOu5ncI1AmARl0fDzfZXeJ
o9IWcYzL1baWWNaFZpiMCboTv2tWpsyjZ+58nYLf6k766ad1m9ipfupXdOtcb0De1bS43TVPvuqg
sepjkCZ+Ot/6uY0ZRkDCjoI0LbyR5CMwy9Vx/2Re7h6WqNbAVUkDzM3t3ab9wgUBDRSJCh/iUSJ4
1ZzDwnnLDZspvx3S5B2Ga6P0wlqM5PvHdTWcw82+xAS96zPXzRKJDr7zUosny0NYb2hqaLSqxJhj
4tu7IOiKyzrkp6yzMAjuOTAoYlxMGqrbIGMOUQjv6WsbzUNOocylaD89xjHP73oleUCZeCfUTOBn
uMYoC86a369czI5m5PVGqnXcgJc8Jvg7aCHgFA1bnPdI53YloU3rUAvY4DhU1gm+MmRONJFJCse/
NFY3j89rzWyVMdwh2Qg6ErjIpsBUzfBKuDCqVI8Ku3l/kYNEVTV9MK6bwfhdCpt2m8WcaxbVeWOR
h8hclcIbwqeVbyOEwhYtuM5DsDI8T3QeTmjHx2twD9IY1dre1BL7e5pYyP+aU27tspXFDznciOXf
Op1K2ndw8B5zk5WFu1JfuPmTbqrhEa9ArnesFJNw3/WTElLI5sxtBtnUFZBRo6dC4LFnbQVFZIQY
6hCcqNx4GBAaxdW/t19qlkTUIloL9FlLWlHCi2AgtiwgqFPd7eLMQGXpwOcnjG5QAqsxg0aUlEGa
t0AFViGb7NKZIR93R41DbZQq0z3JPF1xckw4id/Cgn9V7zW8QCYfYe8azV1Tu1nBtFoxhaoERN8Y
p3KWU7fsCQdBI3ee+o59+jhQbIxSQteCtbiNv23ltQNpylr74TFGXcq+Rovrj9GiiyZRJHsUn2FH
3bxz/6W0x+mMrzSFTyAdLPLj/xkRQfYiKGM0XHLTaNtVelBpi/BW6IErLPCsdxyDbbVa1GFW3kHW
R2uRnJdQv0mW0vyKfHzoRshb759Fis88MQ/MZuS5OJRqCuTyfFItjkOih56p7MzKeE1I/wPCGgOu
Mq1Z2GcX5MmfXue5pPFxYJWwSWZPzygEd2ZbJwvAn5UZo9ebGJPlov+NIBBK4YPyeUyb5heY59mC
iqgcqPSF9VAsUPW7PxGrmqjK9m6VT15DdrGNRPxroDgn0ktOFkzSBv7dCMVUSe2O3prXX200t7JV
nN6afNoy7OAgz4/09RHZQlHUIvSdahsYWJsJSIT5py0J+rPnNJp7R+j+qrLzfv8TbZSLvoXch2VZ
R62T9C9uHkku0ag730hDsUUfBk7/TRAonj2poBDFpcRQkF2vJOTyu1zJUUxcz5oJuc4Dvmt4WHL8
IkK5ZtVjn4yuySTeA9baCYOt4E4eA7igExJYd78gDOKfSl59WoKwnHjin5P+nSZQKL3zW7/SFT/j
UEc9D8c4YGROQxYzVxLdY95t9U5PUk6MLGGeBEb73OS2uOHZdDShLBKmXJ07bkyQ93UV+2b+vQ+n
eyCIv8vNj8WIeUNmk12x4wXB//5dRFTSzRLJ/cDgeXyDJSQa3YY+9kvx0Q8MJDKsiTb2CgBKslnE
cXgEqixhPBw+oXhf421cHbWhGn787L4mi4Rn3BDjolROzTQ35F8O1I6bIdwY2OiHgNZFXqMjXNwR
WUTm7yAJ/ZGNoQQS21jaMgJljCer6Dq1lm7ICfsLCpS8sb/eXkeU1jbu7UYAKiZ8Jo2DiwB74Fxe
DpFtkbBYjnvC4VtSmEDWmHouVI2LYCJOU/qwBLJXRBDdw4/gZEt/+Yp66wTut/66DWYL/BK0ketg
wmaXTIhkr7Nre+ka7lKK415mmUjIkuW/ZbMYf2GAIZ7B1suqEPssWVdpMqZVqIDE5lwe5sfjYF2p
zi9TsfPCEUg8tjFTMLeJ9uNC+4eUxEU0nc9p3knFtelitsbFd0oaBHRSNA2OxQho3VbG73rFzlMk
pBk7/UZaA//Tdbupi4VsnfzzvM1EVNsjAUvIukA6DDkTJ0NMJh+4f7t640FVO0iRG6Mx1iXz46Ub
uSEckY7Yb/AL24Xgp6x4wKWfVIj21eGihY7GFSUzpaBurW5dKH5gioHti07Mw1I7nVYGfYLBKIi9
SaproTbKWz5QNhOAhlMGqmp9swqdik29oJm44vpgAAancNQCDhfJfPsD8QL+Exr3k0wTahCKaQ02
yu9UlTFMrpke5qQz4Zm+BlHOFpN12d+UdHRvJ4rruTplCJP5Q8/ZK5fi1Y3+CURGqMH8dPJxjzuY
BINgt6155bprFn6LUPKkm8Gt9pTQip89HwMxyjn3oydfrXLqvKjJttzOP4Y4UGBXob4fJtDF4Pkm
l5CrzKZvZ/DjWrVNZJv2qF/bOgtC8zKUQDZYq1GT+ZXyi3JXw+9FDvBIUJANFJgF7MZ2bmp/o7tv
1R0Rr4HXz82yEIB6IzuijZ0p82YKukq92fUOw7cQKm7NVmcSOq3NT9QeO3hDLtZdDx5vYYYXR7b4
c+i4o4CiYSn1npQntPsKz1l564zTjSUwSZ9AK35VsSpfXoJY4K8IeK1xaTMzaRI5GUPP+bt3o1Ui
xx7nv1Jq0MmuuSrTsgYM4VY+bMx6zHqaVmprAE6IkeQOGIlHa9dbFMYpXlzORUG/m7eGP5Cf2pU5
2Okh6UERVn4zM4weFhrtVHfXNnP+MUq7fY/X5j0uNME1FAGNQoComHPTedEtvtOjtWX4PSXt/ocf
c2MTGh3VlJIt+wmIYkC7lt3TKQELTrwOGn1D+4Xj45h5Sp1Wzh5f/IDmx0+5c0VxW9FmflGYBnS3
ZFkRneaHNOPqdXkHP3vRiJi4S9yv+1XWBAioRLxwApzfIu/kY/Pj8Beb2Iv13oS1OtlgdX5yYS2q
dLzsZcovw6/yUdDenYZUwpnDCvqiIgm1dDp1H+6UbG86AMsVs3FZ/hO28SMymHWrXlvsMuBVLQsX
FeR+L6KNzkl1eDidSb6Mn9kbkcvBqhq1hihwB/qfcPtbvB8k3lgrKxMb4lDwnpaerggvybVokn1B
1lTwq3SJKtjZ3ViTfjurLysCYxhpqSxUJsd2o61H7AXQrVB6KYkVq5aPuQ36n/jeyms+Rf6EooQw
BZq/Md4EIcOpYaeFVx1GZYKFuMuWNzX4n+v/iVW7k/S+BBSbWTrIv+VVIeAhPlzvvVmNUJKbLR0z
lv+V6jpoC7+LcXd2CkSZNAvQJ/DHd9l7V4Jjm1ejDqkPX9EqMNEt72ubk+95CwE+T52GQnMiKqlb
VYoIW99Xu7Wj5t3q61/mL0LObHa7HAngSipZs/m0gBxlFOyPPPDPHiFKQwc1ZdOuPbPv1jh+YYTp
Q+ycV3ZGcT8OwHypeTNzVj2OIGEBL5TmNd2HnT9f6w/3U3e8knMcE0jBcD/i2Gf+FV0Sn7kY9VJA
B7ZCmAc+KnQl330A2Y3oXGdTpu1GhSxmIHDtnQytfBJJQLZx6YIhGE7imHbavp5uJzvR8P1W6s6Q
K75lOYJPOSsO3rFijLfWNeJNqpU1Wb2oRpZmF2WtwfVPatTaWhM9C6zzvk3AsuOmnlzafNPTUqtX
dbLmZ+ChMEUbB2/FnZq2SuTUydTnTO40xMQ1DK7t0PfhU89HH3jBsrvBXM2cbg4IqevpbmyZM7E5
aK6nfTXoFn/oet8a9wJ/A/QmMjwonI+g1GbdJikg2LJ6A9w7eTLH0TTuUwUCFe4rAxu0LPE07e52
XwAfD1xpuWf5rvH6P7ARQqwC9IFpl/SocJo4ue9tOkspO/HROI996hLQIBPnNHqqIw9t1UN6L/vJ
KzZ/A9vNxb/QC8//SmgJcigRQt3Im7i/jfMB0+y59wY/k9HpNYhGkB+pLf+p33bE3/b8BQl3baYZ
ffUgFPlBi4POfkt8JzTZVViS1vF4kRyOos3UGoWR3revS6w3jBXaVqgY6h7GEk5He1Uce/fuHdO7
dM8GSHOB/uZW2Rfdp+u9ZXhMahuTW1dLS3/vxpq1MYj6K7b2uXPhpwk0/PObQRpeHqfiEnMYDr+t
0JbkH4T4+JmEwz1mF7ldZDdnvRpqG2zi4CstvS5GnpPDSFwcbaQMWbORDakIYyN364OKqmxAM8VJ
8BjY9rRrR71DaKZkDLq6G+ZUv9MvHzor65kdPUz18KzJnoLb+rQvcglC4vntIBSq6bmaAOfPiLk0
FP8WPppOF0iVO956+k4Mv8CR5Y1VU93WrvD9O2ukYfzKKGgttPoZZ0t1K6ZQ9nrhJxhpJf1kHDw0
fJyIoxYZnMEm4NvbFqeSgGh484hdA5exsfCbvUQoGLYTEjTiMERRx04l7QWXCO9AHE95P388aXS/
P7kIQ7+kjiL5SX2wY2VcLy61LIuWypa0Iw+eiYk7TtvGz/22QYiFAb6Bs8BRsa+ziW9bJAmLQJ0U
BT8F60fLSNCVxN55i4u0CEFy1fxnP2qCYpIA1Uqu5IVmJBrlQxUURtu6hZLF/v0kBGoIIyNUQu8n
Qbx4M7heS8A1YzxwCy58tRVgMNIzsj3/vHCJrHD6nqRzjFmpR2YOD8+5D8hw56BYVn2cEnyttS2K
DFiMKjNohDq+v+q1XInqTHHqvwd7k8m9kfE9Vcrdxjff0v3RRy9fAI3+yxO/I09eaGL1Ha/n6HWJ
TP+ctZQf0abnZCHggVvyuSwEuBEmBNn+hKfca+P3APjE+Dyov+y/pmI37/yc18JsNqkImXcSv93c
UfGSuRh1R/K7O6xR7CLIhG0xx/dW3LIGRPYG2ArHNeAU1ktSfg1pAGbtmt4k57x/cWK8NgSojCF+
1WlU8YzeOQWosGpcUwUyP5qRw9nL3gAAiwwrAc6eACouPLIfGah1G7Iy2uskM59olAYdY6b73ZkM
Sy3GNmCkdHuIlclotLDudfDf0S++D1NRMBZihFchOl43BqKtjtp2/8ym/dK+O6NmQbpcU8VwplGv
cYqNqiaytpKUOVpepUX6xcMDkD8zKLvQxIw+mlO8K9d67YxY3B9cpBRBLlwQrBZZcgOq39MQFdJv
m5w7szE4ZHyvgPQ4K5i4h0g6UP2aLFOcxHtZAY4tFXHu/nTO/YO9102OFy0KIIp4hdsznuyJ9+qt
yIx21+bEB+xy6Q0MQ1lGcoyh8O4qTFbsNawrenS24cn5u7KZ3KGVMqaQ+uQeYsJF9cK+NjCQ20zk
ehcjYpNxgFmZzG6bK3NQI49l3e0c3iL7MznP7Dptz4843HVeWW9A8Xb4T1XsmYjpkRnY1spsouhU
+8aK4W4aO+ZOSdrxWd6kdX5KGrNt2YMuABJOUP2RPy8VCLNuyrbDxGWCz56z9JnrOJWkbQfE9nMW
Gl1oq8G/Z+501kxUwUxKpbaVfoQRwEHYWVEuNUGbm0s8oc517MJmE2dskv52kon9AwQG3s0KSzpT
oG/yK15WzWAmVj3Ka8u2Z3JxaTJ7PU2edIIAMpH+Hcs2zGwbLGoCN+w7LJgaDAyigRs+JShc2Ozm
wYdZZmbxhmanXP7zfZoUM8jsjsaE3BL7xK7zxm/N6CCvd8AdPV02V9kMWUEz+viKFnlvvh5vzC/f
44LjhqkMBQthU69jVhMMBztopDxylg/YM0hpo4v34ROaZBrT17bkTHD6XLiHiVnW8/IjZtahKax9
kY7jXmdtcGL7PUIfYHnjpFawwsaSyzJqI/7oMEzvIfRDIkze0+ZKp0esdyiQtxWnPaTpVrbbigte
BCHNzSj5wGVpyTKzHuVNExgWZj6tdzYkZYnmnsPBGQtQEOE9sifX54fDM+XtaOGtLpOknuFYUUFB
L0HRwa86aC+PBiR6W2rf8FqWeziWZ+fwBSqgZp28p8rqizgzWerjlj6I653JiEBhlprxTb20H6KC
1rAmP1hQekdxRBGql2oDycO/r7+QmwKIv/zswf+0KOSC0QXikKirpy69TA0SPUTwBdVCOp5F79Oj
xDOzVJqQ/0LtMCqgpTpHfbObra9S2tdosmsgwSSinEo8HddecHSv/IksTqcxBRAOBo7ebHi77T8B
PWZoWNPk4Fu48LzAcbNfXYxbibQkE5kPnVqD2KLrDdKopV1p2v51OoNLlAVTi8ODmcefGZRR6S4W
5pVqeu0rHmnk3kL7OMUt4LgXgxL7IZlwEgz/pt8WzJwsYBLRm5sUa6SbzuZ/1eA/6spAEiwOZPNM
TD2OzGCuYHWblY9yzw8IkXSoziDRo8P1f4sJU/vxBiY8hFVgSU5hiYSrmymmYFrDTJjjYDw6ubRX
3g49Da5qJ9qo9oPIt8IhyKWyAGMCDzyyzABfplYjn46dPOKm3IYYEwgMRWKPhi5pNvKJtlLIz1Er
fzO7FkdZRcGD+dXA6BxFryWfMP+/h61fgZgN6E4Am9JbwZbdMjWjTzDJZRH354nphM82qNPPJwrX
wCP/p1ceAc1yFTVRlJ31gLl+nMhYa02dkokUfL0p3HXg/YhGz8O9o3K/wguTZWV0v6eA6cLv8Tfc
1ujqYrrSriyefO56uLQJiCoZ+QJjxMrHeUZ8F+39cd3y5UiAKt7/jxUxG6w56gVSpFY80KrmnUAA
0L82MjZD2DTxTFcEpMQkMNRM/LsH0UzsGV0wOhGx525TYzJf9bYy38hH93DP+77tb6KUdjadO+jJ
HBmugAyOc2fxrDc4oO/DAKSROfS+aRFNSZFWMbqbt6xbB3LOW46MmnM4coF1WKjxmJc61ErC6Uyh
jEDhnTFdjn6Tok6qyyy3rRb1Pbe1XbRukvWfTTGzBi8MgBf2eUArvwO5ulHOIoxKVXwAOQjuxwPX
t0qLcp0cW3TNr2nQYVjYZOaTc+VlRS0i+y9J5NhGKj8fxl+9qyrvnbAZEot19tEhGQc1maQCp+1D
B7dt2Pjc61+tJgplggLOoau93fvlfmLLQ+8RR1jisKCHmvre67T5UHq42ClYIqMU7BjGTK6NbDM7
7LEsy5eoPassVzGTJwWsufM9+Ls7R7UKs3goaQb/ZxUeDedbNvwhg3VzvqDuF1VPGWtYS9Tv7f3Z
jRiQcu9YZ+li6cNbzFob+ETcRovHpNze79dzJllpQbFttS5q8BI88WhsCTgw08H1sYXwoeHsGf62
CsnYsCD48S1OJ6zSyBW8hbP+pRXH3vpVJq3F7HOWO2Xb8AHUpjKtrczIEBOYRk/zTvTGp0FxfJAm
+O79+VCHeIWvB2Ma64nn9eV3TuB3wZvtz6VhbJJcrNIOCMXo2Quyl/mqshIQ7sqNulpmqgCi84iC
GJenPWYMeIGubosvi9XuGOD6/ZkpoCXQOulz0RMG4N9bbeAu+1ieSAY4qSLRNUNbZ9RUDM8UDP+L
7a1uf9jTpfLHTQGlB2bGLp/xOCJ0DVjcBAJ5mabXJBLQN3fDcYufoZ30ug+gevyrVmF8XufBaZXA
uCOJx8qPChOc5YvSl+eKqacSzzwYjMHkT7wprDaVEMv/YnO4TN0C3AX2rRJZj45wN2RMisXvFmul
zA6+OlVEa9eemCyyH7lkF9AN4r56iByI3rUWH2kDSOxaElACyuyvHcINKdE0a7g7AeDFOhXBcNiC
2t3YuF65YTIvEYlXQ22d9qR8VLZcdnwU1owNnusx18G5CUXsHhsLPpEZA/vmE+pH3FdR+w3a4IU/
PXcA+RhLOMG65xj7+b7alj0ptQzW8EFP5sen6e+csmknU3xLJv/+RpAWO2Z9bJEvv58RZmbDXSHb
KdH3L8k3iKwzWtk/e/1z3/7AXg+nOAD9c2/31U4ImE46/xL5+pU3/fr5uskiDBRfp3uyUJdetwhK
gsLJ5cttfOVszTxFE9hK/hMsAxMzXpfXEyqkau3kLjm8dXtODLkAjiQcgxy/oQVFKsUFe4j6eJEw
yaDF2NMdLkCEfaPTCnEe4vj4VAuUANyF8z4duLFF0H3vIu40qTWB/Vljzlf8uoiTbnMaFVK9V6nv
lQPTzbAfenK2PXxBM4tgCM9Re0wVp1pc8D/lsAQAmu2pTZmusfXcu5mGO7o6XZJfoawRomRlui5S
iLeAhihQKDKo/f9gt9RbOIA/LEWZsGRyIlgPz3bwvZvDpLK1VV/4U7mEZHlpu8hDkVCX+mjVwPAU
qz9FZFj7BkHqtcik4hwmeJOKKLvracc7Aap0tBdrLIcVQHKDOiKL+efhDXnMhL96ogTzpcwX9hCX
YSIJ8wgcrrhp8vYF+QIq6yKyMDJiCI9LjOlflDOW+PsOPgxzwm1U54yKxuvp9sozuJPo2JbSw0pE
P6gjxfFTr0+21I2b4wSaI91L83Z1uyB3A5Sv1Gn8Fnx2cj+SlHHOmR+m8dCK85ch38aWXCa3smmG
SREAk7JKvOEQYdQCcUMzdR/P59vxNJ3fPKtbX7In9tFUWk+zEjcJS094dMBbCRXrdUvFLCUiIYO2
UWCwV76cHQViTbdauQMIf7uiZv0NgS1GpbFl5X/LPzd/dr8Zbk+lph4X7FPhYagmNIhoPoQiozUy
TmZ4LBwXE8wQcqnS34HUN6rCvFTK4ra9ffCjYnm45RG81Si9+jvBF5bI8X0d7r8LFAU/ZVWCseDI
DBgDwcQ0OdLcnGNTqw/rNqY2v1WYPgi6gDwJDG7+JsCVrZqriBxAus8Mw0yr5guxH3EQtwo2h4kO
d7/GH7ZOHpYXBDgnx3nmFTdcd7mZeMEo0NXdzOQ9B6KobrXXsv/bz7zpUaLa1+jk0YGeUvnOH5oo
CP0SeimBYjbypAv6yleGEIcJmcC0kIEfFyDgr9O2s0IBxC8cbhYL6mBbK9yq7ryqI9+f6dej5jan
cOWfvDoH0LTFdu3IxNsyDHduZ7ws+vFGVN3n1voGFd8qt0VoT5f4r3XV7A07lk+eIoHzOI3ncmNz
bGoe66qX6TP2KvRWoDzohD5j3LiauZBHrblHvdfxl7obu6R2h32B1g16Fyx+G8ugwYkffgHAnx20
vAEpO4vZ0N1eT2UMZUkaFrRfxhkx7wu/DbkeVhg6DXrO5FpI0Mwer93hW3xrW+AFNahM3hDooLWR
++2RXOj8yImdTAfXuVCc+Gs27ekZZ3xfB6ytPKMZZHHZ/iGnvEDg97YsjCN7qjjejjzeEU1JxRX3
ZYhFA2vRHi4A4Ifbjbll+jkPJNZMXWz2EgmcvvG1escAJ3VnMYAZV6kqAkYy2dDwPOe4zGnPfgPv
P/iSqggl2YQVIRY4DaFF8xPJN+BeoyfE0P9mG30Wmlrr3Ohhii2dy63w+/3co6OsOuNK8sOrAbAs
zs0SHY1qG5RzNryAkr9k6WNDVPJ/xixNLANQCvYGFoakOj9xoYtxUxIrFsjIuYr4ypN5bdq5hntc
PojiAoyw5LkfQJLkVcV3AmNAa/4RyUlQVrVOxCgkkmJyeMd8z6VlbfadRsYGFVplkHyPSS1/j7TF
xBEvYbxLM0TryKl6mNM13AB7CeZQ1nWOmAELV7GPA0RovSRRFyrTiOUrIYkOefuGkh/4ez4p5tQv
i7P22PvmeTHSf5hVcMPL8249+/uAiLOzopIJn2liy2TfRIzywmdwIAUhoINUvm6QJCYicxQLE5aj
eanH9Aa9V9Z32MFRlPX/P+E6GCWvVb0mY1kz2snFTPj98Wnq1HdxfPIDFz8J3UlkwtGUu8fVPvFK
j6FCaJVD4eFCZadySMsv5glVAbIJryEnv5AwRCnhQPhB+pw8JiTWxmp+gAIGZtKaNIQYOE+aXNYi
fb8WcjaeM6oojzlIpNlSoNzYUKutr63ceXmq12CBseS1JQTRTCODghG8DO37Nw4RHQizfyYd5P2+
Wd8LmtfAHtgrsqTolNwVI99vJ5aeuxD0gaSrID9VAy0lprSHQMyPLUnUK8Yn1MWgrt86TzP7anqu
tR8BOl4ayh37qJ8n20RK+S9a8ZJHimkBgl7qUEzJRZoC/2VJPHYwjY6vUpeMMhxur64xqGBqf1bz
j/6xaxYdzpFFWm4Kn/TON19FBSV6BaFF3v5aVdNRftKgXCNW4G2l26oVjMFNvY7KgkakJzeBKv4e
+QG0VZeov/3Ow6RdKwPjdisNh8Tc8IojEx40Dy5/4UiG7WGkKF158bgfCPEfdnvK8kLIgblC1MdR
4Qy1kony6Oaq8SMeHcHugu2pZyuzymGdlqDhA6fqZ2xLIogBM41xZwlTcwniTaoJ5c9QBwJt60C4
RDFJ7kTVzENtqA3bDDSzaeqMO/mBM0wxCH/i/ciG/cKxVno90C2PNfCSd8zS51EGhfgXEJZgi2cz
PzE2vAPWy5bXDoU6t65KtMncInPS0w+ajhTAWL4pjCKn1Ku1JHWSqb0CS59Q416lBLWLR1PG6H2n
VlzowZmnOBpvNRMQ0IkxACc8E4mV3mExDVVjnpocRJeFMo7KbsXgTYYO/cPOxk/DYIelWe7tyS4n
AdNT+fGpM7rReFZrSh/D7snuYCkXkbvv11YIfGsPYx2op5NYt7zz4bTF3ir3BKVQqB0zFRxUcRRd
WjrV6Ij28Bq5R/OjAWz4KVbMq73oB3nWxXLXr5iXETHJjU+da4TcyOihBCuYzGq0uVwiyyD72BK2
NqDCKpr5ZNNCkOyRIpAOxt4qZdnpgf3z7gBn3GSg19EfzZcolWr2W45TKxgVvCSsXUA7zIeKJd5A
JHU633O4m4LFDOJwC4T3PesobC4bzJpysOEfcvJagIU9CWaDFFCbdc7yKYHb5R6G9MUverXWjiSG
rN8StiVLKyjYc76K+G+PMlzqu/BfxPRye9XQ/uWOA3QSDSZwjyJCjPBIT48n4r1ruCEl06Sq6E0A
+kD2lk45YHPwqyRxDHnHpJs9+GiTJ2TvlRX3YINpLHjJF+jIu9O2ZupVD6vNn19yxsR3CjF7VjVm
Lgkm4epZdgUBRjy8vjH5SJ2ExOuxwdut1aO04sxPadxZvR24hhfNmQSlW1kDdMBIGElafvdSG0vS
7EAnCA7R9kYZlsMp/yvfz3SupXSWWRIQHABu7pQtPEM7pcU6DWpzxHZOwWIBwOk//Sofn7GJF/Gy
LsMlsJtqvLoEYajEQOjT+vPR4W5OuapdHRLlqubycOS1MR8HoT+Sfk/fqj1wefXAU8uc1Sf6I3J7
2Etnj7ipO+0ilWXp4Iux+8xRrNok1KBZ18gAmhMQkemKG0kfLlt04O4puhQLIuFGmM9su+cjc7Le
uK/JpzL9VeCWV/OfqESG9vsSLW80Dd6vdgPbOZR8R22fFPGaM5v9lWZHrW7G1pzYNuXkyMiOUp2f
91K+CqMw/RxTaBSQ6ZLBlQMCPiTvVmvBbKGiGhWkziUrulhyVXhtMhxtPfgzWwYpq9cypBhGLZO5
yDhU/2nCwA8DD3rwMwu0fb3l5RwQT59Myja6Q2VE4ssWCSeoYI3K9NXCmN7jbLePuMrZiVUJN+S3
GcX11PYMRQHL7atiTExEs0GRsiUgcR3Oe9KyPdEyIARcpo5toFfiZMhcPS6X6wre6CsouMK//GII
Wl34d9vwWbI2qeNBX6mAyZOG0E6JF0kkieXu+YorKHUA7suu3syl7Ukn7Lfv6K0LC+84UGetuHpE
FZE5GW23eeDOzGOpi0QwGCpBVzF8jWIpl6p9QvkWBjPd2I/f/cDorM3PfzNv2bAZGUfQaLFyw3Qi
DNoqS1t6R/CedhxJXjq08cHqpxh36pQqfxFO39150rCIs36z/AV+AD92XwFxfk5M/qO+bryoQF2V
KZqt7iB3NJvTTPMi5cODfVy0z/slC6Os6oKlGkLDT2USfM0IntKxepQz9CTlds095q+zSLpHA96w
0KYDi6UpNuCa+b8Jkr7SXeNYsFnZJ6+vZ8uVYJK5xTj+EsplDxj0zjNqw2L8g80khOTfi4X5i+9I
7lIjkAtvuYl+v6qqSWvUMr9CqGXhhqA5F1Kesy12AsdyjmXai9wLUg/uy/C6A2kj7dh6aaV31WR9
aPkANI9qbOE9Zl52O2euKHu9Z5oI8lwPaCgaRGvYrnVa5NMVaaKFzYTbTjFwl/NzyxKr2rc63KpO
bNg1dTBiFkMPfCfIQXKF2HFO5Ntroz1MYxC0G+5et3algGpU69XX7Auu2vBE/hLzxuVyw2XrD38U
27e+xIiFIEGc3tVEwrW2H+c1g8t7CCObBoDknm3n0RythBab6wxlJjt0ZN+W3DNqW8T3BgI40L5n
OxpSHSEPwuY5dlChLyI5xioHXnCZSGJDHE0CJktZevOSw95SZN/Ch6UVn5H5liL7wlKHS+qUOqnA
XzJi+GjRJocOzMsYOAsIdv0mymh+ge44OSSUhEqUFLEx2RugESKGDEyJXKroX2D5zwReF+4S48hu
COwD/VkmIm4KGepqYVNSX5jbqir5NaVLM0P9nAGHqfCySbZmstb7cURPlVJ+ZaO/Af7qfz4OZO09
VLELS3Bk/ReLf4mib/F19JKWX6ga3tI/XMI41vGKJsbOF7ejDMiURG/deM+5SDQjavKvb9mw4GtA
zB0KZxIDQKI8NhRfRCGWS8sPT2JOlFzKo1Mtz1s8+HnPj0GDV+1ZisYk+I8Ey5Sm1WKejFOKdQxB
81wR1ji8h0LUFWZtzdQhVkRcz1UgaZxF8k7EI0kpLfoAiikyXmM6QxUvYArDdfVGSo4+pGyTVyMd
jsC8JR5QT/Hl3sLWxCtajmZVJ5NJjMZ7gOpkD/RFQA2Agejs1rtSiV+Rw9yVhYhtpoNI+3HyoGCl
WEEGGsaNcoRce5cdHlOGoX+CNgiF1c3u5/ndYMZ61FVytldwfUI1zo981XI8+Ep2TPTvqkchdgS3
OIUHN9q9m3EVXLAr9sJZKosGkMGhy5Zlx3NT5KaLV8VcxHHBYElW7tJkCF7Gcl66fLRFGndHn4KS
DVmbxLqv/G+8duhduQ/UNuUiTrzo4T2vWjRHRYf41ma6siOborN63wbajyc/iqq5hoCfLKVyoOLD
O/ahdewfQZAS774i9AO7KnVh0VdbEJcDtF9QZdcMxtu1Z+Ougep/FYwNtjnms7t3DVWZuzt/IydB
6PvM2pL5ZWzjdqGw01l6fFC0dO7LGfVOQujSJguAUxcBZvquoFdeOVynN57EBTGtIixgIGRdsCy7
cA0IqXRZF4B/0zBpU+nLRBLWcwTB2MGxnq9J0HgWjQ3Gnp5NUtpla0/RqQnAZbcqw457On85WCay
1Q+7+w+1h+wTLS5lRiKkZwhPG/YitUQVF8xm/2n2bX8Er5T6cMCUyDzYxCCnBX6560Bh4wVF7+QE
1pLsGd7YjU9OiQRdhx2mTtqY52nQne3PoaQ58mHAcPNLuMERaLvMXkvkn5x4Uz06ZJjfPlcwaSMO
P9zeu/JjRz0Zgb/9hmvykdElnRv7dNaaNMKASuf3Uq8LpHj08M+9Gd0SNVqRKge5Ckh6x/SyjsHM
dxe/qRG53kWXlVgl9vjSWjZ/Cbc18nmk8ifqwdNW/AlUZon/Ax/HSaEknhgUOuIVhEJTOHEDCsuZ
I7LWsix3pp74vbrnqmCmdvpYsZnIeh/JXrYwerDy0a4eGEXxc5icaw2dQs7fTYDXVg9eXW7gWuGL
4zUZgb5IP+Xo56bm5HM2q3mpQo93ASa/OHlIWbm9oR+070/5C5viaMIRoaxfOw0jG4abCFH5Uu2v
/d8Ca1+kRZrGI8JUdsCQT4rRUFo6+P3wN57S/fN+vhCBhIR0ZHYLO8jqg/bq3lUra3SfvJWHPLtz
H1cfRCQaa0IslTKZnfDDxyZyHHwm7LUmccsHUuAYyeQ4P8fJ/ibI7YOm56kB70EXuzPgx+OdKKqr
xE+SVRzAetoaKZ76vK5bcimBTlVjLDNgMUKmykbc4U6129ECjDz1veikmAmUlwtcytWHID/YJbZe
PNf5Yt9U7tKNnDLiKZubAMTqGC2zGKydGL0tQOw0b3de7/28Y6tf/HqqC4Y9eo97GfgVeUBvuBdP
AFI3quDElYMBS0yXBnSJnVqYsIa5k3lcjndAo9Qyj/7XZNHvT/r2g0wS4UaC4bNAFNuGe/kr8KkX
Kwq9MAYLnbdzQoYki2NGSQKaGAB8ZIflwE5eREMlDBUpP97RBPSUzFnu3xNECtqZCSV20dBPsntF
JgM+goukCcJOkahToJSXq3uATQ49cQQdao4/4wFEEi+Vz+XkKl/1pC7ejv6P7qXn+wW8dSuWdrjR
svcw5yH8xePrJUI2K3GFQOPYmxcMWN6zGMVG7Mc2o8BBLbNJfEC7O8PhFMdypD5wa8sqoTMaoUUQ
9VDaWquS+jtH2g7h4FTUpM2JH2cqX3g3yGsCHatc1LVuQeP/JuYt1zx8uZNdFUx08s623OkD2HG8
Rt5otw6mRYXDYdkzXbhPNm0VEi+IzM0mBNs2mKC4woZkD+v17tMCIRpqaWwyPAfst2NYJzW98yVs
/HSape0tyj0RVroEt3sUIM63244SHxtSxInzrrvq4dA8NvdVZcJ5DXEHFcNIi0tuP2dIdzKhCj8x
fqXwoyGO010tkQlqn2VNYrgBvyvz08tjrm1fIXDL1xdZMBufYwwI1yx1zJu5RjkewQQ/jaDE3OI3
2gzINOIjjYbSXsw60SH/psr91qEOonApksfCNMX08RRbT8jQKKc81I1gzONYn1Pu03ioB02/aH3U
i3BP2Pj0gpzKIB2sFO12DoZCEk4J3XeILgvTVWUc8D4e/YV4XvepfXsHFKqRCw7VyqgBWibyNQgH
wVPube5RiW1/bkBsB0tjcw9qhLCKm2kE6g8iX/inFpiyTMqIEe06R+NcBqROj+Ikgb9zmDm1Fsie
No89TkwQ4Qi+liHyHgNrrDyAAkcUSlbhSDTqQWJQFllwKcAvk7pmNicIe5MOxTkPpniy2G+SgeE/
CEj6JWOj0IJ4Zl4qxEX57prfazv17Yq44oJX9xR8uOtsIhsLacE/qkUUBBbO4uxJLKjDL9lzE7xW
bcSs4yPHD2+GlFExuWUA90Dk5EBnyYZrDdy6beV9xYsLFMJN9GRrHZf2widvsSOin/kFckow1ZTM
FYIe23LQop4HUMEalE7qAmnqfQkiyOAh6hilsy0YZBlFxRW9hEVCFiO7VkQegNkYadFaF5Q5MYks
kDvYXEGVcUJj5AmGeR4ISvifcbLoQUqz+1hy9CCVfGi1PRKi0vXyYjIiXx1XBUYHe8P08Xb7TcxN
vTPCQ2gzLwl2pTi7J8+p+231ioIjli667v3nMXMcckb7KB9AW/oi3sNOBhMNsUfsM/ox3ZDpri2Y
ar8pOYUwo+uR2wUxLThxadJW5x9mYF77ZpdZz6AS+Gv5r/mRrJ6itaDBlcAnsUvVFyISLnUfgd5g
3JhIHSzgqE5h4I0BZQxn4+v8VkQRUlY0AeiIWjg7fFqr6qTn0BqeLB9FMicOAVtuc/f+iNe+k8Jy
THmrgeYSw7OJ+iVpdiEe7A+7yZ+0UjXwzYmyDOwFgLw5Rz+X1fqkOAMc19Nr1RyprnmNt5srOp7M
2Mi50rl8lsxh9Oy+jzFbabfEHL/AP0nKI9zplfweklQXhlvVh/SgLPJYWsEvaRD4C3e0LnQAI9qk
9xM8+8MKrQ/WysPeahM6fr7UzvyQ1kK15j1Al0nvFqK14PaJRAAGU+k7Il+V6UPpnUiDS/FVR7+r
AB82PjBGgGNZ3l7Afl4K07O+UYpTpDYVJnmshtPjY2NGgCdliscvWF3ZP64yX2ZVjdB4Q62m+NOs
dXEPrJktfubyILpxeKOXpGggMurMRNwNmGtN3yBCK/yP2Bdfy0lS5BiCIUOGrvHyvcpivp8Zj3cX
p66i5U9Il+vrT5+8O1LXzs3QC95WmfciM1XOuoMW7gwtEt/lMkSNlQvk8zwrgxSGFh5Fq341Pesf
oR3VXd4yhPkpjbUJILFniwN0Co1FnV9Plz03NA3XSW1zqRYz+IeP4+4LYFz3yyVWCGnannQjnrXO
QAQmqXtYJ1CuC+vlGrZ5SsION0QtnH36S5SDE/PXkY5OvEqnUNcbNgvAJhylADICpNae9OXb4Wdj
VB7ZG0XdQfREOXFbPf8/Ihk7Y7vGVdmk8kGDisJ9snus08l6SlUbIlMPWa6pa8tA7dq4h3Vuqeq9
nV7+Rlq9pbii3uTXta7yfmmZG2q2/is2JxHZJHGEU/h3G5lCcu0GCTOd3Lt92fzRzGkv82xBjfGn
mZKCHx1s0tHkO3XWIX08QHASQkJ4V+ftAvSQYy0pjMrLhxc+FXsz1oHKbqnWGf+FGIzU+LXTaYLq
qJK0oJD5vHu0MvqREsy9Hz4/+PRh5QsGU6t29/lPO2TX9EKkP/0yOtYfy4G92sDhaSJupfWsZWft
IU3jBtBheTF/wnzRdX/JNWh0Wp5vYxs+UhLLn7GOEVFnmrLReIkE+ftNpqk8wJZ2K4/WgwtemfrK
gQuXA1zYM2eTxnqWD2nsPxVPHJkvP79Q4DYkg8HJPMtombJ49Sjs03tpVdYaz0LS3SaeZojMJ5JE
/kLdY78OsY4Ma0ziQ1mtobkeQFvdfpqqCs1yxgRZ8nCu6zzAVkdST16Ba/zsOyGhrTpp+f/J8MfI
hu5RR6Ksen1NR24oq1r2y83VvbUZkRkrPs99ktwDJMaSIfWvmER5CYLTUxT3i5LpptJQ26bRR55/
siFW7R4cEOh6yMsURKtW3jcfSi07P937eRt2Q2uDh31T5X3Bs79dMdG+WCECDkwGrHcesoc2MQHB
1HhSVx8Ejdex/5Zo0duj8b9JYj8tMhiHrnlLTW/GQS38sLRTzQpu13W36DJxiCRuDs4jjxj68qDS
3BxYeKHur6gkkhQvjTb+ynEH7/1bDYZl/05aMeLeIqx8Mf6EoqHAO+Pgz9Y0MR8Racfda0bdPnHV
5s2dmf09kKOI0FxhZDrPd84aNIe1oJCMJv78mpgRuQKKitzn2DUOHG4dNb+UquSkXCoUXjar0j3+
UfwD0p9m+M6aoPmFWmjO+ejZDHC/13LDUoCNrvog6eDfrRN0DYV7xR2brx3RYBn54NV5xubBtCCD
7YTu07tGjv2lSy5IuZyIq6iyHS22G5GbvPTMaMAU2ExuD3ITIqn9sPrcJ+vELEdeCGtAs2iSGHv8
OmHEUcQwCI9wf7OKdNFEb9aDpCsFa33rQ0rflZRYrX9zgzyzCqiFRCow7LsAC3XzIlIi7nGHsPtb
BfoHndcZ9OVkE5bxLuTNoT4AeXmN95RATDRwHpwuBQLLOCOhcBAyJOwCKjeeLPFlxSyhdH0laLOG
nGtI6ZusCwzyTmWl5YkbV34LYCccB5Fru2mt89uLMEB8aZDKRu1vkVatQYBrTY251y1ooQjtLUiW
mKkYhR0ZiXVSOaRuKRTAvG5gc9/qBRUhft7y/3Ld6forloi2xjKx3dyK0epcnnImY42guV437YKT
VDASfWwFHhMUxp68VDGBdlHvP9uJpA8uncVPpLLSUbKek7dsGksai41vUSYB3RsfR61ZEB56PVxZ
MdOWJD0Vy/3xtI7MJUVUTH2q5r4SvLh37L1vqxah/j/lJPapcM7IHAt4hHohEGAKxfYwU2ZdNhYO
1b10K6/M05MvTkJvrlbzKidsgTh6zGHUW3QMkFgJeulkQZ5PF/5jgOfWTSdL11MkQCBi0GT59v9n
mmxu/BIey4Ik1fWevz6XdREj8nl0YVl8fcoHqREO6QT9EiAl4sTSp+TMFLnfshhejF6LfWL/MEvv
pmLl4fgR7dMSaILZfLF5e3Co9ZlhThpYAh74FyizQWEKF46KqfzXZOJHf+gIIggPdWjZBTSMOa3w
O1YRyDsBLU/w1xjzOgDhUqJSNFP8SJ9kBCxk4vTnhk/m0Ne2G5BFO0BDXDGu9Oc6rYEyB2mxdHNT
WGIrmn8iRanP34DRr+1UilnhWEWH0+YzxbVUtyVDumdunTWyZ6xNkIx4uwv5Qp+CzhOmWsT1UYiB
6rOjElTsr87rP1gMbD3V2PP37mcToPCfEUBYk732AASas7bh1WWm33FxGP3lfmxFUGQP/mP7QaHz
iFSDr1nqgugG9EaLiMEoJfK321+Ojpz8v+zxZQUAJRmdjBUxWOjmN+YX0u8mHlQJLGlA0fiZYrSd
a+yepcwoq7BFPHW4G1N6fyfJo7weYhGkRNi6nHonVBr61ne+75+WVxEVdsjioNT3uU6HyW43eHLp
dr1Msf5XseUVq3urXtjtgwlbm1+hExrIntlKaQ5cBN/6F8YQhxNK3w3JmxoK+gA/U8EI5/KEdVOz
fF7m9ykJX7ssWHNS+rNYUbxd1Zb8H3eFKqh4BSbdUhEE/gCt3zBAhZTiijkIjDYGMsc2aCmsFtC0
ByV/dgCaw1kNma8wHOQ/POl4l7qHyiMnoSVDnO0BAQUOzIq6J8eTU+ZgqLmCv38vu3yXE2Yk/6z8
01edavjov4UhVViT0KivkbpTP0PVR/Dt8YW5AwjF8PRR+ZBkyrnaxQSrKroicUZPlhljKS0v/eWH
8UOXEsOiYLhJTTjRyQcnWDjbS0Xak/XrOzMZrD0GFxURmeWVYMhiIzdv9XKrdhTTlqrefwzTC88Y
S34JjgFaKLZDWZb2LTxyqx8YgO1LnEandHrHT8UL2FkkKquls93mpq2bWhXiLyupSCuzXeZ33eWt
U3A5FOGI1Ui7cH5PzS+naG7Liaffx2ZmazKZA6G222gHurp5XDVgCJaQxI1tj2KNrtnKn/QZ1K7m
zSDiKswONbxybFxwsqslyQLEP8g3ZTGsS1JpX4CiRmfK8OCYHSJwrGeHoaDA/8NrkjQ+HDQ7L65Z
bgRNjRL3QZR/GBQLcLJGNc1X1KiCZP82VEXeX23lYuOo5JFUjnsTC1WUxnWEwLqL/Ph9yFqAD7DI
cuUo2Fsv42RX+NY2zqx9JKpZkxIieL+7aDtMcdVFx3Dqh+x4q8lsSZ+hAdv/rjGhiTfYktl0IQCD
8w7nH6qwtDE3z4H7efQ3GKER6KyFXYQ6VJYLcAopcqBCP12c4ps4tDuoUWLIPOwlyWky3Gi3kMEQ
+3azGADqEmt4fxq5VTeFyBaXxW2bjt70TGULgtm53H3NZ9gXClE5Jptq49QkJ1wtEKCz4kUWqpnL
K38hpoiUyQf1UClLu9+blsdEJOKc0iLx7vQ+ZiAr4X3EvLM7KW/GhW/vTH1E+zjH2XU0e5ohWptN
ISpbnzFGcsB4txvdlFBExMrJQ0LI/NntuasEisBpC4qhsUv2GNB2EHp5hM7qIBoyiovMknf2/QXw
fIFyJpHR6DKAeWj6/zJamaGKLEYxI1hyFEdCiKdYJ3SEZQr9FQQ84GwJesPQK0Kg+ZVTX5ONMrhq
m/vMn0wISAgFz/k70SMOmJyQDvGbvZinXDj00pwVaDODhHi8HG5HbBMz9vSDR66zNiAhZJQXtqub
i6TluiDGyCe4RZC7jjebUjmYjZJmxMA5RUin5OL6nLdkfkyswgtJo0vDbmP07YtrefyzvsN69sla
pD56GOKsdVwQP/5KUT/uJeooUKAr6Lhba4EZsi1gc+SR+EZBbebLs+aZfFV0h1W5eaIYRdyG0QZV
dC4GZMW0h0CXgJhY9voILXOBIyrY7OIPJyWV6XS89QlAlN585EwrjUPHaoUNOZvyRn/XS4G/wJZh
8m/Sz+WMaGvgtxkR7qCviAyrwGxwg02u09Ixyr3SUcn5Qh7fDhbrc5CXPOjdqHQjjuWrhmX3AkPZ
jRmtSaA+CLUbPQT570WNy+wG6ZSXDGJGP6H089TtW8UwO2LuYnHyRyhnlbYoK6Wfr8Wf+HP8Cl6z
IOiEjZdvJTMPJPzG0soEScKEBQ41ACpz57w35htLEMJl9eFMM1p7bjMQN/97Ee4UOBsOfVIiKIRz
fWZA3THqZP+/QIIxqT4AtLnjia9SJq1BC46YQlO8HmhfCLeKBZT3/Lfmo9KiqoFUpsMZbCR91tRD
SsIgtbZCdr82w5I5xJFLAaPoWb5hrCCWq7vFbm5Ukq/i3DGnSxAvXnCgOJAiMEKFcGgoW7K4QDTB
oW1sPspVPRqfg/yZB8KZpGEmUNmr2sjaSAr3aDXg1JJWrWMVq8bV3YczG14JuLYK5HXZYCJXnyGQ
QrMmOMIqWcKE5bQTQjrq1JSJEk2JYe6hlsO+JLsX2ZRx/vuI2RIRW6PiNtsZA7SB0068pFZskKRG
W4sirqzT1gWGQwjS8rj6bo1JtUNKOaTljKy4x6jRaYF6gvgKJaA85fOAnFbpsEe5hOmZZIRdkpHb
RrN0nqNM/rDTuC90DZGmzdnMaBxgslX6yd4BdxePJQYXhVCZPUwrJGxJqmdG2weqXaxb0aQk3Q2L
hPjx2CqzqT2SVABmhYvVNsCPZHXNajYnzxed9nSkHNQ1Q4SQtB5Wsc15dLfY8qhUzWitZ6bI5wtc
ORoDxrkWlJ8rOV0PI1t9nwVKKbnNHAD1i0fYHsI04hBg+G8khauwOB+14q1fe1lpfLL/J41h8nzk
kI/V6KOLZ2T1L24x42rKyLGzEZRLg7KeZD6mZOW1csWdvOOWAxOjWaUk47atX2p1H3AXqxmE3cWE
7iRAGqM3Y+5CNeRsgKvEznZL3zH5Per/hMS3rJi7Rz1hvw4UhxErgdilHxtzaCBqHRqa9dKbjgYn
ILgqP0DEOZdR8KFAsRB6ENzP0PIBqVWjUU0TYwyjuEFz60EFTt4BBzGiGbwoebRSVNecEGXfEibO
ekgtUzllxvjbq2f98IWmdidCojEG/042tkb00N+7pK1Q2Rj+ZSl/puZfywiShw6+CQybJ+SOZ2FT
Iuz6Xo+wkrvhjjS4/zpWvk0SFyUXR6kypBJbUNxFdidoEUTcfLoc3pnRHZAOrW7mFwr1feF5RCDc
Bi1Z2cNeaUJoSKoZWJ+pmXvRgsI9g33xXzt8FLuYcK+fxv2vQDgO6vXKd1lvMvd9YkWOyhCJsVVc
5xqEHUOBlin2mdQHSBiphvHAS/xzrVVMmwnnHoQuSfQRKwCtSuHl+OSMiuK8SKPygy8WM134W0mM
svTBBv7ReU3V7aTW2oBWZ3s/eZTfxEqf7kKQ1RJSOnnpm5xdXMiT95ETbZRHVBQ318RPGHSvV4/U
CvqY96ZQAhvL9LvzCtaHgR7IjYdazVZZwMIwN+vRkMDMn27g9ao7tKhSoVyuU7c9MGbQPUs+9yEE
UbapAJjiHQODwcFbe6aWgzazVeG6e6c4mLOpLJ1AfUPDa5Ly5cfHBxky+MNP/JayZcwJzgaijc8Z
p8ZD+V2/KA5VETNfV57CyFlon5PcNNb19BVpVVX78+7HkXj0rfD8QVdJjezIEhJnu3UkyviUZQMy
Qizx6Opg64vCrskkQn3A0sgJBNq64aVdiFcev0DpdNrzz/WoNB5zzxk8sDlos6qyZV3bG52FXlrY
OYxnJiU35y5ryL6WbNzfQmGzbhSsAvwJMYZE/GK2w3tYDZvl/cyXEtNu8YdNnu9CMpyrjk6rL4ek
zCdWtME7hH4f82s0fkaOLHvN054raaspHuyupzv2S8cvd3s5SdtMcJfOf3tPnY8i5jJKbEYNuNIj
P8FMTQUFdLojGplxfdNRlrjjucmt1ifpqV96Rvd2ytT5SCrzTuZrT3O2UXs69l5IkuVYeEFN7Xvg
Jw4X2BmbRYHwk7x3L+T1GkVNM5NPmot0AFi1XnePfz2ZQ8EmlP85NpXXtvNE0SAzfEkvp1dR7GoS
BSfMJrgeDE+dz6CjglPEQrZaOpl4oyoVO5ccovKy/biZ45X3vkl7FFxYS/QG5jVSCxowV2hwv5Sg
HJREPoZ9kkwnEkUb89mFqPE6ktsGzQp+Exr1Ql383etG1y7FMAiZBMbjkENNm512j98noA/6LdMw
q/iBso6V3c/BCjZ9mz1HWw+nkCZU6/5BCruLAByPCMPwrIiUaptvTqXMWrj3Mojjf9B5eS6iShxR
uh8okmmg5EF0u6FAK62gCmRcaYr2sYz3aAoxPYZYZpwL3J6puY8V774B4Dek9KRixwY9W/tBDBf5
xmLO4X1FcUf7bwe1Cv+iDYd/Qt5quhLj/GJjdNWt0uw0vDDxsI/xoarTKmNwONQkeoxTCiyyh0CN
aJmFGDPIHOBcWlhXaprS1jbgttzJ5d4ATUCF6hSV40I/u7HbI5cC8dqqdY9i0BcLlgNMCRlhjQ7m
57stUd1ice7rt3AQYcyAP5kos1ECZ69IKo651AK0F/klAIzTvHGrttP5webr8ue77u3ot7uLL8wT
qMBuAHvOu5TRwaSnw16tj6h5OTsHAwYVNEUhU+WLyGVHuPJlkfixYdOD9KTS0inuK1dydny2ziDF
LPciUksLgI5GWEWF1k2nuLbZ4zEx1uxSByW4h3VsZKUNzAN7E+h7jvu6yu26vp2nuTCob8e+wJ6n
qTvikcPjg9VNsS/fEGxbHl6hQOUY2jzGOKJdlfQAjTGx33CsRiFebiM5ooOT6BhQCQhz7qzeEbdG
c3veWcSqWXtL2vwU+U5soUsTqR1l4upFK0LtZbGQTQwo1NAZRF2RB5s2gwrfz2XKtiXiHaHxSZz6
H3oyme2qdLfv/Ae1AYIXlHMZmN2IMkaf/LEmMeW6+OK+0ogRi4at94Nc223CPVaCVkYvADesp7Ge
u8KZLHo5f3H5BYrqcX/NFpON1gts+u6vz/VnA5pZ+oN2+DFGY63Osr1Jm9fNfgzwdWeiPnfo9FMm
d24ZCIvdeLtBHw6Xs5XDXdlCLzucZiXmA+Y28IG1xzN3rN8JGghKHc29dy3iTW8KQundRdE47W8T
D0nDGK36PSpGZjeSQYJk0BgeyVYGMXYnCz6w4as7xJR3spoJ5lu+n5xspR8gQ8yyLtHTNpwdevO1
PFRYC8sTrWD9vd8tcIX04o6Uh91fYT5gBWri5r41RDxMLHUzYXqkb503xU2gsg+CK+Ho5zWWDk9Q
PBV5iiPnPaEOdLmAa4deQTPZ/wMgDD07EnE05TJr8XPpIjZXtsfZPzSrDVEy+MMC0gWzI0aKoXRW
Qqwv70jQ6kogOSG8GYz4pzvdWHlSwWzfGNFIwedd9aKK5STVZmpezfq5MrosxwHjW+5PUbTAG/fg
z4siOPc8Wddc4OhuDdqLzGyzI7GIZpPa9ngdwb6z8kM0dMsVpjVuNyBryeDUH7/g2HG8vEe49R2a
Npg3wrskiV4azhE96HxZrcAMkNOrjddRUXxWTFdrFjq82/qpbrWAHgjAh2k2p8saYHT8B1PbmOpy
OpPGWsKmAIdEzuLsT71siwSPvL5oooYY6vDAjF8nDc74CwitV/bvtqxWjAs4SZvGMsEa2X3OEYAA
fO8UqY19Emx+umQotVbuLSheUAQT5jyCMvcjwquZyGNd9+L0k3ueSk8PPxsQbfq9qapfd218t6I1
VjKJYcq+F8OxhpckAYkx2d4dwprN5aLOI7Lkxpkd88bwNXFEE31Na3nrMEhSqqyhmEdXrJX+ToNs
ziATOszDd7GwogWQaIegcoO/2/edyXY7V/jMmGu02uXJ4WKvvmeJvylQV0/uZupkzpLf6eOBa5O9
vnAwLHq9gukv9piUDR1u9sXqYQM5N67UNUv5Zg1di90v9iF3qHFnjYB9qyvcTvqfq0jqv5uBRbV0
E3cgRvgUrq3qQzqEag8y71CcnnsrCUN6uhf8xHKZq+ZVqQD5zKRksAnJS0YUd2ZCfPKPqOQ2DscT
DM/RoYgadZDt24KkKK4H5SuKHfpj8TIbpBRAzpvqaBEMxM+7sHq5FWZcaPZeQZb/iFugCfifSiWQ
UkietekwvjpMDmJ/B64VxasGYUrfnsdl5Qx50ggmJScQ0cp7wpmQ4MhVtwPa9AQgOFMmUgTsiCu8
xunHIoQaLEUqbsc4Pe4CxctyE2yPy0jmHW756IM/7dPeDMfumlmVt1lfKugE5/5NmeR7yM/9HCDq
J0SbvLj38oDTJzf/OTNI4DAaZY426lqvs/AHy5+ZfaKeBJroPEF18dM4/UfmDy+KIPHpIqTXyaJL
/VHL/eE1Bpe7nqrZMgE2p9nemQpGPrUc8h+9L8Lcz9A2djePgQae/b86jFUyY90CQU6D7U4PdxcK
qorLfrc5t3mMt8HtIvQYmoJiD4BX2lnv1v/SxjL/AMdWoYPEF5sr2s0hZVT+RIofALUdbJlavaCC
ntnp81UoO5Zb9812GXbM+5xNKuyaI0CT4kHZDiAlhJpMSsOE0zLaw0IVqgq6D12zU+br6SBUd0M5
4ljdKwT+U9FRRB2UaDGBpJco0KOLRiPNisUEFky6yEZGvZgp/W5VsSNmxXhXJFKI2kYvHxoIe+ju
V7XixtNxlwT+mLp46jeq4DbdDzumRL8Zo/btka9NjZj6vZq7BwstebUxnfV5VEk/97rMWJAHO5t1
+0QnpdBFmrtBqrKBvjfEOfqAKbv3kyv6CnmwkAtY6mchjkh6YoV8i0d5mcZNDSg3yf5x86lR4R29
CPzIewZQRYTUXAmgPYNOMB5rQaNzqAvNP0JelihjrSUvwaWYUkaHg+A/kFR+omBZLJWIWJt07dwg
24EjecSRtuJo1PGrK2xxj8DXgZliViKUvalTzTAu/inxzb7liFhPvDM1V8zMAHPZvXAGT1i/qinZ
XYPXLD641J4TleaHsnPdvo7uKbLk3fDF336pBOycD3mg1S61P7+8X00Cw9HHQIyvJq4VMrfHn45/
mgaUWKgv7JSLWiZxMtgWh3Y2LwwWY2q2OkA1ueaXkvRVij5HYsYGYx/3X/NsBwp8kDC4/5yX5ZTF
MDVb8CDv9qDSDk7e+uarZgSGGCMmd1Sgy5Xb+xGp/XCKTf2ys8Pwz6QP/0ql7sepntyYNc8XOFzO
PGh2C90pf79PLYahXimnxqq2tkmA/DemVyIRndldrAzRs04maEseDstrDvWVUD4Ci+sJxB3Dn18T
tXwhQAf8ZUh3fzcfwXzy4wbHcSmS0tcI+NWEcmvuj34BYpOkeuxmyOnkDZqOkpPOSAPqNVfyU0nb
GJv2IeQlbb+wCksDgcEGZMuX9mrKWeASbphNZuIQdM4y3fSetkYHNYt+MPfJ1IMSK1TWa8rXN6Cc
o+vIiVaGxPb0cDGaxLadbk9+fpEqecPPBku3Xn1F86Gs938lK3tsFPi4kJ+9J7okk7wtdfMnr8V0
EGjoRwgzvnSXPFsIYI2+EtDZD+lSkRAyQu7VQ0WR8FW8S9A+FiNJNzOTnfxUwyip7nWsR3B2/6Xr
Zrv6umnVRSyj1SXJgBa78+hilJsvCUSasJfskf+1Z5DQON4ozWrs7pC8rqm5TYda6JMFxn84BkGQ
XMtHXOHosBNbKDTX9mjjpKMMMIs3JTVDizhNifC7dwuZFFo4AEsbsKOVVFMPjGLX/Vj9XS6mCE8B
iYP4E5L3p2hqTC3lDPLuhw9/yuRi6WqhTNhoL9GHJyGTIjnEcu0ySoDEm+A0AjudquJBRxBPCIi1
OO3hc2S/1eB2jU656xGcVPHyjqnGpooYdnaTcumipP1EoiWDM/Kzge+9VqddFFr/w9TtgyV4MkpN
35AehXV2U3q+poQ953z49hRD0+FL61oQQTx38SnPH9zGN0JRiZeojs26R/neG4uTwWd8Soa8X2lt
wNvtAfOm9ZyWYwS9sjrWyvHhUgd9vNf+8E6diIUwJDQiI+b9BHiQi28/qVFGQ1m+oRKuKCze0Hyr
AfIeUitOIS6wHH8tD1c7DoQu+tz8Q5gpP/ZAEWPKnEN0ZOfwW0GFG0sCX3wAHszVdusxZCTiexjy
XnzNQyZxE7tocJumr75WFNlpq6f/tGGqJnXYlxwzb1fdVqIrrv5lLr2Wupfou8OiwFp29wb4Nxii
wMUSq2EGGGbJLxH0h+/cy7INzCar2wCsQgf/5uMhH9yIe0zmcQdoBWSNdwNUBcu0pWSeEvf2Q5Ro
XjXjAaX/kyvkl0tqQJK4EeNhP6nR8qTTsIybog7eEmR9byJFgHWnkrElULLJG5clN5MdMpgD1asV
g9kKrXxoJPOwAUnjk4foQ787oUkrnRNerPJrect08/rLJTDxuXipUJS+z1rAD8bjVdIMEl50P9m7
KJtkI6B61+YnX56tF6iG6kRiGIxbal/98RqYNt5beveVaS3byu3Yr58OQwUu6DFAZ4FW2T/+y0Pu
/iGiBhtQCK5XugWPUxPJRigLG0277+467rRiYwJdoms+AMQvdKRIKpgSbREjAmns14Ra9BIuaYF9
BqCqvZJ9D/ClRj6j1o8WkHhvzSGu/RGEcY2H4ZvRvmrA60yWA7WVcN1m5S1EhaQ3EdfdjTs2f2Lm
B17LObhHIyKO6ZUfWAsrWAVh0wc6DqWUpac0b9dFHNCAjz8+wp+e2vuz9EhDV6lF5YgzR3qiTCYQ
IFoLwQdhim/XSxkCswXdWFS3bWNWEczRARAt9UwFJI5WRcsmXPZsyrGq7ADn5g8XbDddGvDAHUoR
grMeGjeG17nGdudpuhhzvT4z4Y85mAh+bgPmHCOBFf9RFxkrTZ0v/8fGwb8vJ7mEJIp6+xjOFWvH
j0LUcK5LAi/2OBb6B8ntCx9fvv1OAgksUy3ghrMSU8CjMv3ZXCUFGqozmqNJ4cQ9d6imoc4xuRSa
5jSd1egbKC6A1/3IQuZ/hIUcDcvmoeqyjRbedW/gXvh/DyjpCntMMptGEVjmRUScIaARt/DzsIYC
3FtVxm+OBR5hCbU3gN2O+Bb0N9mTTtrBryRjDBHEMF6n1F1tZqGy/STCmKzKP2q7NaSQX8DoMvDz
U64jAmE02lXADYdwqQsOnVvLdikPD4/cfSxcOqTNI1wn/YmjdKE474JhIzhnIDfBzl6sLmYG4ofG
HDUz+E9SxvnCxwFihXIi/Q8T/8G81pVqqPxNHG0r0FiW0rHG9VE41NPuMNyDcnFKhnQlq8LoveAt
2UovfKXmI9LJSjkINtZICtzq9plnfJqHMxkJMFaQeU+dzDumlfuiq5Cov+biXGtEnUE8JQrkYLVE
niAsuRUORdLw0VozWe64xf15LhGGk6yI1P2Z3tUB2pyYZCCq8dG95GMu4/gY2r/IoQDOFxlpQeHO
mH428Ix2qzvSSk9gGEyaRGet37athJ3v+BH5m9SDKhrfewM3+pw059NBe1Y72yOncnIoqb89VSx8
5rrbEjJKZ/JsimU38D/gpbtDIRQ5Y3FG5RdkzJ5AE2wboTRLOWzxcCspB64nzva3RElofKl7Kf+Z
4ovzsCNWvHrH+N/7Q+wx3hilpMPBX0jElkpJrSfAJCvDbPL5dWXtdAjC21XCgx8lteoY8E429ONo
BNsIx/P1pLD39ZlTIMniwxvHL8efLXWCaE6RChWJ83/TehOKEVCyMJwbf7FR0E0M814sUWJxn7Lc
4Cym5dDD1Skb4uglWyncsg/njfGoUGWW7bdOOsLOAyARmO0PoijRey51oKtoQ8azwNiq0AeLR2ep
vrr1oweeBNyBgVdYvmJ7FbeSZC+oqFXUklGg6VFN0nBBODTxDv2fUJbdtdoJW6WLb1ncgT/vaTh6
cPHqY4Kin/G9xDdZxRjQO4S0yo0Nu9WgHSyfMajHjp1nqXCNuU9SX/LuoV9RRovrQG9FFJ2mbcQZ
CpBhg5IQpCPiWOuCsGb3c3Pm7dSrTOMnfYfGVjyEzncCSZFrtJiwTnlF4hkgoXaxwXOw+w5GthrB
P7qd6LPQJXMEi0RxNdhcf5gGAL3gwFgQDnramaa+67AdWAsuWZkHMMomCOgh3aeS8a2yC7nUJ33u
8byW8MzF83mC4430S+h3dNjRxqdXDvnzXN3Pl7QgIvhn1WAyY7OEGNGAwpPb/8GhQcsVez6IdbV4
RBYJrpDs7zZFnLKu4i5D5n/sw+oQwSmSCgFAnivtKramgt4wDzqn9UoOkixIRr56zkzl7kdHZSH+
f5+xkk3/E3pPr5N8D9esW507ykpaAhQslOS5y5K/x6btMrUYL0Zu5a9cVrO2rLSuMK7j2bMDOpDa
4ZizAKsSdDLajrABzvGa7Sx6XE+XMupt08VMV0M0RW6NrMqUsd4aUUSoroTvF02mXT1X0jzjgolw
vX5JHsXfiaDHGrRMdmTfzttdodN56tcgAApb7dioulQqIU86FT+iWHGk/YJM+djm8RJzBx5vxLbF
v/HEEg+VfqLerRaPXp/xXBi4s1JFGyF/y76Qz1ur6B4lr7pbUrgP0JEdCaK8Tw+0wsUX/TYKo82+
UbMNszOj+tuvM8cVocyBI2IyT9bYy0D33NTs5IXbRBADEz4VvL4la6vy59HRFwT4UY++lt047dJ/
WokKpMYmy6BfS49sScOkQmiLQTbw324cgsUPWHLec7MP5iChC9BMkD+Wx3pWO5dl1uqfbwbhRH7D
KfzcewKCeC7VUg4kOw1gTYwmRYcqFqNTLrqZU9EPlfmUTavZdS0XFJ0YypxGDQAlfLs4VlIEL7+9
ybQogKO2hwPym7tZFpJvxGSGGu9q7yRiuEx3OfjgRgDkpi+cWQBbe+NpK7hF/YCyV6TdkAuDoZ8S
ce2CjAp2E0gZmTu3xr2X2unODGogkiYuEGWpXdwP4/ed6YN9AdsJtiIcds+XSuYs8VoKC87g84Ym
RWjs/UV+jNL10/1EDX+/P21zdImLu3+T1TQYq7Zqx9gfUghzb32cvdtvaBXlDnBG7fRyrgiBIrWW
ffx93riCxvoinMH/Td22VRGEOBc8olUTIry9Z2oeK86sYVux2XCHggtKDwbnjwKk80rYuDGq8FG8
/+fwdZcAHFDwm1mtZGMgGFn5poIZQicujODZntaYWcJznN0BLePm94xheEyQmZuE3Ll7pVjwdTWF
gN3Pnq0uRWhcrLpQ4JuIZP2CvLgqIELuSlTppeEYFfVACQAQgMRSVoJrwPo+rFM9yv3DwMpqTIfx
piHVd4OchyO67PDcO79kQcwgaolmiG/k97w6VBFOHw76mkBT9wyaScBslWWSmpVWMH0IVMhTRDIw
oS67vXNa8nRXQ9npnSWFFldETBy4+l4/1eC5TcNQ2d6XhVnjy9xgReApz+A5CAZYYVjsjT0C0T5/
995qVYic0HZ4ay7NxysFeeVnXQTlfGx2vqv3NFPzxeDDaT8WNGXmORFdNeN5UnEKzHfbLMOQhbhD
3jdMNYnceUoyvUSDfTpIybKvcxqEfsTuOT9b02UBmOP8vZeQI9FTjpTqRWCRjJ45RmGyKH/+mou4
WtNqNKulOW8zhiFAZ1y0L7oN86w/H76IGxPAAv9rFucxnmiqmoVEKo6PA4gc8rBZiR8XUmSCSbrE
eRf/QSADVCJiYRcsA9u9Fhk10zjWdwaIWe9q5ZttzgR5OLeAEiCD69fAbANjV7k0PC2txzxlbSHo
45/Z0s7fSRzVzmWimSUgMcDV6UHjDX8dG4vPMLVmOqkYPi4kFAINJ0R/ZLWjugaboV6XI2Zh1yAb
ym5SxvH3yBuXPqu1WhUYnVlKAkvTIVq8w3673LYZXbQIlTfvTi6qEZgecHDx0W/GqRx1bsyPPu/K
BCOSWJVY9ckCtX43Px8GHzVsNrNiK+RQvoAKCVNfhahOAO8SkNfM/EB9rzIvsszDc578ep+In41S
mABXQZ9U4FccBQDIA7cxqk9QrCDcJuwd8jKHP9jVzeXv7xDL8y3JmbzwXeL+3aaAsN1tSjvhw4p7
pvizUzPyhuaArYCI96jLOQH2FPw8cU0FmPeDebh9UmbaLUpvp/Btf53qCJot0LN/9si1bLhfUjVF
XFoYu0q96RDS7NYL1sIHhXraNS3odbu0/j9Ex6q8oMXMpH0W20jXZfHvB+Dt5HPOjTexeDZ8YUFX
BOIGR9veuOjBs0s0MG0ZPZio2qoBo9W6EitbvjjjsKrYYwv4HdaDbWwQuQldTEvXEEJCOrzMEHg7
NEmyVCc2NcRzfiBw+vSywfx4zi4UkmZi+eLSuyn75eI8b5+AG8ixcQLJRVrYVYpX8MabAsd+ToKu
EO5ctWP7Y9rBftKhoaZ6GfyE5dBa+nN0i6po2CXn3Pv9c4ggEkl+cfY5fw5zeI9fpoYG6LMeKF90
Vqn+8dcg04XfXk5GOYH1u4WiQf4D5n5scSfzK3PgSRGgZDK5dj/a9lE8Jrq9jgXRXDdwkA3HKwTq
MaP50ETjHuLIFlB3We794vZwQ5L0Uc5QxoiGHymvbg+032n+TEYlsozZlfMYWDWr1uewYTvdWJHu
NC0j9F8DJd4HaUlRf6uCnG8747nbf0dxbNXF4FYc6zoGwogkEFfnj/ivnxMeMnqvOo7BPd+YNhqX
ubyMxZJEHD0QfsFxgSe5zgBRoEum9Nf9hK/MEUfgwDaheXBGXZFgexECRG4DLCgJaZatdqbHgm36
K0XYgZ+ffY1cX4BxOHS1D9nY8e9/neQngE5VReiES7MPzkgL2L5hEGSIZ6zWDfg6WgUe3ACRcPQd
oK/9RRmhWX134HjGGTNOF4Dr4kc/1TOPWYPDuertm0xFFEcx/zHHj8vwPe4IrXDaBpcQQlsjxjwb
VpKXrpLU73GKfZ4SX+d30niW19EybPkJ1J/jAzyA5WcGW/9H5dpCvSgVrv7U/MRkyB/S7M/Jz57r
x/E3oYcNPxVxWMuSSn6dG3FbbMXT5us+jaYsh0ZfQpaoH4PkBoklPCShL6AV7KZwMVfAlu0LUZC4
Rf4eZ5cyr0O2AN3bn7ix4uou68s1Mfc9XOeUSyWamJ0U8oL7J5i9wILKUe/P536HERw0VUgljYtY
9CrRKNNVxxbFE7seGaZ+cTcmLHYP7ChR5gjSZ1GUS15om2LdnvouOoB7+4jtUQ96dAetN2ZRcZYE
4lW0l+ebjbUovDEPHHhDXWKCcZhG1c0swaXFQEdEEpLdQvrvOzLtN1Zr7J6ccF23eMsnKMZEp5rI
aQs1XFVNLo9lLcsNfhleaB/F/Oq4kXCL8DAgQzMxAOm57pb1iTDzUsV/ykKhFk5UABcjDjwDPJut
1n3MhL4rL8zKWbPhH72gRul9j0O51X79PgEb9MwXW+8lnH6+J7wMq9V2Q/ZEtTQMVI+h7Cw8j6C9
dG6N3LvYl3V7qsKoHQL8ijdZzie08Se/S/wU0WG8sglNQLe/7hM9gP9X/KSBqNFLeL86+aDFCqpl
Qsw0/N15ESa1KfMlHsk7SXN8cIRW3K8gDDijvJKaL0zcB5BS9N9DXMdOcSxjrvSg6u8dqton+B2W
a58vk3+0QmVy6ENDDQQN/grMxrEDTueug8lTqM7cB5EvrudDiISRInCF4s52iua7VhXCK9g3MfMs
/X7NHELE3hf55nD048g9FFsH90HjWyNaI2WZqtjk4c1Fi3o7qowxw2rri3vDG37DtAN4mAreI7ib
fAIRH395bPTpnwQGAR1ejXXYHBBu4kfZveqshpGtzw4rAqypIwnsNw5ZZ7peIXE89iRKaJ6ylAQk
SJYStW5R2AR4H76/cFy+Aqvxd/jwPPhjts7ajCVFmqJMXU/Sxu+IzGfCm17/OHoA3OUz+IW/4vuz
t4kpBMH0S4YFOWeX90JAjLXjpuml9z0pxQzX5ImFW1ONiWEp+KYfeyifzbYHIIheNwvPL8b+LVOL
U3CE2MSjqE1nqf7agaEE6j8UA4K90JRId9dS+bkofASBDVS9djijWZURWwYyDFsZNEp2wCzyrPoH
+mFUsW5qKCzCIP0/Hq+dZsDuGIcSPNn5rx4owt09K4vcpqWmGVLoaNKvTIUnJ0VNQfzeVF0Ub4cp
C9vPUtBIz5Fx4F6aXFsHzbyRkWXhb6PyMUgwC8piB+aj8uFn2fwiIFXtQ2ulIci9V8uol9dr8H5o
IVX4/0xTrw/5oPJ4dpZNTBeXEGQHQRw/9V0vrEwiYydtDMmVhgCfxkzUHNVmVeOwruy3aksjf7Og
mTiI7G+rxewq4iyT8pnGGAck4ROwqoKmuP2P8i3mQ61DCaBizF1xjZ3QTt5NFvWnA9g4RN8UHctp
o0qSagk+wZjsGwDnthDOLEcDa80LOVPi+7USx7WkRLF9PsJVeQOXh4Tj7gvI/Iaa7Ey5P1n8r4dW
PKQTDGlJtdAifqEV9hlVrCCY6eDSlcd48V9aNzW4qbY03QU0Jdx5EP4M77mZde091zNjx8CMyzJU
fmbWmJT6fMXzbHD9FUzn+w5WpBa1tKjBjlR6WhosG8cYmkcMOIh6dODbjRm9VTSS+wu5i5JwZo90
WZJxQ+kbJgsDjC58BKgrkXcoggwAZB5gWO2xx7Cd2XEa/KlL06qnVIhvhjOFePLp+eWn7mIwpS+B
T3z8g4/vrvLDkj8s8q8m40c3SnQnwB1KTGlcaqwk8hqMPanLRM0k+c/3xhzsYaSuu4so/rOHX8Y/
aEKNcQW2HpeCoU4jVZoYSL3sUcock2OUdNgnnWkSbQi42JN8C6s72QRVHAZ2Nlxmqe0W4PudaLmM
NeWe1QLFHdA4ovpbbcX4LmU1EfcdcREG1rNDB0uqJjvVxtfFxiLNEVJ5LG7a7IKj2GDXCT9vGJms
9R5+QyE/Z25Mzp+dGsR7FG93xyLFsML3/vjZMtBkYuVDIbr+3qmTcTCZtHcTx3uhupHatvzyYaZI
rJcnsO+DvKc0lDjrJS7RoKXyILpaSK93QD8ddBR6LzmtmBuZCExTSnka34S+mCWScqU6iiWurjqd
Gm1ZalX/hKDXemoF1yUB256bZXlXvbyLAkRo+4BgorjNRTaGyIOxvxdvTzeSZPZIpgjpWDTltJLQ
rWFvA/2huZ6iovItyD6VKTkknguZ2LEqhqjnfcXxLJorx9vUpoaEfn0r4XfuLr7rMff5V+rjzUxM
/4qy0LcCOQD5gcJwPWWYlat9Q3e4UhADOHkdK+i08EZflJNH4+lk8DULK7QO+NoZWcbCtFgR1GbN
ibIfAhEyr9DM+6nCblB43dZI+VmyJhVtAvWN6AkI7oox1C/4ZW8n2ato5TJjUJLsUH1EiGxtLh/u
ttBBoV3vGg/gDi8sCalSTlfx9VsGl2AOHq9Ra94Sqp2Sxrc6VAtf4KbUHNMf0ygudnK4N15nSZxC
mVFBGoX1++u1sSHG7RJu8dQRbRd3Cibsa8u16Oqriyge5LQJspEnudeq/uDGIYc8gMB2yJv01rIa
z8Ddw9T/2WaZHzSnGcDGcOaDMBr56m1dDnQWsCeP5z7BGEikxeq5eQxqkTLFxa8sntSYE29Wa3CH
/IDYji4VhbHJzR5O+LFIRkC1Vqx4kYOVBBTXFZfMfWlGMYxHJ6j/o3S/5FsiXzE4Y0sM4RxZgWgU
GPZ8D3ElXisVtpj36oNFdkWhqVeyoBpTVBFYWPWSATfrgWVc42uhjQaNOHZY2XEwaH90ACu78uq4
yC3xJpLNiz/xgBpKjc/8qP0WkLsW/XkqouVzzbjEEiD4QHEYPc9F0O50xFntvi5GCIPViyHuZN8D
T1chlWOrShggnPpdQxZGxHtTjd/AICAdmxVmZVSD18Z77hzurTWZ3nMELS0FhQbwmvzswPGY62kp
DvzGjLT9komV01l/XrfBXWeu6zNwled9kElDMl0pR+SiHff3yPU/Dvt327Nvv7fZD5O7bg1VOt+q
C6GRiUbGMUTaxKy2BNlGump/LHEjymGdXR7DNRYzYJFzjB6xsYXVcK45zo5NOIANixe4UGcItcuu
A0QJPO0TXX4eBW4GmMDZbh4WNKL/zCKXOmfx3TptX426SqzbL7OB0aEQ9nYiNzhTvVoJn786DEvX
5lr1E0yPSUiyAUIcQIVHi0sM6VbExQQLL2ZkOt4aXtcFhFpG8O02zwEwdbs4YrdoXAig/zji2pbc
On/+d3ogdKBelhsndNMJsDO3oeiJJfu9/dT5mlnzjUjdai09AHXgSCnvM3fuDl8YQYTDTzepgbcX
8FU1fZpnTA3GY+t+6t4cKEBjPib2nFL8ktekPsnTk6ZB+GU0pizXaa0guBNjbp8ow5gFv4h0MHay
kduaB3mbArpLPi5+d93TuACkcIbFAEcxBfUfue5oXnRmhtLNiuOjdCJOaxXH+SEOxtN4RIyqiUgd
pG/VA8Acymm7rvnEkfEaA4BPX0bL9/fvIFShp2WdVqQePZ2C0HLC7iDiYjrbsLS/czEbLvLSxaCB
Ykv0nnMHvyjXogKhN36d+8lfp8qC9zV+Oexd2IETlUtL5cqGjoqBgJ9jhLE+SdBojgLuK/Urn1pc
Hy+j1/sXREQtCqOjaQnqvormeKR4/5/Ua9JHN0v6QjMGLuSYZ74HpfHg7tW470XFUc00IPKK5NgT
CYHqb7u+qBYlAJNMoOQSb9v1H5MCi3esZGmRQpdGBBy+ZGWdqoZwde2lNPMyRLMUyJzVrjKsJAh6
M2Vc5F4cZB3ZU73bzsEqZt+/AzCs25IB+4zirviJlKZuBtHFr4nFwREJooC9WDvTp5n0Jx89XdhU
fzsOISNhwN8ZmEYjTL9Wi5KUXyWj88r35nC6SuAiWJzB2wTlmeLecAQ2uxcn8tNGqrumI1ydORMC
y1PgcM/G19BiCp/azAW6L6EvsLigcYS+oLl+c7eNNyhLaJAwSl+SPXEy3KcHpKg02Ijm5w94KjRP
NI+wj0Y7xuxA8gfoQKEvBBeX5mauBfQHabiOrVd18dhEV+j6jmo64QscOLOMqd1nA7qLKv4NUx7w
xgUxAJfUOuXnge32HCyHaQOxSZ099Z5FMxvMLJUm8zbBJHJbwna5HxvZpWzYMfMqAtxuNP2voudi
MVo+/LHk2Ouufjhd7V4m8yRUXrT+58vqGevlHKLytQbZYBTxcsIVyNIungWYMacGFw78dJafCLFv
E1+N8+F10gAp47HyOoxwut4NRTebEQh0DXgoFHKy8EJN7w8EL3+bJXKOfLeZgxsImvSoA0xnYH2m
xaDl0q9xnTTrDI/RgWpgNX755f6hMLxD0wMEJV/igTRu1PUHR/2a2bP7Q4dG6Iy4PYSsgPSBDTr9
3TfJ+tG7/YeXj12Fe5oJhvOLCy+RqLunjGLOTyXAKvxBmgHfj3/4hrqy377dlwWf6o8lswKt+d4B
DTe5jSMlXdGP7syYhf5QGi+nQpXW3rFY+Ij/xI3noRt/pxk1IJoi+9zTjKe72PCCXmHjwofmpO70
4NOp9RQcMH0WoC30ge+6VVOVcmTvWVktjmuTOzuLcUIYSSca90QogQZJWKEaTQHndyMzWsGxCsG9
zZelDTMMGMeepe8U8Cql8npYvfHybR+V+cAgtSzyyMImA2qLvkzcKpA4viGyBhjlpU4p0fzPL7nc
rdc3G3Mu8g+XswvUIs3ESF3fUf17bpwmqMgqy6MGGcNTDhmI6FejoxN1ywJJ1jRA4ZkStUF/7vWI
nCxVBblRxHo/VVUVk885GAEHJ6LCx7aQjsZ7OLOTy3eBVPKT5pIegIk+rqpqCA4gcDabySL6erGG
+/PE8SxNxUDOD1ZIpEqwYtS6598HBipT27tfSoMC0jQ7xNm0/hNfEQg/PXhM/ZEzWgn43T2I1x9X
8AIRPpFd92lE54TnU6fI6aIzn5N6bwJ317cfgK4CcMnPSL33HgoZ+0mG4SoDZW8N5PBy6jhZR9vd
AxIXSxMsI4v4VEWn/o3PXxqkFb+izRSE8CLJmmDZPlbk6O6K1bBgDw/Mm3ArlWUkTTvd2p0aZvLe
Uw0Cg5PGpJ4bDFB+q/n/V5NtSQ+onguOdkeI7KvwbqGI8k6Pdao/iYnmm1mlkJG6pNmZVL64uCWL
qE7btBWL4Ps68SUapL6/sbrJaTQaGLIicGUrjQuUPaKJkxyqk44FeRneSOiTD9Vr36addTu2IWBt
oWl+glHTl3Aj31rjedhIrYxjw0XAIxTzgJsnCDCBIr8KO7BCG7n+fuPZjViFeSFgqo1xc1Fgg9E4
J5FKvN4mLSD0X3YL4FczJMnuZ08uZtSV/SodooXNUx8tO+119CZSUfDpwhbzKLc+vW9wvb8GRvXX
wbEJmGrNZcnZmXTb4hYO0p018nmwfNDpdT85ZfhdHBAgVcsHnYkR+xioLi8labSrKcVe+01EZGCx
RgPlPZPrevA90cg2a7EGILJeluFwArpH/pUEfvOrw/qnYGVVW8hYL2GR91F5q0fd9TmOgRzRLVgb
FDswFTgRD9VxXTgmnCGTbyVegzVVoQuusjaW0Q8U3omLKsa7P14mCdq0CG0dNtIzKkkNHpnwoW7V
VtCSFVZEBcE7SWYyoSPAeqlCXWmnhfrw0rkTtvvxpJj4iAPeSoGcLWeGy8ZgVjTjLLka9O3RIf9Z
d4wEU+9by3tyqNCLdzMDgkYiluV1rK/qVkmM8Fhhgr5GS73IJCwDwu8e/nhdb1UZgBvzU8s1L/6/
PN/kMstldQBwQb7kwPhrXw8oG/bzmP7RssUPluaiRWtRfW/nH/T3P4k9zGmv6bVSxQlfmh/rflch
6tE148zmtjpzJT89jl/9+xsrvg7FS2fb75sJCgi8CqIxvhcAyoXmTunx9EVJgAUw/2IBFoGLbd97
s/VDceHRalWgDHVAMvo+loAZPl7wruKnbzPh1z2OLJhr4qd6DclupWH2L6nL97UYMJ0E82HujCh3
vn4nOoF80rOu+h+ekTenqi/Z8ZIjVTrx4Qg5ZxpTuLSX2OWuESf9u6L2/qCNBA5zGo/bGrg7IQLQ
asJ9522axYzPFP+4Zeu03x4K9CwBqVEL0TobdYerasorlgM0XzAjQzN20lmHRssL5O7O8KtxET5C
sIEvJ6W5u6WBKwumK8uGIjjJA5omnJV5P9TWo6v1jEECA5dHeOziVSiBf8XLj3SvVXGeRkZD83dC
YtpoQdQRI8HJRH9pAvHZYE2BfRSRrlFDgChzqi7RVqVnevARmSaoHCb/nvkzVkKNCyCBv56pBdNZ
kAbmTDZGgb26ZrK1eRVzYBFY/6IbZbuyNgd9Me/XzMt8TgrgkHwxzwd2SnzMU6S/Bp0XQ9q0IDLP
lGlE1ZL+PWvdDynxwh1VqcKH1NuQ7HRIqcgrkZ4LcVUKQMfZMS/GkuZJMEDigHgd3K6yfjapXhc3
aQ7TFI2LXdWXfo0nxG4VDmO+eg67NZGC+Gvp40d+vkiwAtlLpsogXEHySQFqAEJOLX7MHdACnJRM
qeKHxkakHdfhx3xwqw/FYtsn3O4ohzzCXjenrT+rWsgMSaNYyV77qwozIfTp3FeOSAQQVqh8mNs6
8G3VqFiiUI9BeAT0RCzAOF8E2yLVshCnmoP5EooNBx1LV02T3p8QmPSRUCU0rbvJA9aZPaAmwREi
qbBkotr+2wFvLeKpCcm767SFIi/qyKbmjINyQ4ytHJj985fK2Srp0XJjjNwXUldF61tK3pOj+7La
JGISljGckdGvSEa5swFmK/w5+FnOOPXr0O06/f52kLW/gPwXIzrKrtWlRGoH9L9XPUZgkiWeZQKJ
hK930aMyLrjeVRTEMDith5trn+o9Ro9JbSIJO5S5+tv+Jx/0jn8xrc5KsunBqLAh84t1KcT+JSHC
s4kUTtQVbbkcu4g/JJeoYuGeOIE9lE+W4uUxTifLOQfRf9ewoL8vlC9kZURCjN8l92vmZKfeXApu
EOwMJXoQQgqmjvQ2jKrB8fdfhirWhjJ2kgyDuhhGjAykgNAhS+RaN3c78dXAREBdraCP01kW9ZWK
tmJyWuReI8BK1SZHejQHMLVxUU5mYy/uWe0Pzo0aRs+d+jY3rmhqbPVNVBQQTS8NlUIvczlakSM1
bsMlns5XPzw8ul0zuLbEvXhdhdVKHhdSNLrq0LFxHbsKE861+ONRQwJuHd1eXjvayQs4CYeR5Tz7
+0+JvtD5kVVUXDMsFT0MbDXDHVoAmDnnHgiBsqtYX14CHEe7ozEYCx9yu85ygB0WTOHj5318dKhs
QRUi49goZVm0F5nclIQbyUgLzA+NVv0dA5uFtnHlQSee97vUY6Lk/BxUO0tl2axGrBmE/BGlADLq
WIxXcRzjwUdaiqJcYV8ajeQ2eZP/C5T5I5wHlJNxxbzuDcJMW5u9+z+nu0PDgeQmypw9i54nyzsq
P/tcUBc9xolOeqby88EN9mL9ui2rEeeKPyMPW4PjrGbLjKllle520+hvAjw3jqelH3GtWCjt33dj
cfWh0/sx01TI70fTXbPqo8StQPCl5V5xXHyRFGyagmaTWBHVhcysonchQXCTsICGhYrXdFEdmZHU
5KRWwVjn8uUcS4Xtnurcrzd0ouQvx4jmOVXfKNzBlIIXnubwmKIX3C+1s/i9VEyqzZP7Kev9P/sN
Wi2ps14WYmARrJJ+9x8AZ0YoTzQRc2PJDk0D99AFzWnRYb+QjdB9IG2pxuCdOw9IS56tY1z0KEwP
mItZ+bp4UC0vm+GWnZQvaf7EFsK/RYsn79OoBvpGLmRLKK5eSrvv93B5/j+JEg/55jfYzDyQJrsa
2go0niBaWmTExrHwCJtUoYZijmRK7KqYk/7uvY/ShPg6qfHuNMUsxkXGU+SkIPrlUbq1jkPAi14B
51NLWW/FQch71MDhOU6H3n0lkjCsvjg7wT7YwnT92k7n8NGl7sUBueRrxdZFbBscmw3lVmVS7NWu
YHYcnv/Me5gRLV+yjeYK/Wtx1brTWmyvxmmOH9UKItWMOb4ui5QKt5Zg2Hv6aZl6fdXJJMU+XX8Z
lZyIt87RWXxQ8f7nBa9nzKCooiQKH50kJBgwKc2bzfJuhQTfweq/LWNvfqiuEYmcae1mI5HypRMx
Ji3WazqYW2an2fxPkEAz8t96JtbskSRd4/DFa9dxSArlkjdFdNMOgI/Gun3fWPVTTn/lVsl6y7TC
1dcWWkle125a/uAhcm1EuSRxI/bLRzX+jEcpM+0o6+0Eczhk4vWhqfZNvT95b6KpqEtkITqv1qkC
Vj3ObzcCXPjgLZdn0C+V/IbxBqhFSNcSoKYcKMhjCjM5uUVGgHw0lYIrWaHZlroCuZLVbI3sMGJu
BKNo2+9pLRSECFf5EbM30j18xMWp9UFQRMC83PuZF5yxIdvraeFFGYc0Q5sQ0KBzN0DAi3+LXBMs
4ekh5etI+Gx6uLMfum1zHoUXtByZmJ77Oi8PFra9iwK45DqrcuzBAhvQ8kQvev3202EYX3cRmhEb
PR56jMQRy9O3kIzgUpjG8AzZtRGM6u7eccxozCQmX+ACUkgf1R3AlGEroBxTAHzl4G4Az9lo7Jnn
TWS0TsE/JHafFhs3BGC+4GX75FUl/T9cRbihuqWWLp5wr4fgNIrwjZO3k/qJx+qX9eYGTSebM/Io
/l0p1JNHimRB/XVQZyiZVq7UGvQbA0qsbbbeQO5hWOC+GqNVb7n7WS3XBU5CUVpRNXCKTMSDoDYe
uJPCmjT9rotk19HHKZH4MJqPF2+x1gnd6btgz778P8gcPenQql1J9sByu1pbAYD77fwTddWjMZb+
iRbgiBu0QFPZZooQPEjqaK7RRiw0obJXDlgV6B+MNW12/s8brhFTHYeR2/Wg2DwX4AvFt5M6WyFu
d3Xj6arpbLDjob2gm000iKBo4WT8pOc7nPURMcoO1a5k6xsmmt1nBW3SuNQEoqwyfBD4xqlzKiWd
mDK36pOwpeFje+DarkMPlfBGDN1dkMyMTRzFz+EkxUGj8COqHqoGeT627g6XFTwFgUIavYgxlBMn
USSE89T5twIatcfFYEtCK2U7nORlGDddEQ9c3RTaE1HOxuJAsLqkzeWGYmv09ENRgxEEAx+qSy3q
aT+LejPBJH6cO5XSdzXMP3+VayfEuzAS1qcPBxQnwM8+SA0XOs9cL4DAoWFU6BBYYKyT6nlhvUcY
skaOWaSblGiOu7tQETFnlj+NRoFK+LLb5SZRluI7Dag/zLAzDtMXlMpFTY4isrhjUKy0AAVDhp95
mVHNglkyumXv7uiW5V6eSaux2elaeffALJYVWRzoHNipuz7KFKjssYmz2W1MmTcpzMZJK84C7EX4
ZvULGUh0bu1tUZ9uiaQcCFG95Pb3tPfPdvLFM2znjn50iPVij7DkK7kfAwfys70g4koXuGFJ23nY
/otNgrE2JG9SfRrVunT1Vv8tva7HhT8DCKCZQ7vVYTYtj4hMykxnP3rQLnDLRDSAWw5Kg/97T2mg
RAxeRI9mRXvJreBp+m6e/cHxlCD7Fp4fooQXiYjp8k17l8A3JE7TJpLItbQREAqDoLRhXd8/Dkw9
Vq2t3SGTtV/zBpaIH88KLLlGdcZnOxVRVQQiEwjrJGCbWJLEt2sK7jn/bNMO5FX+rxbv8+3m7Owk
6yk0Xrvc+TQ0PKz+cwOmMnDZod640ywiyvBao3GYmmXSVuPtB8/hdIpQb0UIMyZpANvPgqO2hYW0
lEnk/R84EjXeHfqLycJ/Cghfr571CuZHDHkkpUcldub1QeqkjBfOy6drGdZyinhvkX+wdveuMlxE
n1BEd54v50zz1u1AjPjbxyV51zHu6bGlP5hKkqOuMsUAE/Ezpclvj6bWpQc9kV66EVtElmlxHHgX
ZHPnOfSBS34+En+3gEQdpA5nU7QsrBNu4+zQ4nsAzbWbv3myYyjv3g9mxRfok0uzQRGjDn7/uLaU
bbWKBeyxUhilc+DhIN99ITl67S4pQR9wa8HtBczEmCrDG+3H2QVNlqACAlqeFbF2+NtyMoczdTUG
/L/eRpl/KZjs3EF4SctEYmXaEphnzUgJ0dvCGpCgKPCgJcJey3mwvEccMLxYnGW9V4Tn0uGHsAPf
P38Mz2lLLnhaSOdvuuIF3gDeHbJ8I081KH6a0ysJE6wfHvEx3YkGsLx59zpDKhofDcadTXmuaxMV
x6ZHSCOblKq2hPrzzlriEMciqBmXiCC704U8Y/TI4MfhDyGF0X7lcVZY7UP0gCLUagtaTZUtxpcl
noA38q4g7hXL960Y6evKMw0HSPmISYIvBe4ZaggIhaXPb///epbF4kF6Pfc/rGfuXHVbIj75ViH9
7aArDZ9qLjbf5Fp94yJn2o/5Ow6Rp0Roe3T2uMX30M8WF2lRq6ymOocy1aMEoN9VRs6k2jet5nvE
HJkH+QpuSDnnpYi9BgdNT1qYzdVl3LhDUyM/2MPI8rSKKOl0UIob2AU3fvlcoYeLKgCj73/njcHV
Ue9nSMgyU6MxqzPcIzeBsfkCS7aqOAVLvwhLTfl1nXbGB4VF30LMEP2FVKHx3VaBuG8/6LiAOgTj
MUwT5jpg8BJ3sFY+MsqL1WldVET6OHqpWuOElhQGARIig1VyDNM7k8S1Iv2bOL2mBNan6JstB3kO
LdiT5RvTCHXXDFgriA5Q3cx5AFNM6JEuzeXsxMxgtQaAQLpE3YiHqy9zKt1JNKAUBN87xkzO5xIm
uxAwFHdByVYJQMfo7eOQgZ6KdCZn77q09+GASx7AUniqED6fDs2aS5osf7Ifnd787Vb6cHpcoO6S
Zt1JyQiWK83zlWsui/vbS0UmePm+CgmD3g3U4Wg/666HCjELqDOBSRlb6DjDZBIddWlBkJLWLUsB
v93Lv96ZiE4OmBnBWcp33LiovO/WtRjy1QozB9SEj2MhKg/iG/QvxqC8NtsE1yPhyeb8btVJjLW2
mPIYRj2/guBJrsYY6HA72HA1n/6yFTojtyl99SawRDGT1/i7iocLllJ82VG/3RSHwJyN2klagrUZ
3NdP7m4ZfRmHYM992II2O2pI4Jlejz+TaO6nwARajwqABqfzgYXcp5kSzF4kpwxLgfrqJvSe9Enl
Z/DEPiLP+GPReUX0jbAwwrVUY5iAX6HcDTDx8t4sCdt+7KCf+J8ZxwxezczFfb5BT/9cd2xyxKd0
fSthGkS1ou7ivZr8v5cG3PibuNfa/yIdF50OlLXE50avWcOMv8rNGp0Dx2h8G8UFg2XX8TAQRX1s
5uihqoEXmy033HssGUsfMEtk+OUU4XnFLpOqZPlS+DGgdpI1UqbebjVqAkgDB5X2cGGe0kS1byPG
+ioKcMJwpClBvmrOztzB7RcHdbrT8Z1xa8qXg5O6ipcMqm2WH8HSsGh7HlvnRKlag86LaKi4REdX
1avI4TwUXBb6ipZ7ldCFmcRdvuxXc1MbFEh9VFexD0RQmaMLtoDZPMPZ0UfADVI2OP2MpRjvBVvP
4QhOneZOk4VUXwmcUT1c36QJ4os8h0+xFH37/S1Ip0WppfwbGEexnn3y44Ct3/7AbzW9TRwdw0MX
55d+8a3kiEimpj4kYYRq0uq1h7E9zcGMG4idaAdTeppo9Hiz0PJfupPSPAMI2gl7IvIH30MhXdsh
Oh3KINq3p217d8zU7ZcIfM2sHOPGxk15NfgzQ28cQAtkOES9i/4fyxJuNd0sZcrmU+qgUprVmPg9
9RV+QYGny+4yMkSxnAtLYV9V97juxrHshhyCD29/rgB2AtVTUgHTsu3uFS38NXv8xus0/IQNDtha
d3trWbF1YUbZ0nNQfqbzLVosNyERpKDeOYoHkSEHPEeTjDlsgsYcif4xQ0wJqDiCXTE0OEXuVvCa
UPMlhoYPgOm+n5lytyG1m22S2Z6mTG9DHaaCaXgBmI4k9nkvf6e97Sw3fdGWt0kSm5npCbCCSAA3
QcLudNKX8NvCb72VcEmnTnRiC0Xrf6r1Z6PUekGkrtpZAjSEUaJHVm+Me2x7nveHj3FRKNDso47y
eTCZxAuD4VdFOt23N6TM4U69EiYui0/cVs3X+Ci0Wj6Ks+j3rZ+xegDic98yvwGOFD1c6isNxUBZ
0HWrAjIF/fxeC51zANTOV2jV29+9bhSFP2nF59m9Hl4VPOyfuTxd5aR9E9KGOn3dQZAQoweq5wQY
pnYCL3sJME5bVg4yznPcY2RV+STGRodlqLoamEF+S7jJ3ub/q8AIR4JB9xGAQ0sNoko5xFY6QQ6i
BzHA4h2aEwBBwnxE7wEvl2267xW8ihekYQv5S5+EfUaDiBjfq/5JolrMg7z5F9EYEUac7lNPabd8
U9bVf1ciEYL1uD/vDfmjwsJaPLWLRI3wRWbKYvo6L/Vh2/tygSYdmWolcb2Nlub8gnn3j3XTRT36
VEsHUN/9O6huAz0xp8emZUr9erDTz+SKZ0ovcH2HKnljjr6aP1ObvC0KEuKlBKPi5irLLDroNESJ
RSDhzKEyyS4oc10i8IfPdD8Nn6fTGY1S/w9eHdH2nvZdPjNPTNZxvW40nkUJQw6a5Bde1SbBO+O7
XQpaXWP0NHcyuApxg4NYiod0IggdsZHinqHHXYEJ0rfdpzQWC4pxUMnOmOBMc6PX/5sW0BBlBOpV
fKJnzAjdktjWN8FrhCZQnnl/LR3ip5rMRbJ3Jes50cXqsfgJHViVpKtB5c6eJSuCAESi+Uq2hzSJ
h2d/vGcVyeWy1+xR4rACFfFsRUvzvNZu8WDcjqiZK8NLacLXhMh8tQuvo3HmhacjN9CNuOPRPsCT
+UoXjKFLB8aTXtTxnrqhv7A1TZxb4l2GModcq/1MOWzb2LkrVXMB4x4eDNvYOrO2w6chfUZAoXhl
IxcC56gUTnfG50ErGlTD1/UtJk5kRdFQ2rBMZp9mVbB5+S8ggOAPgD9gB8TE0y0F+qHjdOAMQyy8
j69/tKXcsLeFVPyCSs3vUb1gUmbytP7Fn2i/U0nMxNOpdvk2TEhn/a8hTyjkV++rtoma9vw/z2rP
prfOntj7522QcIrGWXi0T3iCIgQcGXf0PDeyO4pCOLG7d6eSNvFGH9TlW9gBFQkGc9oAISh9Gnhs
JG3oYBcUS3qd+EwimakyHHIW9wnwS28BkVYDbDPrXKt/3FL+X1OkXd6Lb5Js5CbZRI/3kmPWTkGh
E1GUozXufQibU2ViWLs6ANYcvj6ayiXk6ztmkQzeyIbrlZ1aPoEdL7Gmty3rVEc0+fRaY/7OdL1o
Rss6Epy4mDoQYlym/L7isrnzqL5IVoF+5Kh/dI3iK9ZfW7NFEcQb8oT6OJJGP3yRTOqQRNLrOcSN
YDgGszVZ1K4/QzQFrv99utwEiQxZCZhD2ROiu1vONuhbX1lle5uO9jjW4pM7InZ68F3gUIPpZDkr
nePEwr+jXDVbGerfZjdgnKpLJFWXwStnXSBTqSE9K+mSQ21xXqTmQ/E29VI8GFTGEe2wZwkPKh40
qkvEdE1A93yItqmUavocDQ072A/x7qGT43kRQcVlYCDa/zFKGmtOtE9BSRmKxQIYOkI8njL0sUPC
1+TN2f/1czI3VxtIH2R+wuXitODWpAIzz9xi3pW/Rdd/KTFcTcB3cvHcz8knYcNHwtZ4Mncc3BBB
4BAud83g9M2R9u/5mifOduaj3owajz4XkW3BWadYIW9eriQCwuutF0MwwFYMZVxKYWsMTu+jBKjp
wucr3ap204IHyFrspKPU4xce/YCxpD6H2POa64vg2OaJf/i96wjWntNiGSjiFHfV5vGvBunFYlO+
PiDddFxuuKgyJKihhRWJRpnuPn+a+fQPT/L94nwvfd2bM4dQFQXTV/kJ9G/Oo5GAM8cKDuz78pPD
q9yfrPIPe4cmL92IXpjlwskgotlJNql2NLyvbvcxosMivMdX4B02ed3qgTeeJqyEeSiRtjDQxGBo
iYdIjaMzTQCpkbKjxYdoWMGf4XvasGzy8XNPH+kfqYdmhOhqiL6GBodOGxCqQYpLsNgEs1vGUe/S
4A903mrUTEfJ3/tNcmkzBxjF7aT84z+wB26+WgjZOr7po3SMe44CceU/DFhCJLlASmn5hLY+QGlk
5N1xYe0S7JcL1v/gKlnnXijTSYutJmmpgedNtxsolpjs2nLsOxbIc6TKU4h01NjyblxnisrxkINX
GS3NpbFnteUwnfRd3rGtZFH82FJ0ZY9qRJwwEQuuQf1OQ5GlSBdrh4hymxr6wU3Jg/Ji1yuzJMfA
yS1UKvZQR7f4goVjpeMS0Xqxjjnilp+bFR9nnJ1ZKLBMO7bwTeaT2cFXIPl7HT+OknPw5FFSQEQC
eMSATmovUDm2N35Gl4OVLpqUKWvCYpjzY645D/wIsHeB7jDapFS1Vd0YW3mpnNvPr1xfUDUSJB6y
klZzdKrbrtoOfMsYMZ9uquSjVo1ORBQgQEz3bUfKb6JW3cKps65h/dtiSD5+Q11Y/CVs6Sb9OL3o
Oozkyz00OIK8zg6GK+Lf978/hxWelLXlXstcNvwnUHdrdSnI64Io+7j80OTG5cNFJQPoyM5GotGP
niBjdDpQxgo7e59LvQ24J5leTsV/rmuLc+7PLtk4QLhQ3HfGhxZEgtelAlNcWvQlKGvwMgzyNXsn
olD+f6sUrG4dr6j9cbszfv6NhXzbK12kQ3IL9jJ7ZF2+3cu6DXeLI3pfPhCklUKhMlAJ8d/SkySf
YoBds+wxEAs94C4V9I6ZanmHOa99QFiBCEg5U2TLtWsD/a7ytyhk30qEfn+DjBTbL0CnnA4+w8av
To7Jd/BcS2AXwQLVsf04wJVTXHg4Kv++HAvysd3Y1h+ZN0tm9K6/rHuilCu+B6CO7vWdPjsBRqQG
wogJ/gJy+81MppuN+e+52GU+1NY386Mi9SLHmtgfLeuUgUT5ulr93N4vvgbDckznBJPQE7LJHHhN
aN7pPQiFkkIW7JCVoz8mbZ7zztXWi+6l8VZqeZVeyPMfXKOccTfn62rvL35spZIS4E3MKloQTI3G
ssRk7Q1M+UeKKjuUqScPHV0Lqy8KRPB2SRh24eatJH+jdiQeUhuMNUjbIBELaULziN3vWmzHaqkV
t9UHxp13oOQ0iJY7TawL1xxE0Rxk0idMVnhUeDGHDuH32njPImtP6nTZxrSv4f4iowVDyt+UyBot
Dt/zoFb3aJl08jdNWB9dCsQIr6ziANbndy38/NMvI+XvuA42jGtAST8FACG4D7rAucxHLUrwS5+a
GBX0/jftAgqh9vmAajCljE6Hb8FEnksWCkDPjKc5Ja9UuLPJTskyRRp0WspNgl3m4l6EPXLZPshi
bZCVSw8k057rcrXinNtb8bZIRGWc+auO83YvHyjmf0o6CKlMJcZxUcuYP+c+JZFDfCuc6WoKNJv8
IgNxO18Dl0uzVO9PTbHI8p6d/GCgA/49SJSwEkkETZFKjL2TZp08N0tfFQnYYrKgDNfrdfNoDlsr
fHvCBrJX18AmUkGAE1WRZJdbL34srFJC0KSerx0b6+7aTpMoztczUs7RYqS76w6atl265Wm2Sl3s
Uj3q1nYsxdxTcywTORQQRafuKvTmQ1/vnDY16m/cm91Pfin3AQErIC1xF2+/W3ek15UXxHZuaPSd
GeV765H2+J87isd6q+7t1aSVgiKICNVRLf3vudQkwL38sNmDIV7YG948ZzevFCALiv0bD9GlyFkh
BonM8Oy5DOdXxfpc+WM8/81HNEfCjqh2GTvTl1Wxts+p371VvCTjjJBYAwksnDwZAzxDDtgrC1Lk
Zk3+6hC5B6sBIKPP/3eTRAVK0WlGl1ejsAn6Vovdlswsw3Ke4L2stU1ftCBDvS+zJGfC6rDtyM4W
WHfVWadnPdbeVMwOMvVqkWd/B6XMruo8oOl6vi8JMQ+SFEvt+zUIUKfAyQzu71pV8EhLkO9epzuQ
hIUDVN4BEXcBFtiGarNzQhGthvkqlPpp9AUvGRmWlKRqlddo8Ez9lbzH0PHvcUFjdbwBXVzlX1f/
y5P5V4HcnLsw8uqPja6MSPwSYB9Da49f+sRaWbKRinnWuE45tiCLpTAqHjvc6JhDqo12DB4Sslat
cpzm73Coq66QYU5CZyGHfkeMAOe+xEEdcNcH9eoCTsJXreHO7pN7fBIRYf+L4njZ6fp43uxcOnfq
Qlbf4eQBK1R5zeT0VZzBrGFiZDGw4TKMdQ1ffqrd7AASOV3+QQUBOa8Ct/mtgIaT7OExBvnhDwyI
16GZH8db5w5Jp9WWIidEYvpRxECUvMAxEsBRxjRpe0ooPHK+cr9Tcua65ikP+wMj2n+ZbtmWJIhu
2eWr4WrtNPHwGDa6j/E9KtxyDdu4oGpiui4KSyw8UW+RqRESU635OtRlKLOpCCHtB/4IVZe4VEXj
fhdJ6wAC3X+zCyhpDiuFl7u/E7qqZieNJoAX5TGcu0zvUn5tHgaJ0jFMZndaaN2BDKb5LKMOgNFF
TjT4QegaoK1Lej4T0lgL2f3Met4vRaMj55YDpEVHm+MNvSPBrhN05CvhFJCTwe4KyyHbgVcr+HPk
twAfN6EM2MgVaL15eyc/w9qep7ZJb5xced34/4kQ71NMMfjAY0lhamZ6yIxggQLebCzWvuTkqK0V
ohZcwU797KrW21RyUQudCR11jNiyYTmp0ZQySnkSXNJZ+jgmN6ET3YsMOMLdIxV2Ckd1cbxEmFsG
7BEtvnSviH4ID51rnQAp44z2ZH051Va4AcxGy+CTfBDFi9OBpG6Lr2ZlqyAB+5b0yuLTFdCnirfH
vHzGW/QK2OZUUoypGVA4pZoGN38yvUYYIwNur7O5MFCGAQH04yXhGMVipsvxa9rzSpNBWJKWK7LH
Mw+hsET9giE+y+vpPVVQ7g1CXeQ6qzyBiqWDfhWvkPeSKkbWhF+0Minkn6C5owUQ/YVaU6wR/5vI
23v8tCnVrykT5c2KDIHF2mBG1eFmnG5KCVBrvCWzzA23Hmm7S9tmtKexVoyqUsMei9aEPd+7Cxc7
hqyiyRwM1cJSONi0fjczjhC4kuB0XFtJyLWKrkqcxi7yByomxt3PZ/cPRl3P/+StAsf6CiPw5lSR
3obn5ubJaHZ5NN4AJ9QgTZCQpHtpqnzdnQfjaaJpfVbtL9Pkq/8FAs3WJgnULBLU+xijuPahEpbv
Dq3tsxZJuna1FQ68yM6DNxqKzns8IvUAf7mehUUvTMnyN4ulInvrDb5xG2XJbAnBHSO/2iT7z6Ni
dXhVeMXnbqB4DwOuSic7QEGf5xaFGI57FvfygumDuF6Y9WdbKMa5gmItA2KAFUiny3XYu/YkRa0r
14QauoywUz3SzD4wrmEQy25t1cCNPycFh/d8boSrn32i7mqp6rx81Xy2xGxlbRcDaV8QQCGihZUn
vTBjDOoNT6cjNCfJEyV7tK47FgbPPX8EPzLATlWzVVNeDEr1ZCnFvPcna5mCdmWxP5R84LljBR4J
YZ8HHaQPNKd9IwLxhhGuZGybJFhtmKaiVjl+xyg6sKqPksfMstlYl6f0ZPxZBOBAOkrQiOQOfjj2
3h0OSol4HnDf3TFVH5bNijSxX0zdkxovx7mzVodYq/nn6U92gCsld3QhjqqLWYzFuAZ+zSrzwGBh
rPQc1B9+Amx5oOaoEjGWLEtxpe6f0pLOoF85qz0S1svs9Gg4VPIPqeVcPZcEmtDx00tkqCeRXHcs
okaWuuqboORPZTNGTTKlrMKit4tKx2+ugLUMxN/1Tf9lwmdpCcvM7RF0aSTDkceboyOtS8Yybt01
OMmyYXGR4w+sj4YZxHiB8c+S/+MSoynWt3o0SvItir609+cy+KSEv4KBa0weQt0LYYcfemZI93f4
LQAQIo5ZZkqr42/SLNPMuEE9eOZwDomsExP7G53l743jbtpII/00osFFcKYP06oOMKoy5o7zfsNF
dMqN41FnHoWQRqB2j4YRqhy+9OqIPeapZ43hSNkjkO1KZHOS36aEzbTqS8lVmAe4vvxUdLzOTD0o
j0xU4uluo5SIwy+2dCLAC52SLP6dv177PHJkVOf7fOOjIbbGLaqi3LU3mVfgDMUJLX4Ow6wIkzPv
zMZovmuO4ACcoV6OEWjy9CCn5+0Hn73oPG8HY42Bf7cDpLs1P9Iu01jG+J2IZ5Jmsv1TiG/ftC1n
BQFJ6xsxxJEOMXPcYuY+CM+L6vW0QE3of1KvMjx/sv0+JlW+Jn0Ef2YyQF9jIzPzXTzSfVphiyzB
2ZxDdx6/3PvoWnNRG/mwNj/kysAL2bAt9m3sl5B6jJ2yOXZk9tGG44j8rd71v0HuQI3kEZwJWCqx
jMtYqlphFePYD9BVdBnxoMZdpozi/6rvdJbgCgdTwn3jh3dNbu6VCU1YTdNyGHzKofwR/cQye7UK
jMwYGm7hD3stUK0ul6iqG31FsILD2m70ul9Mh+IwrefIEDdUQxk8XtxNKUaITV0fyhKSOJ5YpamP
Vi5k7iW5PBYKnyaOMgfMkkFSJSyMjtmobWobUnDRZsy89JgXopeP92cxlbDRy+1kNJewiUuqR6FZ
uIGQ/TTvmQuhdvrGQLON/6c5LrIGbnod3CWjvN38icuzfLBhl/nuSuEJCnZHpltNmkyljnnvSTU1
NlcSXmpxKd1IqeLKqWwrP/030E7yUpyV8D8QNJUwU4SfPh3hgTTfaYB6hZ3T9wEQ5zHi/9m3wdPX
vzpk78PUoxB1cS93Sy6mNNqNu7Qbd0YE8V2DFizKGzThG1eIhpiWcAHmXOM5gT0ACHbloP9ofLPJ
ovmN5W2gRxDoIy1wgHMtTOypWxjIzEegSPcQlv60rgyN46bjfCRGDntGgRrL18YPt+OkGmMhF1dc
AhdTcExLdIMRSLCxHJJLSBaKeXvfsQTbNObeXxtdPDpQTohEapWq229cQ43JyaOX6lRv7P+67+P5
XBXgoiZt8SXRSbry7onpUFppGqk1fRNvDktyBYo0GYzuGG8PvErQTxjfjXb76dbCwJb3WNpEUk4/
E3bs3hbyc2H+IuD+IqeyCp63gx9+QRnxXManELzAWFoHB0kRiE0vFx/djZpDj4Ud141ltS7Pa7al
2N4JjLiZ66J/LFyjn3QgT0jz3J0CHnjNx5fyozX8mB0ksz8FbRephWTXru4vmkpPt7BliTQHwPiY
bVkh3SOStVPOD0BUMUh7pVoXHgo+1euBWcViw1WHoeIY+ZPWqrEa2lPwnLnSQVBmGRlIOwTTslGp
eaC3rsMUQ86Ff7gSxYet94k3lhOEbPdq0Q4+S5JvSHKpxRt8Mvj4rEOgAEAB0LWkdG1RBiaJR/J5
s0mgnfRrxqr9WEob8UBQAOBb4gau9ZppZ+nTIzL3LKxMghV5XyQow/sCNC2VH2hE8weQfw6mvJi3
RQ03gQb0cFNcvufIHpm5Kz+Fv/XdF5lrXM7rK+G/cS7BoadHt9YLZ76D6wUc0QMHF0KpD5vo3mY8
mxst2mq2pXt0rl22F7gUR9TVbOnjaXoAL9HHmoP02B8ejFehZ+hX6CUw6Be1BG7gW1VTEyF8Zhrb
YcyxhyIAMUxOaL016VFq/g9wPtjwMRrhsbKN7Fc5YRmlmjJNCImDiQ4CAHQF6dEUbqEmQIrNVMxo
FoFrN1n7rQzhUWc0W2IDZ7Dy7QA9XKZYJmgNS8it7GE3JC1i16fzQdFlzzU9xhu1Z9i+18GuSd+u
qecG/iq57CqdEFU32GgNryIJl44/PIFmK4967zgfkm4xyNKiDHCOFC1Q/L6d5LUTrnyhtUq+OmSn
O0SGOc9QFt4qV8AGTSCNq8EnURkyyW6fJVC7WvFyNhmN4D2TNWZEgKO3GgK4vY5tr93uY/2DkxYT
8M6r/ieMWTObzVSxI1YWimpej+D6UJTKgApzderoAzKq63p3UfvMYUotBqp7EW/Gvdd5gcxO6Er+
pSs6DLLpksKKbzogClK792/RLqxnjX5LvGawGxiisixWU+Nk51POs27FXkrRlnUdwX6s9nYKAUGz
cgwojgCKU/w4MbuvrGczy+CbD36St6H2OAfpIky0gJP1OLDBsaNykdWNc8zevwzezusEw0ib5u9t
v3c+IYr3JRAsf8QqRZjj8jQdMuAJEaYOkvaKBcq2lrWN2BCM7ewhqgLQOWhkoJCN5kKubU/mtRJj
qiJdrjqyALvR5dpOa4lRl98J6kRp5GYV+v1OmE3ZnemTfV7RZBVKO8cOZEkwSYo+Zot8sJtDZStQ
mI3Gn8l10FtDM++QKaUVw//y+Q2ht4cZMuN8MEQgfUusID2td1OQp9uv+wJMbLeEmGmUj2ibIUCi
y7yWhFl2ZcEuQ1GtumfYGPX/BM/mgFflP1RRXtAxgV9x7ZygY16+KbaJ2eMsIVhVlzey6iiLeJd5
hKmgdLu93weKCYvQg6F/O4tFZXcf2hPEVN5rFGQfKIoBT8ydUQAB24wrcJTV2S6/osuHTAGLivP1
giTEggbLQ7lkp03Nk2VwdJTmeqsjIF0tU9uA9EHVhUF9NI87YJ0DT4uzQy1GqLNhmfcQiVvj23lu
whVkF2mzwXB8cHBQEToSHAlH345hRnalhQYiTCfPJS8WGbzGSct1iIBHW/6+oFYZKL7fM+rfhgw5
XzYvOErqwjvlxlSRdL5C+m91CTSqR6JXdNEo1q2EnYuEwhqtnA0M6+bTxp5zCHjYjtMMillH54X4
vVDa5O+WrfzMUoTWqMTM5nM7if7BwImal89xnbPhYwaaaJnAJUup7ndkNqv5HFdqT2Sjjk25xCPS
7OcIsnnxMK0H2NgMw+XEUQzQcs5bELs5Fc/yToNORloS+v48jZY1XAa/DoeZQpVGAv2uCKyTnfal
IQuAcfywKQR6AxOMmrQhEiwebX7ARdyA9HchQHC0HXLWkXTJYqs0LF2l4kvWELm2HikWx24zHIY6
r7D40sLf43FhRC8UNNN9B9a0LLUqJkD0T8Ft7Q2E5hkVGlv112/sdbwaZe4456YhWsZ7jXX/W0CG
5CwdtLlOULhxVIC4xgcm3BRJblHvQfH4IQCNIK+KR/UC7JD+/gA1rO5JSSUWErIGvs3dva/Lwb/+
Hv2AwMgZe+ptGz0eYZJtn/4wWRT49VuG/tjigXaNi3itA3fedfV2M1nkWKGj9+DsL+4kCfLbNoj1
8rMG2ao0UmYBV940zRo502ik+C+M2WJIpD8KoyZROeMFnMAs/g2xnzruE0RKUucc31ZnSx2Y5zVW
k3YfNycR9xbTdW0/PMUmFe8PRSi91zMMJH81Bc0iriptnMDFJCo7v8CQcz++E1vxfTq01Ykmz1a5
Wa0afZGk/6H33YLA2khml7J1hdFP2niWZSeZebSevkxF0no6Q/nKo9LtFqb3hpF+3QfnpMcC4acj
eK7OyD7HpNukDZRV/CEyhZt8BhEocZi0a9yM5TZOPjssxCyDMF6dn6d2X//wh2fVDvK+cU6cEGwJ
En9NkySM8gxsKKRD4LYyHYR/rstXTZh3b/Qe9ynyv+40GXkG/3P1+R8zCSUjRQoF2k1W8M0vlOrF
Lxr/dFo44EXvzaM+eblCWnzKbXrnFtTIGyQ7rIA5X5ffmjAJXiTmKgUxGJetedPs/fRnRsvi/Ku8
izXWyd2ZxqZxEkg2dlIauBbSnU3F5fDCXGOCoutfi3viYOtSUO7TMzQKnyTy9OQhk4iqXtLyB+GT
PZM9k0xP/7dDZ+QwQoF0T/bk+wf/ICBHkSIAM9XT12QtoL5H3JXy8kXHp/sWO6HCy2dpcnuSMxXA
E4mmk8+H9wewzoYUvSB+5W1UvQNmcT5FS8LmcsCIydNHiHUJ1x4jXztNBrKDH9seeh5DHr18ty/n
qGFyUA8w3fYWrVE617hrJYO8Fq2y7Y2UXQ/h223nxdnwDnr1eLQPNph5sFsYqy/Z5K0qrlDNmF1Q
TmGuauPEw7VWkNr19KAUFlPF4CNnWZxDZghqC2IuOZP2dKPnCgIPkcB4lh/7iV5BZCt9B+9dSuyx
ZgplfJoM1UoMUgf6g0lVizdq6xh+uyK054FFBM3tCAXDplZdLCjlzVXGkaL9yAA3/7Pp6QvrGojq
m73g3Z75FfokCQAuXIpf3uyJPr/kdoksi9VwgFR9sudu8flgAtJn2+fkueCGH9N1nN4tpL79Gspd
P5LWqVnKUBOHi2kdeWMdw6yN75bNd3JgzwuZXDwJwVQYnD3WE1RY8Ys+70qGM6mq3D2LelDP6MVc
zQI0ZMe2wQ7HasepzdjnKRHGroDMXb5ldjfNawH3NWkRIRksAIn6SRljaavXfmbLmhrc8mVv4Qo7
QN+sxSjr2vDDeE7qYbVhG+zdLckkc5njFJZOnQ+NvYwKFWK8udAI0z23hhUicqd7RT2635q4N3tI
oTns9DbcWXOOvK/Wir1ESreELC8G+41fPijrVFaYBaPaTW3pKcdeig4z9iuiUgfoGijkD6nYJN9p
6WXIZdEscLrvV9PYkCAgdlV6gn/fRGkoum/1CcAb/Cix100oQka8IYVkFGRaAQzRs6lZ/n/NpIlL
xL1w5wasV5ZGTaDY81M6+jPT7YovUf5uwrFFog3WdxBLdbSeK9jDPtKYbBciZAYg8oKIhKLhIfdu
xTYGIu1gu18xSwBLWfSre7WZU54h5Yx7layVMNcfOX3FItakAaGkpyF7wQpjAk51ctamIMTXHmf9
vCTTR3RzqtZJ9AY6+0HEUCp1Gy/4LFmaQv/0knFW5ImWrPaCtibpiqnHQChxzA2KEQb384vSOMtm
xdWBwNyrZM9+0dqEP8lFwMUIxraY/kv76BEWEfQVjC57EpXQZxOFMCPKlc0sGZfgRRK357oi0Kv5
tEe0jryrWuT2ZFApxTooIdFgfNq+cc1Aw0T8NwjzBNMHQGSAmbMdoymDkv06TclYD8YpTLXFiPwj
zgEja/KqhvwkAQqExWmUBIuDREciquwAMvQwedNqG7OhdFa3TClpalZk06f0nWspmpRQ3Z1dwMu4
pyCyJDdr+XicPVprUBJdQN3+DEh7T6fqyLUr01LjRv55TFvUMpttAkGJZstuHYwKMEysDPMaWOp7
vRyNobij9HaSi+pVI0qVI/JIpgTrwCWgdtV6BVWYOuzY/FqxjZ7tSHJs+3EmS+O0a64NDrY+TX9M
0vmyRv82ytGWw9IhFmu3+Dh/KkOPeYsgrvpy2FOu6gckCzk/YjXz8VSWZ5SO70R1LDb1d0f0ItGS
LJAvqfOpGvkHrYPOWydYRq/gKmP5ET5Lqznu7VJV807VZuOhPqHrtgwJ4960ae/Q+uuSYiVPn687
fIq+9mz/AWJdy18ytUoT4tpAVJj4gBP9tUSwgAZHQUtLnDekq8PIaQLsb6rFVWE5scBNcaJ/tC5w
a4vo0AG+NCPmyRw0a2UyeVXw7Zgooi2uMfMx3WI+HsZ0PivOWfTY1Go4d7HeiVDdCBhZoeQGnG6/
U3KdD4BT/a/BSFarSx7dPlWYnLW7F8FbG/ryIqbZ0tu5pwTMwFmGz7Y4gpn19GW49lAoUJDNycAV
ZBA/GV2D3AyvucEKeBjuI1Ywxit9kMmuE9vS92pJD9nMo/ZHfriBcRX4z4jqen5LA+vlWpC2Rfr4
apLQ5ndRa2Og8bDTvgHmHlD/ljoYIDqkQ8rN4R57lqq0caYClc0h2xxFPiZbGHwUoQ5oOmhWnX2z
WwZEPVEYv+MMnPIgjkLdR7yhxEiTtf3UyUC7V+n1VXV7Kj3/pGvNWJ7vdOwYS9/0z1kPjRtAt/5U
BDq//ZQcY4u3eAb9r8jhw9aj97WT6MPRmNzhIIzsgels2cRct+353BY9CMMuwMV2bN7evw+NfO1u
vFszXh90VyKKJHRWQkQ8O6l3+YSf4tPfwxaoHZ9IXcCoES5t9SqiDlDBec9eEFIJWkddL9lwGL2m
jiX0LSKh/lY3c+rEZyK8gOMvn6GJ9jri98og2wWhXZFUiHIKBQOe2pNrqi/cFicFTAkY41oDgaTm
m8FDE+wWaQWyMZDgcLUyGkt880vSAl07FMqk48eaKYMzJmmxSp56UfkA5jLjbf1PHhqf+6NfWAgf
nekTExyCq81LGD+zdxrdy4vIg9PzUUQgXRowYRKFrAinJu+o/+LJ/0QtyVERnAg797IIg4Z9WQOa
Bghgs8Zsv233oo6fUma+QLu+PpyFK4dvo25ipoIsGVIlen1PAbPa3uGLUUQ9iUBZ07CWshIgQao3
DBinYXh5ff4MwyAqoI3ucUeoe4ScDGcwR+diT7fndte12c8fcXipLoxk1Gun02Hc5JrEFcJbbqTE
4ew/M4FtYO2ZgnkcKb+zO4aRrPOjIcayN6KWMxxw8BplsBOEJu6T0YeUJpaz8A6GhAak5xoAg9gz
4R3ANWTEUUs64RJQNMjIgCKaxKMbpVtXcSLLDsS9wG39ta6VMD9xpJE5utU9CAaK4Vq+byBwI37E
nEG6CvVceAMCfLOvjyp/6SsfQuvmeldZtoT5mJBstQGfSrpUrKUEoNtnodHD2xjMi2xPqy4AJPxB
ljAf7Hax/B26dR+NJXL6FMxvEs9+oCFTXRPB/ts4XMRtft4qstgB+MWLQ63hKtNfT1xyXYz31clW
sRgRETWtepHHnF4W+oN6FKDmxWL2G/VVgQMWTndxbZPCBVenaaAHDP2gMGT9yjx46QRYeh0KTAvE
ouhXNNn87XMrGlmsg5qu4jWehyO55noo9PNn1SdNGgjfAcno8mvdOsBZsHrP1G9NOHrhCnjnsDLg
kHXD9A0xwymV2nCGIsBuP4MnlrURUTwoX1N2d8/w9NV9f+7M5jChD4H37qleJINkF/ECgToLadqu
mBLn5wBK79MgvNWMMPhZrQ3HzjWrIZtsDzYd+pKgGFTvctuTbCJRAiJnmx2sYVVVatcbX2UE3MSw
GLw9yAWsjncfoLGXI9Mbr5bHMDDZKozfzHHu3Cjlox6iz8X2OREj/qB2tSphZ7ArEzzKG8m1Kgsw
ZpoLZ96hLCjlnvXtVGutYIOaYrTu3a9wuvCBlpRsx/km8W0YkX+2JzVa1tPiy0yjXaHampZWm40G
oTBax0eIKB1W9LStN6GSWDul2/Sy7/HquT8RuKy7zPxKrmSh2+8JKEPZ3RhpYPH7Szhxd47YlNdb
zdqF0CpGkg/QJilYfP7FnNk8r6uOYY9nDh5QNK8trQJFUESkavQv5VYcHKccYbaQ7yUpmFZmgl1b
i8MMUciuV6WKGESgX1q9dqqpKeJKJmqBlDUCI1tZEJlDTyjHFu4BJkFJkP8zeJtH2HdV+YMjKEAO
KY4/PxvqBN/OG97+AoDqgi9WbMDeuX/0wLJSdFaWonj4OdfcC8lk9sFcOSHUG/nvLfJP5iekm1S5
qq3NNFzELKZwimguxP7LEo3abdv5FkTFh9iXlCN6BRZzjajRESlITx45Au/wPXpbcY3vXBnrikR/
PiWyiGsxCp/JCT9zDmx/gjJcaMIE4ZiWJYbrwjwlo9sryAdDT7d6oS5qu0dXtmatVQh3yv6FJ7m6
2kNCIa7o/h+GyVK9X8ydZR4i/BH8FdCqEFsd7UsCAsLPTlsZ61uEcsjZJQfneropIfE5SQGwbYuQ
xzL49m6kXU8fBDz0tD6hy4bkhNoQXeBsUIBFk6BbP9EdnuNZC8RS8crP410f6ksf4QKbgO6w28oX
kzHVMd+FRng4PVG6LHrPLn8hQNoLAn+S3TMSaQCB1jcWg7EGPkHARCkKie2IHQ4uYAe0/EaxCpTH
H8kn3S5wFzNjrEjbr3GsGyH61MUaNr/MNGYfSstbiDr2UJsjwbybQvynEvfTgCNDpIs2MNCooWRc
L9Gr1b/31hA07PVrhVEXy8oGVsTsxJrldiM6rkGMEICilij76kSahHjxwQq7Lo7e4/eYcBujm57+
530E+3SrpOALLMT7aT2Qr+VgY2K3DQfi1VFBj47ddlmbLqvcW3rEG+jgoPmARLrD0qK3lpbhi4VU
8R0CItPRLcJqClLCo3L7upAqpYY2KQL8/9c/X9GxvjVXJ3TROINUudLrh5BOfgVDWeQl/y8sYk8f
B9dkbAJaPXJVzQ1lEn9vly/SEZ/+eUWx3Xe1HysgI0U1LdSflGXnGKuJVrjc7/0Ur9wwnmYi3iyL
QnZRik0htuyIn+9zSf36BRc/iIcibl8MQwmiqnymVJ2VcO+lf3X+iseXvQhxBXTQUOxKd6LhLL2G
iLIIPZZgs2aWLnIB8wJMu3ndaEy4YIvgv48Nt5bZ+bPRWHuqayCvo31mrdZaKeZiud+CpMElsltq
ZfOJJ9hSSE+hCWmjVdEJIYPLKleot6DxF8u5n1gUvmNGckojuKjzjuB/f75WC7/57gV4wqu5AXk3
hDre5o6fY5sIaSBaiRIQC5MJDT+P9CtEPqnt3Casd5rTrMM0IrGFg3tizlGZC1X/s7JtnSPRBh/o
U6sFzLPedWZ8gSVOW728pzsmbDYgyVDl4BkyrFSdguhMKNLOrf5zpqh54gjMxxgirNYPUlIutrz0
iH8fbEPIu9MlS+QB0pHaOGz3LidJF6yXxdaNWY5XAoDvRSvJK9LofrzTTnWyWX7RfVDmmjpVmIdv
LP9xvj/PZf0bwVoh/QWgj2nk6Yt0jpxTOM7lw53rXxywRR+qLRBf6NUh1MvwlrPMVQzqmz45UxIA
W9zVCHnsRyyVXmQvjWJ0oOkft7AagtZInHvZeCSlI6ehrwicq9wrakEVcaKWP+0+bgso00X8dwRu
y3cpxYQS+LOKzHA3vf63RqNKHBpO+bmrLVc9DnXAq0zQS1lE7o39P6XicuggV8sUYj45oitbNxl6
2s81OgzrwexHZZFw1VrCvZZSubB1HcEkzDHfbpCmDHVIAKjkXOMoM+8F1b8M41KtXoxYC3uXCTRw
agy4sGjC08AjLp5Dwxg0CFaXsTTFDFTJGEVIqzCpp8jNhC607TsaKsiitE1zGm7Iywu4n28s2YDC
W+wdqRHFXmkd/pGND/OSvs/jHgBqNOnHPjA5aNSHc+M7yK0Pefe8LCtpSk/txXR93SyBUSRs178q
yMlu8s1pSPW89gGhLlytpNtLD6a8W6r07zlYTYl6sLGT3ffIhP6UB9EGDv+1VU9AjXrvrx4iHHrQ
z1NAWiwvkopJa95s34g3nuPtQkeBaFFm5TkKtDsDd1gBP72eblbZmHb3L0BZKktQHo0ur+egoEcO
/H8SoprUE04ysc5sKVkUEbHttQziildpxBaaXLKBEWyPImHZSHSFjQoSFE+W1GBwCJb8txrPz1MJ
VEoS6RL1wbsilHr6RicPriZdRcu1xR9NicQW+jxZ/UJtswT8INT3oMcS3oa4BcppizN3Aa89DyF0
V+mvhfeQsj3jozXxMu879/fU1GaK0JXF3WAps6pIvrzazV2Obz0r91hSFTDok7l3pEDa5U+QM2vM
ZvLN/76udiXmz9cx42OKx9D1HkpmswQXJI2xuU19G23RAN+bkMJrF42XbHPLYM0ZlJZdjUxP2cdT
EIWyeTEtE5z9Tciiloog459LEipQMUeHGmx6sCeMKQpzFOzwhDD7Ocgby1F7ZJf3DHDBS/72CANl
m2O3FlavWUMNye+/MT0e2JNj7Afztz2Kphm2hKSO5rllzBWOoAIRGuYCgUYeIUMpJV7wPNuOyoDz
UA8Ut9JvTOKyovB6fYP5SAmnWYeiSul3CU8XuKRUT8AGwrKn2APlTRVHPTyMzLuAqIiyIskMjAse
7YA49VA9VOWV1mhynHvE8/hpmtW4GYVJNODlpg/y0ojcE/ETbmQdpy3xPH0SfNM5yaOQ0BH00Vw8
LxC6cU65NWkXbyv+o/0JXPuLdE4JEb+mb60CoiJnob0Y1EMn9ShDYTSYX5wOqmFqMFUGi+hAZWxW
BkC9LouaCNOVIyX/j0ZkAm+V+Cj639Pdblj2DH1nFxiJIK+1yL+hJf+o6Um/tCYGNiRc00dKOro6
x+DlwFuhMailiHJcB9ffJ+vD6eWOK3Gy5B3b7Tv6uwJWfVT4gjNxx3KqQ3sW39U9A/eTnLrMrBzu
cLGE8+p7ge67nwqOC3JyimneBmVY6AC+XPbc178VS22WOyvNOoae1PrOjQz79gozcGfpHhz1w+f6
gN6cLIuGsp7LIwr7eiIOc2re6AGAN3vimcZ3ajqXw3aUZvOX8yoAsnAQKLKJA24os752BYFnkA63
rVs6jKsHRT2lmeU3giY17wL0LfZyBY3An+73mbe5t3oWnM5K1Ouh2FsIoYtvLEfpQ8D88i6+jJJo
ChVt+eAC0EE/8/l8ZCFi11XuoISGZPZ9YJUbaRg1hjSyAZavJZ6MjVPXhea6pB4b/Yeg6Dl4Ikif
Hy4TUYINrcCypOvE1ECbEPKym+e4QsteYUcScHOz5mz8YXs1pHp6CQKJEeGrua+WHsUFoXymRGwh
SZxbX/e6UfrsRRRT/OjhPvVlD15gDCQMjFZCzQjpTzwsxCT4rzQVUaxky939eIqPSseqNC4QKkWt
0Cpdk91vd5i8303WedQh2cgzFOi/SdnuUUUM9ygFGQdjGR84EpXj5rdkDLzAfZNQQ5UHGAtonAyY
cPBz0HNMlsvaur8Nx2b5mwMWFRPDBlZfpzm3m6SDxbErhUPkGLxgvE41RzdVBACmKtw0gOVPbcXa
/9NiXhSU42x1WHtGPQ+AXt2JvGLLfbIpc8Td/s0xvXgmRzw4i2ECyE3vSnafC1RXHzDB+nmrr4XZ
DJnKRoYiiqKmqcfHfi+bnC8nYdC1gox7YLdR3CTk602F787pJO4mchppzT9Bj31xkZ41Qc3IBcrI
A/tOjN4iUXR2+bJKxqefPZar+KKLQTdvmsr8mqz8E2S9dbEXXpr9Bw/NsN9+rBLxZTlsvMjOguoO
damR6C0j/CbQC9YL/Zue3ZPvphDokJX0jXUNu/Nuh/57OOQmcEUmIyk/gk/bvWXAh2iVt9/cKUgf
GgoP29RZ3PeAFoPKexU8aJwDunCBOSU428tSw7Neu6+XE+VlJJQWkbYFYDf/BYpFKWPYNAkwF9JE
l8DgG03vltcvVooKibWokB5BbVBUSb6cJMdDjbLoRyifRDdgKyK8n9M+quewTlksL6H+qmeoGo09
BofgrPmOfZXg8+b5FBCi822udT3JAhAXArkrowBp5qv6aE9GF0eecUAVydHg0o/o10dI9pgkfML2
2mLJaWi6wFrgO3hOUowbji9OHBR7bTptTtyz2stAvsZF0FYRe5K17y4/VUq9STwlHrokVF/wparj
SclSvO7hdgqrcTaTAOgULhx/5EDEAthjIQlheW9qsv6ZWReVeAK4BV0IRh9a0YsiK9cCk111i9AR
vvcFP3V4q7CE7eJyMpX7L4HXBuY/CZy2Mw+XDF8DBuztKg0EYSbePLWUYT9cJVufbC8Gf6RuiJ/Y
TDq4dA8Ofjx32iNfCDT2Z6sGCzYmb2fFFsFFGqJoEpWHlUqxV4e7DtMoGTGzfBlQcKbpWWmpz4uH
GWBIwsIzGvNumhYbZoyOW/fsDdLH/Q1UO25Gx5w3NJkGhdMDc/Suh0t/BzaezQXvavDPLZ7CWdyr
ex7JXqYUZ5ueHRDH8+h4GBt8l7qyDpEOCjeyqPrdOPKQKhpLOk7csW1mfADNBHNLZY0DEDjlkf9X
J9vGJ9MQzTKd0nwrAPEDgx5auwo1MTz9t51WgUAPOKtd0EBv2lHpLI8cvCg4o6bMw6OqYh1WOLe1
aMPR4GgUymItFD9rZisJWD/UPT7KwOBYjmQYa7mGJaDxkQYnTznXZ5MCKsGUflwHPYjCSG9JMSg7
kFzsOEvisrpafieAtrLzQ6uNtfx2erubzFO67rXdAIoy5rxf6OzCgbvgFcOg7VhAFgf4bJHrxhKi
3ZGhuOHG342U0HVaUrx/xzkaxkCJqHMV1nSaKxX/UlaQb5slzPpwfzPV7758qL/+Q7PKOXtd/Q/1
ZL4IS7e6h4TEmUywVRsMqN3miz64IVpsdIBJHePePJ3fCmTK9zaR9NLn9e8rFCJPvQHXz4rgp0f0
2ngAIIBwq+JHW/gdxNt5Mad8e7mf9mAw2agOyF3fYVvB4Po8FAfqAhTLuTwJkZoBbsO9xmoTC0fv
GvydQR/H1VafNJrBJLQR9hztbit9hPmVG94FNBOHiXQKClZu+c9DocOLXHcWZ1GiIOgbBhnMBAuh
GJMISOQM7DK2pDYGBTB+6fiQYC1RKQAZkxgEugvYCAuF2EWr4N7RoQDS1zG91dlmTOomN0kgkH+K
U334KxPCQnKLtl74Tc2c9bIgdDCy7jHfwkoj4jY+FRfTd0PXcEKeJULsJGgBeipNgWtCfbQEVz40
NX8myU7drC98hZwy6HHmjp89QYXy9v3pT7387G9sBmdnVDV+XYWlAb9X/5fcrgSzVjpL/37DsLb7
XbnDwEqXUVx2NwYgDenjSWHC4FBtjwcVAGa6TDp+JfVF+Uzr0FLP5ZKE6hKIgh8Tz+YJTuqpfECp
/c4uE5ARCnvlRocRDmK/hfVjFUst/fvpdEgw4pFqYmOM0UmfVZ2YwG8XkeWYqvPHW+c9JNcvWH2W
pcUhmgUTjIQ9XvxIuHjxg8L4GDjy3IgUjR0lgyVhvlMkUwVRFzKMmO5gcNFQDhKeHMI02G+ysaKh
R13zEjo8ExWCGsq4nZNI6aeHKfGDZMVQOO1ksmBK3u8F431mBdck5eD9HyZeNcj2ica1D95vt7PX
f46R396lm/0MUgnj0Q9kTWD7mBfiL7hkGWH7nFOYdixlBjdEgGRONbN9XNECffM380dK7upIP+I4
dFLqOTCK0WHURh+zRJl+67aDTppB0ptP0/XyJV0b8uahDFE+S4MF2NbYOhqiSopqc3SZWK/XycQi
8QkL7lmCKPemit8pPNAXIntv5/aagyFczWHn7ISKjUu0VZfezwLQlRXjcZQmmwEpqBZs9UvK+4/v
kFgDw1iFP/45Ej/9eAZmFHx768D/eBDN6TBHoFCSbmhoyb+s9n89BYlW2O4Ul7buwYmvpSsvLEyd
TUQaC86ucaQzls85TEG8p5Th2yPlAT+2gqk+VeGVJ6qkicszM3En7enqsQHlQBtf5JJ3ZH2wNswH
Fiqe6PH5gJdfw8Sz6EkgOk4HDwXtAnedPPZTVTBz/t8lkLegzW/QLU/Wsg65Kb2NCVkLQD/swkKo
RXw4l/xq6gbqnomcExeFazc6MZLrLOgIDWefz11Sg6jGg5lN2rndD0oy9JrBfNAi+gTL9LQak2nq
+Dnrx6AqIaJuJ9/XoRMGLQAGIb4cONuhITCJDMsNDv6L0Zudhu3l/q0SAwjQPytK1DQKsDTi8bVo
24IBu9RB+4K/nCwvHQHcjoIFnrM61L4utKjNHGFFGCd7WEDWYmJnJF27ZA2/BNLAq2DxowC4ikM0
s6Ogqp0/HjAucG2gp36HlQQICarQMxH66QMSKpqW6wSRegx1SDRmuNb9blyj9JPFQkWKtF98ddmX
jp99UtN29485mbz2LycMYsIxqm4wHJZxzNSqkXHDHLzMD/hPOIaCWGB/jY/gBFDclkUNMr/Al2xX
+1ZttMHs6DqqEBk9D8UwntCwIrXjyyy+Guy1+LKU2twNoSvQoCzXunfI6ExglcL6VAAvdJSp3a+N
c1mgeItLTOpFijXhJ71uCupB9ntf1hP0myeNQpQTvhVsfiP6IiUMbarqifk30q/N2QJp6IpIFTQE
J1CH8x7k8eJ8pFqmGT2Xlq8jUWdJqPVNK8ZZ7alsyykjfbTyUJAruRLWByHUGhw2KwiqvlWXtzIY
XeC2XBbBontfVSGbBQ/+f9Mo/+cqJDuRCdGHsTVmjp2ZVT8lttz04NvhT0sBjo5tDsJUV/xHwqp9
fkpQ5mycnr/WorqAJwBRX0G57JQKjG++rQX8T+asDQ6/9tzGjvrT1fwL2YhA1sg6fYhikCkB7uD3
2WaAv/PRFBV0v5TrSgTvdmHuLF7xYLn+NdHuG9Qk/vQRp7iaszeaxVx7qNaaBE5KqpIHKyMWY6bk
uz0oWxxs45+mo6LeJaFJP6vnRK8+P2t9FNevqf1eURRjoaSmEbYHdMD4hvil/6I1xAG+Un3deBnY
c/49RpCByEg2U5k+UC3QVFCXlGWZMtUnzTmApByp1fWNKoY89uEUAU+gRFJ3pjRo4AktKBRvW6Gw
eHEZhRDB+SCmQKYRb9nRukQsTEhawNOaVHwQsPw1dcI9sPs78dFtAdtybM7fIsuS0KrMbb/R6aQs
UVqLcUoR1/dzILhviWyNBS6ZRd6NPFdcowCUngrQztpvOIdzVmSctE7Zt8BmPCyf7Y1lC2Oryvzu
pk1jmX7AweFKzvzhGHoGZxTTVCr614SLKzjhJeJgh33qfJ6AUxqdCX0LmeFKelhAN5MEa92FIsKx
LhpvrveTkfUVqSfQU5T0+q/6W0YJCcsqsPKkvEihjotnn8y9Q0S69dqhyEbSGF6md7UXjGGQ2HOG
sCBI39Z7DlgeITvi11ZeCFajReLunp1wF3ofl/F9XDF8ZomZZJihzuCj8R3RTowtl/ka8xWhtLtJ
qRaFvZCVXdqNTZ8TOIJb+Cvw6UFUU4z9WjHH6xMYzKcZKrbsXkAR7+yTGRwVdRs8NgzSvRbSK+q2
6aljMIIk4RKo86mpH21LqNKoZJq0OJW5LzGhsDCn7rMAGihUf9LGE4YdSrDaxZM08FGGwS67ADje
Ga4o4rOEn5GhJMubf6bwU8STz9uPrnWDvXO0xZz7/ZCYZN0Xye7Rzvno/NgAGrGHEoOgx7hLaJgQ
g6EQU2IxW+R3skJWBKM2L3zFqtgvy97raABcRqNUfRPWk9nueI83SR8AlYIJ+SoHO4q+9FiSRn+c
TYlgjPXLeB0WJKoGpqrMFgMKRYFFddyGte0WC5Xm7bT8OuqJ3EaZKKSEwy3UIDeRWmZKUQipw1UQ
6yRAbcY3DWK1JXEGL7Mu9TpZUwiW0WCu4oeefLRiIWbCZsdWkt0RszKmlfv4qSm5Y0fCCrmvdRy+
y5/9lbq2WuQ7QePAfz9FK5Gt6WhP428RLMHpNitAg8/zso9iAf97h5OhjNwAOnySwcnW0b7EwF3C
yKu00Gob0W/eaTbHhKKxP8QRMDlR4SIR4+apiUXna+WKp33vFl9opSgVa3/3vfXBAv+w/TVEi42p
Djw7IRehguTZ8IFSJWEjY1I7z2FCT7V8nS9KEY3UL18abgJGIIw5viABWN3ev8gJmaeImfTCmsO/
2LFWL3ca1rd5XQBp/tBn6LdPX6SEoWRNBENxHWSXMy6GoEzxM1AfDwN323QXTsaTZZHtcVrszyz5
eb7MU9CIB63d1Oak0bMttXDzAb2JSCPTeBL8Y6BUVoz7Mn0rhD7BIKOPz0X6BcewmKxLxQCXR6fX
LuggoUMqhLjq6zGnTyFVt0vqSoB2sBRkK+DaHDw1ozVamvmGGeHTc/kmBjKhppc5ATRCTjp94/6s
4Q03VZh0C1JExd+xW2nYAPAyaTGce3SNuoyjVm/+jVVltaOUS3ZhV3679Xj+pR0BK8W8Kswrnw3x
J0nm/yhfF86fc0E18EX9MhnDEJF+kONovz524Z/IYf+K2tCONv06kylygULLsF23TFwtjb3EDN5q
/opMFqnRWW4mgjexALl9vcCEl6Zsb73l7PHtoRCCJF2nt3zIE47vVPX5vJP4ey4I0GFnMdFLOt8b
trW0ixaixTd3+1CQj/5axLqPGPYecM4zj6+lwMRzmGaR7T6KJ7WbDEbOLYaoMAZNfzDyJN3+Ro2b
vO8qhYV8H7j5Kul7EaxiDRtZ5j+PFXOLil/SWXymwMq/VUC127fXRa29y1vkdqYDHvAfo6mMj6MN
XZ7m8TlX4dXPy9kOW5JQ8wryFB+hT0UmD//EdXUsMb2v6LJP765hNepvnLn7n5DZn8D0zfU/XgMv
8r87VrHgHIEgR8pnMSAJj3W/h00CVKrU0RcyXezQRvXBb7s7vy35Dtn5lIa9lVuH0Zr18ko2MEL1
vvLwX5YMAnYvumMLpjMPveOP6F8pu8SayYopMr+2qoSC0+DbYhlmT9LZC5Nb+8aA7BLtvG8FApUz
aZdn028XNjdmtZAt0zQi36ybnl0kWs3iu/t8i8VmWfAJXKwh7Vt2mWVDbkJaasZf6dFCsZW5o5Fr
kcq5tWWRyZPK8EaNJbT91SfCz7Hft7IaaZooi+PJqZtZz4vw3izUUU3eIrUk2kZWzsWyqYMi4bzR
DXsqVZeQDeD9P2krFEH4aFiM/d29qDpwuf26R4Gj/Btrw259MzsQSsPRXO/1okCSghhDa2wViL/M
rt3rDndVrrsyf1Z5YYFo/3j0p+tCNhUjzyHDcakGXgU7vIZCAfNqBr/LdAn+e58z+qtaqs5GtniZ
c2+1nITStTxAqVHmiZ9UHFnpZ2ONoMEaB7I9BfiZIOYPCfKo2OngIsBGAwGqYwHhJyasRDar8rKl
+VGfoaSRxoU7++MQGaNS9px4pLzj1t6Qb4zA8qVycuQJBdf2gZ2qFz0MZEgxUKmegM7tp+iCdP6T
COSGTUdmMaxWAszk7CeX26JfegMTLuI6Dos0bGwhgY5D1m9irZbs9EsrDuoZEpOT8eV9MnhligLW
2w/SjImchtvs2lOI0v0ivDCgS2VZ+XzWgpwKpCP2uPJxcPtDPSEGYMi2sFLpqJp1j8myMngPo2NG
jo2KnteX1cA5fa0UX4fDUXuPHNf/LeG9pg1Y7mqPDvf5M55A9S/96WbmA1S72HxJrdV+zlg+bST1
twd+ExOf2tG8Sh8oYXNGB7cHh5hykVVJpapd5+ytofq8qLvubv4pl/ENdyXwffdhgBB4q2fMG2b+
jCfhY2qp4tTX6+2KT9Kj+ytGW+OI/uTr0gj19zSwsdszu7zYy/PY5TWImfQ7758YJdPpy9uCB1EA
XA+Lz2zLmMsoFH4HPLU6zufqR+l9u+OXPeKyGhUn9jwjNr5xtjCv2v22W1dga1tpZDH/aMYCzerB
FkzBil33PWdZcTHpGSVKEdrqZkSllEUP1zT8xvIm+Rh8HmdeEbaUYmbrx1hVnsmidgtREuU9t5qr
GNXg99uGeCUnWQD3lrWtoSQ3h5Ajlv225SVY6F1pOVKOmxKTeQsOrJ1qpUdpS9HkQef5FK0klAjM
VNyZ1ejZpbFyx7SRCVe9nSjg5JK904kvo9stVBJ9r997QY8If8VMW+oerEfdOnX8kzq0fHvfzBv1
jY45UWPqrMVUff+o/vhPAffUL0RSxqr33QLTSGuZKXD3gndiLjP8GAVe1Tfus9pEkUiic9dfXD6L
MOoxkAalYmFDj2HsUOSG3zXKnBHBgA3RKPGZB6O0aBq1xxTH7DwxfHgLPKNrDVj+JDu3iRlHwtXe
3eeKe56pqDHyOBtZC8NZGaSBPzH+tAJbyIf1YSAY0kRQodptH0YpYfSzydYNKhtMII0ooHOj9uqN
1d0xpzolyTCE8qcJfDdjtAtD5jTe32x+3djaxwvjaUNlsCqJWMsRATIEPvnhYQ/HRN7W4Hba1O1r
DsA5a07LtPfQ+FdkJRll7sNTWyC/L5p6EqdoH+I7iRSA6fytMb5b1MLyjuTY5Oj/gWJneqPK85UI
PHA5nHKEgTu/k5juCNxvotFyJJhWXX9G3bcoyqo2UlJw0IWlH9vQ0tE5YRTzJcgCKsZmKa8p0BLj
zm9a4RdWBbSIOYVukxWK1kJJ2EaavB4WHLo6Nao7sCtFu2c9ElRxovJlDDO/m3/OLljL6WNnffLE
dk4H2LbKEZTUrj87Ylpmk9IC+K8uAfEZQNZ93B5cJDTBwOj8lnxZuc/F+wPFyVMUtpPWB0BO4EeQ
FnUzV/Edq3CTt8YV97kqWfB3q8Dr2rOWp+kZICTmBn6xQib6cmZ701no1G7kCmtXqsZ6ud/ewHck
Q6qQsygy80m/2HbHU7TImsTbH7LGEH8Gy5q44oC7LpxXK6QOEyQyn5jrlij7V+mA7a7nWNo4mORm
lIZqqVKGAR8tYV5bRKnrIqFIfGEkwy0gEwq0Ed5+avWA1s+J8prmsqURjuZzZRiiP8ivDdPcoj4g
DAJ0+a62vGuJ6kCYuW8m+U423POILbFeG/mRYUxgCH02r2VX6CFz1Ei2c1aUw0ZReQLCR+/sOAzm
V/cP6rr1yWs4r/yRTpCDYHK9oM9bZc945WCOyIMx/6lNyV8UD5g39cO2w2hFOy0QomsQY4cEXT5h
IZbXo9vL4F/Uq6nIBL19JaVywWNJbPssdO4mlKgrGpnSY7bhf+rsvSpI5/1UJrVNHEUm1RLyEJJa
b6l5C7lw+tWRW1R165ccRpfBV4aQgh430qofmfXDKJANLv0b7RMnkqMYiQdJ0XOTfRPiW15Z+VEE
cQJ5SbIrr7FUTgidiZlDNyEy4ktbXqeBN7pzVKK7aqJsiRAfyaC2T1FWHsxrdrfWP1BaVtQHRwC1
3yu+1kU4PILIZv99oh82vHh82dKZxEZdiJHjaNxNk8jj8nYTwhF3c99ToxR7Di3DD37gUtBuwqSK
t7qpgkY508YYqOSM93ouzSq2iEhenjr5gqQilVNN6z8ETGvEh5hgGAHUhr7sj29Nw1KWjI0xJlZq
INSJYOKHP/RW/nxislBQzZeKlkkZiRA0wic/MsYh30hiNdYbuZI/I2hRRfdXK+2GV//YKdjtG+H/
xB0909t8XcEyhR6s0S8RiQfr/pk7FAQXxMWrdO0Izwwy5soJoEDsGQBWUAMFMR89gQPxkkfN9ZRB
hbvFTH3BX7oVO77p7cPrJrQF7KX6B+lWCWo/GfPWeco5/tzPAoUI4ssYbpxBQ9BaNDjMP5ot2jt2
DDaQ3DZgO1NT2QBytpgTumvIGd3O08j1Q8r5l0lkHJBaPs9A3HSnrHx4ZwotOeDFkyqJsqj9MBI7
kiJC8bWDrFH7SiKe/NTzuzORMTcXnhkj5+VWx2VXjlnKwhDvQvtW4HxA7Ump2syavLZitCM+ruUr
M/+QWs3WbG9Dp4HKUuAXlbVB7XvlsSrnSZ9NihcU/omzS5SEvyjuqsSpNugOMTOWINQSFlprwYmL
6t/rZmaTGzJnRSe6UT8vdGt77TtAbRdR0jd1lMbS6uOVTKmuXR5BEwMGkZn8qn+w3wlvveztdLTk
mbncbI1C58KuwOR31w8E77kvlVNQeQZkBy2sE9ZUUbFN5brHtisda+pnKLxyYim0zLYs14ixAiDN
SfpW9//KvpEFiwUhsLYeCq96ysxqIK1mAshfnH6otbwlRUmWojgZq59l7nHGtIwVTfVmAQ7WEd2t
62o7M+HM+bpP4Meei1VzScfir3OBZ3MlAU+vucAy1+8UhI1Qk5j/sOZt+y2yo2K5byweHgdNesci
PvWANzTPtAjwjhfYSwqSXqEToqHvQcWhqFX5Dv/w0YU0qnqEKHTdsWqI8jcsuTJhohOR+s4q/IWb
pfbd35pkzl2FGIprmGYo2PmI8GfMjHnofd6pkCJ3ThrUQLjHqSJHQpFQLpGcLAHiyYSd8jahoMJg
vnjwRcbbO4L6SNkp9YlxUDvUPwPtjKVuG+O4EX3SH8s6ggXbkfoXt87lh25n0JAw5qerrl5K5xYF
qynKMpblf7/O98vkqHY5tUGwN+o6UJYPQREFYTXxw9kAUfW0QGRC5SvXWJKNHyJKODAFJIregJbv
Obn6a82tIcV41GHf/785JO//e/INI2dM6XmUIAhGVKmcKGOrBWEuuyKCXpu66zUo2UwuMZqdyXNW
xkPRDjSlxP1WCR+4I3+a7L3CEnM7S+M/x7fZRqZE6pnl480EVTFXMswk9WjRBMNZ2fbLUqhusIjT
hj+BnRSg+cAH7Cfn5yt2K6J3uPEeAdBebL07aaV4xbtrWma4vtd0ynfvqQUsPj0ZCgwrD5LQ874z
W5RHAfk+U2K34eqKkt5Q4m5yiLNTYh+Y+nJobWZzPkD3lNCNozXKDY1IhP18Ig81ijWX5sP1HtdD
GldlD61PLZ3XgE7Q6PPpVVxTC41pMW1rEPQ7DZchRPEpydvW4Yvo6WvaM93CFHCW47BE+nUx0LKD
Ob1ZbVj94nD41xxswAVmnqU3SczuvpG7qBUDo84366b787WQv+afl4UBCkmZiizGH4C/zi5Ow4z+
L8iOS3v2dpODZh+y1nFL3Ou0km78fMkMP515miM2DgUFeePLPQm3hQmwIFlsMY+RckjsF6FD2HDh
u/H/IAuXJjeHHXPCuK5M8xmEXvHO+A2RKEA/WEoueHqJOE3KjyAYH+dYpzywHeO87yEQInZxVKOz
cn6auCYbZplT8iHcR01nVVf3GOOfqZ/6zWzUirrezyW1c0cAYMoIWwfa3ETk54OHhZeWMYDB/byD
BfSPHZray6m7qdmvr9eQ2S80+KfNjS6ewSOz+sHwq06lOua6WB8ZODRL4amrCLoR3zRJ9gBG9lst
bNsyLoU5Ml+Q4pgA48VGie74Ed4780lH09ihJQ3BL8Dzunt3JDYIMdi9in456qJPDpBq9dvN8/TE
+6zf0yFucpm0VBD7+mZBTOR6/Z/e979uo9ac8ZyO52wquZN2qgqj3Y9QBT9QSyqObBj2Ar/H9MuC
lR9VZpur8DZdx+GTyziEubyyrD25hFCg/BUxfdedODy7XRb3HQ9oyGxsyb/WUy8Cd3jniLM51DC2
IJLtx0zCDi51AVfSlIr3lLnvXIW2nQ4Y0f5PiLJnzCdncYT9oCqtv64pIbMQ06SsQWK7yWadzpev
iP3QEMsm1920oEAvlkXwgVCDBTJy8gEmI6Eb5rNp2sF+ER+kf2OWnrv9iWWowQnCSBo7O4RO1Vrd
j97F6nHFRw5FCqigZNPJqzClW65cji2C38xuV0AkP5GQgh54zWwnNjAeFm+dvLHWjd9Q7GrdMZ2R
hGx5Sy1abd7WIL1blHN6jtxAp4GWc1WEbjr/QYNbou8txsCPD/c5tRrlUDpZ96Isgh4K0x76MjRe
P/kyPwAxdebZ7VWON0AJQv8giPFoJvs/odMI0sJzyGD4kCUgHGR6JnDBmsGyhgFsvxgjXi5gAdh/
Q5Qsz+hDD0+7JvCUpKXBariY8zLbG0ZfWUeYizO5X3nHCfNpBgZE+D48NEBmbL9mA8Gm6wK17xao
P2teLiZNxt49urwYAkf4dAxbPwKTTqRnmj1fw6YabuUkvWaBFT1DwlnhCVrrbwOLHlWij+j/F/sN
7BT2uqqMEUVoiPPBvlp7kMCbLX08ZKdUTE2PxphYVsu4lAaAj2ivicLLdNgFa4vSt+KV4HXftFQV
gDGTQqYhCxusJikyzGSjG31aax6tfP3qazpt3xJXvouwSjGIsTOatDPSZrEjDQT/zGVAiphcc1ia
ujepUDyW5I4uQKoJc1CuZSatObRio+CsR6AQFr7oFTOnc07lpuBnHTYB9syezcN43L9PNWceU0w7
OCGmFEHxcb8Y5tIkBSJD5SPYAYYZVdy5G8ZpqE3D6xuXJA9bNlolBDo7bF/dzjISnHns0BXtIRxK
R6QJhuCl2o4jXu9RMnwUlo51GydSv9mrrAnJbRUtp/D8PDybrZixMnYYgozE4ZYXDFYI+42cdyyb
Et1xFLSSGpyGYzAR7oC1H7PM8AJ+yDwZr1j76f/wc1uE2w/hr/G4m+X20G+Nxkp7cggJUzlQcHlc
WaaiOEajqBqOPKtXRbEnI0KCfiogdw4TKwDSckFXE1jSE0fwXiFnjRnPoP08aLLgnVZTO4tyjCXJ
RVA8meAzDlqfxIBtv7UFfC6vKk3qESAGGfSeq7ftNKY/esEtxG9OhCyaigEi7C6QQOmB4T4WZlYv
95N7pnC/Z5YqAYKRa9+u+TVraBDzwVm+4CdwesLOyJecdeS9pS4jkftlfyXRYFGQ2h0oA3hDunlU
ymxPtJWxdy6bFcj+yD+MrKoXygXTXFgcnQrMuFJzRXL2r147182tUkR0mJ8+tLyvosgdv/bi8+qh
NsggeryaXwANg6J7sKjX4TZW7qX++jPYYx6zj1puJjkFZM/HFa3DpRb6PtxVbEUMhCy5zbRKE8Z0
U7k0rc66br5z99pfgLRMTGNv6Qhrx6Mmb/ydexQGjS/1VUS3YDvzcFDRx1FvydNB4N2axBNR8FVu
N58tUvgAJBVH+FVfGd17pJnu+nkCerFJSONOKqiiw56t21WFbNDI4NCFtzAVjD5KV5JVuiiGIgp1
98X8X93BDLnd+AJ4f0SLgIfhFk4DGHAgO2jZm4EyAo//3BytaUGzpCXJw1ax23d6qW5HppGYAqa4
mrMxPxQMNGbsQcqHZ7EXxMeKmR6afcnIr7R5kFY4XrZdCHQC+jb1OhEtfEJ5QwgsZnEJWnGeY//P
mYPssPnMCcZr4xYItdypPO0P4kz89/BP/65DWD1UKYzanT4k4HRFlHWeASUgE0bCYbt6rcpEYiPc
8qL9NA8dZ1YO7kHFwqDyFybSxuN1IORhxuxgsvAz7axiLtQKfKaBujVKRbctFkb2GqGyN3uca7pn
qcfAoYNWGuToF7S5UA6B3ej8CBOn+IjZdolbXcmo/feyZNnCdl16wVFnVGiazWnP35BwUyZEox5+
VRZOpTX0IJw/eLt36eEl3M5jNfjDgFwN8DSsgd5/Qxm3ggbgVuzPSa6ChNKGFUSjp5TkkrCA92So
5IQJsRRnp5sDPipuXkQnwODactex9kVSBNWrML8jfCtbZA2ISloG9Jm3E6JuKJ9WBNBbCxeR8GxL
2rc4j8e48sqKBiGJKeChjSqaWdYfWsx9t1Yh6sHAvfKY1pGGoyvfk0gTKyHVWjRixVvJf0kFctIO
cohxBTLT06Zzlz3+JLX1SxFsfuU9GPizkT+DhMfpsUfflze/vNSEdPFh0SemLXJrTwUVZ5NGNfeF
h+HbQIOoQwoWBl2obA7alttNfy72SfqwRFutGM+rssH23JCImXC7B38uGeUKZyT0A9RSFSQ60NFQ
5Sa1lMcQeqOOkKUezncMeOSpVDOBr59AhBYNdPR2c/MQ7RMooDn6BMNsgBexMjwnPEFikCLIl1pU
2wxkWftMfYkWhoKNxcjGlBhm/jgeHXw1fNDzmua0Iuz1/lJXOjs4fooQL2BXbs+iaIFAcS/EelW1
iod6Kmb67QSFmlbM8qthm1qSwYsUylqM1i4EVPLRfPu7pMhPBRAR34yqJegKcgr/HFZ5SNgQdjh2
UHaD1WDHDZfq0iiLL0SI8Ja90IZdzFZCviXMJCV2O3EYf+ahHaJ7SJMp5j7yT5T7+447LtS4cXlC
2v1z2MkpGKcdGNeSrRkJ/1o8FYC/60gG0ZY7cJx4G1FutUiSLqC9xKY9DW/L+mu3vFTQ1aA5v/lZ
9WOArD+4Ym/Qjla9G5HMguXoDShM0kLumXgME/eVgNvCZxNkPa9zSjz9rbG+YZI9KcGKmKN5Q1u8
zpiTCcdw2CBkpd9Z5Zdd4WUkg9t5jicqH1flasv5kqWNbCp/Ibc8cryfzBa+gPlQyW3/dJila17h
6m3sEOcyvXJ+bD8h3smxKrlgDGdhTpsP/AMaZ84QnJsw0Zn7hwDoyppZpOOR2xghHuMmWV29Oik3
ouIJz+O/V0hGpuqp60fYFe12MNLjw8DRHWSXuhpQU4bz2dgPBhUyYLEyfsi+WWorQuRkIleAWrJC
RXBpkN8ME3zk7C/23kXqnnI1fJR02C5mHTumWe0HKBYIqscc5a3oY9ny1kBNKyYIuxlt3NJpVlXA
3u8S0oMDZ2K6R1YVWObCD59SWXeBh43BEyia9M7WlaZXQnhsXou9bAlWnezfJuiYNv4c928uJHHG
rwWmaCfkyKJwwjsUC+yr5q993UWCylUCbAWKcjULfI7Vvp2c1B8KBtC7uPFQPoPp2RsWMcLpOZDg
ozA42ZlCaVj3LkxCrM+ZpMGlNlVChP/ahA/IbJCxFckBlStTYauAWtzhyukNVK3XMSZfhAdRKR7V
PTqDohLivDTlw3ATprE1Txu2CQkA8wt7Vr0263EQv7x8ZqZsH4waznUktWtUJdIEXMDzSNWQSt6/
dN2Zh1TllgXk32EdrthgMERDHS+BmQivYchSZu5dyrMrOAaZUbSvYGjgy15vOyita53QwCH+/L35
oqlB11/ZVxj+jniWdmOJSgwE1GItioJ3YyKtTDUrCFuUwR1Y90Sj3BQUIZJubt1jBH0oGOwToAnG
+jbVtAg8rdP0PORjGcQT4t8Zc9A2HEkbUL8KRrt2ZEsm12F53C2PHtNtoz6of9VgeEm8gppAbxP1
ZFjkdcGddzQpTcoA+stkQQ5Xj7AemUphnszIeOr5Om1f9N04vKWujzkik8z978zAacTTlrNs6D93
WWArK3SQz2dVsJEicR68HpkSgFr9yEAuPB/syIgkHFW0yvxyHwJl7wrDfKqjT2mELosrcITumlfC
yZJbe5FgeSXhHrRAh8H16bloPioQ22N9HHKfPj7DJAQ1luIa61L+RJ+ynbdzJ1DmyMS6gvZ3UaV9
O+cJyGrPIFPqfPIgpV27Lrmly4XXJ/bAm1lKEaCdFDXxzU8/6AICotzIEwKwmv4DKM70Aaytn/q4
jkp/VPbQLuQA15vH3A6LNXKf8/7b5QQH5IrCwUS0nj0zLoDC8YtpKMLV3NFcc3RZKQZ/VxevVyXD
iC73OtB6fARxUbkZeN+ZoG8RYd/o6c99FxpQ6nSaS0nFttm8OKJhafJ3shJmBndFrlJOri/ZBbSj
UtuLUOcGdbQFv1baT3f//zcN3gf7jlO6kLNr3wbpScNPLmFuN1lUBWOZQm943IDoo+LSIiupQaVP
YYT2SyKwVu1EEFM8G4mY2npR9uWePvolxjhQ4JT6H/+utYx/dzG4J8tVjuQXhlXKKa/242TY8gnI
3lsoAONDhxWBuyU6rAwrJ3HPMqB14wfM7X1ftFFx0BspAKpRz9Ex6jhaqHCzD+FIYjlC8uoN5Zvt
jDf42h67PnygSMiRsRD17vMZXUXORs37vRfh/ZePGAPb4LUim+q3lzMcy8qb7amBzYYtGMNZ53J+
D5vl7zehuCRkMPJmTDOZZquDcLrX9pqIW9MA0GRoJfQuKwD3TWUymTG0gt/yc05XhuVF8CWx9saJ
Khi/coGMuul4V8KgACZssoP5PtGg8sJKCDcDWxIApiN650XLhsJD912T6rQLiyjfO0Z0Rf2QPM67
Q9zbNUpUhbGANi5vixNMfrep8vXy0Bu8MD3i97hlpXSY5ARbACq3xAG4Dk81kF8IIPR6+4hWX6Oc
70fvFD5/mD9er04PXSHFM0zQZyzh9UR8MRehXFk4nlbsvUvy+58O0nMrgMDVriCNmQaMIZx2lQ8b
jz7tIPjab9dJtV2LWQWn4exwN3Dr4LbYwRwM0BwCcgpG98OLRBrQ5J18IYzqXFELM47OehCx+ayE
0iiJXR+9kNTsKkvDS6B92DLHhbq2f+AAz5qsYa7R5d+9brmRWTgav/7yvwpzpi8SjMqTVurUxzmi
djpBvzb8dk+KXgeL1Ab7S02v0HzUjX8UqRbMxu3PnmR0Oqqf1sbx/sscJYV9cWXVYMlzi3dXXU+z
ZbkfpVjLztqyj41Ygk/WIPqigrTRK/ZNaFgAy+Nd4PJpsq3gtiiESeHO+wN+LxVaJOwQnOmjInLc
fI1tQCEl7K5mfvWFMRrj0o78e9bCR1B0of/Jdn81vBjBAxt6n5+KqWIcsdCU11wk5yxdwSWIXnXo
wTw9/l4QIQ0D/ZY9hGWpdFQGdaHu+N2LTHJRtrSDjCiP06bN8XGdg0Y0CB9HOwKh3l1LumXQJCHG
o9QyFF6krDYOKmS1DX0dprlDvwQg3CsXgMqwfW9uZwScusK+WPgbd2za1/sPg0TvK0ub2IPe59mz
UZmc/NqhFSHIUKpCpPPp9NTOeY2t5WD1DknfYUAgcJBW3v16s28dg6pDftLYDwpQvUXeGGoVyOb2
M2ZnLV44k1d/eFXCuSIhOw/EMbrzFe96n6nT5FqJ/jCHMMlRYc/Fx1e4DdtSgciuRRkwFKOhjsX0
g3tMdlA9jzjHOzK8SJeUCRjx5Pbtqm7oOQ/kpGEr1kb6wTZF4488t9jNiexJ7YdBZ5v0UrH0f/+k
18sum4Gvrh2j4jp3ODTW9V7BZ6fPpr1lF4sM7Elc0D+DEjc+jN3jjsicy7XNm4qi1wQaAYFhcqIt
UT1LvY1Q24aLwYyOX1CJKKRdIkXmwXZzG6eu4Gcln41pEZ3byIHFZE15sbk+z773GJ5G68guSGNg
4enncdBpobwFD6i1RbZUpxfcLgZm5MYp4CvzNdxCzlVL/iRbnJzv1OuIMtWfAPvaXqQd0FwhW6We
ghtHaQBtPXj4N6s/NkgUOoXpjk77TbiEVDakQZ9M/9jjXr+WBDeNvaUbJhvX8SXIsRuae5RTJH/x
4uKUpAsAsoHn3exxp0korwG/gh4fQxrPMeNDcj6plF65Gy/YDq9+E2qJhzxl9jqFVlInxcH/XWgf
VApEY4DMfBjMxoPnD6g2INsIwqRWiTwcU6ZYVOe1jjxtbF5kgJBUtIuXVwnrm1lV/EzJeJJVM4tV
OE1PS38oOdZOfAxWmaqbOLOxSqP6G7Vei025IQkf+3FOCF9RzR+wyQuPuqgv0pF7ulqvNBqQc3mV
OENFivJ8MbDLqVVY8lfpQSeLvxh0UYH2oiNwPZl0mvTLwv7I9cJBbPAdpMOhIsAhEKGMFOr3heoi
0PCEj9Ndl9oH7hXwMHyV18/p0wYp2phv2ooFQtEcrltAbub8qUEVWp3U8BnPKnnu0x3b1kaEfgBX
sJNgHRt/goo/AKbd49Jo7o6uE6IoP4xAWdXTytSXcLGOGbaMM/WBx4c2z9ki5I2h9DkYP1UBISH+
y9a2ABO8/nMISH1dH/0nsIOzaJZDLp+WBDD1T5esOu9aoIZjJXj2/q566YUczo8eFcCds2QUG118
2jI9Kikx9aGPV459+Jm2HDSGrIONRt0wmDxt93QwcCkJLvhOH4SyO/YJrgbpP13BIHaIBJkXAm6M
YYAhPa2/HO3i9hDaUrsvjcBkzbx09JyVXSemIi1y5KuL/OjQslc8xD0o4LYTs+5k9fa8yi4mT/c+
yIuEvS5sdQnsRMoC4NCpyUec4+ENYnc0A11TpPepIeO5nNnXasMg8ofiviDd2pOShtS1Ke9fINXE
YMLLnQzNkjOtlQ+OvP+M1I4ff1CCBvu2n1Dy2g0KfM12MHRrLGxVPDhPjXWXDjotdAD4VxoXb/4v
kagHh1dVecmftYXlDLKkUW0KmOqeN2eRK1UWrc2Y/IKMBMmjqkjGFU1EZRcJJc5au7BJMFXRbyKc
o1nh4Jfp+lZ5q34rGjTptPclZB3XFa41LbA+MHXaR+7R1PDMa3ovcgFGZRtDwNelBbIsYm0LJ/Su
x0xvpOwPyR0bmjCGa2j9iO1XAtLSfkojy4rOAuIkjzPyQ0BriSuqnksY6uhgdNmMOIh7R+OK1MMP
im/gg1zyMHRm9sCG1DHxlKghv1Oh6JTM7uAy/g8Hpi3xTNxnFFvWicIYCAGHSvp0RiX4aFo/Gxz/
/M/7C6yBUZQVJseYVzBzBZoqKLMLVUFnpE2Lr4sei65plyE4ha9ETQikY0DSZ9AsIHidNGixNGW4
byFLhKC4IXpRxvLbevkIgr719S8jqDEfYxIuh6Q8tkSD9o9LavHjVOzF7ZGRaQYb5cdnDAf9Fzev
ihjVwAUxaYBbB1RJE9bZ5iO0TIDiwQKAN+uu9mLQT2VWdGET/tnlFn2XuBBtxVwh+SUq04Dk2f8I
JnPZkcKZRbtcadptdxSjw81u+YLCKTZ4dIohURnCxW+6P6dOERBlPxtOQ5MfQsOIB9nlhRTR63ky
cOG7lw+CCtYhmWGxhx91MBUEFSvDh1d//RQK/Puyy15gcE3jTnmhIQEY990z96+g8Oi1i58vf1Qf
I0IWPsMYDndb++bNlAAYHHIVf3gZOMgViH+v4ib6Bt/Pu+3JBB/MFUI8KSG34AFyzB0JK05mhfBQ
EKIEd7CL4ypFOnUd+JfEOJGlkFhGm6XBWtVpCTr7hQjwlLFQAMFPFl6Uo1QlACPZsMGYHZEn0C+s
QZBQNHTUUd+IynV/CtuZZFETAvgu4YYd2xf1bCRNDxxI8sA3gdmmBZIVGtv50wQbgCUTlAPT4c08
cxxHfw8z9kOeRjtT5G9HzhTYFdsdyl72zF8OL4hXWmOT8e7M+8GKHQ3USmSHjpgL5cGhno0dFPi/
ChG6QYMnz2zkzrA/dEJTyhHBT/+39Bvte0AHSRfyC/FOIh2uQ8z9bIClqRIJggqADoMJ4kUw3Y6q
PSRRWOtcK2BMQx19j0WsCSlD6QAIxemh3hnJqKzzZykfmAStOMKhKdaSPRZShii28y6V1bWdK9m1
AtKz60PlKmK0xWGMlb4XNR3i+eUF1LE1eYfe4nE8/VqatsFM8TWw4SRdqsi8Sd6luWDDC8EZrvbZ
DNUhMLE959FDCXmlLY2EfdO886cuGZHJ+MIa024b4WF3etRm/7/xevGnWCSRdlMTK7137YGex30U
+i74eqMYbCXL8rmXafEdYclsOL064/8HK6cm5MAFm/x9yNNEKiwUEXHoTJvOVrftzOd3EFhMLVQx
vyBZDpt/BFL3qA0I96bSSXKmQnH4nBvc0XIW/XbYfLg0cWLGzcosbFLWkiXqw+EbqK0OBfMgb4am
/86x5kF+IH68cHZ0+U/N49+xS1rABX9upKXbAUd0usoRUPTSMZrU04fkzP9DgHaklDZu3TuIdsFX
mWO9PmU6xmxg6nA0a+s2B+leUWidML1l3RlORa7YpaaR+O8I8aLSvI158LFRHL43JBF6IH0qIl6p
RhDWizCIU8mxoZ7E3DxS4z4IUNqIZFnPGVzbppXuiARPZVICBI/19Sl1WSAjiJbyUPz5H7cvEQI4
HDmOqNnNsillLiBBz6rX7n1kojhpGlupJF0Sn0vB1AR+O94o/IZvG00GGXrukiOcw0/t/IQPSjlo
2gjJuPS4g800L9peCvaBXLejMr5QYg/kBzKMPIR1ck4t+CsQhiEB3eRl6KU/1Vcrwqm/yMGKMApY
JIjD81lqz+hmp4OaBOX9UfHU2kX77H/VXhctde3+Nz3MUXNS4e9mvwrwWKiJnhsuxNIqC37vBop9
GxlWx3O5I7Z5Nso5MmUZ1aDimlgrXEN/JYduYI3MTR5en5FL9+0M8QMVnIqOyJ0iHMNbmhyrYwnX
sTsg3gqC+RZ/f4NVVDSxGuPLN+ZimHK5R1OS56Kglgu/AgwQSi9gWbUzIFexsMnTNX9HzZN2BOXJ
iFdP+/Y7izEnKL+vTe5a+TzW41hTYXPavmgYPP/rrbV+grdlb7z4CTXA5CZWyxuK4z0NADxMGr2U
Wgq4qIO3DRRjpE2IWAlCjm32a6T7h0sytcv09gJVK5EfvZB7wM9dxvLh3edr2F+QlUB8cPKccluw
PXnXFgMmaT60MMV++SP8AGqOPgWS/iwl6QWdPQ+euyi8BoSiYrIkxseLIjwwkehoKLKcDC9ltgU9
2t+Cv6t1zozFnCAynXycQZRzYEpce/SeL37XhTSVaSHC4DHDS+u+Dk4eMefZ2d1lRdn2l05cv8/u
lXfw3C2wnWjBXVDCZWojQBekKOTMfY9E8byLP29d/m+dz9SNXWC5JgJX2QG0X+aGmJIB5YVvqiUF
WfCsUK/oG0HdCBBkjDfEhmqczb5EI6o5ExzwXNPHNRRkHdPDXs4Nvi/Vr/M+pJeyiLeKlVpe4IGm
3tibTGej56xRANrG+3KqVvASxN2J+mRM2UfRM5xFqAvQoneu7drAycT40K3RSpVDk8BGzJIaFQEp
mLdcqdR1TVqG+5yaCxzBslHKTeUIxPnz0GWbyXqbVtjOipplXCGO8T5HAGQpjahTA/qZezCztBM+
cyOjeJfrQRMR+0A6qkrs5hxi0Q3iObb/8pGOcYAF7lDWX4iBeobsV/ZJVAQkoFvNSJGuDoeqjFiN
GUEr2uC7QnhGpwexHeoPKTATXmLYD9qCUE9B4O43OrYqKtYIak0R9iqrCFomwqbyV8u449/pO7fM
7PDqWdVFgMr1nVqW2EzVJGZgwXxDjU0Ku0WF5FbsnFwAF2ft55SiF5uWvjaUXVa1Xk5ETYp+Bx5W
sMBxjNbQmeUDrRfaFXsFqsMyvGUF+xMfV3+iUS6SqDdZJCoARMdY1HSJ7FFYZnsz+uIWFMQ+mht1
uNlNLe4Qyp76Pyrwr6hK4MN1PYvnabKcYqMxaNSH0uQscOSs/9yGQX9rnD+fTRqV05RuArcUfe2g
EuZElL9FVvbuwNuUmOFhZNkNV2/DQ8cWsNLbIj6CPejK3qFpbjxZLIwZuBmG1vAyL8/1EoMfTVjF
jHz83GlLIeOEI9eqXuGWu8PeYf8wjomMjx6Cf9HswHY5Y9TvgdwGKI+peL3WNzWejEoexj2Eadye
+FW/adpAmB/oZNT+qecwS678gMKnH25E+xegn+riOGr2iY8i0sziL3Yl4FzTdp9WJFOuOoAJchur
AJwGNJVJcoTPonwyjSPc15bXV+oR+bJtGFVXrn4hWl+UE/0jxFA+lfW+N86xEKPB0whoAf6g/9HO
218L+7DI9LsFSTTlhF9i3DW2Y8cLXFwpNRBl1Re8BM39vY7Cv2QDt39yB/b5KHUfEX8ga9NpT6jK
63goQxnnuR9pIzuVIQSiSC7ANMdqp8AGyMimc1MDmdLZT0N6tUVRP39FHDU6fLHHoXBjmNFAF0fL
uzMJubfJJziYi/TWQwbqsad5EUfIeCJsjx+uHjBJWAEzNxIT3ARpFdjW5N+z8s+gyz5Z62uUH5+c
ORNsol76M5OM4pCGeOPdRvPhXMC0k3HLsqMZ8MYbgE5Pb3pm/qdbI8YoLG2EFZcrZHmrwlszsEYl
q7j0g5Hye3t4Pur1+mQCJSqPs0O7zNxZwJQ1GyreA0LAC9pPtvr/9bXo+IeSC0GXvibiB447wxBN
RIWL+z9D5KjKCxD/y8E/WnvOnAjI+ODNf/5ZEHGQsDdbFIOdaXfb3YwcDd0ET0EoeBtQqEMXUD6T
+J8jg7NOG53pFWOMLEJq9Ao4zxp8FEcNwnp48DnYc0Ezk5LOAA21YVpd53h+Mv+0UiHSdRaLalsO
l22Xlk8Se929kfm4/uB/JFNddJtjm0O00nxjznmKL+SVBO8BuMXIqBbsJ/GEVrsDcoLD5UYz2rpr
FAklwhVo/om91lwvMoa3JptVD7zgZPZdCewhrArdukWHxVohSY3oITq9jD+LROEsjuTa+L3DsPKF
uVkTp35ZJifPIdUXMMNaJgEe+j36j6biweeSGw9xJmnwD9PvG25v/XUQhcrAMNfnE/iTn7V955iK
L7Kbwp4xEmPk62+FwC+PvpEv6KcvY7iHCjfBr59XcEmszShi4ec+XSSnc7Om7a0IsSzeGJVp35GX
VPM8bnNZKvxeZypcISOfemWJTiwCn4YfoQdahEWntyAheatkpC8fHwwJWOEaFXEA0LwZvgOKIMi9
maUIRSyVxyqCaHgbdjMFlf4IRyHFQQPAa8f1Pa2W4111yhSAouyRTcsLBoilO6+DUM5Wd5KkOajd
riD3HcmaXWUkgsvaGBI7+scQCexr3a3utMiyUIwl4gbE6L9xmzjJY2hP9DoiVL8Xz77wdm2ovtgS
MwdySlFmWE98LFUueN15mLYBkbmBUNVeCPKWK7iIQaOc/aF2vIjuLCNQjXlNzFoWH1ELsX4loUUV
gDPTjDF4MZnIAjHbdBzdnqtjLCQk9KTvilY3ADCGJ4WQnwlxQdaQlKkEPAWs2q9mGKfalFk6ohLF
lriloBy7mDaefnAtPb4KTR4yu+hCaWzwe2Mj23OAsx4ZQhbU0yPx1KfBY85SBj+k4WxhFBd7q+Db
EbEsfVxFBbXBfSigadgcko46cXVBgGtzP8Ss8dczJbWL3hOPd8bI5JdMHl35K6RuHWK3+EZ66rFB
RuMhQOXvjwlt4gMuLmxaMcVCL8TngEW0kKP5HEjkgINQvnGABPxAxRhXaIFHSXAPXNQmrAwCQuzK
w/WxFNj6PoWaG45DyQci5IJfYeoCh+1+PsNmfiss0bpBAvDx11l/fEWJLzgGvTGtLmWddMwHKI3/
LHU4m1cGDbBA5ZK+Om6aAS063BildQVAEiwDgsPWmbM9KadsoKMK+U+aZMvOVhhUpQmz10b49Fnb
FznM+CUy0TZWvIyya3TNvJVCWvVGNMNSTBzAmwuz99ZIUpDhoVMtndIWze6ybh9e0YCGzCggUfKP
loNE7++UaDViurZdMAvmQ5gcwLSuLTyri2lz1GSMDu2vXvsfmySpk5XH65e7H3tYeGsnudItBCmW
rIGpnfNxok6eSFNvCxOgUr3WpKZ0uzufguC3MQLnoOO7e9oLRuSg1nz/fieqeZwWksMZAC8admL+
giVZwAPFuR9zYv4nAFR03G3SWfpHaTu1e7Ssoid0aN0UuSyNOBN8CIDDq+MXS6atKk6JVx+/rL3l
TBEph+bbdllSZLbH4KzTJOEfHq2ANQOr6qKnYU1hamHOyiSGKk5XY6j4oCBW7qJRz/M+kputkDV9
L/oXV/Tg1UAtIl0eTX7wKPgEJbsZ1/7ZGFQp+nrbBmfsj4Re5kudMNHex3pevuscxxj3g+0lsOnG
MRCVu4fiXt7bKT6YOdYmTn8IGGoXunIotvGumMVoNut/9Ld7XUKPdtFElAt295c6y1YxYPCAi5T+
ChCkpA4wY9MFD6o/8P3Xw2uLnQkhNkpUDg9h/2FGjju7FSpfFyL7bMhOl/TJkZzuzobsy6LgiUXI
G/CT7EWewqr9YsTuOuIqeUWD5ZDMUjv6v0J3FYyry0WTvgS6rJzqdrzSDXy9uAuJkR8ljSfYRK+n
UMga/r1bG6Ey/olliysM2BydkY5AZkxAUu8AGDbM3l3OiFDtH43fnka6DcM1GjdpdXx2rfnaXNs/
pYfpxVc4k/eZ8IRRQG8FnkIU3Hqiy6NS/l/Y1hR3W9HINbvJq9bnZHh+VqaY6KhBZSq1XM+Dgwyo
2XR7KaL+5ox/H8YnuPHP+xai30Cze7XJTS6U+hdSRcdSu2pTQlmGn5XxIMmpmL80bYcdnbf1YbT8
zBa1/1sFGI4C7iRAUQM/Pq/aegUaDrxINU/xiG3rmz8wYIVSrmAFarAXXSjcX/zikTG5++RN6xlX
09qiEj1SjaChcfrjibnMbjFt5ONJR6jDMwWayk5uKZyysD2Kpj7iXv33Pww2QF7sW1lV/5/uL/kH
6LEn/Wvk4dB1xs8E6eAC5jHAv0ICnqjDoXNmxcxImiRXY0fHyGgWT2+8iMXj8yq4oJHijd4/Xxi8
8+dtK70fbAnuncaPK5QJevYuf6uRrmWUEGuo3ev1mFMj2Rufnsq7u3OglLRpYpUfuR+Vuvz+D48z
VXIm3TUwR0yaIgHiPa8jekYqryFp8H+3j2ZtmGdBwgN4r/0bvtOpqJgHJCgm25fwJKCybnCVPozi
ZODng6b4nNIrvnDlDvMU5T7Que/HQ7krR6IrVN5EBCt9gbAAkllmb8ikDq1epTzm9oBWJJe40hGI
jmcDhp92+jmDRM8R6H14Wo+Wa4JYUO8eevfBdhz5SK92CpI8kGgFk2i0eU5h9Aa2Va9pzblGHJ7x
fWeVU+mG1WHu/hYuND3ecC4PPOjnNbFFz+vxl2r8u8AMpheK1XaxDnI+k6Pkn3uML3B2gsy4Mjpd
E0zrGUEf8ExB/HuL8HfXV9vAdrTM3+tBIPOq9iyOO7efgZwAnyTaQLkaPop/Y8zWo1N1vapH5o5r
DK+uDNvsrm4VkFh8PWJmrfrJPYM6AWunoxsgvbxIB3d+IWDjPBDkCULVctoXZR1nPuoUARE2WKu3
K/XN0HVQkz+ZvWiiEMHkmMO2A+ROUomc4v1hZ5/rx675JeGlgTCNe2NWY6oOkxOHq/Meo7RL1aYK
+p6sJ/7JJJt8ACELYJ1MEtcLbUuo5acy0i4fBBQJ+n8CDXqssZOwGpv7rR+0hrfx86wIdF8hUxwq
9ZyIlLQdfQPmiWxGwD4F+GWnCdB9Sfmw9zL1RJXC957kit+Br2VJx4vG7qEj+zdPXyM9XPyhMus/
bIZHiYDzjOgIFiobGw3Nyw1xgk/1TXgtAo7gY6KdHsPpGC8p2/mO7ZVZRD8MJIUut/p6MyEfWXUY
qads4zstdcE+FkAtYmAUGyja56xdv08jG/vAFasgm9sNUnWaJr8iEJQTGZrydNn+DUxrahX0br++
XM4WGxfzVOaXny2yIZ6xmowz+eXWI7Cy1E8teb3E6HnV80XJIWsiUAPmLl8oK9UmMVRFEacgVqox
4ZVB+bm+4wkxGpIxbL+tktsBwp/sCP8yrTIia6SgVmiu6rio7rEQMNdMqoRly09eWnF4VOq0+tat
v1xxVjeEnA0x43+2CYpQcjpVazqzdWgDV0eAJbWOv7aZ/G1YuW5rx7W4B/Ic1AASTpdmgq9rQZbM
uuPUZVpPNAiM53yvM3i16sOHoqHuYGbzRRJDhTPKVfMq6P2fm6fATH+AN8+YqjyRXPrU7iG3cMLd
AN4ht19N2fT/MrU0eJUXXo261qEwaeJyYebvOk1NsKgFlAozUtlgXBqNzECAgrimINWnQDFhLUrR
eJLRau3SHUk9Sb2HmcF4vqGI6Cs5GmfZXIZSDpuZ9QG5Ss0lI5uLjVBw2euhfObJYSTAOM3URgFT
kIiFBanJTdR1MKQ8WaJV0DwkbNRzHeFdY73rw+Cv0h+8T7Sl6ZN6JgXz7jyvwdYrkHrYMOTdoLD+
2PmmFHQWDoKI2GpLnAFJLu7JtudAzzd7zWMCuNrHiym4JfwxkpgHdN7r35ixYFa94W+pJtXpagAe
JFGP6WNwz/GgvnMagDJoSWY1RnY7lkXefZE1tFCfQruBzYKou3iZFBH5be8VLScJOuL6dVJhUJMQ
HlyOeWu93IJVxR89ly0fhBxDnHMYe0yPZl5iHph80jqw8AOOBbDqS6g0ECRoVy/CE3Rt0uqlC42t
tSmO1v/OLNTTay3AEVFhA4btVnplR+obvL5HwVsYRrcH8n+uDIufyKezVfb3LimhKOFMlkKBvNmw
vb1eESu0Ge/KLWd/s3cm+DHgJYwr+JGdIjL/QOJOTRcvFGla3W0xQOvV6iLXg+DCPh6fy+Vn7CAa
1GRi6n2JZ8w2ITulUXe197FvcIbYvEaZg0KgqlwLCurRUlQZUk0+qxTmYRYP7LzRYR71nJd+Ut2t
JBI2i5PlQdm15p6FFYDToi4pSAHsvKjNP4vtgQBDgGs9uo+2KTA1YDqYpUaj3gO5uNs4Om5O/ht3
DLZvTNYDlZA1Thet3ihdVsOCdPemtKi+Oz9LO55CajAgVHm681cWTL7gHSUVR0CoqX8M1npDCCen
0raYQVg49LhpBVA/mgMToSYDXOOWIK8EmNNmuQoVXBdiBSldUo2X/OEg6YoUVVejaq8Z0zf2+Efd
ub68gl355nYYMWohHsDp2umOwNN9b7Wnxb1uNP4IdpNmJbqXupN4JRh7ku21OGIesnKNU7URqeAq
GrTPRm8o2GMVdGJcfdwoeDZyr4kXCoJSQBOWyWZfNmVdoHrgNG4+KHooFmcXim8FzCf8TZNscG32
Vx5tn8q+lBOVgDAtp5hFHZwZ7ThHL3vkfJvaeGRepfwqDEWx/bgd9Sq1Vejl7isluzSwv/pdRbXq
CQiCwiWKaWQjjcoIANif7Wf/UQyHI2nIrnsrXZahF51Dj1mGK/0Ma8fh2PfM6RAoHKb+zENKSbg5
/yVb0o7A5MDLkXgMfISl3PLyaRNeDDrIACVNbSX+hqgwyuecjjPUMdFywCp7RooYIzTsvUxTeRER
tM4myoYPGy4MPRpLEzaqWF42D9DvcWL9g2s1nOH5EcA+KOJgxB4rntugrmf4R6ubpLpiwybKdXGK
UoavUVQP7XRNQ0ci0siPMuuUmcQHv0C+8G1y96jgLzz7AqsPnGpJtdst2GyiHvB1tF3H0+vi29y7
kpuugsgF7sYT2AHGytAar0NnhP7ywMZiih17Fje8RzdEZVojQ2IiiHWA/oHtj12iH4svrYd1r6LG
1NmcNIDVKXTu9PDO+xh13ORvkhMAFh2fWwcquy3dBI4bns59mpSJQdce9p0dxIJLhPB45Lh80K67
E6yKlPhnJCRU/Uw8Ejyak1f7CVVh4wd9CLLGyAvXq31iFqUXYa7UQJTbQtGNYkv+85SsoL4KfkcI
07d2cdqEZPW+6a/PafUjqqhX+CbyvaHYOwE4srhZXBFvwmOaiXEDHO1Pn3+1txVYROAUGpD4JXo2
3E2dOyvFp8bRCMCsdzYlVmBgbuO03Wme7D3lDrMnp2yKzI49hSqnzypBKju+Yan6q0s2nWfgwzs1
SUFyXt3r/+4AADdCW8gzCXKwQ1C0Xs6D0CiiLXmFSdZ79Ktxu3e0qpAOj0qADz/HSvaZTc8n62vk
/l3pW6KcKK5qb483MyahuA8dcZ99vO6zW8zm8yRq8the4hMMFXUj33uedF3wIV+GAXqB7nf137RF
/jtDtlWYr17EQaJVp0GpjWMXaHIni1FoK2GVpK+T7ZELEA9eMrT/iN348RNby5aS6rhGvLLdtmCB
ggsFq5dBsK/LsqCLOuI/+YWs+l6v2U+MGLH+iDGVt6iCkH1MqdlOMaWMGCHMWIZmz1mE/UYGiXBw
LHzwgEIRga0qLQZ8/pCx0Pr+A6R089bCeO79H/5orMtDf/hWLj5VrOKj1GVvUvGykCDQ/lv+2i2A
ykRSK3Y12h7gfFij0zI0Jhfj211FLktLpZvsrSRLuMTvc4hyVLdN+frxq4/biXE+K/cOyQ8p9Jqj
U1D4Fm4JozFRfgQRN6feAnr+ZpHQ7PvP+jHW0CjAMzfDcxeUZ9P0I6r+nPiYJ0wXDqrAMcaWRlpE
c3M3Nym9fll+nydRDPa6VbdjJzTj9s6J2XcrdkPxztgko51nPzvZm3mtM0bdqaUsREIIrhwqxwGT
o6WbGNPRnosI1pkxCpjiCKYVtd9/vHhNHD9+t56IPmH1fKuiQtYenJS33X5UhbWXVlrJKsKP63hT
Mh07T4WqNOzodGF35BmUv/6B9TwsCfmOz+nzWnlbrlPypc1yopussTQxU4ydJCLfoTFLqQSkLG5l
1WetT9nJwQ4OwPBymUYQJ/k7uK40Deliv8398RpHRjbBXmgwSY2Vj8lgSE97WfnmdilaK3Q3SGsB
AvajR27r9vIS0zDxWRDc1A+kurJHMKR+eJWtv9GsSEPhJ1lkOi07yKfFNxf5orlhlar537JtOjyY
A6XLhHDe/TwTXQmQA7v2IQVBYOa29bjdOrsktOSG7NjrhLbFcleBd1VjPIQqztYr2ivx5uj/9tu2
+N0LXt5DDqyruU46cCo3c2eigHUZh9F5Z11KVUTCCwoAtKlacvPCO0p3dt5hSOtRDfv5pXlqErmR
MrgNWHrTsy/hVpkSxFdCuQTdU0wm9QL7RfWxuHsUMcX7w4zOgtbNEqei/hKb6WDc5g1GkBrYkIxu
o5nhod2wWT/6sznwJB0uHdnsRByoN+1cKvAMErssnlMRHDTgvZerhFOnlfKltgCR+q2vQhLMCQhr
oAGyrV6B4UPnoEyc00V7Mpi3zuY1k9pZyWQy/fkogBzHvihc4fQepVnwDlS0ujHpDfvDBqqN78s5
mmQEMx3we5dH3DW9X6n1Z/evu7pna1/pkfv42yFRwIJJYPdofU2DtEvHbhT5NTHrw7HNmmFjMixq
IG/eY62ayC1T0kd6EvSHdBPSwHSHB5yPVGIoG2dwal1XbaUHTzNeSCuwyH+79l6zdJUGjmx1kvJI
KOdUY7YtcD/ZkKvFvD3iM2uwVWiFNbWvJWZGV1+fUWzkAb28jNJ0yfxvYbziqb8Sjd+F/puOh0QA
eFxm4Cp5HKpjfVV2WwNzPG9Ef3vg7XdYZHrjGR3prc1PJoamPFId9gAD4w77+on3P6U04FHyXvKY
eCCQR0HjPq483hdKhJxB1lSaRDQeN0nTFQ2Qz34G5BMhQwNfCdPWGWyvSvQSrssfsw/JspXRwLZO
MW3+twe7Hyr3FY13NLKSIu1hVvbAmnRUHLBzCRGiY8KUBWtOUDIuPvN8x4+ufiagX1vcNtpQd3QF
Nij3wGJbRk8dxfqmk2j56F3nat1/x+iGtAHUITEkyafv69HGJMhj+x5PsibtS/PDM7PbUFwSwA1a
yVuedFzQWuqs6kYCtpIwN9p/pMByE2In3CQHwTKuxG5CUzNDXBqW7gmWgkzT8aO8v0C5KgtSwVvI
pqOZDgjyF+WZGR/slLSPRtyzvNXNKXO8t0lw/YjKP8jkX8ld6ndZSfIarlf1A+6dnPuCa5tIAAOV
7Z08CYqP9JHP1zZTCA1J38Mz5uL9IMK9xnRkJjBtaZei02ciQZfaw9IXqDJ7MMVOHfY5wUt20u1/
R2KRTqiLna1gW5kSTG1GPYqsVtDdm92B/+u0IppUFM/eI+BFpMotKlPxJhWNVUwwk8sjaMgE/llX
10EV9myCmoca+4zhkXktnQvCaBFNqDYplzGBOxaqZuEp41st0Ls8hDZrDvJqgqTqy+AEwpHsoOpR
3+HPPoQychXS8ZjQDV5j1/cS8nKm9CFC+V4EeNoqKv/0LbN1CiRTTy0UqyoVmztdaibN5+t4tuJX
aEq3AcinFGwbd5Qx45DgwdFAj0WN8CBFDGEqmPERIlPRkfyWLlOrDUsX4L6YnP77fY5H3c3Hrj5C
0H6Xvrg0yTAc59RzDunD2TZ6ceBHAsX5jtIamowHHzFr8PQqopvdYmnBMsHK+mvkSc8wsP9X97L9
J8/IiObqypFsOlVCzBkpHhKH4/2bMtG5CBW353ICjN7LrMsDobKkYmpumGg7fVP60/drm4bX9rhs
IjQdwSpaldtg7EHrkVveR+kXUr7T27709XdhLPVgWwGwVmp8Q3IzW3ErIFDgBHdz0thoDu9dVOao
2heLKzW509aMjnAg4oHwWhhRapS7ROMiDLgDEwmOeptzu4IUoFrzOrRNBbs9j+JAODYD1JZ9e469
EakM2W1zXqBbtZFi9NDrt7cz+m+4iVpy8adkjaAVi8ZNCbIImQJ96fLEz0MzJFb+1fyQGM4rlZbO
mrIdxm6jqST4Ef8yBolcuzOEUNpfiUU+zAtG1iIytWWByWLBkqrDVN3OL0NBYsyCUI88bHzXkOhc
SxVMp4Di+TIU2dfjPGbOYJUWWrfEMIkWJ/zDY3zwYMxOW0FKVdACntGAg1AMoPCwVNjgIzZCndLt
rDytAkdWT3UIFxVQCCy3yoUZRxd80y7r9SVhEhovunDXjzDtzAZklciX5HyHBVtOeaMsE0rHbwz8
VIBbmDVDclKZQC5jRgIOg60Mq7xCtMAja/GVJ1lJ+mSd3HVVpCZzaXvwPv+iLmBmj4+1A17qqocH
/f+8m7SOgT3mCUHNMN0arLl0b/WFKJeN7vfN2lH6kU108jJ826LxEqqkLZ2ZTarurl0OonXNV3wL
aV2nLDwK1+TvOK+eBuLpu/wISQsOdRpo1+zZ0HmcTUT3XFIpDooBiO98mwt6tozjHfqWPCma3AI7
Z1QlYsZTvhBkh353Ab5zvhFW5DZ4ygobzaAFOuefxytFfbGbZOBGNrgpNS2O4qvBDFAYdLTKaBzM
RzrJKRqw+YByADOhJrOsXH0rq6iOTxlknHFizZcl6vdnioQnUDRs5M7Xujqi3I82SVYRaVySHoD2
v4plLDQx8UpdACInJMnIhOD828O2DGRNX55hE1sG6szEirLKRlERuOoZyrFun7ruZuasCpzx+Ndc
+qaVff2QNCuo3lxrLMPDLfn/ZwzCCdEl9sImyzDTV96oG1bftIrtPTixk/D5F547UkAvohEA9N0I
PXo+b4JjUjbCWGg1VPUcFOOWOFxxaFOO0lpmLvl4HpdrtGGetZFfs9qeg3l/ESIpjUfikPExxbtG
bQlGdJq2/kEwIQL7LNVmIcLVDcQ47zPM5XyOEdivHmYSRctM5fASlJ01u2Dj0bV2bPh6Y3SOisWa
4ZLSe3nLL//j+Hcn1HDQjvlCFj2GkDGTBMNcypbVGBcUMs4fR7os6S2Y2FB0NqGdwYwUeaWaj9ct
hGsXSix+jJuUMT5jKAJtuS3Xz3Bi94my/B7zpLTkkJ41GX6siLcw0u1W2MDuszw1jKXswwh6R4Fb
/m4yW/55+4t7FM7Ae3EAeHe8inVi+0dngZUjRFpRCyqxX2fbdKK5SfDqcXqhbclXUpVzaRJWbNIA
awfx6MXTSOy9EnICi5DKJytjRC4/PzSHLfPjGtQBTH2/cc7LANLFi74+vUFp9Xqc5CR9mi3kFcCO
9Z4TMwfqaJpoArkgMwjLORiCmCQP1g7NNicJ50Rzah/r/fHVjvC225IrQe4X25IyFIDebHVP0N22
wANY34Inp39NirIhVqUU1SxExGmadsMNhzC3sAiP8IfhqeuBR/e9Qw9qK9RGsF122WcO9isEq7Zi
w8kn29SA6ImneRclnf7xtZ3l3+t9JXxgwYe1SJsW+vwF9izIjWvBHI/IaSwmnRbPj9O1e9aEBVdS
uRlLMHocKpGCWs+l1xNN6ei3ETnA+QqERmtu50qeRKwH8BnTV4P+fAaXTmf0Br/LNw4bxEGf+dw2
EqHuNXmChkM5zX97tWfiMpEmRVJkrgAWZzxIsgfyRiawYpy3r+VSOoJ5tY/DPC/aRAF+QzYveExh
6o8mvX33J3ACVtl8ohxlm5XOzgKVGWJHkj5A2cbtNtXyJPO0YsGOlFt6Tkb9c4Adl0HcSZeDOj8r
u9RmEqqCjieBQT+bTjOyEypD3AmkFXDuTgXek2+4u7t6wEGSzbR57g412+rJZHuANOpJBa/xI3Wx
MAYGZWG/5E+hfKnjsSRZmtTagV7RnozCt3ASeOVFrLhRWb7OIDC8Iiq+vxCC4iAY9UOG01KgleX7
vUZogmy5sL89HM5vtA4DtaxYICTOJo/OYWEHhpgHLY00cHFGXHJwwdiqiE6oiezbJtPe0ReK9Ltb
w8SLQOV+f6RqW9CFtitmbIi7wwxL3cxc0xEpDQEW5oQB8uNA0eCGopbZCOL09usHlztp23JQ1yX+
sySmGrzTeC8VbfJZsu/i14VqWsf0rg6lfDxw3G7SyTEo/gWUbmkcThjoDoCx44JuReZzFFRJQdl6
xbLRXHeeeE4mjjtsD/z9HoA//KjB8ejBDY8/MwoBXMG/9hg7mNq2l3wakpziQIBCy1YF8cgHMUGE
S4j6LAOr2d0fdffep+xp7li07KU+EDrQtPcIn7Gp1E+Kn732CeuV5NLG5iRquQwrZIIzd/hoXYkZ
kRFlZKki02tDYq+y3Tlw3HHhe/7xXom/jACo5nfJSMoyx6PU+TMqNigB7HJ3xhjMKJGd+5jmMT/s
99eao5fqCoBRzcs2ORU2ECdfyTI/s8a5W/9FiY/BHSCDZPk2lHshnITX2Ci6E1QrNDPtzI1dUBy7
pT/TD8a1P4Su0qhl/E7t5CnE1SomwV1yqlh2lBOvzVyj9wfj92th7c3qb5xDBJSXSciaPWErnfQz
xjhEBhShcn9k6v6sBgLaPr9J8yJWD0WQ2tsynpGerNw34pP7TMXIIaMBbwziI8z8mUFdVcoL/y1G
gkEYwN30MHx9SRVZnNIPKMa8Tev7P2UE/aq7nTSlLSVRohbbr2MwoQYj8rBGTOBXRxc+/ue3i6ar
QF/7ngscUC7LqHwbXVTN7KRFa54ICgZajleRfEt4xACLokXQb0Vy1IxqAnGOqMzZBfk3Dx5HTPw3
a8/8h2E+mfXMLdrdUO5ByK9K9eB3LtNo1Rva6UlPjyJ8hhUOy0+2di0sCARtJ9UGtRzDfBYIMSE9
J2R6sSaniIQRQqsfzZ1E57eh2nCOMQy6ukXUCXab/ct4NdRW5tBTX8orBAxeHWv3ePe6Rth2vma5
PuxfKdsK33vqBKPD5JnazGIqUyTT9KmdvtVYj2jwtwUAhwmB2hNGfa1MSLPFrs/WEeF83eku/LgY
Nr+aMi1wY3qykybY+yBvQGclmxoUS2uAWowBny8OTGAHshoxnN9u6B/3BBvCxsVSP3Qk1z1Oze66
vFKPHz+vdpPETivxBNdpjQS17lzWOm0bIaGqCyK/ACueNBS+41lTZtibHFtvMTDUJitRbNT6y/jE
kJ43/sUvc7hY9ab3BS+Jitg82Iqp2cBIPXDp+xAi/6+C3LBeb1EplGFVeW5naqRCpU3uxSf6oNKv
Mds23TcEm402AkJ9F7phS/vYiF59Tp64Ghy5LSStD0dnQij+214RHMedveydf//Hm63/FYMpu4N5
EQ4KhARts+SZXXKGOED3X79nsX+M2IM/KuYhblp+43Xoti4fOsoxUjOqjFERsNfDdFLO0mXbE9e2
pmWSd4iHowpjpJteWFbRu1TlppoiNGDCGFdKxDxyZMjcnxUyyn0G+SNhYLfcH3NFPHFL3lWbOFEH
hoe97DRAyEuypJtj7TWYnSWdlNEq9yCWDxihsYhqwTjY8rZ2Tj8MHn4b2eeYIBWfsM9tLLNay3yI
cuJzxKLO9hzqHxvfod5oZrSTF2SMXh8V/wnr6o2PRtzdob0nrGHxj+50kAd/cn2l93lsSJ1QSypR
Km1zcFosMSEw7TxnE00FnOVcLiKz8nch3Ecor8Mecb6x5N0gPaydMboV5X7+S8uSWh+p7dh5Etxo
lGGVUrmIkmT1xkKd5HJjd/Hh56V1pzsqhDsdcYTxOJ8SMztVW4m7yTEN738P7eFO+JljwsPLRxoK
5F5AMP52rgnQlr5BHOTeSIihANbSgi15r+tbDL2wkqvyJwpTa0FCVZLJqVz3OFWeVAYY26gw+3OA
FEVA+3KyAfjoY/H0fuqDYLQ+bvnzsF8B34u/E7QBANFteGy7iv8gzL2Aqwx5L5Tg5N9yp+HaZyvw
2ODi5JfPekmGBN11f5CxTyhtWQ3J5CiV8hPTGuSztPbSOmmpZS/Uj5fhq+wmUnsXia+iPKvihvtK
WSP99RGRzjPXZCNUr5jBVylImIP0BgLZ5BDOxxHM+rEy2Sm5oBZo6sCWCZNMG8Q0vVdpgLOPt1RF
kr/Wi6RsiwGKEuRNCVG/ON2wCWKrS7x0Hlqqn4Kh4Qk0G9oQE418XKtPuB0ddjxP4+kpTZQo+Sxn
0yptDJOF+Y/IxLjzsC26pilNqS+SeE8FImfchO2cve/S82Q7w/BcnvScgpB/jJc9zE3t29js8gUy
hb+rN8X5rSb/4MEMnAoVmXh8Kwwtzpkd2Z4ZaewI3wX5RnYYFCzg7zzKHpS5DNjLm+LEmK1CCjQ2
RB4YOtlgngr+6N38iPK/2jbbC/2C6Cti5eMnG3E1BjalXASD//FteCs8Xf8o2mTabSz8Hw4OqTQN
BRG/R0r/74vMAVXS5BelYL8B9IcwXtmGzFzdjuvr5U49U/wsDVhTjw/C6YCsRm6+xmhEdbvRpLzT
TFmC6TRYC7HWtdORI4DLQthLAOdTga2s+uk7I7/yEjRQVDUAohrJlAXr20c8bx2wV3qrdt0hyeW5
VsaSnun3R/d+qwjjLs5TIRsbSPu1CSeH3YVAWwfee6Bh0oi1lNE4bsdPyCxIM9ceMwKa5NQ9UzM7
smNnwQ/znApJC0rNHKPGfQSz2dHp4md9BJwQCCVWAeyrvHd12vzixlNsOlgzrd9Dvtr/YfedA755
w6mQEaXlWmO4Mu89cwudX5d5hn0Po66yWRfPAXJCIhJV6VWiYpE1a4ESE92L2j3y8vLpRuE3qAi1
MASPVqNHAor+LD5vmthXVwtsBfNklmUXn2af3D4EsYFHzqDG2aJeyAW12GbxDKtQfqqnDftqkN+H
ltvv7jPgu2zr4VVy5hmI0ceURdovePlmCDZI8dq4wgytTIp9iKpZ1VSEPqOkdb2TXyMpe0voazCg
HqWAsHSw8syPCPVXwFnCM2qU9VQloRkwH4xu6o9ZxYNvcJI8i5bmBT0GK4oVhRPuCrikjEBc/PzX
Me39qAr4vCaiydB+z6AITFzc8Y1X94WIplhzPLn75BI5szLEm41owz64x6ZQJPPf6FcA82+twuuq
XVDmvi1eFbKCwVsGYSZESnPBnLQOgtUEylXlWQfSt1D15RXNo+3iECHVUpKDBg6dMcz6dNNBeSYT
bp7GdkclzBUt9p5dQk6aztZG0MGuGMJR8YGK9pwkc6dZpMk6lYvB/80W63qfYqu3iisQY5hM/OGq
Y6NGtFEaceFgueJOKVduAVhc7H9Ejq5Fdg1EHyUvMPk0vz3NsFmnzxecEvYttaidFYXigrQg+RiD
ieqKwfz2+JLVFaT1DzbDJzlcLsAxqv1bfXRH8cCtkTEDcdPGs+83/iRZ4/Sd36iS7j3x19yiFf9n
hg4xun5JpdVdmg1qDjmarjpLrZ2DZ+5Vb/PD5WsJ9Z0rm8aF0WR+39yGLroI6IAMvmbW8CAwjJfw
BCRFK51b0LCiwnPrUuzsCNArvbrccf2zdYK2vf1XUWhPOcz6axgj8rm4HtStXnYq8UvP8okrWs0s
IsQPA+DPCBSq2YMBBqjhxE8C8vwughd3A2WMuxido71et8ATqn0gBik7VNZdSKQracy2fXV7yy7g
TtT0PKKRBVuV4U3IPwYQbIAr8p2znZH2PFUegUdyL4PfE6O3UbgflGN+X7VfcRrhxeR4IZx+Ij2z
sSdXaxoQ1kSF+0dHOU4WyhInWLZ9h9sTay1bGGYNZpQ4JmCoE1WOf4SE+LxkWRwXZNfkqXJq4hVq
CxzgnrhrDBCVzdPDX+SyQZ8csOKMvfaItJ9vVfADxrLA/7yfXEsT0ji/kUPeaXG88nlTvuk9MsmW
sbE7iv0WDLH/NjtpcUTzaM/OPZVTfohikpsKoZaUHXTTBrKYj9n8hcOkJ8RqVI9wOvLBRw6ihZ2Q
P114iwmvMizFfD/a20viWwp6czbTQ0iWdbEeK4Acvt1AK7jIN64H9ElvlgwQujBRdmas/4ogW+8g
V0Qx17mm0494BzZXKN49HVybUa+IddLHbTfOuLVtzphG6fmODvYVRee71WrKf5ocTd5B2O9LFUSl
hZce4osrMJ76OE5qLxxLKS3UPJ1jwVPt7bi3x0fgDt2h2yG8qwXa1gO/1be6wnQ5V1oyHfoDFhO/
UBQVCQ+ya7/ZlKtp9cCoY1Py8y8ibC53+bYoMnwWw+eXTlXVvwlnrwgWAnTZe9sCUopOu6s11Rvy
TpwWbs5hy3jFG/6r2ThDtck3nIXsrAALs6G16A2rWLYw+Pk7vE7RyNoKyBOIpkWMXdv4+jsIZvAb
9s1FcH5d5xK+0moj8lMBM3lLJx6Kdlje/Hem41qdjvxJ7NaONncDohBNT8Yqqvsb4inmd42sn4ar
TBDRtqneTkQ0HLBm77oWzD41FUWb+1TwoYrqwo2gTwB6BYNHQpq1rM5HFH1rPd4BUrtm9D+MkMZH
N503vLaWJmWf6DHCVRs7WxXKLDOD34lrQ7zxYHH4hjbHwZdCs8nGxvtv6WUe9FhA8Lx37jZL5e5E
RSxVirUA6hq9ceibiRaknHK/FaGs8IhH6RitLuls3ectMf8/M6TrI1KwUB8MDImOIFRx6j5RDkAT
XHkyTxE/jzeBLvDyqHujZPs8RdZvriQ/ONV23vLzC96koUCBAAy3HLcF2NmHkWkDeJik9LXix2cY
np1n+2BxyTFUsamoF6dNd8amePHad9Q8g4sxoldNhMOWyySSU5Z9NWbVNJLj/uB51qAIB7e7UHKG
nChFLXuDf5lRn9ahB/p8orHipjlvBVVe3MGNaR4GNQ3bgPy/5LYuxMQH+yHWc0d8ehSdh+E/tFmx
oq6MA0SyvGQSm1ZDgwvVYjwbyZ5RfIjGML5Wdi8lEDpxRP+Kjc2dGeNZUNX3uc4O3WltSbtKeXtD
dkoJUWgF2cs0R/hj6ckxlxiqHmQR6AzbUx643rnIdBNFfTrZ9bT8HFknI5E1vLnlbs85oPKSLC3S
tMwUTAVlwYD0HiXF02jzlDrgGDr69BvytyGyCgL/kgt0AnPkIAuulxFRWlpnJleBQIIRsEhVZMd2
ZRA1n7WdTTrzK9DVr47jKmH2DCd4LXGYW8yTGLd9tNdUpjCSuMDgJ1muxJnw9ZyeyN2L6SQ06c+U
AlIC894rVNHpgk+dlcUHYL2PtQvYzWbTVG2BV2Kw3cENgCk1fkNcy7IlqsZ7ktTsZ7c2IvGNfvBX
kyNqfDQAFYW3ZlpgPLAUD4nQi3ovKBdSJNGRl2EWGKpRpoAJRZV7oFUF0l/8c870oKgOPHaelwOy
xS9OuVoo9FJ56pFE/yCRdCT+6qGwTIOQLZGmLGfcaZEi9luxEsuGKrha2wzHjGe1fK1OLx6mq0wS
QjNdd7izMMeAZtKnhItCze4XAf9axvklDORxtYneEgXXw6cleK/Wfq+epM/ELMdN0/VVRiZ7GXul
y0lRwi66Z+ZMPezaTS9/KYJTdOL7ODtaaijUsIYq7P0PdH6KVWIaq3iDZxW0jGTS7NAbp2NHnQ5o
g4sH15k684Qj3x1pFi0KBVyXRfdCRSaKvhfuNN3DvhiBNAzu+k0cnlxBBmeKgtcpPXJDyv5hhBY+
ogRHsLQPexC+7bvDUCpc8LtbUUZ7TMfMMcjfBzs1KQwkVwvxAQWgVd0OlIMPsNciSYduMHQR52MV
yPYc7Oob011WjBDv3ad/F9oVz/4vJEEVirPs5eNOZllCDVcrOeHUtfhH/b/56kJD3FO15es2aKPf
gxaSUe35JuG4C+0WdUdqVqLNMSermBWSxszIkvGo6LvfoB3U5sDe3wTSpN9QHv16f/n3n5irrRx8
5j561cqCTcWbS0DhH8cRtaZVyUq4TNe4A6PiVm2URDzz+FpeZTi20FZVcqN2dGKF63axV5zhMg3w
U3o/xUtFBqT2yICE0Y+/B4QCxtzxYrNYcG0D14b4jtAMvzmN4e19c4lCn76LJb9gFFTyw3qTvV3e
KShGAKmGaTbe1MJfqZu0iEpL2s7/fB5bsb6dFiK9eafl5HoZLFiHmgxNY7XM4zYUxOPkYvD2AsMU
26FqCjQG6VWl25O6/4HeNZ+CG8sGxIz8DnKF58DrN2Y9QMetH/7dDLzV2u5sbSt0vEfPYf7TRO59
mzofgQXoNQvTmiqt4gqJDZgb26YmUosW6PzKFghpmGwb5omZiEQM7gDpRAhYy3XeSRPKJHzA4PLl
yGC0kecX9ZjWK0dqTQsavx5CppKBKqCtlV+EE787+SXsMCe1iX9uvXrWWlRpXMp4Bmvk843ANXNd
gTptLmqIi43yt3YXontuo+r6JJ2e6rnfA9/kVb5bmDz4KaZoN1TsuKtzMxpj49RvJTjyeZmB5D+V
AMzDALqPaowanXmN11KxLXBtn/onxti/mZZ/rkFNnKUckViZEun7+Tl3JfHZCsHvXeau54qVvhnq
DkvokRkuVO5aP3SmPlNvhJ9310trNzGvs1CXic0i3ja3xsJzy5SKtz9TdVypefE3PSNYlkTVehp7
1QH2/Jb2p6ziXqGgxF2SBFK/1A4sdpfyr0syeX6lB8hO3PFkOQTl17+dIjSzTIHbZzbIU//UuQkt
XxWusEz3RTed3C17lgGC0SXLvfXlZpnIJ/dtGKjzxS9Cz/qT+6RXiwe7IpEgsfLxcZCnQwm8Vmoi
y4+/Dx9aKBbpZZHJCrfwGmYRC+aiuUjUa2OqAmB4zVtOONHNxIkhoC5g0LPl2SB3synLyh5U5Wmk
eOZwGUteeaSIl3I1LscpEP+oQBwCxd/FdVAqGnjMnwzUuvdA23CJJ12HraHm9jaJ0TSwrrpdLEBc
PvthW70CBsZURFhNgry2oqf7oun09CmpAY9ws+UlprEj2A/uYXLb/qOQyVPtiGq0q8NCDe7bzULm
JjeRmezvOAL9dNCeFIEEY2bv0ZcnoxfRy4236taYcADh2id8KiOsXxcSZeOO6wHWyTXn7SRUk6Cj
+p8Sc5mjsmE+GEzJPGQov+/NXXsFTmLX6bLG1M3VXPlqFKOz8gRrFFojtR7uc9Lu71NEUvdFZ/nz
hi4hiFA2dnUrvZxyRQy3k18fJGMnLb1v0rq3SVBb5edNy26EucvOAnO0bkgH76Yjur3hKllEQm7M
i6h6b+vfhfbjUO8vE5PSb28HSWpPt5RcD93wdqJk2IlpgCMh14gML1ZISDUvsPbwyZufTNBZ8lBk
0lpLxKGWn9C36nQGcjFEAvTVRStE1S0+KymoJjswYcvZx25Yasc1tEn7VJjOoQvF11MGJ85Nr9xa
xnXCRvKChmvovk8E0mL3KoBLa1rHIX1dLoYaMkXMvULsZUoQ1ue9vDQaC46M0znUujBZrcskL4bH
NvoWOOx7YF6TL3bwiSEs5oBxelzrpicPUGsDc0GpgmeqQ4m9pJ3aw7psqbtMLo36QLwbvOXwp01/
tL4yqlISMkB1+cIaOABhn9Gtu3jebbn+4EcpHYPwcrtAHOwO/6fcwRM45AgPRdhtvANu8jf5iP0Z
0bUP/o8okoZu59C/16NZYXjPZ4DbilRWps8gLc/GubeHkavsVGjtiE/kfzQeEgCRwB9LDD8Io+8H
adGGZcCsQz1tqi1vtJKXuq7oz/0bj7X5hQF58Zt4l0NFqRhCG2WhNjn3l8mM6U5PdP1+G3XNG7S7
qYA8kmbvGMwUuTsQpQICKqszWDERSQGwN6Mv4eFKk4rISBpuxJjS2VVr9kjup5SsEjblpGGvB5z6
l81Q42Eh2Efp0gXq95mrZuWbl1eR9E+GecV3wy1mRbXaAd1Ti9iVeVnt93mA8xWnOJ40xE4oLzFq
Gcor8ZOdVJk9aYNhz73fAqir03ioNkcW+RhTApNgi7nk847wd9OpWrpc9+un2Yh1e0kXwhyO12cA
v8grZwpZWbrfXT3iF40aJtRGeq/bDcXWdReM1uYmiq8tP9OaIj/P7OahDxMwcI4HpnCPXo9ExIOO
b760bEDNiRZMhigRcpKJfVeyeY52JotrZbn5vRZ5PmjDiZ10pMu16p4Mh3oH19DPwRKG/B9mjvJo
xfNqBYpLZySgG9Bi0jgzBpmZkWh0iDjS/XFEiFzDMGpiwEuXaM/ZH66rgPicEW43KDj85exB35DP
IbdUQ+Bq4f55XiZQ9oamH1jQWc11IlUXATrZbltiTF08YQdqSeZan/CdmqS7m4PIfPbBHIMXWdoX
1BILbV0+pWkhDszNOL09Z5zwgdyVSIxWTj+9I9vGuQqWmTy6xr2fUFEHSNqA4Q7gPwTY6FFZ6ZXx
SfcDXqCrI0zDc4xxZ5/mf+Zk8tPQz27jusHMWq9rxbBPqoPKjDzCUEx3mDCCtvU1osVsTkh+h5MG
WDl7yxVNEdbsdAXkEHYCy/yqs7Z89sSi30KjUgt7br8tQ4/Fbg7BdrJvT0jWk2AZj/EBNb+7x1u7
qDawu7UL3pvjhVmUCVCSLT1n+bV9xa9JV9oeU+I5pY9g6uRGgqBJIo/dvoxWvLiqWUbMfrEvt0LF
iAxKeCUsFSQ4UlpwOT/qAVXsGsGt4Wg9R9vKrBaWrp7Hg3EgdFSrS+HPt6erdCySY21eB4WZb0iG
sPnn4uoB0kift0DsBMczkeNSm+NxcNsRG3ZjRcvcBXdb1soxL6slhK4X8Sua8DZdnKGwb1DeO/9c
52LXNLJ+Ut89o9wTHzm7T4r20GeJxYEhWjQ4r9wfvozy7V8JOOqc+vLQfcBYKQmdd5srt3aUFRzN
pGRhjNEPJu4STYtbu6LLi2vPLgxiRtq3pu+70t8sqoMMCaCI/rih2ks1l7FtHjCv651ibE/R8oZ2
MaAcT6krG+odWpRit7SxXMqhsG0MAHETin5JFrm5Ul1IwAxrzyLYPzvLKdp3Bx2IQ0SSwMIhb4tv
htmwrttHo+pYhJYcAy8/gtbrksCpC3WPZ2hBdmiCKiEae1LPWflf4mS20kfh6dURn+B/KKnzIpx+
w6VMfpDrNMqYvzH2Q0yl4D9dJF9qWNepWf/48/9Y/PQJyFV6R2NcUV/FGobViLkyF/RodzUUDcTp
iOxee0MMYNab1cx+ry2zjORfkXJJ8dHqXJk5xAzPpxtmGxXNVvVu6QeMag8lUtnMZIJ91PcHV1vj
lHf8pLKxDgdTIx730hwM46Td6hUMTrQClnl17t2a7zDjmsen/qyBdfNeP4LXTEc/pFI4hsVbqxSn
9sq0t/c5AkifOBvl7k2ybidV0L5NxCHb4WxK78AKAAFldIoZPTGNCD1r028voohiF14/DU+tD3tj
TucxlNSRoJs6NsbEaFbVBUgWE0RSQffnOApclMc5ggiH0ZE890FIrxXsLArutsUNRGfBjApgFNNm
dX5CAWJUjO3T5C9UMNJXpdmcyUAOeYQM3FA388MvScfUHkxiLOowL4XCwb/LxdpMLzolrjKUmkE7
SfBmSs4WeDatrpuzfUNctEM2wQSSiUcBxUtb2YjjWoHW9DTv4LqPO6lqxz/C4bZmf2PIn7Ji2Spy
s/xcUJhHQvB7N2aqBs7RMJ9PIAB9d6EPD1PvZF+jYtLd8tx0SboMsYWL+0pjRRbwpn7LtfbFP5UW
DGRF0jt0UKWyf1NyHMzme/hZWc7t/uMRMtjTMKzzKLjQZ7pSBDlv0VsgrHKENLtwiGkR9HLuGSq9
WbqB3Z5ZNGCubvMVehaQENH5GMmcTQMli7Sg+5EIJVbpZ0vveYHNaq+ON+e/ou0B0qsuvCsJfPzF
bq+2xS1HZBx7Vw+nNKPcwTDMH39E4W99N3muS2ARG//uei206o+ErhhoRSUXvGBRhWu9MWe3pCU/
N/geBMRkpUmDWnX5uZ9fz8d24AKC0+XCD4SOjqg268/WsDFB9FpITexhDyZpxjK3x0t3KXHMGOSM
CTWOF+bSMzx6FOI4FQUATy3Kj8kSsYMBHeOfABZh4N0rbcFlLWNoRlf/Vjk2dvfX1IMRKHftY/cG
MSDleOWptjUKVReX2ysTrZUfv6+LCUo4JeJaWoHe2+CTjlrqYzeCTbTXMzoeRyHBZn4sEBY4FMyK
7RdU+ZU0bTMY2OnWdBzfZqF783aiPQM19lWGCfB4W57M7nSVAvD5GIgdjFzhjNa7SQwv3V5V/nEh
FAHH3ta1ZQvFmpxh3GypG6zWWL/1ujXQdKeYF6kg+rcF7bNavipvGAkpsWeAMRWfuaFSRgNn+tLF
+BbWCjTJkxx/OBEqOy9NMb25sZDvUQh9s6YqHODwB8bqpDoR75B1LS3KGaKwM4fortISGB3EijPB
UjCjI8zMgvqISq0mnnu0ZFZj1VHrM1CtMcN7urPmP7sRiuxMiwqr3igQ3Caxd52NKfsMs+O3sbMz
eNEajGnbO1Xf+JFSuowcG6NuPDU/dvT9uxqlVKoovj8Os1Gsc2l0yzJSsZCzFHjDIf6z+suNEj0g
k4yOshcCbjW573uN5hbsovTJd0h9ljBNB2TsLp5Aw/bGhg9Sewi8fC/aewV0sgEsAZLOPdF8Y2+A
ZWfG6BenkG8uuK9W+TRP6wG0Kx8ll3hx/cnhdJOlQvEA4sK8bTNjSLVaiCg9qjsUtDHkBKmHn6Dt
0xNIOayAKrF2PZbzyPhOUJoV1+F33QHIvcAcomdJAJm7/95//7RHxLZvGRgf1bDqXGqCknOZVhj5
jVuAcv80GaCX7TU5p3zab/hXZpQlPD8HYfoxL8t+72dVcm8DMbnxYjfdcDWgmuMaEyH0OWOAv4A9
n4nk0LxKbOoT2e1juJaG5+bSMkjL/SoNIYTS1Nl1NsvHrplG5FUecYclHCfDpNqSMNPuODSjLt3i
Cdcec3FSLXtDN9Y5MLFi7XHs+LvDEQDK0mSez4nDSOf9TWSknio7bfiUnTP3XJrIbApwRh7aOJZe
C/B3tW8yFjXSWswJjm9BddklNAtJ/rlzWhBhWzljk4mhhenoqvnHMDYoIzzxOJFeg1gpt7nsV9Jg
A2bBXuRHb0mlWK53nh5VkdlEj5kY7ShIzcxAZ2ea1W8+fDFKR6S9R7z8fuWMfLYn/T407Wjurj2X
1QPOxSwslx0x1kU88WojSFJC2/eninA3L3L+LjvGPk4M582DYnwY25ibHDJc6S0FORE5TL2LI3GV
niVnOE1lnDkmX53bfhXE/OgAgIQA/1ZmRcq6Y7cL77rAYiCBSFtHK8G156OmLs7BoRahUS+v6fSZ
pqrGTltlERv+FaWMBo0W+j6QOJ3DgFRPI0t82THsHXQ3V9ThW2Q9J/m28RLbYsdukXATyMxAfOvm
Hzr45+Igqi2WOurCsTOyeuJSc0HCv7ksEHq4LcI9S9a1UqwwmUxP0z6VdP3vESmN37Yjrh7rkVUy
nmAo23xjoLozpL5KdbZc4JmhqZqTtHrJQre1sxKrE0fMn6oOZQV+14PIi3nscxru/i7wrivQsHTD
zj6OgVtj7dT/pYbiQh8P017yH8DyvT1P9moambwSnU9w7TJJEaHDoEYFFQ9eWMHmkuaWYFfzidym
1AvF7wsY/ieMxEDjJdablV89QEfJtoI2Qs6voBqUBFzPomtfpFLeU/aFahV4O1+KzU8L4JnqIcip
mrUhsNQ+DsmQVHRHqVZTaSS/46MsL7n4z1EPxcA6lZEQ1W96uWkbCdB7b3CUlsAEAdi5key2yJQj
FgkiwcCjDXJJb9SPcYCizDIpP+dbr3cr63SzBUcr2jBAinqjYRr8jgNaMU3Ki68fohQWrVoFOmBR
MjaATtPtl+uf+R+lQDciKJUhs4eqRCB61/0glYODpaX0shqxAgcM1CUsYz+m4iE73F+ucGhQ5W8J
TwRFkm2TH/hDYl6VZ0XWuOuYfAL02lCUhdnzTnoUl4sf4v6qA7vFltG4WtzTSUaQTwATYT1IlSBr
O4ku2ORoDh1TjGbn99saQRyQxEe4bzKTWhVNWbCADrNnir+W5hUtSbCGFq92NjwCJBbiuvSCP21d
yNWGCa4kQfAD5xd7NomB7LgdhpulbFOsSqWbTI6dIDb+FZ8/c7hb32qBGtBEiF9GEt7c/+rgS6wY
o2rZnqreFjChvdK1nVo21mfNLD9z/t/ih0gGH5xMuonZbR5navezNM/TLH5rNmV5qJzVTF6JnRqc
HW/HXVBOYmi/oKV1lzzp2qZ6csYTlBWwDT5gtm+CelPedkmar1u6caUr8apsymX04o0TaTg+4sy9
UiagOGqdsUqcwXkhQ0ufNQdF3/uZMr2yeBwUduY9Pb6WJTr+96GlvvTmqEGFBHm80liQhJ73yVNu
k5EKwydgywJ9XhjKaChRlCpfEzrKLcbolTed5H/ZXnr/WySazNgG2HTiDGs+NssjBsLB/f90yXyC
RqSkAmryTlg4RpHaP+iaiWHIpAoFBUFD2RZFdfzSEE8ovPZzOzGf3XL/xRBhf0XVX8U72QBfKFWt
pNeJ9XlLwoGbfmFax+zOjQEfYWT94Bt3dAn9jTSlwQmYvCdSol++aNhHG7tOXrWlcwr4S+jrKdZ8
ztz94KdAtraHzTStWz1fuV+YtiIo2I/rb4Zm+1upbfdm4mZH85JZyCfC+ED9XLchOVZTCAYzz7oT
QOdhvhdbAedlKZ6b3QVetxEVwuOALI1AXnbwgJvoGA1PF5XgQ4GT+YsH6TiZZtDoZfJyDnaF0b7/
1vbtmBoM1o9nI2LK6yj79FU57iiVUQIAqQSgGmE8a5MYrP8OuZAnQR7dbisnTLs8EYhw/xnu6LXR
PTfOe5C5u1I8ukwHF5dzsnPPxnleTueEdTlvhR1KAVCJtahAF47FAHhTTWZhCSeNyfkXcZAPjUMD
fq2/82rOvClXJ+rGpYIk8t5IOujFkKZIEsPCDgMXzM1XXXirNiioVUGq3Ri0BrCIdVXa6q3yH2yp
fsvFc5G6QWAYo/2rlZNjieH7y/UTTKgEEtCCMlxP5mYdy844MRICYorM6hMLpiClxPyDb4bRVqCk
1jamitzvWGlW2xSTaFYWAbzohQ8Z4iI7yWBKb4x1r/1gUekA9tHJAKv5n/vRSVeUuvvUnFQCJVCo
Pr7yKPhFphpUP0iOGaQ+DUH9dg1zNsgjv0idUPu001kDi49DTPIVOqZqx/23Sq6I3oOB6fI/ELRI
Q3/Jh1jCXZKILgafEMhd/WKfvhtR/Ym14prsk7wvfR4fM13nHEnwUvZhlzScvkb19NOpdiEqmWde
BzZl5MziHsXbFa0Jn9jJTNTS68cINzsLdrkqnwpYaN6JJBrTEw729ztNXsPg9D3x57EVWNhTr/mp
JmzZKJPixqZQE4brOwW3+owYKX8Ruu/l6zBjmhunNQacX+FJpVvuDE4RU61rrolrLwjALgLEHDCM
0mkOA0wlKqyub6jrD1UjQuzyG6Seu/n1lG9xsp6SoQAbLiqUFjEImYLcLMt82HqHdHm+mmXuHsdt
NBTS+3DDkdAoyiEsjeS0zoQ0CrxsxinbpCFbaXYDRI/X3cnvwIv9eWGZHTCWXawLx6ux73EIZKmw
ziRxHxMXsj6dwepTuLsrwEczbl4FB31wbHM5WbtPqQ3D3cS26mr6GNyQ+9knfSGAhvnD+1mT+EHo
W2wNWcxUpeNK8a16VBl4dFoo5iocXSVPDqhU6ZGWoQ1bY9bLhhQIOiwvtEBGh4tDxTO6gB6WZwxq
fFTAexoyf9Q6VKlNIYuaVp2SoYGxFNLV9sIbfMT9WaM6P/GIqLIyYvhBANDl9tLO1mtiemMgszxl
XgBq8pdl8N/XQPaEWw8kqKLgJ8Rd1U9nQEa9jrLTR/sHIocBmvY9zPKT2usYkbIVpKShuJoBgAd+
YHcfHjvYYPUkUdeRdxoIfvQegh4W5bQ4epdCfNaLITt9kZDyfnIGwGMe5w9yDgBL7dnpkA5+F/b3
OrKYeFmnCtGLGxAMFh857vdTXj/+wPHqzsscfZhA/rqM+X+e+a/lGH9EfFKX8Qk79c575U7O6yZf
VHphuf4TEsBoz7yscdBMtjfrtEPzRulnE37pAIs2wRjkpix2qmJS4DfNvqMeTaDeY99AgWS72o5m
pEenq6mn72ldaPS5j/QPM5AxTnJ/KHfUOKf1GDQJwMNXHl3P3kSUnTU2n2VkEDQKzEjYB0T1l/ns
xFg5OgE2lvPVScv0hDYLDRoCohE3+8maxEvezhUcnKo5F2f7qC/EVnQo7LS566C0rQzgmCU3rOpD
I6fHEZf1J6LGf1txOOhumOwi2OJJYarpSXJ99t1Yz0FwSRUpdIzepF6VAeZ+VPsZE4e71XyGXeIE
Bei7agfPa54+cuLKYK87I8Ce9+PpbF00rl+auPkXpAG56Bixf03fbRvjztEivy//IZuJibRsJ9XB
UpJcuNQVqvsxAAVz1NjeSfPzTcTwDQ8a8b1xf/BFdmGzA0KuFLxF/zgtr3nRxBm+WY8m0OKyOxr3
0jNlyklH6qcPnFnatppMtIcZjsw9vTPiAZALTNA/ATOXFtknsvhwbb30RMmQRWieOvaxET0F/A0j
hhZqb5axP4uIIiHZ6/BK86JAg+sbTQnDfRPiR2upv3QPDzPVSo802DP3pkNFgdKe1rURgo7+qVFe
Ap6EG05HJ39GPX5DRlf2lwg2A+2dJ41WfH0fQjCKR3DWMFlaFem8yxfVSWCz7MDr1+4vgbIaD4/p
umz5GVeVv3BXdeRXVjk2G5/7V0tcNYdoyxnEP07T0GoVJis+D+p8966C2g0YRf82ooUYhRFw0c5s
8/EHpXFFomGl41QyeoyMF9fgskzJhwTHKAhNu7hG+sXeLh3m6EueeU+1DWeWydRmQZYeXGHENUyG
xujwg9zUsBsIX1Dd1IjAYPYk8pp+sODqOTlH9gSA/fyXB5kIrn4NmNxuntLXMv/y+DFctQGdSjKe
ytXqQbV16SNXfnpNDthvwLGcBOxOaeM5/oecNGhpaHIR3sToX7q8RE8+lw7kUaRKDuerWJ4ma+09
kHqgKmS/VQv6mMNOBhv9mJ20GFUvPaRhldgBA+C9ZFKMtrc8tSVtmaz1ZiWdfk1ICSeEikJ6HPrq
ieodDlu1nLDdMOWRZOsNLRH2NzXgh1YVhPqFIJaSXRHlGdE6l5XojTrZrVe8qKA7FlMoEJNRdMSl
fiRlkS2xEuzhFvgLXA3iC5/gnRuZRPRHMxZ1uB95uLbDVfDskh33SD0PFxGoj8VIJ+xdnO1GMQPe
OOw8u+jigovPQl368hW+7DWyRtOfBdPyOc6HaRCfV2hzuHzyALGJIJERQLv6qjRMWBwUoZc5EAdS
zSP3BT4yhQfDbyNNOfRs1r2OITAvyLJz2GT970yyAtcV3fm8LHplZFjGpzRgqWmkdgfBzxE7bx8R
OGeHYfrEdhdeaVurq10Hf+m/2NeX3bLhNVrPCfOLxhYYp8HUt6B0cQSfOhtdoKo2MTMtJ6rWSncR
8h689R6M5miQtEzmGevqlnmhrp3uTOsEx28FzTZuIYYib5Ta5EvCQSxZaBM+j2mU3CMhq9WgmSbs
UFT8XYMudR+fIMOPR/E4cpK9ElLuU/qNvWvRt8zrAPkotTBEinvyHJXF70xdhCcIURjK8BWbGb9U
ZtdFiaBQUlcEYmzGgWo4TTdIwmafkoDWE9jwdrDKV51xv0ROt7RB+ccUYMEFf2JO5ApyfT3QCCM9
2R/xV9DYTmHX2unNNtQF/k81KtnZkYsmB/qvJMGZec4WUkr+aGOTBjMuq8miDEjg7Vkw9GA6Jr9P
1Atg8atybTP3s/DEXGEoEQ4gu4XNEZ910pair7xO5yD+hCKEIhdKzsyYWAcmcCXfbV1u8fBq+yVI
q9Qs+YxHAlp0N+5uSD9RIFSv/biZckuOKVqqikGUI34b5Olg0w3WPYUBnLMbHzTp0yB3EdZEuDVU
VX/qiAZT/UP3PxU6etoiFWw5wg8SOZ0KdvsuKhiHXb4nxWGU7EaKCxoVJRApDu0yDMS+AMSIIupD
53OSQsBhMV0jYRzmGYUMUxBjxT7mPh+LW1lTDTgtRCLU9Xq4Kj3gMUCr+z020Q3MSGpPWiAg4O7y
sn8gk5qtJOGHAV6dUItbuZDWA4jDaoeRcoacQ3+Vi+H2kV6AQr2Wx13R6hWlAJ6F3eoODJUuB+vc
yP6fobDtFphCZjZCDUlsD5h7KPAmjWy2m1zRNsBVKq0U6yV+XBtQyuk36qBvvC7YeKla/OSEvdzC
LiE9ohVX4pecYxu1RjBVvO93s6ndqqfBAVBTL+P7MIgexTWlvfI4H5MlVac6ABTUCk18F1M5/c43
ss/DWxyhZH2fPVQuInQfhjtZssAYXwdnx+ZalTA0eksR3bz/0/MENBdSWbfCcIPVnvIKWterAh6X
6hnEcjZt//gdyhJGCZGRRtTdYs2uyj10cV2XJET42gwM4HSX64gGToP4+Lj3/WiI7BpUHSDOzL9l
bTJP0MQKzlsYdvGXCiNlWM5C+E5CGBoypy1/mnNh6V3AG0h3pvYroyfGffuZarh1hmlexQIdtc6o
AqpEqx9NQVWcFqBbfSToyl8C3iGBf+A0ONjQolq74qHSTPxPTz5CEEOvtaYucWoAf97fcN5GcUVE
6GDXRnahxVdnkqXOnbq5tVe8fygB4aw4DSI1tG/p0zxXThT27RnGNrW6sKTsbO0bF2dN4A2zpGgl
xzet7Bfu53wLvMt+98HSPGlzEL1l28AvrA8FJwslYmDmxT7Kkt51JNY5jsPNmprUuCadYlJP1e9J
IMH5xhcxlR2MffnUmC436dlaSuDnb2+ddk8YwNFiD4amOv1waBPIjiZQxxoUvNQyk7gqYCRH7RYv
lL6EXZ1FnBwz86jss+QOeP3x1xg4IHYlfLp3MlxiLcsEygBiKh7kcT0573FWZ2o8VxcmnhFPfcO1
4pD2k6MMfYBGOnXKP6EtdzJS3/rA3K53tdumuvZVm/D/jiYVN8nod+ffp7iuzdRF8SdNrTgmIy9r
SCxq6KEqLYLzzGr21OfRVhvEdxqMYQyC2pbWSjsJD7MmMTZKbzog436071GtdwwvXSJw/obLeNrP
NnQPTyruHf2c05N5MsFHac0BY/in+ErbKNz4EH4RkHHLYlwk/j9paPguRqqFx/RY12NRbX4JFqEi
cU+Xf+mjrTu2/GNaAgEibsrmjpHcZEWLzPCADoG9T6JN+3Bq93UlK4mimwv/UC9YPmbF8VP3+P+2
jHP05HYbcWG/RbxpqTY2Mr5SvBaQf0sg8wCqrpU7PFkexJKgTvHZisL/STDCy+Yn+A2hCn34tiat
C2iCyz47OOR5i5wylgY0tN4t90wh7lakfpeP5P0p+0pPduWsBjmQ9Q0zkBOAUt9n09oc00KCz7gi
FB+oWCQ4Spa6ZkdLX7zNc4JfD2Jj5PcDDE8CUAarbd5wLt9WqtyhY11guArzMd/0kggpcuu0cXbl
iNmu3mWLu1h0V/z7cL/ZTxxceYidhK6QjaOcpH56+Bwmm9LPOe/daftkE+bAsbpiVKbFB7ndoUOK
MvSPjaaaBZ972jwdYR9lttkpz9/mnGi4IdkWFylAeqnu2O+VeOPM8WHgdF3ZrPWRgZrDdtRBBe/r
e8UAD5t8DtbyCOsvmCro7yW2pZbh8zfRdUfjQfym0qa6Q1HconTj/j2FvzlhQaJ2MQaJQGV9VTdR
637kpOkHdZK1NztGflBVhUoVbBqsTmkiDVZpuX8r+OdxCoEkgRdki9uu+b12s2susS8zdmHcNKKI
POU6JG/gzY1HNAn0YJ2RD1dqJntQgpEY5aWSWFNRv2o2ETYj6cRSp0zcjXKnMmKuw6ORqp+AacFD
JAvYeR93aVqzKobL6UhjvPlDddnac2KDR8QW+PDjggt7ooex1nhzXxsJ7O3fbFBm+CmobhVsxMfG
DUZU4VLWcK6Hewcb15XwV6OHxaSQrBGnkErZN8iB0VdHd5TD5682v5QmOQao9WjRv95IsVxKboxB
9goIFwm8wpQwrUNQOl0ef628PJ++8Xr9SfNfZdk6axLcIs7XvJYabSIIcihV59qsJBRNNE+yrkif
lTcOswrdRoWQEzlE1V22TJULDverIZMDe6k9jB2Y7o//FYCWaK7l9nvpSYhpnO60SwHLo1EKXG48
8k/9xihOVVzV6d5UaNBlE9xen2mzOC1corOgYROcRYBGXxbJ37VZYzR0SK7fYzOF3ezrPrrw+KdR
Zcx8PbDOZr0rug0bV+xVCBdepIVGxYv5NUEA1Csdd8iqVl/1Vu3Wt+sRy6cpSRy1zmzJzQn4lm3C
Lt3/wwRbPnwjg1mqmZ/mb8hHxIAhUxqRzYEOdUQEmm/C22g9/aWp1pS+J9idj0QJ2uHhyxmMicBq
9em+dgtWS5iOBCZbDO5JQadXcQavC1V+Oz5b9RMZ4tssrv27GjhFW2AI6v79Ri6d4PuH4nl9o2Sy
SmNnJ7//3V4pWD56nz6ad83l7r8GQW8KgE8+FEKuxa8XveKiBnlNq5MidYfOlRGlQKVuKjdoFXdU
voCAe1d7i08PDOq0XY89C/zwE3LDP6JIJWmMnsKS+/hw0nBu9j+kZzL1/KAJtgt5rqtTwQc9zX30
QM0aIYK//25xdvE7NFyd2IBNnPeFAFv/7svdvKbQnYLO+eUcH7ZHMIVqUVggjU1rnI/aqQ0E0lsb
B0P9KC6hIZYMFicepFJiUgqpDAgOlukmyDIQD+yZ7S3qKeTv0pCnvh5y1q7sKAme/fOuPufEWJ88
ig9MLC+ErBR2uccflqqyQSc+E5LEG7UmRgisCooJ8kKs5hddXqqPDDF+6ntdHFesZ2+0D0Vb/pUv
vwQPZTRi/ss2AEGJSmvVDnydy0wUOJNZM/I5BFLQ2wRDgp3GsllkhiGJ6g+9iAylFPCuMlzH5COH
pLROgqsuCSKBajwe0eOJF1IV5kSu9P5Bs8ChJp/ycyF3Bw/aCfkJKoF9C83omRiBBVz9cuWxL7E9
5ZtSWlWGzxzg5B2VfSiU//rSYx8WlTCbqWqyiAzcGjGxq9vNIim3a1QChwu0NVUdyEhYzpRR1pN3
ROp9FOCKW0/e1Mi4vPEXnL4sbQnkloKCv2/GMQ3fyVA5rbkZvV8uei4QQLp+uTxQhBU03ZK0+S5S
mXU7C9yBjSQRtVhiTI3zxBCs6PNjk4WQ0x9VJQvAGbqsHHmm0q/TtBytVtP/w+E1dhxNsVU7/Vik
FE6q1WI22bENwdL4aHZw3Lh2aIgbyWRh9imE9KIe6ABrSSf1KFoaUTZpDb4sjrZNxrHqG1BC+a3v
Zopf2dqX/4tqe4DM7phnlCOMMUs/FgnPU7FbjorR6qLRYe8rHgBm8UfF6LVzzru47SwESWncUFYY
RvPkl4Bo59/GNBZ80Mj3ISEt7gxn5vvakh57RDLVxBwm/nNaZEe+u8CFrBKPYSAQN0ILf0gap1ak
LGHBebd34Y5uUTrxBSHkGFdRHwV9ZQQP8JRcSzfOfeL7wFh5k39TYMxlfax0r5qYAWLc3DlwDxZ5
QkakQtaW/6OguDhHncVQ4SOVFR6khHMO/Zv/jF3HkUFvDpxZtvVuL6DzPUC2jOr5hpE9ia9zgKM5
IOIGJjUCupPpRanjhsNZmcAotxxrBthDHFFnq2eSqbtKK+9bXJMfYKGS/zfk5ZZQQg56YgbdGxNu
muhwwIKVqCN4c1CFgLTl6KOWShIK097Hv+cmIQqMbbWzdutiyyiCDT/wztRsroYtPMXQ5VZ5GMNm
Hv6ePVyOk6l+fvLwSC6KcBtNS1Su+wI0npTy+wR/Fh+y5JcZH/SVMV3matd1ahK00vhvifoevSla
bgX3eaVlvxQH6s9ZDiO++kOw5VG54/ksuhAAYpV0Q/4gDttt1uEx6Zj3bCGS2399REwnNMXPSh6+
ZkHZFkyksnzhgbRqN+1GNTWbpZ/sl4R6bjiIaSF8VSoyZTLJOr+WSx3khRVCrz5riCqVwv6XY2EA
2mnE+FiAR7oWPytt2z3ZSWrJl4mh7AxpRJSw5cfS2ChXFM1b2KSRLCa2wBTZ7b/Q6cFp5rsCsfwb
AcHCD0cUProsRm9O8YNoyV7inN9S449tX9PTvPvvrEVz4LE6j+Pz4hQspGz4AgCRsYtb8LDPzS0M
v+7o/UfIjO2YSrS3zULzdkjpH2BDgNgF7fuF+eQnYxnFmfioLH296UihCxdJcA2rULf6+QSTg4kJ
6zc1af0QYobk5yKnr9MJgj23S/3x631OP5YEcpyFRfi/fefUlpSJD7O3C2sD6g4z60sd8xKFk0ky
8vjf2jXO5/DjweLHj2xu3Fi6oAd0sqtJF2UoWryyJHQmW+4I0rHtrqE7G35NUpN3cUzjpLAMvhgx
JxcJYzpnbm67IXCa3gcAQo06B9VL3TwZPYRlZvXMrmk43WLicm9e9uO5RTGd/98XE536Vkc+lTkJ
E63We7q/hC7L1I6cN0Z/lJKmeeZ7+H7xebmPpzaBuvJGmv+DvJbiigprzu3cNkx3C/ZC3oXCAIlL
67Yyzl7TufiqnyNt5XZ+0wA7uK5RqijrnvoFHDJeqCcU584q6IK7dNlI2segvggfgT40kv0Zjcya
AMCycQsGaiHU8qAfEfoDbbq2IpSCDvqCqsqEF4S9VxceIAfQdBK76aSO5zauDhHSzC10pu4EChrN
SI18jwHtdC7N+nOs4xFLaEF3yUzJ7uzI19PX4NU9Oe0Keosh04V4L2pM5yIsA87JHngPTSrOI6Gz
ymtCi8DTcHTzfc1RN3pVJrLd9FUiq3YRaqjqsKwWi6rzshusufko0f9W8hxbuXB5PXL8WWGoEYJG
bnkqUJV0LCEVYj7vM/r6T1mx2uMra21wyg6UzahSjYxMK+VttEoZXdijxjo+Ptha0CqzjDc3WmZ9
LcQbUY917+O0kw4Tj57fho5MqDjv/v7ia1HbHM7Or1Bq5JdNiPwIxSAfRNy0jndu9I8T+sr3hOHV
3LVYjY7QSeIm7WQ8yzdfIYEQcgqSgUmK3xZP7LFFxJKuLZpWrjJRh7GDa5szc+Wi2vd9QYKTN8/j
xuroWZaw3q7W+DESXuqABmpA1YgidknsuFBQx6AoEqc/fMRlWHVwGpywIymO/vAYo5SN9Nj5osJn
VblyNyEQjC+N+teh1W+jTQuuL5rNxEdxMzilozr8IPpsBxrUaGXkmIrYkAnMaFZHy2tE+9diDS30
+8v1sJHsaNZ1DgUCE+YE4bQrY69h+vE1y9O6BJN1RAUmNs6q44vgVjSpEwioQ5hIyDB/OPh6XNBf
EGCq+9mhCIvxQ/CQJkjHzO7qLS8uUW9EYkXlzXwkPud7y3vnb+RXSTzKRDoStCNTgdnNWjFDr085
iMMiCHDtsSl0KDdFGZQ0EZ+den0CL37tOGx/B2GzK3zwh1MoDkq6IaWRZXuFFuoGmIrMey5sB791
O3Vk1mGoE/OYDTqEr8KPgXlVTZ/jeINrRCmvpmuHXBcia4oUevlqHGCYGpiZUgjGVhW1K3Ye9l+S
3vWqq7UJpONuBoQX0lapdki0A91kUFkbz8+lz/3i9a3VoohhOYFbZAu/avd1psoJUeNXcNEUJnfX
nZ9z1JDI77G2kVBe8Txi3vpY91jGLxRGh2t00N9AqK1cgi2AU6TH5hrtbgGwVf/wiuQnsmcwT520
2noDTYWtA5gM7gcce2riTwQfEreL4t22uqjr4NwydboikPvMFnWAtU4aJKetRqzi/K+nAWkzk8bY
k+DPsD1KI4q0k790QD793diixgLxlNFthn7UCaPvRn4luO9Qgvpf4UCyNe3fVfavCNduolZfrwFD
2cnYDPC2d49XkGAds3mRjIpBUjaBqfXx3+Sq6Yb1ry+qGayWSLIJPSQvmcnuGadg0cC1+z5PFRiG
Gkpf8V5N3Gaw9sdaYUPQHWlktaRTGVAdcZgb0f0nn32YDc80tIS+jcCDLBXecUnXEqdNIZrTwfYJ
hNpPf2/wxorAvnaurWvcQ1PvbxfycTnuNVJJ8Xu+9+wJ+K24DAl301rzi78+1D9F73oVWFrJKPew
0mOj1o49eGMvZfKpLR7YPLf0UXpWj1p4OcAdPond+5Y7REgUXBpyY6RDmoeTcRRjDvS0dB0FDu4u
qnay4mgRXYY5QGhT13WwEPa6vLXqGYNfD2vbnS8JXgQFeM8flatsGaDevXyG1W5PAkC/VXQ68Fmo
NoZdYg08ycuwY7PnmVvR1Gq+zeFm63bvCYHMlcBQjUy9GvR3EgbxlCw7c4orIpTFL3xS2yoCYiot
p2sfv9YPxf0rohhHQm4/r5TYlgWYkjRL0Cz1gxRQmkgyzSaVV0scHNOkkvRm+OR1deJa4DqxlfJF
f7G2gVIta+hxtaGgnmJY6XpFUyir6TrVpJFVJLbLNFzk2jQfUwSFnwEPRtXNdmrcKkYLwbdu4rEI
t/LbuVBBT9rwgsJ6ax1wg6idPj8oOcao2MvEf6ty0KOOal/192GBvcTvGIqIxbIXXwx6R10ob0yt
TjaafzXAmnWIoTeS+XhfDaYQy2aomlCrZ4mEZpS+BVY+8yrusLxhjdHRk3EVgoDw35UsFkYrOm03
GZYNCVtl+6tg+9TDVmP2Of7SWY0PkHAd0F3l6MGQ/9ixe3gOOhP97pcpIjYWUXz6V/ihVeo6SU1z
18+V5eRtJ/xhGS6gjmUPyClmQ9ImDbqt4C9dT5++SOjU41nePCqG11OByq9+Srz86y0l+KcUglU6
JSSgu9Qmg3jhwnKDSzOOimjL6skhpgd6RLmmxKqxZN7WjnJ+YJj28h0TFDKm78jNVm+d/m33XfeE
aXRGvPN7x335+iB6oXm6yE/YHE83P7KBe+T/mFnvef+bBODSTw4bEqCQGCUdMsvRiGN3ZInzfcWd
f6UHmVfvn05moWhal8xbWBWxZ2PxzMFYc3puFnYZTg0WnOLhPeBGaBxeg5Yfd/0Jx5xuttbrHidL
Ni0XOK33/757WycVMmrqNH1osq5JIh9xViuH4ZuKiuc7BIfNmV7KatbiuadSGS0F6ljR6yMP0VVQ
dDS0ywMqnDbSXMQxBqsRC1KjhcFurC9Znqh7td6SaM/zlKWknl40Mr10TefV6sddm0eHE07mHH2Z
RSb2Ihc7OGI/HEK0XuN7wbys/5f1L7wuw1Z4FnuvkfUzKXjsCZhFcyfcsNnRFh2YajstjA3dgP+Z
paWtw0ETp6018+M1kddF+a+/6tVBQunqy8JSBHuXzySltfXV1DnkmgPFlJrIGImurLYOjB5cZ1KX
genS+I2RcH0me0f4Xo1jtCcSYdCqe3HTXUk9GgUHnUN8trRbJw2KNVNq2K0Gb5/0vHUKoEYHSVkt
kXfD4HxaQSUINNYSQosooo7DBJBSaSaDrq/9LFjy2g52jqWPiS4j+HcINYBI/saQskDEr4o92C6n
dWQFXKqvmEQxm+s/PwcDAqrowLgscb/puPvY9oMFNwWSNXvCtnZ0Y07GQZGfFFEstNLZTLw4upix
xYYKptI2IMqh+cXaCvkiLomejhIvePnbJIogjfXcU0K00CLRsFoC0IXK0Sf1KjYYmKB78Q/Gl36o
fMmejheSo80qWPdB0SCt3JdiaPRiDXh8HHsCaRMBJfdadVccHlCCVVYntA80OqbvyiSPSk+YvV57
EvfTclRx9OVjydoE8mEuv+/PmVQgv31feQ9hBCKu7LkRDcWCMoL1CJDvmmvaU+8grIUENTe2gcd7
/jPFrRQYDcU/KH+rY3tasd11TmYpQbQmQIXw2hWRurzjU+9IReDZAmOLmhlSmC2ZFN0J2H1STh6x
VTWChf/kcV56jX6boW5udGk/uFr1K/aWxP5sjiSIlT7rC5bdGtClxD+A4JwelMhyIoZg/BKiGxiL
pHaguBU60hA9RfXPnoGvNPwingmUhXV+zVPqIafDjAEpfG3dvFLfnzLr4DMbn2bqbgpDUKWh15tS
Ir1MqLoAlv0MLAAo1vpzjavrpBynF33lXbPFn5VgIAsXrXnZUQHWRfrqXT9Bm2++ECLlYj95jrIy
UR/Y69+PquZS+04H6LCIgRfR2jc/HhKdSS7tGD1Nxu/IS4aeptdaPSHvaPtVfO+CPb+5sOiJ1ybb
LBmCWC6GywilX6sDGrlIEBIYNMTmpx4YFjkDNiOaxLn8m0XlHrEIxxJsht9zxOKaAxKm3WsmUZvN
T+atUlQTHP5x70ijENMZS7nV4JKgo6q4DNOY/HnBLO97i3mes12raflc5XSpsOsjsBDB61z4vRit
u3m1wW+PIYum7OZJoP6W0QaT7IVGS8D8/dIiSGWvYLmp5U1laooJUc2LwFYXywot5rUnSXqUr3mS
LaVB1c9UeWnI56rCXKCC56kCPtvLMb1i5Mkn+PZjhX1cLTS36YF3wdHhjWVrAMsJ4UPPHWZ7HupP
HvUAjLiWgNGiCNfsT0Tlivv5LSpYy6i1gBCvhYmeDQ+lKmqwAIQpZh02Kyb3ZznombS5fgtiLiME
z0zm2wRlCVgukZxJNvKqcA64kf5i06Pvkqq/EhX+RAjORCmgjLAcgeyUN+I9E4iOCgrkeGCjD28k
uGaz4S3damp5WzoGEbQhf22xM0oHdrPNISOYhDsUn6EvaGI+aY0yyy+Mq3zZkZQ5AJ6LWC8RMu8n
+UhxZh92oCMS6EPYthKb5oErkT4g2kOeeLpOAaZr8EjIe/bUh41Tb8JrJKfH1vuZ4tlY/EJRwrtg
pMGzV2mbqIjJeRMDAFRahJHEckMScS1kM9UshU0/l0+KJWPMdc1nTZVhRMgRYQb3iFKdo6PxKgXq
Zm+LlpHkO+AEsQfpMHTdNFlvyvArvjbKEudlJhwYah3FqhdjhW4cOEdLdNyPXCcAcnycfOi0MMVL
0Q3Cn8qt3dv+QuVRmzwW1pUdT86G9qvDh2pAGDo4cgi5q/wixKCowbmF4KbOrWGrC05/mN/54QQM
WmC/l5RX2gn8FrSsYLdWOqaCa9yMa1mEb5kKvXSDFlorHycnb0p9H3mAtOvZsaoSyx8/7oKXbGTY
mJdh3QDHt7VfnkXIdn0HNewilSoIAHCiHTDqSjPX0qmT0Zran0flCZdhUFDwDxukOWHBxi5cwyuM
/Kf/UQQYMrDA/2AMOnIWs89SHNH2WU+LnBULLbVydwGHYKnp+Zl+42oruXFWBwVCSbYDIXPZKvJU
Vra6ixXX7ZZSkHdCexaTNMW1U1w6LJc58frHQCsVmlbwQZeMSGf2OXhb1pDd/Q9/am87BiWPoqYy
50o34tWq3cepPOUxv4KGOFeGu9JWQYW3HIdq9hUaActdz8TPHWWkAIItgvHhgKNTMaGPfz2rdPuc
7Lo+HR1mFHmg5A6Wv5t3sXifhdGnQaSt3o+7QkkfWMCtia05dhyySHPudYjx5RwCidYPtgPXM2BK
HfKbPJyWbyquc+Dyvo0eUXSXLMig3zloZ6vPqGC8+QCmtyVtt4lFX7zt2Xzv4W8t3nLrzL8vbldE
M1wZtIFNw7ZZ8BBfhDEEq6pfJ53VTe5enKTvPJEm7fvXY6XQ1/LqklVmISSJfIyZqEXDZtmRBdyh
qlP0bt+4vRCHhlRemqpeJ558NOpzeAEA2AR0K7Xv3HO8b0hsIwx6PWZcZ+N2NoGrTfTjIrtNC+oc
5FQyFXYNshSzrLjTmFAiZyxu8MEs+2N5ME9hUgOK3FLKXDNM58JW4gEnMoUCiLnRPVbK3kytxtqZ
VC7AvPs27NXAHyMIVsB3Jfze8iSE+RbsYqzUkSiIsQbNLrn+1dVtaplu6hr7EIy08OdZNSBJx5yh
hOke5AIr+u+FZB1EpqWSu7LCRal2i38wbGzQEC1Nt2v0iH9k13n6yrGJvo/rsPo9a+IvaEveveWs
TxGeF/S+NogTccDcmQNWP0WsIYry2FA4qtQOcpWKOlXSR17x/2zvu6EfttFetZ9dpuH1cL1wtl39
NMCwwL2zdsMghe1MUsaISWTKl726QHmqUA1DcV9DXEM4g/xdF44V6suFz7kYiW/qfx2EKM9Oa0qc
5jkFbhBPh8SoIX686JC5KPwpLGnQ3cR/BlRkSWuTbhq5TJVi49woBJ/ggn2JTtp5ychqP2Ts1esD
6GYi8uYeQa7GqSlHPD6XatcuYChRjU3VYSiVMjykE9fV89WuRY2SS5TX8Sm5kR0OcJB3BvIA/uiK
3w/rqVNF+7+1jv1eA2n9YLb7VxqBxsJOZHwKp9L8hgL0lwKwOUoOY6o559fzvpTtA/jMLg6LN9Ad
a2IDY22X9tOpyFezq5xWldZgZQ3r5wPZtQTyZWPMWyD3nhmS0PgK3aVawhoywKDvwRRmv26aCVkj
d7zFO23VaBGbdVErOQFQOTTXJQiEHEoBVab5M/THi8UmQUOwnOFi65pX9GlWvAqGpr7L/XasgNRs
yg2yFRspl4EsyI0p8r2uC+HVjnnuVh8U/dBM5xMsry0OlpJhhdzZhVtV6pFEKSAOZ4nE/S0vQVpd
ZbfawnLS4ocl7XDSS9wOSZwVEg2keeZSG4ZPRxxLFNRE8LYNztG69VTa3TO4OeJ/ez8URMsKL1cE
G58hlMW7lnTev+gI+CrI4D4kcn5rLC0zg4OL/p+moULPtSDF/5Ef2z0Y70wk6rwADnJ26Yq5NYJl
SL2SzawZzHZn/UtreHWyhmWr+lIDdTkxN7S770IJ5GII6RMmVChcKLZOvXS5lpvVtF9lcNwI2LqF
rrelXVWurVyTb0dQ39ToQkcbWn9tUCkhyITGEpgWxOomNagfB4FcTnzqjRz3lie9N4MqCm17L0Vm
2j5Fx66AAWht0CRLtSOtcHo8oZDE3DuDsIIJKNMzlVL22DwWLHw61RPlqHIt7xKSC6ScHwsf1oEe
NGrEtdcfC83QDVtSqudS1oVJbH9/lMovA3pTSxETmRZC79E9A71BlZJGbY1/fNhfcQGlQIfAYy2d
lL+wBiWP4OwFzat8SxvVFBtzw8YybZ33Dpb0d0M9gJBC18FIwMiniXj2a0X869NrOf4tKQVUo+O5
bk/Safvb6IcnjE811YfhZ6MsY/KS5R8Y/ihpJYf2zO6oG2DBOC7qljGXeU0av6cOb0e8hZ9vD4rW
rJgiaPy9sCMgN8VYRaHnZ7yUFvQdQ7aDdAPc7xfIdysvS9VMb9xuap5IM+0PCxVRnzmn7R27fy4c
L1Wr0CgL7XYIN5oDFrtUR9A1ErT/INoGGTxdtGvp/gF7K4bLpNu9erp/RX+QtemIlMsa9V+RNzVX
Ncl36vMZsi2iZqCYLbCIqijXOOYg7xvbrRhPG6CyIE+8v+44QHdu3Vh4LI9AC+SXsDm+Y7eIkcl4
QnB9RpWlM1RXSEvqzJd2jrCrvz0rygN1AZ5YrIDnoPkbCdWt5Su6RdBWdksQL2uG49fBdTMC8mRN
E7NloQNximPKcozKqEDzXLot5G6rXc94anK/6CiTbn3bhtt+eHviMhb9UtuZYQZVFyUwaYjV0PON
IwnD9igYc0TqqEa411ujLQabX/zncjTnPlUWlEZ8H4I+ZLarXsJ/v5QwGY3urN37Grn/G4oS2x80
d4NKmv7KqCSo7xdBw7ejXbd7DRo2AEOFK4AbUNZMvSS6QJNYPI3VQ3vwHfN0OGiV88teA/6Gj4dB
Mh1M7iS8bC3Q/n574fl58w4s/yvE6Kmqqr6wiDSzLS5VnAtU3CpTy/fObWvluakJk3cX9a2Zb83T
hYcFVDdTkHVlGVLROu2UAvB0rWSnj/jXxpqIld4NSwwqoNbXP0X6n4xvA1ZYUg9w59VIYgBZJ/ce
R4/kQjxGa01bhRecXqvrsna5UA+e7pHNYnNaCEcfOtkKCdtZ0LRuRirv9z3tdwv6wHwu0r8P2Hkm
ZS7i3cuk95LPxHfNky2e1vYONrCp4IuikUCORerw6fEBui/lq6sUTz+/LrgV9U56jkRtQerQx3Nv
KyFMfYN/gKfzgEbXeGLAJRU9vXyCtKjXsWz6UhguUqTp98kEeDmi/UFiI01/HHP5UmpQ41yAz6ER
JBXckmtSgGTqImzRF73obiT47FtV9wVVIwKTVrwOxbBDJs7JqEVD7F/D9oelDwKeRLHylF0972zE
AIEnhYbHODS/P+16zKHh56w13TkH25S8k7f8QFu6MawuaDYjPLK9/K3YdafEkpn6JvuaXn+RQMCJ
+IszjQwVH0H75Xmi5PUDXxBhMODOjQujJ/eXOgJ4u4+JEoyFNwBHIhbcuLUXd6ep5bZJrbrojox5
vL1UK0gkC3tCQLIREq2gHIs+p9UzbjH26cu+xRvuaVnOtdXdWtlfk2Vn0+LfndLCDN2wOD8nC+/w
6uJ8ATMXpKH5ez/uEXaub/7cslcDRQY5scjfAqXf+OsPmX4bx+xZHuuMb8ZWKWgC/B1zCqttFlrS
LIWkvm+mj5RlStBEVCaHJB1Kyp9Rz4fjj6XjaCSYhhSqcXyqt7vImkJmOZGIBJyhh6QS9jz6uMP6
pXO5Wu7Wz+fqH8LoSK4lSgqzaXo1WsPF6Ar2TYlejLi/N6rl9ZSWgs3m0a3kUq4Uc4Vt7C4xVh1a
dn4J1NbY9Sz5Yle46RDyWROhgtnk2cb06GnUx8XoGbgBum5ISKlKPL6vJ6FR3hvq9Oo9TaNw+LL+
J1xJbr+FAcyv6DkmXDu0w6L+6taVwPiHH8Qf+YteC7Vaf17GeVrE++9ZiKl5tGu0IesePo2xOFhr
NFAhnxcopKQGJYpJQFsaMo23QJ/ZQ5RsLgqNv7To6ohAlgPyTBtH1ZZ9mSAEQpAt9l5I5weSZNuZ
AnMmEi75jiduqmZpiMTRXIgv/2uvFUeIOGWJj6Pq/DwgflSPGGLJZYaRfFfQ9YPvTugPChOTz99z
dEq2ix+c7QS+2/q6yI3ffkzSCN7ySvSniqNCoM+DY6pinE/xMIq+KTQ6EQMDDVeD6+1+Uw3KyX+l
ILNnjo8nJy7tz3Hnz5FomS0WBpHglyUGdca5XvTrKZzjMk6ipD+MGpYb5kZRqsDW3rO4WxyVh39Z
+WtbMGiIgwHmNOWJFRyItCVOkTzCdGBCjd4g30c+QzRkD27s9G9rFrn0GZgPqH4O6He63igjBrba
lcD56xTznQBiIYq1GDh5L3KoQzKZbnOZHxN1seZAgG5xoSLb3KIF6zLoOIRZR6sKwgHt5rNRki6Y
HwXKS+N6ecSC80PnksqIWXcm0AH5jjbe1Us+o4StSjdccP3EPnQ0HugWUVrT260yc6A333qLqmqw
3NrajQuRs8cDJ7/1f7/5OzdKdeut+ardszqUQ4XlJAvue8uTK1yrXZ8lrbqHD8VShFjeUDZi5AMs
MAn0wreLJeCmeaCBOH9oy+MGHiSkNj3yq01rfzkphq55ry809ofPOXuQkIZyWxJcEpNfunIVPn5U
RnSTUt0ff/6aprJESFf5iUfm9vOcujaaq6Y5VNql3/6FJxHDP0vVjfhVTEpPjhD1BX0q8AvTS4bC
JLpdVENvWiDpdwhz1Fj8vUmdMf0suRjKF0OCjPbFAP5bynmwwzkQFHEOZcXkDhh8YXo2TRBw4x6d
YmvDLTPAHBiwBoHH0O4AUZs4rfsA9wkzV+Q24EA9wB6q04jzLRQ59zvENDQO4dpZ9IFPC+ckgOVv
B0Wwqm+k7osud6T+dAa32VPZ7JGj9w4yVVnNzGQ8WD1RzOAH0m60MD29PY2JBizyBmFNt7LNUrR9
mCAz78x8rQWJEGgJyxTu0heaHj8xTdolvU5UHrDRhoxLlMTG/Q9wGPxV/CcgYNGI7AJN4jxQZfW9
eCKuj6ngjEBVaY/kIUKQ4QJGKkqAhvx+kY68fahZcnJUA5a2+ObpQ0g8eUOGwsq/pDDrIcDlzDV/
G3c+8y02FZqDHti1m2Cjfn+hpoG5FguIYyCU+4rSxdNVQw6hoiP1NzGfr4ocAuWHFqxrib1lkPIO
hoJ9/jSNqbaCMkqbVmmga6ONRKrtQdsMtSuDH7C3fTUuEh63SV0N0PNIHpv+m3MzsKfd3uOz0lqx
F2V9A7eSmEAwOPp1tLQsBFRjcPJ7WbQNG/RjnJmQXI8BQ7A0yMZ2xHvi6Md996WXcpDFC56Z+gdP
hT4xL/ni0VH0IORDcWJc4WS5jQQusyM8o/XWo0kBc/2Ib2oThCTXNlSSZM6VP2rxVBPUCH3oGbVm
bKn4wMPOzIzj5LipWio7fO+1sRdabAeu/aXo7Sl9cFKwg7Cab5/FwQxCR8acer39LMlZnv5GTtLR
WQpTf3p50qsZWSbPwM8Lq+PWypP8ObKuP69RA31YH/7PIfv6aO8AlGZwCMo7ityJhK0eOS6vOrEE
x1AjCsEl+1mJhpix6uK18Fox4QBns1ovS/81J9FZbWzi8KXo/UYSuloXPysLSp+Il35tqwgh45eM
gql3UT6H49ueAjX6+PJti7v0rrSUlDW8iqlcYLQo3jZRiHmJfqNXtSv4Ax7C6dRrVi3981/QQqcJ
gmQ+nvnIBnosl9yX6RYGNmbucwmL4PVeA84hTnueN7808pA3dkCFnhLkNapxmr7tYbmEDTlZBe1f
3pA6o9cR7w4M/8igCq7rQF7Unn/EBGExOW8o3bz7GBBTKLc5F2ZwH8k6lVvbHche6vNi2dA9Vp5U
1/1OFRqtqMED5Cq6dJ/B+vCHfTtJZ/uZOem9AUL0/R4HWClYUnek6wJvso2cEPX/dNxG8llrlF/n
zyMDAxFDIHn2Vbze8mI7XTH7Mvo9T/BbtIH/zId3zcqT6owKmH0eqgkDu/a590zGFENNKRGHTUB+
36dsL2rspo5Hb2YmBzmjahFB0Lqll3/zh/MYFoaQH/jG16Tfv2HtKdsEvKoD4J6ZTydQ3WJv0MbR
tIQFwqAY5C+mwAT45ghFrxGUdvzhcUP2+ZJlUEGjYOlUiieWXnbHVRPv+vzyp9fCpX9FHgMoLEEv
J2ZSGqZM4XzjaZoaIRl+SQH0g1ZbSsq7D1OL2K5Y8N9hvmQDZnnosYjJayarGvWlZ6Z6WLzVKSC3
jbBMqNzeREvnX/hE1oX3LV0+N3u3dzAz519+cLTVx/qppvS/MdHDkJPlttIFLHE4oCnNUY5VNGeD
f2cvZyTpwnXSzdn7YO0EE+XCC1gTf1q+0az6N1cCNloGhPoRQDomjXGtj9NLj7o2Omc53rKKRRlo
pKWi3h3bI8WxSeUQ8Vf9xGCwwfiv2f9YoyVkLGQJDkHO/NKS3CG7ICzqnJWwccZPnDtlsA+Y5koK
Jg2H6tQR5XHa127w38N3HCJMl7eMuA5YHU8JxZWZtI+QWyt3F6ABhxu4YOo08yVYKRA+/PrZ/ILk
kzrmhR5hdTNkGs2aavWD08CFWM/pY7h3gvcREUABQdu2hUFXglas/Ryd4JxVssPLqC6M6mLU/1B9
zK5/+0Z3EtdF3nCaYGOnfh6rwK5lq8QvOZL86wfnQ3Rkz3ullIsc3/z0I4bX+89ozK3vfdZAjj6q
6MD1rCMV1cShVmTRIASMcS9fheYXPu5DXMxMCtkTYj0JD4of/ffFo0Hmrq4Tx7e+Hk/wFy2oU/LA
qUi4Qrfuqa0G7h/co/z0DEamEbO3TtnqRfjyNGTJj/EhyP7utJsAuTQIoYPquAyiZ6ucTyJY7e7B
6s/toQHnPuMbiukhNMUj670SJ65fiJwaDhiG1s/r0iF8+oPPaExgBvmd1A+Yl0phdGGfiph07gme
gHRphYr3OYE6X4XaH1R0BHFQg8kaQnQ4hXsDjQoDTsxZuCdSLl9dfdton923P53pCHv23vcoHqQi
1LuXLbXNAfixACDukPQEWmqu+M35PjB88N0QvpGuCz3TWcyu26sHDxx67cgWQE/0rSh32k9KNoh8
CcYF4CKKgJCzxpJTB9nkKfX0n/0D0FPBqrZoVnXq05L6USgAMkBWGm1LRVl6ZNt0o6fGIiJwP3jO
3ChZQr6NcEHXGMJaWpLbQhSNSucojmN8AbzIlfDVarijwbMYkaBiifSgbltgTpZ1Wjenmc2RmRBh
Jt5eF/v5Yt+hUoWIITZGt5er8eDjJoI6TyiZl+6aZbM5ssGTWwhtyHr/ooEZCcLJiPN/kvh5pXOu
jDAz9lv4IJ43go57TrVkEaXqvU3KGHGF2vGpHzypRsbprqJ/UhlI9ZpkGwKnL1HbRcHXDszJItZb
Ti38Pdeni9oNj94ihGrrLN8xWagkgSRF2sdzTY6esyLy/J2Z/olhwlf58uqvNdxtwAvB4GDE88Ls
rFK53RjQnQLvGraCJRzs1entOvRoT7bVZCUJKcg43tmdhjDiXvepP9SZ9vnw0ztXzXqrPBMl5SDH
QWXQEZ/QUFwBwRzHPD+4og6bbWDsGvS/QNd0YEDjlBcgn+A1STOm/pP3kld8XLX+vBLozHpNjP9g
eN4xkvDabZysgz70+WlKm7ZslsFjrS8PV7BUaymhnmt2ag8uaM3inEnqeStkQ8O4ucv1RMeH/rgh
pQeaXhz7Upv/00OjTTovEfB389i+a/HAHQ4swYJdnzkrDxjbahSFa4jXftDNqxZG700Y4NKVHvC7
Q9gBBJ26dZuWILbe0AwHw0ZTW7JkqZiRKktZ2qXLSneaytqsC/egtLo1UB6ms8rHxx/YVZjHRXM+
99BWPSfo+f4U/hBlHSslAtNo/zfJJLzQwMIAulaADTJn3JMo3vsLJyXPAh+wXIBrrG7OD780EJhU
OKGiw2zo/kgxMQmPGLyq+vqIcGA3XSx3B43VDV0VMWwySJYOahYmZ96jWw6bNdfcAIVnhPlYiOVI
7HINZzq95SNgRdfrvPBFk03nbCn8w/O947FzRldCm3ZU9QAU3rWLHHXhhsgF67/rQMQZ28NZcm78
1IjBGLeDOx7wf+hHWKtkxYBwrS38zyPgX2GUyyH1omX9Gk6Kmv2EHMr4CIhOiNSKV5P8K6uJdH1X
w43Ik8oCfultAoU0ksln52gxkruAUtdsQtFJFobGuct4WgbXC47xjPHxto8NYs4I83P5hEjIqg0/
USVK8xyEBrBLox5yUMJNuEsctCpnJdfK3WqI5w1DoMIjFkagDd49TYdlsermHIqgDARGW5kA+6LT
pX0i0JxN4t+wR36MZZi73xX1lpewhYwu+fPsVA6x9RxN1rM6m5oBySTp+rL96u8x1Fc4fQ/BRtEL
clCoAIJNvrap5JJ4pJkIs1LqG4yWE2TYCDEZlE+mD06lQI9neJlccSFpqmSAQCqimXj3+j1iHq+X
rWylx1e+ZQf3/6n4XGxZEv9oj8SdvTmWSpmW8fob4p82cvYS90Pnev/MyW6dTNSE2lWNjp9wzl5u
1pyKrQh1mnL4JhOzaCInI3V3OcxTjiqbXv4JGthgZMQe07vLP2MJBfbFfjlpZldSj3f6oc8qoj8D
3K6UzVL9Jdc2TBZZUvKRpkzyL0kqa5P/FIfpb2iBCmtOZaVrVakhcFq3EeaJx/xy/i7/Rbi5YXu3
jOgQ47CiHyjfyoN4dmLOfvXlrjnS3wt/ADayLKJF6YCP2M1LzfJ2yRCEqH4Xqkj0n9SOketNdnk6
vvnToO+yMUKAnbohjmTS67SX7vofy/++24RfyugMTmw7j4bAeAW63vtRow4i2jxXlNoTBz3T9CPx
w6CXRIyey3JqdB6c4UH1xMEfL+4dOAe4j2RvfsHRQe+gIEdq1WLAow4prJuOEu5cjwzhxrjpSVWD
ZR28DKRBWAy2WCZygS5vI+FJGfvTekReWama3+noMK+sfRWKWKCzSH1jcy+sXsVz4pIIixTnjbHE
+od+y1fGR0rt25u+NaDgoNKxnorzYHmHWXXQdho0hPdQknPQvf44jznLB2tcAO5csmFNYW/dSQQA
0tAgXMKs4Y/16dElkiXeDvV9t92owUCx/tY9xY8GqG2c7ROdCKfTyOftVRTaeKRCW7s3q+E/ltES
qeLjiznjFsFLmmgLiwuZiWf7hJqOEmaTRjbsdIcCPZxP0aaDlXYWOzFb0lYLBCO6qgcaPTP93uWF
ZDGqrVjYAUgcYRn+K94hWtYTt1Nom4eWiahvKH0zYm73pDYOr0egYiP5+q7eGYeGjiJCYVebSBbI
rhEhaNKAukB5dqgGZyNYcU+6p2pv/7Q9LjOsyaT9AUxVF2upfLgR/pvgVHMlViFqqe2HQpQGXnEb
A5I+oa9U7n1QLQr1+EsTRB5bic2ReoGRiAaFrmcaBczu6262aomJ6vbAWozzyR9cwZ/Vrk+lzJDC
besimTbTZcdHVocn5Cq8FUQp0iBCOMFrkA2RtYT8TTvB/gBTv5rom84GUlWkuPLbEPEjmVk6swvD
mIK/xrhKHxsq1WsRbsm8NFfjsYBnCBMaN/2blseJgmVAHJKXguHuIbg1jCvgCQlwHtbSTpSD7LyV
12WUBtH0POeZJBq4qSvbg7+n4o1Hwtm57SQNOlTAF9q87bMKNFkz/m6suVK2c44u3eOYM9EVGXbQ
CJ+4WEVfEVllwIoH0X4wKraQkM+N08FQDYEwOToQTx8CTBAuBlNSQF+ap3+kwlxyY6l54LolmN6i
uMQVjqB8brrTpZFP8U8aQpJb8zBaYv15YaLnwW5smrzuQex/FgVmeTUFJr5fm+fq0qjcV+KMbJyj
KdWTr8LcvOKP4nrOHWHrs3+p0H3SchrqcIftDXiPoGavSUqrDFfhjcYlVPHXSSpCkJB6a7oXewVT
7rPPc2sHxYy6Iwe1dQG95zf8g1CKlYUqHlxXDrFC1qadqt+oKOwpAIYYuyXJ9Bb6V4/dDfj95VqT
ZkJsqyBuap/tvcdkKDVVv2AstWU82SInrhZPjezsXr51EV9IjuzQZKLSz2oGgsR8eudVQf1yuIsR
er98z+MwXk7nIgzfnuVQvitr9MCL9bRnsR0bqfAW/Ql14wSdPGFMA9mZmF5zG70ZV5FK5J5FUc4s
BkFIE86XYvFivx/dJpZBOw/NoTM/2M6wmEJKjhBlXj+fFVnqPDD9uVA1TmQ4/Nu0uhuIzs/NedXV
fkqTICVtyIi9HJvx48z3ZWNLOOtSdboYSJfDIdASfeGPDjk+f0/kPjxD+wuf7nACf65AOpe6PgVS
cM3lKaDqwngiRKKSLyOwgD+d2hQgXoZMJg5Yw8kT4hpzI7N+k5lPzMq5pH029IgDWNL6+6iYceLm
8Pcfugln84hrGjVEnV+lzVzmQUuYVUFEGqp51yCAdIl06425+K2mNs2SXfUjaPxa4ZvCm5znh/pK
14yY/AW9UDaPIqUBkWWj0H6i8nlUWVO8dn9LN1uePQ6SfL+vhaxqRfShs2cQ1lIBSJzDn4DPRvdH
o2edQ3ylu8cwnt/asnYakA9pdkNBJtBDNiptRqjQC1u1xXpPf56V11LjXws/MfLN+zhp+TgJKYmI
Si+BuhVm+bv27D/CFSndpFpeEbGEzEk9VP5qDXH5i9OkrjP0JP9lUmg0EbAR27S5wBKdoK4M1R2V
yHAzYOZnCwQhHGkNoca7mZfSyxfg2vUey2xwYfdn2NpJiVhT+a+fLGU0ILGmH5d+XGLHZcpTuhVk
g8qXeq5MJI54vDDvrYkNHsMeF2uiAD3G2rQaObyE2a628jne/lfpDCitJJc+UvrQUsV6PFdF07Hs
T+dv8Wwh02nbma/Xm6WuGhhyENlf2xwak9Uqv9eRVfvEqoZAcEnyMPquoyvXU2NOPf4imr4uh/vA
sd+wkzzbsa1vbX2BHlwlMy8LoBT+rJ2pIdKONGve0jSE1FNJ3Gup2lI3Wlm5vxlg+0CvwSdvwJ1b
NwAHyR+E2JUsPc+OnHJfoo69jLYm4CnXGvwIxJqhulIE5L7iIqUJRKvnkiaTWzl9FINnHKdfWUBJ
XuPeyhC0+qlNsCRC56QssHT7VPcb8damDlxPCcdsRSN25hJcN5aHWhm3cEht0nInoKJmICf07QfA
uaUS0CWwZXLblMPvxMtTClGq642s2lM0l+o/wV6fmFOJ1DAm9WLirkk5d0VK7FlSYhtaIhVnFDeE
uzkBbl+5rgL5D4m8TZl/ye5eQeXIMh98X++OVds5dsllsZ5JzM1T6+DhOiQgi2uwdzBdk3HpzIKn
uKbtjM1HR5rUDo9pf+7o/XhLre9S5Y2qg8W1/kFr0D4A5pKRQ/ZVS+Fil/cS5wShaOKFPCkPrFuJ
RmUsslOjeno7ARHnjA0qDZM7EOSP6Q07Sf+YM2arQKK6UdkOAcy2Xk46gkKmSg2cz54MlEIrHozJ
GG64KqgtUw1CZAVfR47avSwnizr3ETYA+QLji5v0zGxYzyY2rov9OIMXGXcvnnKLIJlpYZXp2+/r
YbM0WA/eAG8EjTohVLXVQfOsoNIS7hsVCo3U0evZUSiEpVz8q/I9n9NnmFm3rt91rdCUwK+1U0fg
dOtNECQDx1N6CtnEdqCHyCwIRLQN68hqSZQRHQzkAroB+2fcRwVS5nu28DPcMzLhQgQ4uAMWwTuV
sUCw1qme0YObeLIJAFyo+WCGmkQF+G3jozCpt0QvwC9XT38eqT1/OiZqw7t7O5aGbFNl32ocdQ3y
m7m/qX4Yr4705aL+NXniD+0ViLbEVMcxd0yCuF2snv3G8Nes9y6WZcwC38mU1+OIbbkgiiQgGamt
n7QDW0rkoovS3CSpFRZ1vNeDVR8G9N3lV6XNGU25REm9gY3nbt+1DofVNmMuiIO1HDhhHro0Yxdw
Jwvwt3kzY0jnwJ39f4p2bmZSxnmquePisGyl/cD2phYZY0vG05SY1a0Q08K6VWfbuXeSJjKLVPvC
eEJpMJFjyJm3EcYabG6LpCfkx72AOVtFHetR91IULKenJV/G+vBFwVE/ZjnTy274FoMlZiOYwbyN
WP9MjRuMTtE/N9ndyqU4MH0sj5uIJ9wmps2BwXFjsOIF6FJ9M06zNNFxq+ynT5TKn4CQQ4KPq7k1
mqqnVt1kyG2gCCDX2zselrslggQUZaw8gc8/JK66fjrAiVufQDv+pniUaaGyMAQuN6vmPZLteWFQ
Z7SGfwOX/rz62VzW+E7J4YYKVIPh4BLS8JNECmdWpVsNllgP2N3ZwRziAE6KMvHY9VVR27RmXuuq
UGUI/z22B3rRDrfV2hrpBdgDNPIfHQH/4MiK82K6t4dvesvN+j9EaabP+Ek4OtHT6256fvTlXfjS
Y2tai1odQwxmIzAyIoAC9XGv+J5+hFZ03jZzFXViCMVp68hkdUsBW+GX4OlchIjndM3SI/SCj3Zx
i2Eutn1K9Lcj05JTa+wIPszGLKw90fk6GFhpha4SY1XAcUy+fWXQ69XaG4RVKrwFJpv3M1uVgf2G
/QiQO1Lr4o1oLADaaLXxoiktOTppY3WicfD62W5yEs8yB5bvmzG2FuWylhEAcHvnHc9xK3cW8Q4G
mBlPaRKIkC1KqZ4CcoRuuc/WUtV3uqn5ec7UT4tBO4HV9R3qR+YVjH9wQ99WgdqG23ni6n1XsZSm
qVN2vMdsDpG99IoVJVSp3arprs6H9ts9xnziJEKgOlYlC/yts5j6oAIWEx0Nx34kNa33ViyM/d75
D3gM6oq5Ax0zUl/xItKT2Rg+tXDzwURZ7FlOSeQYOE4LnIcd3ZJ393Vah5SrsHO6odYXNXCihb8S
hk/xV3D7dL44nfPO+tekDHUBSxrQSCK0s7+UtuQ/wgO3L8n0+2CmtqQSEKGNfCQYDKFDjY9EYPQ0
sKW0ujNjqzdkUWfkoBxsOnw9EWKkBncOW4Zu5oTE6zQJEAVOar3/wIceVPJ5ys2a59FZLrWegNzw
5ObMDU3kiqjCJ6iktAvY/4b6gUW17ku8jOqHSMXRatUvEsazUltvmCOXEJH4/wSPHgaoeR/XWa0Y
k3pOwwKuDPRH+trkkdRo3f8QQAePftwBQ+S/ky09foaPy4LVyxcEwbGiZ6O8PZNiVimnROSZDuGW
vmu+BaSMiXX7favPJzH9aesbXt4auMEQ1CBcxSPkoMKQTkv4X9J5EWp06nmzPnLztKRco9ZHrEVd
n1sug2v5fmzUjxZc7bzHUFfHSMnaixmaNHvmmtyX72YqltT124yNz32Fmfg+aBwgSWswFPhRPdVF
vLXzMTMlx4NpM7hVOgetD98FHqelmIocaH5DoyidD7Dwnoa0H6F6s5z9XGndasTX5auN0yShnZTu
K/QeAlEORVokKA8VtvKeBQXYhetakdKR+WMUhfRL0whdcUcGMIJGE0e4r7VI659eLmgttHKHh8Vm
ZwYDx3ozHdZAwjcZq+LpLAbmzmHPLcIoHEbvIjJeLra7RWvQeISaZyENYKO7BG7bWc3icARXhe4f
aSxvC5CdM4YHlWTrxRHliBG/sLI8So5lBqQ9YmiN7rZO1Ny/TIJSPvTF65jHx5cWoX4i6mWKUgSf
Kh9zOb188g2JQE7kLLpoDF/D/LYOb3hhHMZJsz7atewmCsmJCkk5d3Ebm5cvjYTVHsdZ6Jg11Bb1
CDmu8jao55ojT0RWNdJfIgH9gtZsSiIzWW5D2Esk/3GSuXAtBReBkxn6s8gJZ3KvAlR1LENNmqLC
i6Eh7dBe7zpNFVJ+0dltfPDN5tjv+MtJ9AJKOi34lsvMIogQzcLYGqgvS2rkOx5SIKAQfwLnJUdS
X+gC0uibrl6VIHUoY0tw3R63ug5ddgHsX02Rt/d2nLk6RESg1pE/RkC6qr1lgXOWGR8eS/j9hltP
w6VYAAaY/GCDDEOoqoQeRLjULjgPn3OIIMWEz4V6P1yBSnYAKgH4gOPHQikEjEm3SFIPL542GdGg
5Lu4DgFn1Smh9Yx0ROk6fRgMsMAElFJFciuF3rPsKMP3cR80sfpZPHc7dnXI/NkcqWoPFtgnq7/y
NOQTHJJPRhpU6yf5/WTd5bQ0Xx79dmEpVdBQ9nMSdgFVZPhJgT6HoM6hlaCLMn9kLDCVKIAm7Jw8
H4arA9noJrrgknjlRlXY9Xs3cE2j3XeQiTQKsCgqdNu7x/aqzdrNS4yQvpUau6Os+Onk7K9vpl9D
PV5nPsOB4dToni7wNQMODQaUzvbruysGCVwTh4jnzRZ0TkVFjs9c6wePSAk47T7g0y2b1lIcTMo5
WYV23FnRv8fEvv2WaBYnBQyChrqWi3IqkQHfJPT8LLMnlHBu3wmAbtLyrS/z4Gw5z331L4BHdwcV
6LA1CbEKhYnDuVXJDM7oBqCJnLsMmYBE47QwLOLuv7PRpMsw2jPPi1x12Jr7fJsGC5Jr0GCR/60c
XUN9TUINEDm4QoMmegkVUBGriEdRA6pG3I+Q8NDxu11/2/d9uJLeKEtD/8q8tLWHUIky1D488i+S
8FbrxXyFnT1cQGfbFUI5C2s+xZVt01QIy7Qmw8+0Vr4DeC1hSrU3L2hD/InrQzpeV8XRwFFvyV7S
ChTpy0eWnQttnUBZzKTV3xZqcdQ5XdHHRGokhrSKumYZlTdrkZmemyHiPD5WlEoKidmRg7YpFO4Z
WqBgcgcasKDpEUitaaNiSoHVzGVMiH4QaUga9cWq458bKYsJlQ1PO68tFE7O+Lpc921tphal8ZdR
caojEAIKRJehUPQNSYOKyiDOMMQFzGFhTnkDzKxT8ETwrXlhiL2H44D+00domRtg7xkXAS6QVKaN
YMPWD4nBehFMgD7gukUX1coUg5ajey1+SVYGqzdOU+uwt3JZB7MI1B2KKZ9FnHADMn75Ixr6vt+n
Sl9v0KlzKU6ymQqaB8ni8vwkrLryXbcChyKlb6xV4XGPlE6adAJtALgHxr2q5IODbrLTOJ5ZjkK+
2ymg2JxBBtlnSZC+67me/5H3R8w7rV2glAKpbIjBKkb1GSeNrQq45eutX0bDeBGPcbD2A8pjASZt
PZXFuW7sm7PkWIY/ue4BLLJia6O5LagVLp5GALAfJrz8DBZGzSIbu7qhgvpmQmm61KW39r0oivZl
8QQwVpWYLXVIp8j5LHdCBIy26ZYRQM1COj+uae6EquYRXfHlvzWh72Ut5wrndIykNEnQ9vDIMkF5
FsxorUve//+RpiJUl4rwLOap1m9pHw5DirKwCFkJU7MYy91/V3v37z8mUHTxFR1M+inyJ1INThs7
0KrOTbX0cgmd6iTYfddT63oUIYgwWGektManD20tunhFAyMG/C4omZNBuXY3q4kpXBu5GZGwFXeh
PMV4ATFKL+inEafMVWLuzPUtC3/MhhROuBSAz+4bzFrSL/Xmw91oNmQJEDJAm5LjMABvdleFmSqc
xUz8+mfNM6PoZktqTDOruQ8745bDSJDRq7Jp3fHcPzAZDhRNK43tSFwEsFDKy/FrT4oyYVdlElRU
yxG9gGCY8EXGy83kipnQ7lFDjn/dBF1+PoowB4Eazh+VhbuNdvAeCRnNY4YX2B9YhXB/OIRvN5tx
2s9RqRRloKoYSL0Fdk900td8bkp+tLiRByW0afeR1tUoWxEeUsik8aLKTSz/bslsPfJoBskv3MiN
GlZiRoFRfZbNCRhfncpNr5KG1vIuDbOFG7Ocz9edUMkRJQbhlcBniNMSg+EoGsnZDOZcGpsb20uy
+5gj4kEb9Mt0wjAF++xqrgauvgC+YArDRL7IbnG1bgUvQB79Uu9BtbDkSnQPwxJ/Al3fAozrxogA
DzNe1OADu6U/90RX6293CQuiTkJbSF8KgfKPwLDlhH2EXaLsFpk0OlSyU85mZmDzv20hjpe5r+Y3
S0MOtl6d192bu4+bVb3X64Nl81/uCJzMe2pPkeTAUP2l0JkrgTz70jxy4hJyGXTBrL7xDZVP84KC
/UVbB4AI4rlwmq9ghAD5IzxTOqMKnE9XVe/5ygxix98BI/y8NtVTH43lFL8QpEpe2gLlm9j/CpI1
Ti2F8zqBZfBebfZByE74TNYRjI+WlznRXG/fvDTGchY6IaCKUYINN7fVle8hK4er1b1I1hLUvURp
oXTwQ+NTwkja5l63cnIFAZDbw3QwbSOwEYM6dm0Qugswp+1OihvYfeabvd6SXA6whs8gj/7oPL7J
kgdmSw4SfAJKkjE61OmBvV262//qfWYUQ78RQFHfcGPNy+wlneH9DCHKkZp1FyuMawd90a3DgCm1
qqL3uc/bV69wc/a7PelduFjseb5ao1Q3sI4fxWTb2BHJ27VZtRvWznzR567L/vyZPRHvWnzZPGaF
xeveMjNzYC6lBRr2FRiCaHrQxdZHUkg2ajp7bIYTx06iq8wQBSepu4X6nzeHrMbN9Gfovt68MrN0
+QYOCRoQJv9EMfZB41ASd9GaTRxhS5WPKamM36NY7JJZUMQ5wMMBs6f6MFuQgn15IqmwHMBvr2Bo
f/MkxozKFfRpY78b0VCxb97ssCO6Vt/XL+Tg4p/hAZgXJB4Z2a5FjpAIb2xpg+Lf/YLwqRXALeTu
Kqo37/oR95Zt8nMrhHkg5/1WHfGjqLGTZ+FkmSg4QsQL5/05MBxT6rz3xX26UYuoXETcaexvVIGI
uGk/JEilcsA8eOO6Xfj5zcMnt1XdUgWmXFuE1Wb7D79bngKTH4+cI92YaUANQKpmnVFM/r/6B5xK
Nw4tzZtDlH2Hkepxt5B0w4FCZA5NANXiv0qZ1ROw4Q/1UbC50pxohQh2rmK0fUZXr8n8bbVKEcmP
dSZ62rJak34iU2qCOm+CjkX9Uk+kGkdF7TC44HuunZKAeDfOkONEOryyU6ChR89JmXACQwtIWiTA
rMR4YJQAeWkpa0UvyEbekMwm9vZPpRg5dBEZT12JXFxastKmMoZyH/xRpcV0sz4vgovxBbbx45Wk
2tT0Uljeisbr7Q5/uIHOUM/hqiNA5QWAauitOv6PrpjSbJLu2zrMFhbCT7nSsj1H/Wm+IRJQkdkX
Fdx9U1VSd14qU55vkXSsjjJfg5r0uXkLiU8STnSkz/z25b2zkM24y3SaobU8tQ27SMLhC2YdbTxn
3lxqWuaY9K6WoDoui+vZyDz9rvWoBZANwK9MpAc1qvXTP11+NMTUkaafuvY4zWdLVM7mSnWoMvhm
MT/FGJf6Xfxevk56qr3qP1eDekpT8zhgSIYTE4YT48cmSxPuNVkbuhbXVl1sqCxMxdHg2qgF+cTI
4gO2B+S80nZ+HW0pmKNlNZpLctuFFmlI335Q4cOj64FE2eaoDBMUg95oEMPSCPtc4XOtQPrvLTAX
45oOkYF8S6+xCuow6nZuAcQ17syB5hNWLvUIb04NM4ZpOplJmo10GUmM/JP7kKCjLOCSwWWeewID
PGO/oHFYQgymWeAgECVT6aKyFGUEy9Q0/gK32x/A73AdLblOSqvq4n+e7GDN/u5mwyO2hZ+QpnVu
LkUfsM+5+qw5s6z3kVhR4Bc5c0TpgVtFNPhNjnSQqkACOT7hrMZtxGON/GQ8AqQBENMBcz3cLRsV
fJXfVUHqG1RV09KZhe+d2EIlnQSUG2GN7UzZa+/5fxV0DsBXV3tkmNIKV8aIhRgBikxpVdlhaZ5t
FGdjL7lvZGFmeKOYp6hcwEihL52N0L30Rc1WcmDLoYyIg1pcv0lZfY2Sbb/0YfTcJq4G0v92NxI+
EZK5d2LfzRuxTZc4EaxGrVSwITgi25YhzMwbbNSn218U41TlO+zhrEWdktdREOOteJu0CCL+nb6h
aRbcW50kL+ZWSExKRVS4UsuvmZbmIsgmba8w6se/s+Qm7A62VKFY3hfEOvWyaWzRsFqNaNUF1Ek5
3BNUYuv0Eho6zO4WyK8bW4MVkdkz95DP2f726RoiHDKYg/Y05FVPnS0xZTe4lXplECVMkiIK7USz
pUR+hrSICOv6U5TH9PYxKYPojIVABJPPBItDU2t3HHyCEXuhjvvs9sPr3SbJOladvoyT3o2ndUQu
NSxq3kU5UBPBuXjuE1xJ9AYJW9AyU04teHM6hY/748E+rwvC51Uv8xT59C4Syu7hXpdF4cDKGXTa
9hK/YhL8+yuZKgvdn5HpLOLOc0kNrcJUXLMQsMqfNpp5hHJbn0FNmXIqYqvUqF57GeSKCFbuLGxl
PbXJK17ceK8sOgRC6VcyC9Sa29W92nGuujjhvC1+S/t0dclGw9hP1H9xFMpJtY/xPjUtL1HgPH9S
/BwcTOv9ZETj7HECdyvT5tDKGfJ54XUbS2c3mQ2IVHBBpxQ61dgx6MMIjgiK1v6uWr49I8Jf/AdT
u9eCSAsb6+ceitM73h/23dU2mw21HVqLVwTujKAKH37rZdGm3EKXR6gOdAYOsL5L4BVC/cYQ2fwf
mfowZ96ZrEnP/HYdfOSW0/rLDJtDRfpwQnMWclMT78/DF39A7DM9BRclxYdVAlA5bvr8w72/bpTT
0yPWshiS+Srs301/yZGECYFLUhPVoHLtaa4JgqvmbKMx15xquIOei5t5plXnjpCeHEgM0vbxWZGt
YpJ6tbH7NSVTZ6sjTpPaygrvLkzWHpNgRy0Wdq8dsB3wIw8yakVJbOO1kbD9PQzOnK7wj5tsm5YQ
ssFysN8JxYEYFOD98JvftxpyR3TnoiDhQ4xLV/yG1KViUBrynNbQHhIY50rWoeUPr4j0+ScUSHnY
7SlVK0wKbYiumwGj5UDZ/vgIpy2c19I3QDPSHhPrpxnpUTSYpqEA8/yVBruN6X97y0gqj7ufMBcQ
PtrmydHAD3Y60cPblMeVXz7u2hq/u1mCECQcXPwKPH7AA3pIs5UGzreVZyCtL00u6K38fEAWQrmp
hn4KT0VkCDl0pPYpj6KOE4p7oM0o3AhFtnAUz2EddFI6T32XTJ/6cSWe7o5tAM76AOjuuhWT7HZd
Ew91YaWt/xnIewtuND2uRRq5w5EdlebV78ESAmSXCEfk/QLc7rX/z4e2zpHeI4NnuNbdjZdtBsfA
wZysHbFRMsdVl6HgMNnvfnTj9MvyTSLxgsNzu6VT4XcnpuqpxHnttPCLU01AlyGAGlsqpMMLtWsW
ifCxZqAICISxHHs6N3ZfcgU4n1sn/yfhk5lnr7BaFfy2W7WT2Gj18ElMshlO2fIpJaGBm1OA6Fdj
ClWWeP6aGVrebVWrnv7LKNzN4z2ZbrTl7dSITE0bbob0kIC9W+OO2sgbQ+P+21rtRhpqkXDiAVwp
KyAsWGSOdPkv9ferWuRZ1nj2ZHM7sDsPXsf73cLqJPCWlZru2ZKjvXvi1CltQwqgPc0ZuiwLEwB6
3NsoWhHSwBXV1fqd7Cv1e/ZBd4KQJq3YgM9tm4DVzhlWHoC9RVeXfLs61AQYsUFOUL0J8Uqw+m/h
Lh1NUnOoI/zZzCc8ohfoWcYyr0x3Nk4r+/b301BYRdvGGQQBxP+Y6oPAlXh2ddxiZ8PxVgpB/BXY
E7yxcWmz/B4YUmyNvOMq2jNVuhaluQZNN+y3eBDile+0yVQNRbS7gd6tKmbTyOl08aDxls0mx+eq
y/uMm+UabPOw8kJk2n8EzjOPsztED2UHtqQCUcx94iAoOkM9WlRrdTcsEaS5m8hXifu42N0viJDM
4x0h66t1m+NwjQ/yk219qJLA9RNcuGoy74l82VoJBFlNH5cof/bNsxZzK0jXM6ayAEECBo94I4V3
hdQUgahuK1aAasORm1oer0pn75pYCNYvIR2JkpxTOhujn62YXfHDW+CpfIybEbGzdcpR1TlK0Gug
QiWdHEftZa/TEKhIUiL3S0CyTgfzr6ZERGMDdR+KnYI22BZbIeKJGtaTIG+CAkAzi2A0aqMn+zN4
3XHYIU+6AY/BN45gbN9OqyHzxHFWMgNGCCykKyNbgju5Cbq7vFSm5+XrZca+uF03HRxO7HL+y6Xh
4McJqAcmU/RGVDrq6rs5UQSO8mm2Vq3qqR9mFSsvcY8uhajAlfXfCQEJSIZTKF2VDjyYhhOcKzHf
T7twtkVkecLqCVC5Hvh4PX/+6T+vnwFEdnFNrYtLvexYiqfo1+5g68+nAgPoBeLfVaIUEBU6NmiK
1j+kBaIgqw0+RC3fdoV1OYLkwbpr9WwDv+Xo9Scgf+k9xrgqSNFG//f8KaW3CJokVZG+qA5Rt+Z3
02ihcJUeW1Nv+cGsaikpaXTNWjAtM4nFcAAo6pmX+8fqJ59Eev9Ohc213DvqIsD07wHGkSN9u37a
pZcGEZIPXid09pYCJEHZeI3sg4O42KR58gA6nApikqXqgrzE0ie4ymbanWzPGyLNcUbrjE5BodLv
LtyQJxYXJ5RKqxmlBpEmdoUB6YNqhuMJfiLH/ZpyeR1fk05sFXAxI9pgW62BV7iXOHSRcYhkwJ0y
MvMFNe9Zy3RO3fJoZR+V/NEjNvRAeOspLcbh4Mq28mdy267XazcBvl+6f69c1aghCp8ooZjsbkHe
S/z8eHtIWcGyH5GjV0TmiYriK4DsvlKJiYSNdX9Fzt3I1oifSoT6mwDjw9ruHogHmAdz+pMFTsXV
x45RWjL3KFWuvAPPu3quZAt8IhbhYFIg8zt4C1de1g35cGO0bZ4hketMhWVoqmk8JWJYLJEUuf8z
MmVPoc/R7f7G9h5AmDLXfu4KNsgXbWDGDMlm6Gdw7/n5bO3Y0MLRMXv+l9hemnaHiU2Ectk2S8ku
F1CvG0tij7R0ZXLpAlapR+5P+BTqvYOygRnVNv1IwHY/GDPDa+jnGT3I4OyngYquQVYbXKxjeokX
DSo93Paz+L6/r0eQHMljiAPVIheGdZbB3gNXLpIKtADI7hpA+TpxWlhIx8ICd7s3KcDgpmBHklH7
z4a1ldcqQv23rgxgUhpgmIUn077W6FKEvoIf7twJJJlUOD94Vfb+AqY1BdJmWZuNA1t/IAoqB18q
oN5XQrl5/bRroDUT2iJL72BUcwMU4Cffi0Ls5BKumxbuPd5k7SPOrqQ3iCYu7XBwJ/cAZxGbtf9k
hQrTzqPhj4rv2QLgXus0ytZHMil2hCE1zDqlZ2cN2Ld6CNbGK9VGu4EfCCf0leLxMxBZAiDwW04h
U+Dx7HQojcLpoZQGxO0DF2ya5E9r/+Vtdk0PB9fC4PmEM3SbMiEjCnIafCetIn5NA/Nd1ZCsVzH3
6wZkCOY0j4jqUVlfzZ29/cQFg4dq9ZGv2R54nl7HJKE41Ca84R3MRb55E5oMWwX2oXdG9Hf7RdlG
cHH9B1Y/LNclbgJG/DZ8llftH1BKGSKVpiNU/QyjCtKdR8lGRel8p1RHamN9DY/lI5rVKMOcqQqY
b9/kUeWddGqf0bXKjiaKIO1+NAUBm/N/QpR7CJ09toJrtvepy45peCIiEI1BclZmHAFNkbocd45p
9PgUZEgZQooQa9YPOnK2w6aRuclKQeWWkpAgCxZv1EJ1XzaESenyB3y1OndJd0sJQCJB3+SgqE/s
wOA4McKRzD0ES0VfwRLLPcljtcXPFKJ24Ebxmwkz3nVB5wSyTmwRfH1Qz0Qco80W2uIz/k+QjZdO
2zIP/wahgL5zvU9PS7L8umvQyMKQXM98rONeioQUgScWxUFNfOckJuKLrbENwqh5gvKZrwqOs3XK
1Ge/2NbjJ6RDnScGS8NhX8YrGk9hxvvoHza7iRr70kW5v8mQKNO1VPtbVUZfRk3894OouEgOzAbu
TnS0r4Gqjf8EGZg8oBhg/Qie+2QcS1Ib9jNi04HXEwU8aVjgO15TiF4cy0EnKFlgh7SIsgT5srwk
KxTgL/FuJvKRqF5W0yFWfIzupFkCZlQSOnShe9M8w8S+9BiKlbkg5gSD+y2zGrnJKE71xCCdMhN2
RlH9pAtF7aGudRIGL63yv2SIF4eHR+KryPbWd/5zQDB1nkNzYrRp4PbNrlu7Il7r3XgpixnN92ea
p4A1aDZIXreSyB4S7bfnZZ8wvz8F3uwiHOdy1uiWYi11LJgpLh9+A6x3AlUPOTnr68qmwp5r56J2
Xl5+Jm6GXsr3pTotfPDMoLMDoVHjXtOJ+MvbidCTa28BENpmk+XSVmS8xKUjOnStELEX9Y4mW/AT
9zf7wHx31hQU4czmCBf5ncCZUUA0+l+1zhlxj1PSt0L3cYghrHAy1Np4WdAq64XJJNIZeaO9XjmS
D5sJYsz1oFIPVcWyK6JQVV/oL2QnXmIZo0cpjoFiXbQzdwJ9//r+PwU6TCpfp/k/Kxwvyj9rOOeN
n+Z/ik9pudTjBUZrH7epjaU2qj28H+BPhZ3yv/kDsOzou5EdYFPStlQfZzJ2nct6a11gMzWz0TVF
keGAP28cuR1mKajVMlOYTH4e9BGisBn+wKD+Qn7fAlbgoQ4Up95z3yQAV7ZGywJ7PdmHV1P6LR/k
Zospw8r6MgAYZ1IZC8PMYfnXID4s2V7ovOAoGYQ/E3aWUYh14lxuiSQr6ESUdhrFqQI7OXuB3mJU
Z70xTVmOgG5roa8HzxJr/uPUJfIqezTsUx0kzTa9HKavrmc+nnuPVWJGzIDLxTUTkqt1c4T59B/A
FXONO00BVJC3PAA4OImu21zDUAiOp5TmkP1d/voixEysvh0s3N4PiQAxPcZK67S+H0qH+pQZbnUj
gU1zT9OqQL1jlg9P0a7765GRm3TS6tbkPJMHDaBlyj9avZNeLXa3O08e3mqN8a8K2K/ZPUxWfEdj
GKbyrVLr4bKbP6e+sZSeg28hHj/1VpRhy87ojcdqWNDT3sqpMyN/pOO/0v77U5oFwMcxLXFScaS3
x+HixesCaqg5hV4H2mZm0GusaEkLIOjsvAKMTf/onD3YwJZddY6qliZooA3RjLxUtefRQLxZpjHA
UPBfDBpHPXEGLTQArOcmlQlF+yWbs2HX9LARli9Oeur9ucFNeVoyEchRRsh0CKgqp757y6cJEbFf
RN8teVdQHzZbp4QgSAyuAyUueulVjL/NWuVddDCtnqc+liehSf/uVQqUPSu4toR6lG5CG+YlhXtV
P/Oi3KGk8qvkWhsNEFeQCis272WWWtSdrPg1DwGorNBMx2HYD+eVpilY9NTCg4aCia91w0Cz9bnp
NddA5bNb3MCP056xkhoLnf2h5FLjPPJDyPrgZNx1WfKygnrOVzi/5xYDPEyQt5Mg17eqvVnAR5mA
Hl/sxMz1CsOa32IJ6pLhIlvvpIR5m/jMcm1KQLjE6S+S2C7A9brszzHrvimqWevxjZ1mssfxuhK/
t3kDTN1H6skf1+8mMiHqXmYYqba7YVQTnKJdPdvEA9RNyqGWUZD6Om9c/rMKLQT1hr15tCfnQM10
qqcUQh54S6Nf+aLXY5HXi4TcCqBPb8zsIwX7YSy4iJj46vEottZWNWvFN+Oj4naPEGGYDqA/6uEg
8Ln1PyJKVJE7P29NY5FlPPuq3D2K7X00H0N4N9Z9nSc3KUkEDjvBDo3h4H19dXbtOPPp1uHvDIKK
VdNJ8OwJzmgv7zgJ6v+2bESSf+LgZQnkII75XcoxltiIdQtTfdrY6zWwQ3pumhteI64mZm5b9E9F
49kXcIWhrwc4UOcUwNQ+3XGOHvnyZ42r5EZ5iw59lJ8SAgmgdY+JH4smLdeiGL5UehHPcFu3inSY
sokZWf9USRngQh4hUvSoDfY6ru1Ok2hLQG+bPq5HCiDCAR8rcVQNQ/DTey95jkk6z6yF2H0pFXAO
7yAq1tFCtl39tIKOGpC/3NcrEorTZMSH4w8vM2vgSwDD8l8bac0FH80doWFMxwfyA2dzCOYqe4HP
FI0HjiBxQhfVtesZXG/6oIVnP8UDDxLFbS1HmvG1qO+goQrVk0hS+cPIPs1duW9Kyk4w1Dgh7Xpv
KhK7EI8TyMFsfMhq2sR6vshLE2YuSn3m3T2cBpJKo8bNYHsVJCqloZDAKDxK+vHj4rtVbFnb9X0m
k20mooole8ppBdzmp+/UlEr07PLI0J7RTLS361Wuy+OfW8320F0sfeMYElmK0bXM4CFwJmLVwu3y
O9KtSS1Nzr9GCW7VkFS+qI2HOAqpcbbpWNhfOeiTn9NiNoqf1cp/6VE9QppscB23ww2OOVZGw8ft
y2MxDPTwQiO2PBGq+FZXIg2iG5+Z0md7bYfksvh5Yf49DUsxsYYPaG7sl9GCAAoRA9yOJpdvGKEz
P1LdhuYGsTHXfZ+urGhira9rJFidxWPYNIl8BsMQcbxjDIZtsHUXFR7TGIiosoXaQGPYl2Yk+uZu
PxO8b5vXsznbZAEaldO4MyXIEbxyyn/wx5sXN6uhbLmTF1FTkpSSyjYFk92lrcQnfRjqXsMARZ9Q
cdzUVPZsplIz5FMHYELBP6A46hRMXWy6QQ3yPnrHq+gqvjgedttHEY5H8e7PazHal0/2FmzFhh5M
Sca90j6WbPPIYyqnwVciqUMJ7JL+Jxj1VMhPLzMFk80FjMKCDRPZ51GjScl/0wkXIV2TsUIw5hcq
/7TxJriWecWTZy6pkeQWOalP1eD55kRwag7MqQmDGqd7XcmxO0aV3lW8F2jtBL5g/dtXFbKrg4pT
unJ2Wa1ic+9SofuPJNZS4MYYJ0gYkl/VyrEGd0EjLOJIonfBCxQ6ZrE1IZe/10bvjUxCttukSHcj
iqaI+kdh0G7y2dWxoMMlt1mGyVZASqf6jvSREWr82s9FN3kpD663x+vZkQcwR9cG3viUKA5C7LzH
O5hzrwF19y3rH4hL3iqlkGQCMlstVFvEE31/jpHsXmEVnQY9Ax7p+L3pET0YyKzp+tM9sWCtCLR6
/mGhv8ztIC2ZvuUXiNLLHR5+Gm2PxHlg+Jmbg8rVcMNPWqvMMgQQCmAJT3vsgwW9lP9BXymlVPir
sxVaEBMxzAA5Fqx4T9q2jC97KzPVBakHyVrP1bbxKTIgrjSCGH3K3oCfnSZR9K34jm+I0aIsP/Vo
aNNbUKRidgXKp2r2JRsbYbC2y6AsbEvM9WW1LJkUJggL5t7xOcvojav9LPMUBfe2Vu03lvvqAaUW
YNLR4aSx6qal2E61ROE264UJ0HZnUbOnLfxEfnZTkZywU6955AwF5iqDnB12RUl9nzLMBu9l6K3F
iuPj9MEv0+t0P3woHdzFEhshriNlEI5LZqi+l5dWyoyFjQ0DOHEOP3OOrP8d+4eN8TknKIfdIR4e
uJrMaUFaVvZ7dva2qlHAzX3H9fp41n6kZgusFiOMx58LkERt6aFim3CWLJteC6ogykFvAsCYh4iC
O+rd3XuQY80Gpo425qhKWEZ9I4Jou4JfAbb9j9LGw261hN7GtJxUwWdgYTzwTglc0emGEzLXZmjI
mkwtLfI9BsbLDFfV0CAjqJPD0QJe4a6sicoVU1STGJe+3U8yVX4uyNwfkpk36QH9nolUMKMKMGhr
s+l6jzcSPudExKq+uDNoL5Wct3JeXJX5y97IrkCl0I1Ars0THsIpgJuJteHmmE0dZbZ+fb1TauHc
Yw/tvBL0+FTfjSkSF6cFjhjGlizJRP60wTLWtX/ujKxc2UQLKTitD0QHxC7b/6aJwxjgoMBjJI8M
s4oNgEQtKhDwTA2w3+296HgjKOT+QvXSDrYxpSxbxA0Kv0Vree3sb0rDhTS6/K6GDEMXPFIr350G
Y6F4+mzetrpuItzUYGoMce0Rrm/koyE1Z+sx72LHXJ9tuSA4WR0aIxLJOWXex0gxfUhGPrv5EsNg
F8a+HFhd3MxOrkTl3GWSSwVaqxf3YNxyoYlRryQ3GQnMrY7yqWJX8iomFWeV+awVz2su95h6IhXb
QlBl4tu4+1iyoWDFlOSzxXmEDJaKHCA6ouMlwtn60BnOwKeVhcayfloqtx0UX8v+MHupKJR93SsV
b7dgf4fcOvpUGfS8Bhe5WEI6oZbV9XObz4W45jDtRx3ogmlZV48Ihfly/gcxFg0uQPXCnqqZaaCk
5BFH4gpXvSH4O6aGmeIHpb8BIE4ZizJijUtm63RYgTQdAyHXqk2dXZjTmMlf+44YDeLBQ9kEmlx/
A5VhtVLee3s5SXYAb/YNmUAepqbgn0sQAzi7E0ZJUNdTzmS3lxo44BCdcdlld/09+iMLhgUcfDtM
ubVdnwieDJOf+l0eNy4/ETWagaclSsz32KlmQWlyzrQfOQCefFD2UtdRPAVNiJ7FpBTLVoZrKWPD
p02P04id/M7htFWtdBbP1pMIYxj5JkSaa2AfuHcMzhe20HRan6tXxpfedfZZo4DI/KiIoaZcC+Df
mIzz20PcA0BgjegemRz0LVzUtHIrF0akGvytTSuvWffGgSN9QSu2vn8JPzJYh3wtJ+taqz6HnOdj
w1GKucPoSikniQjOkgkP4hFjy6iOfxhYDYdsnvPswcBKvx4zoljyd0IgD7FGWKUc3Ya+JRYNYU/z
EszsogpnrOwoP0MVrUbjv4dxIX1uijJZ22igbk0WI9eFYHs8DBeJmwN/H8taYNLtQ2j/Y2ryJLUe
UKfiXliY48Sn8dVKC+GzN1JlQayNXLAEa5IIhvUqvN7Wjrh1PrznkwY7Xp2puD5tg3zZZZTR2MPQ
v+tBD3qeF9BLWWEGJZNj0d14yIXVIftXzGde2nOLPXOkPqzq5eFejHIzA16PkM6B9TXZ3yUwixOc
9rTbC1qhEWm5i74QB/nkyprcJ2QIzaHX+28fzjfbOUfv9uatXXZrjv+k4hB20suOV8R7UUlOUaRy
yb3l+x9txPBD/sfHzf2h7XmcHwYZFH7BpTIWWlXuJdE2lK7kPB9OeKmV0eKawQRCWR5f6AK6YXOC
HYecC6JrCUYjVsO2DQUzQo+agm/jeOIsFFFvrL/BDscMS5nfG/0sn08J5N+6gUrPKy/aItpviy/2
+rbkr4S+tuOv9NHjrhneRox/GtbQ657AbV4Z5nsQk0SgNbyKIgBLfz0Z9SRw5QAnB8IMdWY1ywPa
rnRwNFPjczbEXNeDqpAMsb1K4GGtlxKbdnnC7qjSFv2afXotPCYHMxiodgUbL7KdGDTN8J6Ubrjm
Tn8ZS+mevkX5INQxI5KtFgyZxl8G/sbIKiPhlIheCI1r6MDqvCy/SiTv3PMGT5sMVCj4LqpLgClu
qhb69mreiu2/JdmwvZKeg5TIbNlVkgAVBhRdguJh54PrEUDwqRDpwY3W3QrunEPcfB8f+j092Wuy
yIdOF8omEJ8bxgWZiLZdi26awHrU1n8ruRCUd0GgSIqSpG3Aitx/5RHypZDy9wruysP6k05ZJg+5
jfZWWPZX278ipf96VPWJmcl1zLyHjq78gDqfxSaFnOaTHfOeTODRjMMW+7TU8j+Y/xUI16ZRjD1q
3nBt2jnatASBwt9r3fb8IvfxFyeKcr/sa68TAOlKWtQD9PLOfxgRQTrL+hF6XsVm2FKovJhzDi3u
ft3VQgf7wE26Oti83UBqQQrEAHSWuCaQxSOckmdwA7MrZja0ISUc2322N2GfnyUFADU/GmOkbYN5
9ukLQywipBKXFs1vVgbyF6jVYz+0mF9oOys3s++2sb8MHw+LLb3r5ue7WrEGWZaHAixsR+X2sy9v
Pt/frbDGZaNfeeDGBAQwMQl4Q6g7jOVtce9PjOpc0ZOwF/G2yMuUYNdswkTaZYAeeAJcv3vi4fa+
7A2txlMggHuJ/TaW+CgemtJUA/QfaVBo0mWW/CfdwVgOehtXnJGVnejdhl0LMd8TvzJqf98oOl+2
WkJ/KO6xMWHLxK+X+RXrUiOm53SF1jyuP4Ry7acZfsq2wgRD17GhFBg5sAsJ0yeRq5sWtVf0pIgk
xXYIJInkeWadIu8eyXvjo28kyUoKmaYu1HGSQl4LqiGyuMGtr9EatBmz2RKZ3xFu1laE1mCSaoo9
lxE1C4/FTK9p8yYKFg7LnY+EyG/Bnl6ibHwtVTZGDbqcGeXS5AlGlJqy13E6KiR+pdWjkOzQDsn4
dfLZHX5cBb+hg3RadB6sRGgE1owASFdE13H+7VSSxME2XMrbTV/TW8PknqI3jjtlCgx5x1J69+XB
uWzqNIM9u2dSSteINEI7eVh22ukRzh8ljlqOyveRGBKj9ba474eU9/heesyrDE3EAgMZX2kVKXk4
PThxmqcZ7DpwSe87NXPZnmzL/utyFbHIrzrjgmi2oz488Xu2mP1vxBZqG1i4fzMLbMkl1Tkw8k1l
DLe4f85Uy8B5UonwR89wGEH4BmHaKmbM83FTAqJOVHOykjDKNtLg44MAElYu1++wXVPax3y6XiVP
tYLI3L8liKp+pHD0Z/38sp09k1CHlaCqsdLi+JO6tTWN8kYnrh+amZ02GI1PNB8uXRys/sNdY1dO
rqG6miLKtjMt+zpAd6cLEOPJO/UUS6GVRvqqGYwNEptleRoihpBoDtk7TBnrOYSV4T1a5FhWjY9d
wP+BAirfNMgySsAZ2YwTIO3MlQ15OZGpJ6GwgZJr2lf7y2XMlsoPophv4BT+1HC/F4iHRW48Iox8
CLvus9b7zeVOTqNFt0GLyYwza80ypYVEUptN9k98CDfhqr1bUWF0TSvmxViTa8Pz87P0r7tpMXr6
BCeRKPzAuxuBZYJecJz6Bm+PMB9o14BLucSF1FfjxBiSi5xH/E7pJyWNcWu3SVMA5UgiR9aW8QvX
4U+qbaOiKkWJvMn/l6OhLgAsKbFj5vvg87RBTn2gMWYPsh2veCtmN7rRlSIeWo6DrtIjIODhPrSb
xUeXJReOsyM33RKp3sMG+CrhSl/4FaaJ92Jv2gCeTfIv75jt8vuy69MSWi1NPUm+hdc5cxHEPY//
kWAdohcZ3FDlpyCWVFZqUqVTtKQgfoV+ZCqqrEoJKEEcprRRkXdY+V//zIKFoOkS4GFCr9LAB3Dc
m4A4gesuyvZXJHqhEYoAz1U9UFHZMpwB5XvT1EgNCTVq5B0rk85QpDMh1OAfTdcpbuqYfSZx8eC5
CVB8pZ7HGscrH3GgibN83H3B47vBy07pWYuKDNfDGbgJwV7wDzle0O4qSDjwDfcOe6ZN0rsAjsut
+U/yBjNfuPo0e7Ox16pcXqw/OeMwf6Jh0U0wOc61wxVltOiI7ZEu9WJUhNG3sPXowmM0Ie+YpTQq
LbGipNIR6kv7b6+AmoKq/pnq3L9nuvUDyh8uMNwJr18SRK9yPJ5J3OiSaTv4NGxtRTzbOc1j+I/u
bd33IsJKoN2h9nhV3H84lTI3e+MIqlu9xHS5hYdMVo4B/dTtM++uK+d0ry2BoPt+kVxEc9Q5jDvS
AfdFXt1xekFrSHqxovGnS6BdbvjhbmPLjpZcpOFqPID7PP50yneqP3ne3SzmmaEkRscX0e8krPQw
HBP0QXqL6jK/xzwH8O+0Rp2wDCZIlyAniqakp/s1mtMCQyEEBlenA+0oYV6Om6cfM2/UGaw52eVI
sLXCyD3qEdlPXhtaDOuASNe4RTRd6EyaAV/d4o5B8ljOIJ4Aeesv2eTVGHlSfG/lrMwN5d1d9EBm
r7uUC4ifbzenVsWpQ01F3Tnqsxry91UEdOiWwbbJhRBMC+oTo0eZju2P+RTdHbFKCFCwqUjcZjCE
jtzf1EKO7cnIeH+qPJtLVn34Z3FTMRrvAxVLVt8pdz7uV7HHpCNjRoqlLDGW2WvXfMGZ4rqxqz0Z
c9YvY6i38D30gPJUJ9gBRitNDts/5ZqaXarXVt+P7O1p30FpBDaoEtdGMYWLLYBVVLLyErH5FBkg
dyDU6W8wpF/IuZyGiIu2rmAt8k2F3VnVoZ1w2PEZIEwJ1lSkWQO8tKdjaZJXDMQGYs+piHkNho+E
tuYW2EkW8SqTKahHeiNZOxXFVJ6TKComADABWrSbYWMFS/RpdyeW8sNH1dJSjvTjhBo74bM6G2Q5
jOrNmiZ5A87XbYyXQTyNumukrOXIg6VSJIb6/V1DhepCwascVaYhVqwvVBsfNpRiJ4d8MZld77kd
BFEW8J+CuPuYcxJwMMU2X8IuKbDUGOJjBlQkkZo6BJTuWIbu/V98jx2G8J2DQZfp9IhP4uSLBXmL
Oxx9zIs0rAGjzpjFDDYHXa+qF1JpGHtWhYto8QackzTq0aPCiTE3QVk0sbaTvTW59SryqU30U5Aa
V/1ZCzzdIgWfcD3mGeljtyyXlyDS3fQgDmRJhZAq3pE2zVvtdwl+Osw3S9U5RhljyS0tCk6SAbNd
xp+zYtyxII1/NROkJATIwLbtbRn7SLy+pLMLCTBgxIolIhz35IMsx22Ig1N7xajizjssM1eweMRW
6vEiRfLslGNKZUBHGa7JbL7kXHSngu+AwNeDf4w6Wj7VZ4DHodIr8TYn1p1P/jlX5rt/v1dLK+0T
pj2qqhwocIA6QabVTXeUbkBwo4W1whd/fz0R/hnYiZ4aOK3Ieg3WWtZLT9dW9QFqKjOlL2Lef9WO
aqtN67jAwkJapRh3gXays4LkiKngomxbA9dPohXffSOtS3cD18tmXpXTuG3TyYelLxYq0XpgzBXz
5xGxL2FNFGIVezP/GOzkEveCI8NVf4yNLZHtHquvcZoYpomkt+BRH0NeGdTua8drqdht0xv+B3rq
mJ4H6Z9KoLz8XNv6Qphww5z22Ofmz9NXzfjjubqCz3I/gw6dfYdK9/E2u12fR2Xm4E+tOdcjmqqQ
ZDc+qZfxVSQ6gddGUqKci/6QbjxUDlNnMY4bYyKkiyIvc5oTPcIGCQO+LFAdwiaiBPf8WD/FU8nm
Xv7UvrmwcEqQDdIrOxafQLEH3k0AvtlCsZ1nJwGSiLuiAwRkKthl9vjEnYaYkQhjIOsuds3M7qzX
I4Yeo1ePtA9g3o2QLh33XjxiC76D2HNoz4i+g1uAqpCyQJyrPDjgj0Xw/EueMTdysCNQL0F66n/2
EWg2xUDzTCJaz/hhNmKS7bokRNqYr/MzZ9StvqomIv6beSNEMEbKBgwlt6gpWCVeILZlCYjtUIxI
Q9NWaZV7wkrk3QtyyP68hvYwMvWMde+IG+iRhaUHYXj0bqZpqg5oDexPbH5/n9j3N+SKiOujuhXk
B979fUNGSmluW7PBMmo5nsN8TkHbdfcPNEXgn+gAB+2nETOQSjOuPh06xNPV3zBmUG8oYSAXI6lR
gEpwnNmvFyjDW2ZrCBWUzp2WkmiRxVpsBHbmH0KNFdt9Ocyq5hbX+A4lOlskCsibVE6GW8HpADR/
7SW3+rN+vjqQkiWLzOqgqvEeng18K3Hd0zRMWsZHIle16o8GeynhXVR6M31+XInwGwX1VNd5Ei2y
63JbT953vcy4MRQPylIApgSwr3OxCbQGFJOyoOy6zbAXnNgP21parPE3SJ0SGU/u39c/HRgXo7Gi
Be3ONS3M+CYVtwt21tDVW0AMMtUHpXIRKancQ03dvxIQuCZcUW25gruETSlpOuum1xDjcs4cELfB
K3ZZhk13K+8YaQQv0IHHEueNH4N7dFEqcajSbSfjHjukei7VslSi5EmsbIP+Piq60OK6XPCOGthV
SqWQJBT+kJdxTkC0q/Jb2PbUR4xVHmHqRBlAyR0dPLgYaiXB1VtypCaiVEv+6qsRQporNlYgXn90
+xFPMU7GAwhF1l4tfx8jCMXQ06sdT65AQp6zoPyOOJ6tmg41m52FEAKle/+c1H3+OxhWVkWPSrCs
FvlMlMPFbx5OcZgemEeuVGi87BlqZzo1Hn+coN9nIKIQeZNlaxmYgWqUToTFnxDdG6KIzcg9k8RV
mbaFJjncFGngAIepu0KDUsMgU229ank+YB2dfuHAEisu2f2aC4gyscfiVIv5x8NCa9QtrHb4jRrP
xhtpm7m6+WyYiYJLxxLB/0KE/qwvCCG5ykJkAokK4oFLElgs0Vz7ZnNfh+XzyP4bNcugstgUG2Y5
BFFX9kwkMBSbJn6PAAnM6SHzlj2ARsFYDqe7sD7tcoNVRBk/gNdoTGR3uMj/nzl1YqtTQjDTPtaA
1x+K4+DT4NMIjYQaY9edKOBW3anu1wHwZYTHu55l6q+K3dtH1f5PEkXNTXPQteD1Pjfe4N6qaUtc
gPf+8V5ituVifICacChVYJNq5ApTe9Qj9KOReiQAd0fzDBvTLmQNBB/UQdzhWl8bmn569G7J39Q/
YKgsF5Pzi2vCHGfhGbbzgvNuA5+UoQn9IQYMpOvgEtKy574XT0J5RjgGECr5s0oBe8jpdR2zrJ8D
ThF097rmPDAtgooDxVV2FMhs2/XmkXQkbVkmJGXSRLljO5jqP4tQMLSq9i0I71X7rct8NB4djX9A
b9icHfwPNQEsVKIjR1RGAiztAsEIpMJu15827ValBHY0FXiLKr8h+uFVttfhtdZ8GSzcz7sX/qMo
34z977MJXEi4N1FSdYwH1r7gf61IKdhxc0pvdgN1yz7gfM8rcTRXwnYITOQq7wvldedxc6eua78r
JMo3XHWdsOF6Se+Dynn+cVTkKcyPfMdJlzoVTLYMm9r22/3biU23FhqerA/CMIsfuh9GDrLh5Lzs
mkZynWDTG+PyuIL0254jYnYCAJuF46nAURpoo9lzcipAYDJm+49q9QkWncPrmAFKcjW/uC61q9vo
g+FO4kMLjESzFmUbQNXcEBcXXeTJTOTRi8M5iJOm/QOwOKBLoMZ0m5XO+4JjRAlvKWP6dgS4DAlv
tcdJ/xLdczAOUVtDPwnEBL4VbZ4RprUwbB/U9Fc1j9CJfTysCYQhzjomh4AEWlwVRdr9ky4l3TTr
6ZoxnnqzXYKhIyvSzOfojD/7f2Cw5veusdnqvTmhufF3sWRQRIfanvzVPiG8LTnAhAyxZwVaGn3n
J8ZxO1AOMwAxS/yXFh648ovJQiQAqsEWGnZbJrndfxK4qkoajZ7V0JGoQYs49FfESeoliMDiuj3P
ax4TzkZZB5CRiS3hpuO3HZTWOCPqNYvMCoePKhBmO5KJ4I6IVQO4qWDnNnVoTrbVhFRmMC44qbwT
hB7ZTTdww4lAIQLfz8AEv4uRUkCcqOcKTSarfnZ8ik9/tHfNq+hRT2RSWXmgZI2WfbFy6iI9Jrjs
jx9GZ+sxNhnjfsONE4Vdy/p552dPDsPy9FFEyf0mj3XMN9zb/XLJ3BjgH/tt9CvO7ft7YYx9iOsn
/6j4LsLxzBRFR4aGRofoVhoyI1Lkl7AOdPx4MDi2OPQozIC99n8eNp3FMI5nlOjvHEdVqzM2l6ov
vBZ/5o/FVeOQiy0LFXlYzP07Zq3p3i/p/C6ULr9Z8V9lvwtUs2ZiC5ewo+DvpKP++ExRo/wDkoa3
N+kJRmv502uPNUTvjRlE24CJfndI/XDK9Dvom58P2XaEK7oyvVvN17lpokkahsvsNPndEMKaXyFG
HyUUevniZRbYFZ5XFieV4NmvwL40vOC3j3mdgZf+fRKdC9P6tiSIg+9rV502yBK3usX6LGjVkwpr
rHzc8w9nlrNgef2tD9szXUrVjXcr/pPmLRYAskmKGmTRxf+34K3/6GsotSS1n1txvl3YKLyLTo0U
6VaRCzBQdst2J00nAg7HZZEEoCxt3QxhKaPUFyczL8sO7CT7t3rlR4nRcv/uE7+g2En+o8taiqVt
aZF4Kmj51nVaYhmOBIze5JVhKX0KmajwJ8MujeS16ejqJsRtPAjRUt3j7bG0vc+KD3fuk0yOPMZ8
R8cDsyIPEWVQhhSX6YMltML3JvoB/lmw3M9e39bsPycZZKBM9QDKZ4pXTD3AWwjFI8GYjAoTAsIl
5rPEnzb6ZPsGhnxuIuuN5aewRHTBB2OEhZM8omcaWa7OzcrFj+J+OGIP0lFpTAbWG9Ff5N+ppp9e
WfOHDnWgS7hiJ9svNJbvfC1sYgr9lrgEDyLhLPhx+Watc8226At62u3pb3KX5oOATA1ITjUpztbV
8s/mEVO+5yvdURXAXknyctdpp6bclqZeQGdqLK6OXvuUfugdkgQaqTgadilbmCcM+w8rThctwL+q
obDGrI0kpfHWjLo8K+a2ctZlM0CPxk6l6X0c/XAZ13zFy1eruuT2OZn71t5B9L9OrqlaTop3+Qyg
/PEnW9BTgH7R4jD3Z9GIhu+yJwHEPJVBNxAni/GjfFkE1IDEcei+7uQXcXglxKlLiMdt/I3wG9Qb
LgytBmeTjYUcu6juNxafIGvncTOS+yHC36/quH0eFY6wa5GG+wJm4I6ziaRmK/wWDTfVbt9lCYF3
x754DGGEMxVxomDasmRLL23jkBWPLUcopa1IWpi9qR9xA8DIXFSzCiymnA8jMgSwOmVhZqOcG4xw
QTqZzOd59e1Iqv7kDUfIMXvMnP9qOSB1I2M0Un/iLrQIx/loDhR/vvkqmMMUnc15NkwaeCl6UtnZ
Eln7xl8qJQRVp/Argj+zH6vTeYJ8ChCOJQJNjE7CLzKW1n7R1KSeufp3OBI9vVYALmP/bjou+LmF
zGv7nB4AxgscA7xizOPvRIh3iYg7FKCOBqJk6SmP6aDPNCbOffa3UrBTniikx8MlXtB9QUti7gy1
FLS1Rj9zTOE9q9bBm8jHcu6O33Qk/f0J/pw/Pwxt5HEJNbBsg5BebYMUrFdOyXERbndvyeisJFpV
vluw5Sqf27Tkxo3hDheuUBrUoZNXDvIj59CiBxRXJ8kelKwxgZvmxtU2ECIo7xgrmmuPGw0oynyq
0wfIAOjZXo9N0JKY8dgA/napGUkUp2Ke3Z6j75qv6zY6njNjWapWajcqymfUkMyta+1RBQGDd0yn
xVsHa4u5MK1T9OO4sSJdsrO/Aw4uGgSAfqUfnS+uNNamNGAgz77OBAD9Llfu5fgXK3de9OBoChwW
vToMJCW3On6XTpUokIY+iP3bPzN0WqI1FkiT0gMcakD3NL33Wl5p8pXlczvbDIKL6U52WTyEsY1t
souQoTPy8DGVM/xAktKz5sJiN/9im380ig/RPAUlNbjVVYH0XfIUoGqjE8AWx3bqt+j8cTbPoiLQ
4D2g2KZH8f256mpy4jfE94dYYBFvUue3iJNeJkmffkUSkS9qrvP6ZhIVa8U8DfQWyL83KoWgTj4B
ZZnEBSm5fc+JwO4ufxt9bsxHIWdS4B0oVpc2TBhWl0A8OH9p2b2uh5bILqWWH9DuQ7bSTlBLusqW
AwAVyecdHEC+1XMjhpZJOdoAJ8P52jf7OAqOjOAHXyiPhJ2PU9w5zLVzn+xiKVnuZhpifktS/1hN
OxvI5bpPEDu6X/RlhOn4sm85A1PjBxg1vryEU2K+BEgf7XEvxqmRdnkcUivuBMOOavG0lJNSgfnz
j1roZ0tHaenynXkGuld2Oto5fZons29iN+GQ+tHXI+J5HnkNLEXRKyg6+UVtOlhGCirP5kLjK0FO
KsSAyTdvku3yAbiEdApF9bdo+4Q0RRDU0vkLRcDGFQ3d8kwCCli79KojDp5Mi6crWwdgDVPhopM1
Rrimfg3qZPjJ9WE+tiiRkqhV9FGvK6kyIumUIuNl/rbVFtCPYHrbaFheOjihMV7kR9H1cYk3A70p
Ffiif4TnfJKt5CAHLqf5KxoutwXJGnr38rqbcCTlVLdHUKzLITrWnMl73T0KmTSaSG5F0Y3iLp+s
Ww8Kr0onP33oR+DH6ITwrAG+r2EmhV5ebYsPzy024tJ3ja30rIlR5B5Z+SbrBL4Z8yJS/8qMXH6m
A5HoMQNFwB2zhKmRVj2SvoUHojyxAILd2BLrfJp+lu31B9hVVGrWe1JYjEMMlw+FjivV/IrDSdnc
J3JxF8ljXbYZoJYmoP3K46VS7c7Rrpxk4aSmzzYJgLi0O1jQ5K5NkgFtFo45Q6lkrZ06KBMob6wx
plcx2/PhWZGYNJ/3kcWGNY8Kcdk+JEJVPJaiI+X+XWb1DL+YHnKN8vrMrbNytAuzoOZ3M5AznJJT
Ve/30jJGS/GjfaDmfpyhgeUOJe5/zeGPKP6ohwfo0MN0ECMek4bkPuKnvEMNjO/YqRwOKGXgauLc
VvYo/5f7j0jIUzNt6pPsqsbXeVzwSBPNkwKskQkhhgT0KtOYo6E8vXjWzWOjjmZAOGLlBp0fDYy4
Ufug/SMDoDfIGnSowsuK9upj0h/wscI46LHa8+q0iVqCBeLKz4MVZXp/JalNmrg9fTt+Qj+MUhJo
v6m4BTbpvz84PrHUNXgeKiSNSHzbsZNCEMLzvAOs1xzld6VrE/z1LJsGKJ0QQi0hHl29KFJi/6jI
/tvOmofY8g7CRr1GQlKVTXjUQQN5D9mNKD+siTPpYIOUQ2OZvUXw17tgCCTuylOG7OlFc2VFmm0x
EaKsBnvYUqB52knVFZwXCY+YZtDVwb2Z795pAWvvPESTjnmi46Y0N+6h7tDR87qBSlSWDxouFVCI
Qv507NdDU+PXDSwYMoQ5MLmorrtK0mRMWBa3APgnATgAo3V1tKsYblNcIXrUFvNRy3e8bPllODn6
ml5+ZFTA5tz4eXLb+yO5qYaZ7kXZ40QV56ftqHjpbikYuhCnP4yMTjtd6/XYqv2QWBSVZSdu958r
Gt50+xnP1AbLDrm5XXc0Yy0JMyoOwhYXKTzq/+2nM7JylR0FQK5hEM8+iCpMY7ix77MEcjN4gDyn
gbUueZrgQG6C3a1LJ8tKamGdksud2usdcwb+doC/v4to0gwLMcbykIQbGBH1ua7IpCrZNHJNyl/n
bi4iZyAwblsiOmeQUSUkq0l0K4uVL/hcT5/a2rOAgKb+tYI9c79eshUc1g7BVhw2nVS5B+fWCzLw
4VE3X4Xh/kAIZFyx4PuyqXl4AwTiqD3RGCq5REpWGcgaUrqa601YD7MiCsQmtxTBVLXwtBucJkPF
LXdnIHe5A70HZwTKtK87zxjFwDL6Zghj4AKfhDgvkbyYy7UR0rgT63S08PEIy0OWrM243hp911nH
2h98CpY96toHwM5ac+J1GQcv0TK3FFmjt6Ux1xnZj0Br/tQQ4oTcml25VdfIkaDrXa8cug9d3B2V
L7qt4SKbrlb5gpmAf+zG8mk+um59Wk/CZ2P1/klDOq92TEWhLXmgpxNonRsS1ktqsEpI39Qvmpg6
4Px2SS7Xn5XeelJ5xnCtNOPfKxrHAqNutQq4ovMXlco5LOVrw/kx3SqfOJqiURXP8KMQmotOsn5Y
YBerrhV3B2Mi9eMism8ybkdrel+d5C8ahpvxhQB5b0G6JLVKrpQHGjxHv110/b9KTbmDFO/99SXT
kymzzNASbp+nP/3DcPzNGl5ZrtfOCRqxCipGjo3AUz2DGlncI5N/GQwghNzTUcW2SaRWrIPIbmK9
lJgGgi2JPKMAElds+Xb40RvS6dmRSWqzHqwGpGt0iHwfT9vPYf2B5iRnZEmKcXDGrftmfxP7DqOt
ki8N6keZmdlP5Jm/3tL0EsCHGLdScCx+tJaEqNdqJFr8BduQ/rgGjUGAjrYmU9NvnonUI89Aw+8q
g85nSbobAWHkPgCEcDsLmVTwlYGPTU+BGAG++jswzFF88zDvMrN0tMFU8EFNyyWCGUdXoeKiYBZ6
Dkl5SYzZS99nrI8uVaixdX07+N7JF9Bm7Iy/M/agtaBsuwMn+uxxVc6SmZstbl3qqIIZi8ZVKwdE
quxx1hFqxNNDTBQgu5ExmOX8+C1J9NT7It2QQH9JZ/8NWA41PqJTeeEWuEQbul13rnH1xIjfDSec
qglqspXQQGbSZFs25nNwpdHSeyVidZzpdTSiSuK61orzNLp5GVI4XTU5ybhbS8f5PLcI64sfo8N1
ojR2Ix7Hc66W71ZLobGDgLGGn0GAWmzl+qM71NQ+sBExrXNdRIlXWJcXhJ0mgVuGXUetQPGsAXCq
3Mi/aWs7Aick2yWO9gDIf0GGoHwcuoiM3UcXKWXR2RjkQq7Q+lo25RVbyn2lo5WVA28c3ZYGiIM8
G3kUdXF9iJ+H0BJ/PUk7cmNSwrwiAamnHL8vZzLFSEuDKw0ymmUTxjCBt41qsDcj7rhPUuvJTGUY
CUlXc4R3WdDLCogfHu+4pnGFVLKlCMWEooaFima7oODvvME3Bp68Fq/57/l4ijRKCZJBxUgegDX3
eKOnvSckZ5CRBgzpdyKqmRxnpGJOv6TyaMZ3mvwvqjEF4Xqyoohr8PoWH1oiweLejIeLEXpSNEIy
cfA/lLuFdhXNg2ktZW0i7wPDqmDnmqMw4MnXiKn4KUpuJFHOYNQWo9EGs6zNio/NmgdxCSzSojr/
mnidLJNuvQB0dnG/lvQxkqXd6a/S6Ia1abWD5BhqPgzN7aT8ijRbTkbZplRpOyo97e88NlRnbU6f
h3El74CoDQLpoaXJE5YrVJCcCE04cZycgFmT2sfM3geIxOTBkFQnzsJWTz7aiQMfELI7rjlXl2ij
YOci3sSOhUx/YufzHU10R0sQu2xnIja8HqttMEMDg/frfGaOBXQGIS+Kxe6UmKW3uuJAMNBOMjcw
5xi/EdWXwrK8SCxLFzJ8Mm4H5koS191AXw0n8E6HUIc0YLhXP4kxr/V4EOyvmEWsFiuKHvwPaGRQ
Fvpa0Bz0TgMg83Z+36ngPSfPpw0HRa2vR2NCT0Szhq5SwGO/5E/M6z5WgkYL1r9sCDd0w4oG1nGt
aFhh4d6Jk7NVPlBHdTvaSnSD8W+1XRTX8o31MwwhmQdWks2K3WOh5b9lWPzRzzNCKSMUn8VdcbXV
9Q0QeRqksafrqU6IrLyENF6X+yodSkRIlk76GT6dR3pgX8kPXeTT7QiGlQ2RSUDJL3FJrHPTSc9S
UPs/yJRXlMY8tWtn+wkhFOI7vOGtgVdIYXMHBKIvRUWHvVxkIoGHVgX2YfNbzWIgTSfYzlPQpJgt
aDSRr6dkt4E2wPISYP2Te01nZjT43qwK7XJGuypIrXainy5dFcqs6jQAiaLNikSLsSYN/6vtGYaX
ueBZqV5uP45lndZ/Rdae2K9Xf9C86+Mkds5Sya/uwfVt7iSIDgUYC3nUaxtWwtPEvHuxzzBFu7c/
TJpK80S88eu9hs/wP4jhJpU6V7P8NYre9epOTacW5fn3BNOhBVyFoZN1M6kOlWeGZSSl+AYkvcDe
Iz1kTe516/JlXJem22Avr59FtGMQYssRnKuER6JNC6l+ixng0EJtOfQkl6vXcdKt2HbxfgfDMlOa
hYJj4O55lB4qsabbwhJtYnIQQXDIBRtUdvOakwO2LsPWGd6M4IrctKjJ6XjVpDB12fd0c60SCq7k
rqzKvWP9YkcwwdmUbjyqNCgMHK0diO/vGldCJ/CPF6oL4kviAE5WSUndYuK5RX6kH0Z41f/u3CBp
cgRmia8YE1yvFY7YQq9Dhfrr1YeOgaL+2DHbZnAtQ0l2YCyJxgsipyFieCJL7/2g4mrYlg8LMWq+
MurFZdR2ucxfRrI/vikrk0OOFhLvjCaqvtumPWWtZPjvwdzZ1fTbrBmhr40OWEfumK8ii5PIzSpb
i8iTgzTM0G4wlIoeSmQ6NKjMPkPY/Mn87emtYNz0hM8mhYLjHFGSmSHGOPAhKwljVJ3kiZN1pNtx
CQpqaXpCoVyw96Ny4jmrTIB8hCweXHyQbsMI/fXh2zxZ6BURXu+6V2lBVwcbY39iYnVT48lSwxPq
7mEgCeNTnzBTRxzV+TynMzDcFcPHmBxRgxZOJAV84eCUtUhOLvQ4o9QEEz44NJDx0j6xQgRjiZ8Q
yg/Dob/oebapPZg5RgVGUeh9Mb+ZXeOZJIU0hOym5METdfuIf3kqVJgQDe3zF+cbwtPDwLk4iBnH
hTg+7hCU6kvNv0o6rTYwk9+4YiDdTRQn2y1zqCTET8WBXl/21SUsJXUIr9XHQDw98q4EeCxzz2T+
zOw5A6pggKlYWioo2pfTSQsm9B10/yL3Aqv3Y/gJW19Q6zPVMf8eH9d2w5Rl7OKvkHZOeP/fsbh0
OnbStXGu1QrU981FG4ZRHPzAxmgrhXwhqrBZrmWwfHNQtMZ698nVTBorFRqaZf7ymfYdl5fXkvSH
Xyf2j9+eoz+gwqOTLViqiST3OumyZPQfV3BtPPlgHhjevf1GWD3WYGCi9PYNDwotxcUB/PFmLnYN
xm4l2I+Z0t6c+p6d5EQyukH1MqotGYIknjb73T39dTzt8AlZrJvc+BsHBgrhhKtsxwBDscPouNOG
1usiPXHD91MOqCT+v2xWgR7TiiQqFETLH075BXiwOwk2ASJngYKUzxd0yBHfkPnawdUuK1o3eSrr
xkgPuECGmKR28TCcmoGgyhACvSqgAaJC/80D84n8LXFmktJMW5OinNCKcS1e1OL8PBcVTt6VjlQ/
xMDErF7ogPP4Nab2eyunMbHMqy5TzPmaarmN5IbhXIsFdWFRfmRnqCqvIbzJOX8xuCYILJGuusSr
ns+MMmJFT+mV1IaNMkOMJqlw2ix+Jez05c5st7nWHh0mo/SS0d9cHK3bDUcOifh1eLBG02ENKb56
H2QjWaF0Uz/WY1+fmjTXCcPMCCtD5k3CDlO/XI/51F9n4UWqX3PlYaFTsV27uzMOtJPAeC7PD0Qn
sM4WscBrEZVMd0JYdD3yFrlK8+wtVITYPmfgmYdGjmUGErvk/WnAhxMfoRWgD+e4ejExNk8eH/u4
YwtIjsU0nL0HubSX5OONxTNymLAQrT9nKHMifoN8BQELq/7LucNnPjHwMJTxU7blHcvtYxUTeo/Z
+C3cR9DA1I4O2J/XuLhrhXw4qxlOfg+Db6KOdocC2SJonMP3OqIj17y5wcm9E+bhmgffGoOOOm4l
Y71z3D7FZ/vqI+IMyOhYByb+d9sWLcjCXbNxP6jmUApxOEubx69UHQUvO645zvMCIsOzo+uD5C7x
zkdyAurO6uFdd/fm7Z54cNY3y+jleIAh3NOMzYYz0YeiFtMtfD2pKzXmvajUllumnt+YyoNNyElw
7oUbn9T3ofjNOZU0tQQL34bw+VcFS304sD/o5PokcFeVVtjGPCulfsbqOW7H4u0LAFpc6s3l03EM
rn+X4ljQaKDVd/V0GN4OKHGCBZGYSZBbJJ6B6bp4ujvfdZvsUtirl3OwKtErWwgc0mfWavveYuBv
1H+sMCY47z3iJNmdZmwiG3Bpt4rKb7jm0BPvtO6QjPgWBHiRQ91/1unFVbI0+ktQpNj5vF9X74Ak
AvSzzEDQKj/agWOpE2Lby2jeF2XVlVQ78s3eXrK1Zl48lembBG9waGz3tFwZKWPZ6EcgTWlXxn/7
nPMSpJxi8gUj/Mie31BTT0DWMccH7H1Fs86vQ1V2lNJt2sKSvqLKfVxkEo1wdyouYbU71ohAcJd6
ascdJzrj36aTinCNdMZ0zRzsQMHuylQvZtWj8v2YM1WFcnCEst7YPbhOM9f4HesTS8D9hROtGNNj
RBJf2TmDDD9duzJLkaTnRXLbhyLmy1FCi19mPIaoIH7tKFehmDSUtTL+l74XF4LVjxi9br4T3WuC
Lkqoy1ti3HrZnOPuueIBPF2A8NH8Dsg8xT661aO9CiRutICkTBrZIa7JXXtYNCAvdhSAB9NKt85q
u3Dqdh+Pkm5aPBMpcFOIUQkNLgJuh3QxrgHF+1RitF1RGY4ygADpB3/JS/cV3LpOJOOPne3PRfIU
wPVQPG7pXO3tzr5Hwi08uvMhmE8PWmDAB+dcLNt8YbnZsnuZjk7c27dPuB3hg/mChy2DknWSHWQ6
5Q7nr/iFYWlQKLN+qAgREMfo2oR4uitxlfQsh8Nms0j9MSBwti2YrByiX462qqdiShuYUBfZ5T5s
GGVyDPbw7+D3tUj+4btTzdAuQqaqTLnsbZ4p4Qk8dSp2j0fASUVKOBrSJ6E59KAlctay5kDLTC1/
cq55+TU5jcAXlN4jwpOplKHj2n0sFhx2ZaxGU04/YengWfFF6RSsPfsDcAa+ggsM05L09neOu3Nu
7mTBnsmJS7iPVCjAOGPxJzxLFjGurlZgu181WamoUV8g2CULQJYDjMXA8HnQaN/3R62gXPlopZD+
XJ1S7oH8Hssw7wGcUoM4r3V0++MkDcuqps0GHWULoJ0PctoK81zh6R/OTPpi/zpZCkTmXBe0+JkZ
XHU8tBaLbfrD7fasrHNpnUDCU45Ep72hP0q7OrmU+XjYNK0fC22RrdeKyoi49SvHloZyTdwXaKmo
453gM2OVLeXJO3tQV8s80vcAQOkaEU+aKAqnt42SvPtkKZvIqqK1X0PHI0m35m/pgk9VrNIjtQxR
Ug8q2k2p51LZQ0RogdaONHLgwmprlWqhSQpK0Zwu/psi8aMxxzJWebPFQFURnCEDluvI5RrOLb1T
BzvyVk/rdqDGckyaewIk60cgOqpvHygSR9CFFn/flXe5jCqCgKt0xQGe8+1BTjgeDl8cnJKy7GY0
d5vsZuDXlhT9HkrObvwvqGhNYmw6eohJ/yw8DVZsSUrd/TWIcGtQ4FqEDw/ygMdO1r/YCSUPctKC
kLsS6nzxLwPw3YN51k4tx1c+ymSDBbuLsfGqFtvPAdEwFmFNwKjvetZNtG4R0pbAqgAwiRECHLy8
mRvLxzNTsc9mScx6gpQuQDOAVEkCtxdcGfiasLaSm0PJm5Cjchze6hPLuJ1perTUhqIJKQ4dsapA
CO+30Ca5TqjNwaeWPIgYS0dXmV+0IUTaRCrwAMBm7+Y6xW8QZdkovTHIBAQsK7RYLjYy+bseS50O
UI8uav79fgyXYw9zWz4U6wPuPcBG8+enNtWQPHEkVYD0ZJAFljuNLIH5bB7fRIT5mnLGjznjEqRH
+NJbvskYd2L/PTJ+Q2P0P9Vz74OM6Bv0Vf0H4l4we+PITNwMdvzsB5RLUSOIyC6ZRIDdJ0GeTMFd
qBlRQY8nRwnbPvCO7rZDEZtsQ3ajQIYe1acTw976TYpkeyWpkbvirIr4KZ0jX+i3gRt1mRvW8Nxy
FDCeHMpp5IJ0PS100ta45NVk9bD4QFfLg8i3btWCDCQdWWh4+ru1N3aBMpvWVaEU/6cRFN9X9ZMg
S2Fd/2QoNkSRTXKLzxK3fVs60EvOESZbarbG3NHfB2hzgH45ZjxglnC2kyldKvXD7775cha0uVC5
NwmJRXffxV2hlScX0uPLF4Otz4iWXyIFJ180ujjdygP1ugNm8uvPlWEJ2Gth1Imme6bcRpWaXESI
buQ8f5+H/Wp55mWJS6pUii3pBlAJNYXJJUbwMWBAWBONkhDQe09d9E+BMphUu9bWqwKimQ/i+hkS
IRPHMxBwit8sWs6LGC0l+vriw/OsVyA6DqyTbObsxDfHKaNI1KVGMSPBXZ5jySUs3749GnI694sX
ZqBUvh0FCNk/xkA8sEeV6xTzTH9QxazwwE/uZgcXGiQQCLQibp2r+EiY7M6GGhZYlTp/eZqzk3ec
VQaQBcnxWrkm3IODPZ1VPp9eS04cDoisJjMiH9rkyV52dmq+F7YyDltmRJgu9S8we5Gj703rv4Du
2tSPFxNCfqWQQfBcORJwosHOUU+frWKN9WAMTbJnd3Mxl27Z6SK/FMFUYyczZzLtq9qMoeOGONMK
gQerKarCSzztJE+9kmVBMz6QBB2ArPknl0vfEShRBewncE5idQK0QQhAdAMnVYfZfcAjMZEWwA/D
5O+CJP75/Id7BoBGJn5SdMpOGP4EBi0EqD45IFwzbxCtEK59vl6PtVS/1TGAFry58y8GPIWxbXHF
i3H9AADKj9eg00pJLa5YGsd0sNn+WnkBlo+Iqqv5hlGZSiZoEnmwtyEGMNVB4bJ6akUY9wkWxZP5
9kUoKlkvBgphSvGRYVdnyOB1OAKFoXtiqWQSDao46W+TbVvR5lAoIaLITIOjiYFT7u2cNuub35CM
rNNomHVStTygjg7OH2XkWyQnaonJDUmHWY3JNPuUokfFQe958sLtVssInB4lGdBwQ2KJMggxuQ0h
NaJL0EBfbDiT3SZ6xZbY9Cu0iALw0V/CYqvmfSeDpLst7+KbEICRfaLeFx2pIA99x6FdssdNM1WI
jnSYAkuKiqhpqIHe2bbRlCnP0XSoa9pab/+33jH9B+jCvEwV3IjwkWcdVBRJnN0HE2oflvgHBikg
ZPA9YlmYdk/UNos517vx8l4ZzmvqkddEUYmopbwojlflIngsdpYbhbOWA8yUXeLYQZ8JS/tehdix
lX7gItjmwMN4hnvXl7pUUS6Ks+cQSEYNElshrlMiwPbGJmxYXXn5af+Pd5TNFb4vAnYUb+XXy/CC
j1MWUaotuNOgj0RSa40f8dHSgMEQM6bzzuLKiVKVuz3xCgZ9zS2JjL+5Vpa6ylVNkIJZH8dHl2Y5
OuxmkLIfuNFAWCxgHGjWEIqacCIkp62s1tK1O7KPq9IpDBYgcr4A3xJftdjvNoUt9aPXzj2jKkY1
sXErmS1shTZfHW09AhJB7/pff+ExNsFN8sOvq5i13Zb8mab+48Xce29YOvkDAhq7FpBPQSZzpcHJ
uoTFTvi2k521LHfRRioeAwGPYwCN+bVliPeJpDOn0Vlqf+KdpQDvEQNGjCyV7ECczYD9Hr79ypGF
oQIw8I32g48QMAROGqcpLrRwWbhiCKV7wQkeLKmusrFUF31wRQa4DBlpGdp9z6pbl0CstkqVUbOH
zyKaXLe3kzPDnnDzL/Pilz2Kxp5gP11qTbM3aS95AsVu4JCNqz78prCoVXwgN3QRb5oPSsHuVYsh
vsFUjBckYqWReltYkYwNbtcHF60FLIDvQS639wWMwjkCPuZMrTe2kEHDxDG3t5xZwqz92vgp6aUX
0WDBNPyh1eOqByv2DnL1d/0NfNfGHD1kpo0AeoOKCnsvOLrrfjRQQ0q2t5mBjyl8mhpL3+Yriabr
NuGcD/qKKHIogWoJrq0mo1FkiGkqkc5gGoOh5+x5zY29EPgsdevbZjzZIWbHdsFWsJPEAsA0Ef/T
93lyN6p/6CUshI1uHtO8AshySMJvW+wi6Hw8q0m0tM/9ZRULdtuFzwyWbBmdRVqM6cH0XYGZibat
1s6u8iIPT4YpLUtqw3e22J1J8+vRuugHsnRka/xwA36nqhkfZlb7y/nkgOPJNAf+gwFnVREyKHG/
zxshARrMYSYVf/HgBGXDGMyOkSeefsiutX+RBIuQGq9QF/mm6Eo7Fd0gg3EcohDvVYWRkRnde2f4
StWnVAVINYB/BDKQmQ5d7bQL8tZrCwaIkYwHhwDhCbg14MmLHcBt90TioM1NVH4SWNYKBNk+Bp6e
3vIJXHzcOfdgPCqig7eW3PWPzUN+BHJ5N7sUBr6Vcgy26/AJDweaw9umy2jipb9NQPmLXVkZKyi5
pO064uR6CatFCXbDjUeHJnOPXx9Bc+R2AaimRcWehPCyikKMvRZmAM9FsPCJi7m0f1XHBD4ZzzET
5O7ySP9NRHHv3wfGO/qVDnXj0W82I6/oj6gI4fdlgHG8YIWK1jtXdYfTyylMZglRijNCQwvMiphd
S1crk4g/Mgsr0KbnHoImeO3UA5++1BXBmqzupf4rlPFth1LOVfj+7mB2VvvW61+hzkyYWs3MDJtR
2a2v1KiRw7Ujhx5aGc82UOCa2W/hIx400z4JVKr0cShDVdQnX2KOte/saqIPCdlCsaoyicqAwNDK
nxeMglGexSMxxnOhZCbQA3+cKrGFFwe7I7tEENcBdwqz9Kki8LaqRmGVWAok2pjXAoIEU3YUJE8f
gRUwmwu/5YMP/4wPjIHLhCv/i3e4wHxOnDgPQDvLsVE83QUQ3xSyQDB6VdI4AV4sOJicAihzxVIS
gKudGsgkjCth6SfCUws+MYkYAEqSZgPZaLxVYiKxLfMOtXYa3Oq7/Ld7sOUNIHDdWqQWku3UCgie
G4b7dTZCq+nyjojBzWqAYpbOgZoFJA6e9L5NFPYCcqQu++/oCsT4WD50oyMpS/kdSjfcB5KufGql
Dg9bU2D2LsD70Rrqjf1xFOXMcbrgZzMWocTtMnJg4Zztzlpi+8xu8WMBIsJ6VZ21nlgKZld4Nt1H
bIFt4MvNuWrOlDlDsYv4sdwqBLEgfhGXwcL9Cmwozd5VbltdJY2rkm5lwJhU6TOcAI0ZKF1EmVGz
8f6OJC2dpNMSoFfQrYuF2s6L8WAydVWt0w1Q/wWbr+xJRNcUkEUIy7a21xTV7lQ4+aNtzgXCuOA+
Wr3HyMric3OXgIDhIpE7xk52l94fDl9pW9YgdsinbYK+cENwtCf4iQrmpNfBzTKuw7wEwwMAx7m2
b4IA9qOpi26DyoW18h+USlDi4gr26WRoEUyBrtjk356O6RRwQy1ck6KnzVx79nFye60AssSYO3dM
pOFPAhxxAZNhXia4ataPmgHEtNxQBbuDste/AvYWdJrtUlXlOJ3Gp6cRuMvpVi/iDbQ1qtLIC1nd
UiubWHGYq9pliokHn6+Qb6Q7EwrdNoC7CspOT/0ZurV1j2Jolqd188MwYePpWZd0irDcwLigemfx
dzsyckXD+hk0WmaxSKyE/zfg8MriDBseZDBYRclKSTSOXpfAPbhBaXHpJY7PzOneh0sEXb9t3Qh4
eMcjYdzsdVqtakjsshRGRrg7VAnZXcqohqeD2WOM03wm7e5wjrlNucFaK13El6qhuoZI6+2lUpiK
btw1VFJBPMjOgUxT2dbYV9HN2sUy7PhskV7x38vtG3t3fURQoidB1hRQR5f+dTkKS46iw/eD0Kyr
BZ/jjPepyWEZPew57tmytqEy8aMoeizhi6offMhg0VreW+BHIR9Y0MgXy/WcvMyoeaSbz0RyRyEp
7zdrJY021ZGiRF158nq00TW8bu6F/whTDN30dpKQMPpCDWZAPZFqv5/BJQbqMcqpZ+EJ+zRQLN8D
vW3xdr/8TZPGBaR9PtNiVi89CgUcffVKKwBvv7ZEdZKKriMwGtOcO1MY0OkyZUbyAWvA4cW35YAR
kbUa1Yn22SzhtCmb2ceMsSX+DRtNlZAwbHMp5QA1REVBBc9Uaf84Q1yNMkYzUd2m9dzCjTu8GXh4
8FSYw4vt7pMTNhPJcW3/8SNlwvWB+72vu8FWku/slw03YgVEtUcYFyz9Lm3kDUQSoFyFMUtzl6Aa
MQFfDJ4/D0NJZnV660FnxWYkcLEqGz03DLnJULN5NhkVooyR8VSnaQ2HuRG3vh6nLEeLjVezKgMi
eDFvYx31gKjrZ6ZXU4m3LrlyzlAD8pzNw+mZ6s+9f5juJ5IZwe7Qu92WhWSt/YgU8kHqzwdoyj/R
Aj9IF8SpY2KrW1G3m/ZB33xmpSZZ4Bsbnqb7lHvmWsFoireysZOz97iS08/7UnchwPmlodFMDmc2
yV0N6VcKDzxeS9+6BLRyBPexh2CVarVmL0Xqp1uky+JmOGc78kv8AVKYgXib9xFi1di/1NUQ+w2Z
vtKcVlReFMP72fcemAJkRbrbD5v5ZIsRBA/cjWtylhjr9JEWGS6xueviAz5CIC1a1fyRgji5yttK
Ws1bBIySUgrncf6K7Dt5PiRypUZTbQgV1kxDvq2CJpYCIO6O8P+4AmUWh9xRp9R6DLt8rY9AMbV8
Zy0vzmChR/+P+qPOcSmch7y7mkR245rGNyCCq1S4/9L0rjnr7NXeDZdJu8Zr080PtRnbfRiYZxBN
/07tXP5GlEEAKDa5zDnElw+S/UIQ4Bg9JxMBRKIsuUDIIeP5tHtpc+vxeAdAZl93I5R/I8dw00ex
CKr7w4unYoVzXowJnpjU7jV1pk2ZiV/uwcTuMQzoA9v3RMpt7hjsV/flojs3kty1yDCQr/cN4hVz
eHXOCd1UZNPpzOMaDw+kt++8J4TTidaQvL56y8SshAURC1hmauLdmUw0NZjCSmBNHbIXpRASLslW
MVY7h9gb/P7gZkRrohqwQHYG/0JSeyHrtnBsmjpjfAxnM+bbpJaoAaZgb8Ko4Rvw+biV9hkjWDPU
q+7Mr8zkmewRAvK9efdUND+fhCOkOM6YneQDvbYjbCN7bocdPuQqbY36mds0sph5S1jcgAvAGN09
oQZOGwO3DL9C1wERFZv0qz6roEPwb5CcukPdiPvlLAjux+rBkBPWSmpopJx+uz0nIaEMwvt0WUPh
3fzkdhN3w5pz0hJcscj+xJGyxLcnfZTpj+BRBvNSwo13b72CuoJ7npWX+XqIouQ83bAdfpzv1fIy
7X8fMhn/PLfOvp/fFwdP/M04CHHOTM7yK9g3nqHxNaxuLf/MnXqg6q8SzqQo4yFWilQ8rYD5/l51
Ux446Y4TKVgvaUpd7vkOr3RRVOXwyxDPHW/PMaM5EN1mqEx8+SOefOv1WEkEbUCc2SGO9r9s/G0r
SP/Cy8/93Y+PbQ84CHinOJI/TcHnLRX1lgJboi1vcQdPVcpbqUo0S4eo8iSILlsx1hvVw4PmRunA
GDRHFxkbU/18zGYpmVA7j+6HxCvES6ruO31yiKAdHrZWgubn+GhkLWcLKLel03W1Whoyr/gNV2aD
MN8LLhDRuJw9x4QbM9ERkRyDZpjcB/GTxWsg+ctGJvBmFz+fFAQz14yMW9zGbjMjxsiVjHFNoehB
Qw/iajkDDZGPmtJ08iiS0/qdw/TR/h5jwfnM4DwexCzn27378Dhr2iujSitk4o5K85q0iE8YQMQ1
sTccB0LsvUvNjMe+ml69GXp6LrYZYDTg7hDbAckTB4NXQEc+MHqF4CXTFAoAODE53FlI9jWG1HyD
PsVLmeSV+g3RqwD7jZMM45LHJSOPVyPbKPwaCmk1xSmPPI2+VGL8X4GKfZy1lZyOMjsUSsqU5U6H
GJDXk4+CQXO7Gc+3FxyvS7aSdDymmA1hlfcVTTEHW4H6+w8LPrWzEImniBS/2QNNqBgb6g2M5qo9
jXdfEDzUuEN+xFg56mf03ZsTG3T4W4NTXkkjpWO2Pp1w5UtxSMzsGtWg5uzPenL4QMP2l1L4COrx
2U4ERSjnsU4AvH1NqH0iZcex+ATrWE+IInuISZnFhxgHX6ENQnZxQHPhnHsq+3K4pOJ7dPWvIeHY
SJQA3vVT4YEg8WB3nk5tZ4fHbngMtthjX6w22kgWZWjWARVCMp8AWKnRx8FWlqD5Pyh/ASBFyRSr
b9qJ/v4g3nKMdQAWKZN58l40jLhQG4YFrZE0n1QpG+ky2yo3IN+Y9Z07EQco1dhpRcawEQD5HCnP
1+50YSBYvXLs5DSWiq9df22ZcNBsctJ8aIhVJgKPS2HaVD188ilh6/SbScACG8/H6eBr8E19Vy+1
3tW0erN3Hfk46ZVsh6/bT4DdqA0pvFl8q7Z7eyek1lY4wkW3Cj0h8T8iFLwTx5PV5QyYwwOvu3Ha
0GX1a00OvGbPzRLivkRKZCti/w2OVzYxcFM2dWP+M2QcnQB8vo4RcDXrW8pIoAdA0qsGDhZUnfs9
PZ9bJSPYIDOkYIrJ97i65ZohfzNjGFul2UW78/LTiDFrt7/Wzr5eqCsBSRRS4QPnBPuxERlNXz6V
aPk1RnLisKgFNt9rCyVKALtbzlN90P83SwPgmYMse3NxcV7NMaXQYwdgrBfMz9eU+NAVvhLY0aS4
rILL8I59yP63ydtFtxGSLHFE0SFO7Tzg80/qG/i7K+s+sP2vzxoiYhsrUYcCp8gDrOoefeTColP2
hAm9H8U1tOorJ5OAzDOsziuEjnQd2TEtLf4qcScyQrmq3vDcGSdA0QaGeFA0+9ON7XwYoVFF7rk/
JPr5ktlCmCBkYosddNWZWVrUnOwDnNW4BNpZ7l0Zs4imkRs+egPU4GS+CFBjokp2ksV0F5Qh0rR+
eO+vno4inIB6jte8NOId+1abql6OjlP7R6YbkrTuCpm5/rben/WPHjGofCfZbPHZWIo+SK4oJOL7
R76YlKnz6ejHfGXuUqepWfDkxmbmyrs7qz3p1s1LDmXovPDGr7gT2MDB3wpHU0Rm72K8MH74Av8S
j3PTH+BABrXtK8PZHoMCT+Qxj7P7b6vRzQ98rErLYpGv8s67uivMKR71H1VoPOSuABZ0zlTxVLwt
hDmQqUmjjVcMwMFcmFYdQaz8jFTB12cqPt58OOxxxaRy4qRLP1Z5OtZ+OWgAuvK7KEGoJU980TrH
5/COZk4spCpFZ8uFEsCBLKew49bWeYtK4MFDiJdVu8KGXnR+mkUk3hDXlZ66g349580nQQv49tiM
ZRjra3GdeDIQa257txgX36d2dCtIlFoSPRhdz1gj+z9hTr5BfYwns2ABmwUstodJ4kls6M50L6L3
IgJZlYPVTtlZTHgFH1N4VUHIi6TkjCaCBGtQiRFAATKJsqr/IOqdVoqwoxDRPjyTgA8Y5CE7Ymmq
MV/BKaHUkNk0mg2U3e1tR9oEEVyK/o38mT1jDhTETNMQcneNPVNQ1q72vWoFIYwg+77wb/9+49vS
CA+naOnk6OkRAImvl3GPoRNKj3AZyEBSgEJFlqq6fkaTWb7+VJMr56CmHwKNg6d/7UVazuevKVcZ
oVYTRBi996rm7g27M3+XP2qZrMXF4TWJMeo/J3rSveOOFDqunpS4MDznt5OUPzf+EiDi3r+5Pqq5
ZU1WoVk7n+iJ0aG9ts/4Rhl2dI3EFTYLtIQi32K/GrPH8GHqFZTe8OLRLo/9bJusu6NP+N7XYrGC
3ErNjF6/xSFPezioyPanhcfkhxxfcBUBsguSOrte0X+0boh42kOEGIpmJroryIVTWUgSaZtNXL2b
/FTXWWsf+5dYdipGv2w9mtB7+myKZ4JpYOGPVu2bysyBn38qsT4BxuSZY6L/boYpOS/67iMn8pN6
rcA95DaSeAYjA6ftIagwQyBpwIyKDrMJFgd9slCw1jW40uIydG/IsgaXv4VeWd4EomQp8w0fZL9h
Gyj72iP5I8YG2bVEvGOq+/kQXGz28NSFXrhFN3MlMie3pIC7/dlrnWyCYAOv2MKcTaw5pGTBJsMC
wl0i8XQk12JH8S4eBKXRVkrUOJ68AfK/zjxgRER2GxAVGFv6HO9DHKYVxzfaHOCwnAEpy3PoXabQ
H2rL73DtZis582gw7+G/UtVE3VBFhgLm7xvgyE4r0ZmCnyh37iCfJMo/UCSSwzuvWpNY08BuZqH9
ABGHGsqsI6FHdUj1COxbJefN9o5hK/33LCcm9ovuiGHiuB09uLmdxokvjiwbFr7JTQfxQkzFNx6m
4pjBFXLqiEZD0URqhgL10URG4/gttQOrOj+462JICHx0Zk83bBzeK/UvVjI76Jy3PHmUL94pekKT
5SfY5yQhaYwLzY+5MOlp8Gy+GdrvEjLyxGJM4sCUfGvlrvshkzWp4V4hZ6aFeYrK2XkTO+4weInD
dlfHHVOpMvZrYYR26Gjt2vgQRYHB6r1lyFVV6OHPuAixPKEyeGCOioREBSXlhCm0ziO6WkqhHErl
Q8sXQ9isUVtaWHcxGHRLOenJwP0D+WYIqR3XP+ysYO4NqIuSgkE4HbMtcIfvbcg5wWBZ51FpJu9O
8bcC2wGTZAg5xnvojWafrLejLyhaovnVnWMg1+IPXfi5MkcJc7dis1d3B/kVRwk0TWPeiG1KAMOv
3zO1Ivtq1AIhZvbrcSHrsiKPb+RPhdVmDpdkgOOyoPKObkEcQetGq2fQ0AdlQzl4396Fe3tsAwjo
Mti/6UYQ4SXcOk4Ssa8drIRq1skSzDpLc2EDfy4zWKtOWAiwri03IGxl1LSD6sCUXX3e+nAMb9lF
S9REJJZVaikP4mQpefgS2UiTpDxf2OBjHl0lMdMfsVmlBCS4ghIi7hTV/a8tGlJqUiJ4a3uwyTwB
uL58bF+k5kDzCSOl1jByygj9kE86t0CPEdVQGjXvAsjjktB6OtSw7mh1UaKrWXA8PZiGw/9NUdsn
hSpCV4AcULuSst5H/NA0Z+wS88AVuCyIPBWaH8uPYU8tDThuTZR0wuDpeBO9Ua4hupnBIteqSJhI
SXeluyBM7+umYTUjbH9uIhD9RjAJcyYLpLuB3Xkvc66HYtz1FPN1wTrWR+gsRZi7R/3cOrqLhvwt
29MCK94ClegxjhE2qGXrT7Ll8rtcPLPBn6KaOcG+u+rS8c0Z7VjrSoovxBL8PgY16lHkcfklHowO
ZSFaBroD0D4S4P3DI736KIjvaGPOyDfUIauUZX1CxSE4RphdfDyLxVyKjnXswOlJaqqmjZyAvfll
mhiuENE5rjUeG864cID/LpG8tJUm6RDWQzKf6csy7HkjjPwTNubSaEskJpYQxlmYF9S5IROYMz1T
2apP2hLXfqrhY/74jkdI0bN2VjimAK9wElY5mPhv8mU+KbGhYxeXjmaplzG8RGIBDMIvDpImrs5n
HcPblqn96lXQuL0+tSC9+sbZR3DlgIy/BEMOjdWKttG3fSI2gUapxPS8FY1G+kBmPnhdTiKf/jNL
ipD8RXNRp+D/lgN830Bq8zbbfbGsvyuHa6aju17uajHcW8B3Mw6fCDab9IURzDgpkhMlgWO7EHWh
faIuzrs4l/ixTv5KZZKj5ocvcFTz5JIgI0ssaLFKNEzzl0uYlPpQUpVaZ/HD+UG3xYYK4nAsSSZD
V3rwGQHOxZOV2Fd3HvdX+9o2SiEicuLGJ7FFMpKfyiylVrkro8Fe2Vl3QO4J6meLTnDBU4kd/581
QwOAIjd1uBuq5B9w9ipiX639HHc+VIGeU5RNGgtRsP5rfO+g1wfkRBGobysQv0YRP7Kk+Oqoz715
xtnja0urOL3UV4m36MssNUGnJ545RRK+BpW35GKVKYXkO8edbMSfQ3gf6jMPVf/YMXETcL5AkIWU
EYfVc04M8QQkZqPWGDFwlFAUzsiPsqsyvWqIjvtuLRHfY21PJXAnw/Q9kO08cPtyM8s3YTiy2kIS
IPAOPAinUUYi9GcLleXAXBmWRaeE9HhpH/TQXf2Jl4CIyU/tr2pUgo5OEW2WuYq2YcW/MiE3J8Mk
+Hzen9zsfTq4E355SMuhm31zEkFByR+1bYn8U/ryROJsuZMRyFsO2Nt8AVCc4gaJQI5N44GCoN5I
9Fl3KJQXuES3N03PAxK+BnJwBpOBHyyzt2THOdt6lr2bEub2/BSrmi8g5yCh6ALOwGCFx4jYReoT
u4bbQS5cP5VtjyMF7cMOlufmmTSLTNbBpTxwlY1Jm7GVWPQL6CJxed2VYypeVLdrbRzqYlPsRsef
alzSu3nsPALYlyhXNQ+fLFPQ9j0Oox8MM5ky5VEdzn+CsMBnptiF7FVnvSYhyRUksiLVuaQNlauF
NYp0HfNK4Qi71QOLjbYX5WoIXL3QeGhMpnkp2CS5gpWFt/06dWHg9/YAwhVMu9Kvdh9Jfk2ZZexV
8oxNZT6bKhNG15oCuaByLHtAJlYC2EseJAWTBd4WvotlLtE/BiNF+7caSIf+CBpVMJ7KtkS6nAza
mzCTG8pGG7kg3d58FcIu7g6y8js96x2h16aA3WSrCTnTfvIyFiPk5uxETHg5B03T6iMg3D6HUHvK
2YAtdmaP3779fs/L4TonVdJXDfdLluHz7MIYx+O0mx3D1W5A0Fk62wXwMe0tXlVWO9PBy2/n82uI
MhkE4ZZZ/W//BRfJ/uZff7h8KF6DaCSKj9YDdVmCQMpqF/1X2XYRJs3DhsVqHuDE4W3SQ9OFL+8d
+EhFCtKOLdkAjcmN5Md+HQZDbSqGV+RlBZdWuP9oN1mI9MWHllQS4PChVF4vHUJEsWRI3UYIAzfu
67HEHYyKiGTfmqLdIqAWNObiNV7MQCid175wXqAmZk4IbQTduUwz9X0KHFc+MVDt7Jx/Bsn4/RvM
eo5AfgCrScC6ffD418AC+K0sfZ0vBE0xElDzMPuOtt+SlBiZAZEyApLA4YHkVoaHhscCOLmR3ftv
IHVidgGsC8xSr6Ttuomy1/YkV8MhTn8q5IBP9IjoeOY2s3Dq8poDeP7cHA0RlDFoW1LkGpaFNFDa
1McerQuwucKBdXnhaGQaSG2fTvfObv3vMDssTUoYFLyQ/WcUQ4HnQb0AFXJn35ieZVnmbe0BOMtF
dZKlD/g4sUN8xkYXoIm4Tim8VkmeW50dex8kw8Pa+Sv5bnUxmrfYZElzq9To7yKTq5DCTd+yMK9R
dIw16Gmkg3KxYngf5dYyC71bREc4h/t2O4p0GX76hlH8dTeOlJEv2o9yQqkzxmJq1UuD0PNU+qo0
wQ15BN4YkxVoHQAIcOH36DKQ66sx8WN+riWiCiT17eV3Sstxvo0QjhCWNmrrfFwXjtn+wdsEVJtG
UKSq1UhiOl/yoHtmIm5D0qd34b+MPX6Ttl1LUrT+31gW3azGj2tvzH40mU/0Uky/kSwKYoJyqwK3
xg9NwuwLSziqU32yoahlTLThdPytpK00NEIJqAvXZy8vvaIFflrbz+sBc/y+DQsBv0XNXH1m9dtF
a8aff7Ga5aJEs1bRvzTP8TKfs+kfmUDPpPzJ4Klf43qokJ8MvrY2WpT9SG+osf5AXsu5yvakEmgm
COSKoNqlW5WnDtYcFe6sEbKugSSqCwWxJnb4YmjxCpWQ/l865n9uzi/aR1f+KkYGTRd717OVGEt+
kkNWIbLdGIWM6za5saBRo1k9i/nf6ZfErD+h/e/Tzu6V3oatEn5T13vwp36KWFnGBSsxJ8c4NqGg
2Ntas1pyMl+aYNo16BtIn9+ivtA+6B3/V9hV4x0MObOgUme2ApUBrek7PUyt2EnPEj/A4FyeUVMZ
sbaoCgnDTabHnVeCK9CBTIpSRrEqO4WXrOsHyMha0zZPtv9iJSRoX+H/xXNWCYql13vFLI+0rStn
+3CTMyoLFljN4wrQ5F5RSF3mFyLGykKe8vFASfXL5+jjithcC65BrzA3GWVA//FWi9DIYB4UID9O
e6QQbUIL23w98u72PL5aGXBVD8u5eOXvcBZ1NXI93T92uz+4aVmKg2czqzGkFtEllYjjjcuxxcOA
tajwH/k5PpAzW04lFZ1tbrr4EuUMnLWlzx3/bNtMs7mweYci/HH1KehYh5ph39ov6sAp/fRtWAcw
I3XnMtIb2uLXy+5nFg2xxP5crgOZQFFUjBpnbSqT88bKsHfz4yKXQf9kgeh7S12CUjGGXvIw5cfi
T7ijdoI1SYn+zMDFpx+2m2RfENtTVvR1mJ8PStt9mjEQsOjIoA/rDGPtxiQvJBlXoUKmmv33Ns68
pRDe8TFrR0XVNguqPex1WYpUZv5DTucFP8SFMaFrY/C6exYLCEzGR7jXZ9XGUiRFqrxMxX8XehpQ
5/bUe+1TnN1ncirp4Tig+St7SfSRcDhSMuybHwoPTq8l8ZnARA54w8GRIlaxyW8t9RlZ7jQ1MI7N
YqePk36Cbhcgveczv4dDNHylJ2ABSDwnGUv0fD3FsUWhE5JkuM0Bt52a+qv3q4cD+laEYGM1dQ4E
+2rPzoFMe3kZbi56pKJm84JeP7opA784KVuTRGImIyzbVRWrOY1NLJwjQ0wJZdBRBtsZsJFBS+dp
b9DfCvHYEmeqVEGDnGaU6D5bpRbKBH6E5bo795WMdXgN4IkXNWLJ9YVjemCFh8d1CKcoMQHipQO7
YEvHQj5nVfsS2FjXhrUEPEAk36TRi2lv2o1qQj+mYcS8yVqJWY+JRdaedY2jIgFPwehFg+o63sBT
yM4NaLOpphKy4NuztqMGK4Ohd561CrLhqKcxkoi42ZpWJfKP+NA13qZlbzQXatGibu2buUknGdQj
lbCzjTNDwT3i+oXVuVu595sm/ceRUwXXoNupPljDnOfVCsqJNJoQQDKAe8IcNEw1a10I6gHEdoNs
unJozPJPpuAmooxyRAVZm9mGQl52pLFO0CfsyBLKjbSJBtVDELsMtAZp3FEZ6PziUrdHvppaMGQ/
us1/qu5SDLquAubE2nbXGMs0kzmtN1rw01MptO+FKFt06k5UxVF2l06Rh0yG9VgrKkzfMuF7PS70
/6zBucPMg1ixmWSOsfC9fBiNEffeEY0o8wT5HIfrvkZa8YUkHnQ8t8rpyKGaxYmxnTW8Gg0Asf/S
QBgSAPf09oIYEHrLHUcSN4T6gbRI4bQPPB4jNz/AD2OEouiE9Uv4VVkCbOzr37t8voohVqNZ0Pi+
FBjMxDyTIS/n5KSp2RzOMZRHStL4YjBjJRTCWFfT+RxNwt6qIlomrLIDjqSTTk8fMK2iP4JGZcVC
rHQVd59MglgQcG5w5Qo0BCowGKzSN6uhrOVW0OCmkvPrCrkuU9PIb3jJWyl7Eynd9tH7czutbEyY
pQaxoiaAwGBfDO5vE2NyYFFIxHc5GAhu9Sa2pIRwDcXom824ZPfAHrZSaGozIxfOyB+Iu5ZQaiHA
DrlF64GjMZGgtR9S+QyILRqXq2UzDzW0h2v0/mF76j1lK0p6fZohyzlMjQSSgsuW27rGdmfGDM0g
U43pSKYsm5f/BiL0gJpsksoaO8spD5nfdV5yHu0m68dm8BaehmYTt5vU/y/2PanR6C/8yi7Iu0Q6
gxv4+hyiiRUkrR+Kk63hbUU42okN3R4v8nMbqICi6Z1GoVNUpDKY+jXQJKBBmmZNvJMOYE7seX/Q
CaPiSlfcFPZszeeG2YWEflnyiEdD0wpSx0Ufa7e31aUkh9Bdpmw9U02+ywMDe6eVg33h2zCG/+WY
RSDHjmPggRTBEGTx97mkdQgN1acXgb/enhYOfTO2ujOIMrnfz0h8Xl0V6kRRzcTBxXpnu8Fzzlci
MoqaQRMW61+oMtwV+7KsGK4cHHH3Mxzb+wPCK6jWJT/9/wtoK5IdURiSPfezlvvlywWxrEYULSbM
qBzMm7rMG1HptPw2/qP5PJXLR+aorMFWUc2gwGtzAizJ+1j5P+6c9u0CFIxJL5XHMK+qybFGv/cs
OnYDGOSesqrM+k3IO74v3vBfV662Xjk7HtDNFfAQyxgzjSJ0et5y9V4E0Tp8QYjy5yYknzdc0Ume
cAw9eb/z33ej2gb9OCBq32QaV4hc4Y9LAqdB92qxdZMXt9rBaCznWja7EwCrCCeFiW4FlYK26fCV
P/C3yj68e12YAejZVaSMcqYsMPNZ/kLJo+svJcPtB4zNkcyXHy7s7R181pQ18C7ZrV/O8GpTGazz
hF1izSc72IPZyZilgfWwdJmYE462jVRmZySuB4jgplzNu9VnuRtox3yhBQmAdDCyPfI3fmR5sSWW
Sur2uazCJ9cIAqK5pIkc6MuMxFFx/0pDPuWvETGI6yyAJ1IEMAmjN83Md2YYexdIr8sqUDRY6FvR
9cXZzUtNjWQV6/mmfNBVpujpd4hWmgdlIZ2HO0aJa9pcNqyytbv1j8X3Cg4x7IJ5u2IBrJrYq/9F
RnElNpdwVKwcd6MbHxkdR86Y+ekNpFjffO6EN8JFPPJ2oAOoZG7jSsBzIL55/GqrEDhQBdlZk8RP
c7xI13Tb0jcCoVFRO9p/CGiQrwYt52WWAAEvexgN2weSxhHKsOeQRDWukbr6wTIwdv8mOo8tK4SQ
AFhPFLnJEYWu8qp2u/K7H6hO0M2HcKZU2QSszwMWpzgJx7I8NFC62IQoFwnMiBuhdYDM4glEvGsl
789EWpM0Z20hEi53CqoaGSCiQfNIaMYHDfnm0Hs/H1j5qffCop/HQYA6kj6Mn4PQkHQJtgAxXqiH
gI0jm5J7ZGUMK3sSnrhWyFWl6UGeROxrL0ie2K0SttJU1keKKTfx2zSW0tEGF8uFN7egpV0zpF85
68fTw6IwspCedyNf3CDa2naA7JZSMCgQIwYvl4LuwePtj4doZifJClTX/bvza2/MzdP1/wWtYtSL
b7olYp4D/efjUNIkbdu5+jUL8G83g4gVey0rFPGTpMHFZINyL3FrJACLzAtPC7Q6mMfgB9PvKz9H
z/52wLTzglpl9lzUVNwIBETnjoiNCRGVcYIy8ERAn3sZTPPO2bW6V764W6jHX5bgVaOE2FgAsMm9
zZBU8IgRXl65Sy94dynnaBuDAI9agTSQcQQ5T5xh3tt2r/oSwS0JEGLXZCDHedrGjFDTysQqlgWx
/fhvdtiUb0IJZKfiHfDGB8WzYhxXeJ6kDEadQ7UxMzauGhZ/5wlXf6DxgqvJKD/upJfFXtjan1Iu
pN9STtC9bNCGfUUDoMEWFOdfEg6emc6p97j4pBaPwMAa9bYCZR0Z03MsKh6Am6Qwim5HznkjqgSI
B+/f4WY2x+brknIvNHnYhynq4v52uFOyQXMUlVb+JfTIsZAYqreo1YqLwKAS22u8hmEKeahco37V
XtjBQa2CLsxZdwGbFkrkT2oevAldmT0Wb7YJ2GMIMVUIfEon8ZgIJg01PUMEgQ7LfckXjDOz8Xbw
4RpiwiI0gH8oeAMNLadVKIl0uNupew5vv1ofkxU8dKMJ+Q8v2IW0riPCAEspmSLp1f2r6ejCkmSI
mFE4Z78BGz8oxRBP5h7KKD1gs92PV0qVAjRzGj9O6iXyXPVc4cP/s5sw/vjp7+LknozlJ0amtAhl
Xyo5JCwCKN/nzQtIGTO+GL2KhkUOaGZimzMCbofvxgTlcZbv2mvj6DhFCLeqSDelP3tASzQ9GuoD
X0rqwkY/vghJ/RrZH0zahBSRX9uL0827UJhCyS4W9NVfslQ84DAGUnUoUElE/QtCSAZ3AunrjUKs
C/PFYHKpWMPPY4Utp7zzuUgN3egg9Got041MWQy7X5/NsCmwtRY6Bn7GCcsyh8Qv60Tjm/t9VyYo
kWpl45uBxxNc4lf49URZkb8Xk8tGiLMDLSYgT4AZwp6atvMTyqJq7dMpfQSvNBg5FcpSD8GQV10Y
ANIca9z9nwGKWHTxOL3S9jzRnOgyzXH4JzA8RCel9yD5RBDsdUufSPWB/X5fFrESGI486x2OO0h2
4ueP3j7NaKxPmYT9cpkdznaTiXGTv23ZHEZVoQkHUn2tdv9BaXutyz77eqFUh5n/Z2tqQxUxlA4J
tK/ShqZnNmF9yMT8JGtf9UZqwf/OGQPEW0RmgcrqnK9xUqeDiLESYTZrRmF8bNFe2smfDLjydGMH
WnQY/Stshc+I4IVTJKIpsHcJPyQvDbPyXddYNtNJAO6eqKW/GrUPXOvxSiGoGB4gd48sOl6V4Noc
FnE78ViVu9ZdveKXhVBs4Ms+A6j9Za9PVC2Km3ie6ItpSDHHVVoRnIKeU77L/oNXR7t5AhA46HS1
megikLWA4Eh0XH7TqQedd5g6PrkJQgkXkYnklLPg2dQk4V7dQqutUAmPbKEK9vhpmc0K8N+rV5x3
8FeVLw74f1Nw2cEkSOMAdNxRysvHEK4X1ysx3feJkpQ4Oa7r8YZZ9D68V/rfKhzeLqyU8cE77yrq
yIU5qhY1BbFtehGSFdqCilUmof6+dPeEEZ8BTNJ++WzWXCWxftupVbJU31j8eJrXb3sUH6Xt4Cya
bQzsXN+6FYWvhX/viVB6HPx8WbtvvTQUV2uq3/IzW7HEk/6RKyR1OhS3Q9xcBoDXNGkdi/rkMLVY
e35IYhHmk1WwRj6loGChevNsGsRcxDT57ui7pw+w+U0Cf8XMdtC2wvj5anLwIkhYCbMFNtfuaU7/
E9MsUFc10VNgx5rduJRsCkC2Q6ao7O0XHJeodVAXooboWEC6Hqab5F03H0CbiT0b1GYtAnapbzqG
dADRCwzAMtBv4xmKdDvvhyvAILewvIsqPOkBs0Lv+KBSWmYDZlnrVTm0p/jgs+/doeAH1k926XyO
Dto4CkN3E22EuT1kKSnDMBCug4qaDAcD05mGUT9RwD5cyvTZxv+7Ga9GwJgmLK+8IYTwRp3gl3Xn
pmBMSsWDIunM01U1OCVj7vEU0fbljPrC9pSQT6cPNr1Wc6dGiDA8a4wAGksIiId1sOQ+1GvPVudu
CKpSWMESbrDWlahmhdQlCCPgcd38mYPikjru+RcWJ/DXU3xPl4S7y06JCQNb6FA50FcuaAg91HwF
YtY7tTc9wSjk8cYGFsg+pyZwu4R7BUW/8Jq9q2BtfaByETJkQvTLW56/Vk/AZli1u5qWsU6piYeo
qNM3qBORQRJfJOfnVMDmUpRTlHcy2EVMiDe9Z4+MV03niwsOkpacmadLIFTTDQ77E09EDsefbtxb
58K3nyoXzvvk8uvAtgoyvd5C3xCR+8z/B64mUKqF68efSaWJ6Tf5Q0gKxYUsTSJBggLekIRYRvm5
ooZvKI+zxJoLZSULzxbAhDytPD1oRfeptGUjiFWv6+gbo+AKSG38HS96FRtCE7FYjpzPlUMAAW2N
rj9Y51h787kY08yaxE7KofCXPeojNLKuZsuf4HKmDXokotShPfCBmbe7E6fGaki7jg1CFqtKoIIg
r23uXmLLZNUK+9DbauNkL/s2lsYIT4rd+TYKQ7Wk9gJL3fI2+e0BEmeL+uZRLTVM1aYfiCP6X3L4
zmGT00xFXq7H1V/GRcqHjuHflYtULMLqLS1ouQN1YvBZYeTBtb2pUdicffk57nOL1mtlO+7ecTKk
j3LE8FFRJKl9gUs46zXKCqJ+QD5qU2grprk1ohAz4QYSrCc2vHupDN6/afvwDXJqWY6PtxKpzkVc
xiMgeKUsxuH5IR6mov9E1Gjx20/JH2Mx1aVkhplH8FNt2uVIzMhwcdcViFELgzQYuwpjJs0ADRQS
IFf6ws/Fk5Mf2QIgtuyGYVnO+ieOpLjuF2yhf3BiI5Yjuct9n5v6HH1MJPdkeO/4+j7EVpdTGA0O
Tj9zF8uTOpE4hcBy4En+tin23F/hD2CEQR7Z8Jquo1b1x2GeQx0Szvj3g9+k9voJ7tAHQUDRcDe+
qi87PFlP0nac7Dn0uk0178+WUQjJRFmDVWzlGXlBkBdaDuvO4UGXpPZc+XdE3IDmn9v6W+3ocq7F
gjm0tpe7OdWN91p3spTzVmzlm9yjOU81EMPgym06Em1TARovvnQC2PVThSzIgSvUCyQpZC85fn1J
p9qauOMoJ9orf/QUkPr8q2IplizPZgeNKmgpitHhJz7dvjtGete5tisT69PG8B2kfPB6wpu/MZrE
M9wPc+WL+Qg9j/J6wZquFxzlqOC0mxGZo+2SSW8ZZ4xJyfMakNDssEwaaYEuvUS4xCj+AbfULtSU
kgt0shgidhGt5XDsVktgkEgrT1nw+7+kRB08ISqWQLBpB/TV5+Vjrdauxdaoshv+QKPxQbFiQVeu
TIbIbLeFJFsXgNPyJPTTEpSWi/bhfhltDLWqhnmCliGd30LP2dCuQ725DmEzVcyPOPzVRtzUnjzj
G9Oph0rn4v/hlUizhVyVZkaxoCCn76dhcU9yFgCnG1Q8A3VkdCCMxofl401CW2OpJRcFIeCOCjE4
4Xb/6gc7BWZxRAef1/lEB6xkJwpoog0er0zJAWBmTwZQJysi5xAfI+/dKgpPONhFo9qRBLDlJgRK
TVAQq9g6/1zvOyWNXEt8PFMKkbZ+6O4ZAQW8GHfim/01mAw40m1dGyKdIiWmYXXx7njSQUxG1MFJ
/smq7aB++KQx1rAu3W2m5ppWQVHjk8ID+qQFUzxbR7P6W194kD0YtSXo6mjORX+RgIBSnqtDsZZL
iPbXOb9Ri3/kGJJENGwPsxweTz3piMrv3Qx8ml792hVzdcLkaabqefBPMIrfNaM2LaGJAuk7fSL+
Dx8bBMu3PDHo4mMzAJKO0zrrgp/EmJDQxlqSqGTQerJeJrkkQQVB/6kddZcESkAXNOwHRpBjT+II
uh8DH9Dskdf554yfUpGt1ODpy0+651qH92Lbz3tCpshNaAm2bMA+8GUpIDLsuZZHbnlatHNe7ElI
1RRmk2uh+Gsn3JRaU5eSpBu2dv2BvWY6nEsL2tnZJ1LDz8XMY27tkEOqcOPRmrx7JgahN4SCv8pQ
K7o3PGjxyGvmXtJY7I8tKn45ehmOmoV2AVIsx+LxzzNhO2tLlEgyia1A9VZfwfpDkT4Ijp10c5T8
2a74XCKqDVOvxR48hP+a6e3lK1P3/zDVXhDKo2iKsurQ59eZGMIblV7ZPMjkKyjADXGtKxx6HO/6
JA49JYXZbJ+tRYIeMnCtQHSOe+uz0jrVXiY6cX304zW5tRVGevcUtWXpcL3uYDRi0oEl7n/dwoCJ
tFRaL6MDFRdUfa5PCoPudRTYRt/OVtkTAR9Xn1LrmxYRXSi0ksdhXCy2r3QVIkQkB3WH5OjIhd78
64VtV2pRVo0mJD1/pPCXWeA3xJ9ub7U0nRm0Un3CjhydNFGs5nAgl6JapCkIJFAdGKyfzmMqQNYW
gfnYyLs2VrGVM+IiciQ3R2EmOno1bvke9ibMeTaAq76HtLkej2r2maB8QdYulyEoa40D5sofLdFf
JXB3YCZIXRIbmJ3CgVMl1o54Fe8uODUO07bDHdKojUXLEFvG2qElwC1OjsVqlh5lrTX3olOyM3VQ
yVN/HuDFqVvhYM/0YF572ZfeqBc9Gk7cHdfVbpC4Qm2Su5zI+gMbqmckJ6atEf7EpxthoatJ2u+t
S8a2G0gfZCy8HcYpZajkRBRzKKqLN0QPUHht8rzb2PLEXCJhskqzbcCvtCTfDNOB6MneIDWTJHpv
4yYuMQryPE59z2DANfAVqpd7HATj+zopIAA5GKSSzlYorDRpUcM6XTjjIMZHXzvgK37/Q8AjI//T
rt8pCU4BjNKhwmwnanaP2Kvn/U8En5iJO6lThEuWql2iFv6CgKD5LzEHS8BVHencaaVLoQaIQsSq
pwS9RzIGw7rnjslIiscZw8lE/YhjXUDWYsQkvf/qLmUOSlwiR84UqCc9NaTRHtwZFnIfQL+J9FAN
FLUOBRJKuH4/Uu4aLjAgtjKCzeYm/MQNnioYFcBlJkNxXTRsERm7BWCIw0U3vJDnBrGAoG7zRDrK
Xz7WZTZKJab8NYUHybZcgkoXN+dN7DbU1itkOkFJg0LCiXmSdRGqLvcG6HMfsHMDv9G2G/Pg5Zxg
SxfnV5+Ur+SJxgvcb+YCFEl2bTy5p7E5+Wh2JtNZ5oPyaW4XNCfG+hMsJEBi8lhWvn3Of7ao5EOB
cGdHpjTheR9RWGnxuk3K2Pfmxz68aGvbElV2ZjT99qMcVsGdkppmuRic7xjD/GrU8uWLnKjVsyvH
FraRdIFSdFKfbafRVJ4G/L15RfZvvCpJI5HnyTydpc4who8qNqEUL1YCLem6sLLfHAc4zCIsWcwR
l+F6xDdWnZdnr8t7b+78x0OPtGLXp9VsYjNIEK8jz8PaASoPAV3pPb9+PFbWCxQdl3s9NUST08L2
d9JVjTP2xr15TRxXgMuW9L07qSMgB/nT/12dBQ2GRMyBv/8klkMB2PRtBZYV9rVSadzOnoyx9XO2
Jrlan7NCQ8x/NhdYU3Es/h4oKHnno/vB7svI/p5EPaKUoF/jc2uTej1loTJsiTH2V1Kg/NH4OwP7
qj45I+Xo0+BfaW6au0JGjzYWxnfTTck/kV5r2kA1Hsw7YXpXSXc4OrMg2DP+B3rIqaWc/izNzX98
t9WMhvgx4Ntkd0FlqEw/7YvCexGPyP7wFrgAyOMchqkclD4cxlM8AXFDwxZUDrxmt3tX/4Hbv49n
T1QhoRlcmgrM+etK/ix7XJoVLaVbB1vIOMO4iDnGmmrcPO4BKiMKC+HBUpMOKbDLZitgV9/J4edL
BvVzEFmPTu16/6e04K+k8l59gCB9CPlqvuXWUGbjkf7vG7vnykh7Lod1KEJfn9JLeU1P26m81gcC
4ei52hoVX1JaKwOxVaFTg590r9h9nFwrotkQ+cw1fQ1gZRJvOpTIGM8bH6WYu98ENUV/7ejrfBoT
TbWtycQzuvrJ03t5EOFj0F3C/4Ps6ci20SX2AkziMxQq8bEgzR5WEKA7/0jhE2RjRbBhtZ5dpJx4
wsgRpBUjf2nI1gqPTGKq3qtLtJQ8qoocou9eTkp+sTZUmTGAuIhQapokWbn/sTvwLvuGmMIxJZ89
8myuL3jHdy3r5K5RhtAp0vw3vZ7NX2v0mKvEVMDlR2CLN+LzdALptHFjBQ3urMwuZkAcGqxlA5y7
9BJt9ISDvTUKgXriS/hxhZwDpSCUnTpOSM6iXLvRrV5UnR4oPs6gUE9OXaY6cPFHA6smVDS3ETbj
9QSuPvRXlpYT3cl1a0FkvXeCawr//TfvBOPDwgS0oV8quXvVf0ySDHyTmoE+LFnZnrhZc5hD/naK
oHSU40Eh3jCphlMarb2DzUbbivbnHyuiVR2W8nokYbR2hI4mhRYpG7Me5H/d9XbjwFk1Hex2Qgu1
KISGKSWCxmMkSyTDw5HGijMGpA1oBamEqhHSqvDDRwPtqlm6S1UF1aQSwm1/L+4Jyj82FiUZUUjv
ATFQCocU1Nh+IuIP8pmzhOE61p1OH1H+lubT2NCeFolvQbiq5Mnp/+knGnt7ehkDkH6kXqx0K0no
js5hvltUHuw+mdX2ni1+KaWlVaeb/Fo30T45Eaocmh1BIpLy0Xkel9TqIoEKS7EiLRgND9GT3TSN
ELzDfl0LHXYdKXyr4w3LHOdsbCplkMppXmsy15oyEBxcavOqfIAr/NKSP45byMpaLE1qc6AD1IYk
28khE/SbjFqceZE09uhFzdGyzj8GeMKBFeMeYe0rtimtZAsNI1nwT+z0bhJfSbnwm/zzkUzTui0f
sxg+oPyiXkVSgXEg/8lkXEM5+C06dCVte68dCFFi+tzGsVUC1aKzyOcpjAg4IC/PZD7uFbHYIx9j
AWZClAcb8iYZ0ovdwCHJkIxWjLlaECm4XXZ1KKKaeQKdktB0XVSzw/xa72kUd0gaLPMXRaJhbXf7
uAOENy4lOhngI/nVomkLTKjLDd6a7UZMKp1PYxbDwo4N/MD162Idcx5Qsxc+8XEtLCl7BMsUMzUw
fA8uc3w1onWvjgBM5Lbw/IsNEyqsHT/CLCP0cl2+pjZo04xp0Ono9pOVt7OvXdcH4T6me7fYZF0O
Rn/YV40Ri/5vY4XWuZSiTU1lYRDjGuQORXJUGrr73GyBCGPQu35SC4iz8/oMf3QIdtlmv+8H+7F8
wl9HC7L+ZHx+Mnl7bg16VKS07TsS1U6TojNzB1cB0WP7ly7c6HqnszuSU4daTOMPzQfSlfaxaLZv
oj40MALLdlG8mnRsEvwI93BW0XjK6Ui90LcrYPqSXD+XjVeD/jcVATFZ3Pnj9/8Vevq6VgnchGoN
kH21McpU+hQD6LjCXmwGyFpqXJqJU2pCVPJp7/M+WbaCvgE9yakWIpUDorG+0FCe4h6cntEywMhL
kyD/1ZphxTPiGct7arp8MPMC1esh6RmwPK80QwcSPkFXNv04lzEiOe0ZYXOWuYQ+MMRCtOobfpkf
3ZeZpo+glkWJORcM4FhFvKwDf7kBc+Ht0t0/1fSfRR2+TRnoEsvl/DXl9jRnR3aPKYsbLHbyScaR
EB2P75FHPOeIY0RjGGdStpY9E5DWI7ksh6Ai/KksU5ITkfOPxfkZetLWfjezO2ySfb9+Mh6B6lMI
A21bMl0vtasQ4xuSIiZkMG+LpQy6j3jLvvCw34gWY+fqM8NMw1LmiN0UXoDSFJ699Yfcq3pGogDp
cTrq1pYtTAilQBEFpAOzHGUdujGp0TSrkccZjq5YCJUTuGbo/M4d/urUxRt+TqHnnkiMvV2/ml2k
LxWb2QxIdXkPtGiLjGQCfQceS7XFQE9YclJMk9ZF1KXNdgGHSUio+r9G3foKD5dZ17TJMhNnKvC1
fv6JTcvlzBGrD1SKwxWFWA7xzx8AoyPXLW0PhgF4omny6SFqfXn0/xxPW1SFX6Q2s4NJ9GKXeRW6
8++PE1w22e0kWozoMMC0hJb2pj+hWdHLLW1PQGIDAHNlEkkpESFFLLnOFCiWOuX83apXtVSIiwmr
F8x7FiFgXcbMV39UUdf+/fopjNCTYijbjMFFZk8E0wxlrrYvc96xN0IYAzqU6ZGMKEE67aXaUyUN
rtOrw9Thci9qLsMbWEjqdSqzaSSRaA1vknBjkRSeIva6f8fBDatPhZB8PmdlGHw/e3Cz37dTvJyb
7ZnJS96IY4dQqV9qy9GVAnWBVAlOcjk2hb+tf9pmT1VMF1lEgktlWfokTuCaWfqGWc0DL843VS7H
7A0Z9x8oAG9PlwLOHdrULaMvnxNo7/5IYuXu4xmApbqCsvgohCqp9zChDig+wD7milOxtUztt4vZ
YVtXDszxFxU2fkcH9K7t6AFixqko4JINvu8IMoVnUK+cMWU1zaNnFkRm1qOPWTRGzGSoGXrL1Qxw
TJ+m4PVFileMFwhLGOmRIUlwi7HtduPNFSNgWpbigRLGbVs05N/Czc7L18WsTlcRYgp8AmewLVJh
ZF6n5a1b0NaUnU8yBWhms7UcJsKyGaMLxR1XtjK9uisFMQjNR6jtRUAHRvmOT3N8XNeKFnv/+15z
8DSKQ6Mm3ZF3+9e5Fv7fH3VWoFpfo2YnFSw7gKlGenfWgk9Aiy+9apub5KznSZqnJB8In3jSH/KK
zUdgXSUDL2L8v8nJ4Ik0VxHouF2+ewdgEI5+degHPvHvnZ/BH6l5E0HKAvz/37zqqWLQVtqdbATy
IKGeiWTtpjWvFIQrysRA3uWlng8Y6iIY3KDlkWbttDa5YInE0ezPYk1JzcAldrczEyMrCy9c09Sc
NRmIDwR3DoumNbWGoHj6512+MLU93RCNM9+kKeYQa/CwxKmz/1nOwqJPRNQWK7APYU4c+PQP07dC
0f3ZooxdxloIxoxVM2VKHKKh9WNQpk2j0KQDR3BQuUIiNS/BLbOuGrAvO/wJK0ruyKTBcYCYV3be
VdSPUcCQh3Xl/5HkHfj+9Q8CXTt2qS++qzD4XrX7Sg6lhYO22lAPw1vETF75ouQUNpKfjPXjqEuu
ayoFTSTQVWRuPrzAEek9JrWsG3OPVdOtTCFfu5x22qAIPfmEuOd3eaSUy0JF69wQ1eoNCDTvEtdd
C8Miu7cSBobBZiyE7okzpBlNHoqHMR2uLMK6L/2K97GJltOhDs7JVpEKuieiAM0nEy4TDDEXZ83g
Eczw/4uvLrAZSuBniXFHQJxc1geXrJoEgmz0qeTAUb4gWdstC7UPB1t5FP1YocrsX5KO5uwA1zKX
Nrf23T8GYw19NDYkI8Fk4kpXoZGkZc//MDZWxkhbcgtjEtfbn+suogHyQ26PRUCQntuBNtzSe7eJ
RvZE8rrCbJwzUz75QnF71ZV/gm+QV8HE40lnZQ7MUMutqfEL4OoUJUfRIKPWGrP57+rsCv6os44s
0hRFVMPa3AAKfgJZlDLC2b8NHonVrMYouiCJuGMWkWRr8eIUOms4+olEC5GWXd4ZNHosI2zg9gXh
FZFoHP5BUl3PkJ/y9kspFAe6z8V+e1rVIx5Az88/qgNmSTyNZ+BVa0Uwhqg0xjEgEimOt+zYuKxx
k61sDm3Z59k53CVL+LII2Zp/5v/1JhL+tQvjBTC8R0+5Bg2y3lyrI8knD7FxFPGXjXtwvbd4dMsT
JRIVCh+SWfAhLkrSwa2/waroTVLsWz+CgRaBGkrcZIsnF74Rs0eGWu3uVshE7Fh6wCrKxw8wZ8SR
o1T2x+0AC77qTwgjWdWr4uWouC4RWbVcub4dD/LYtIdblaKRgitMNkJttkLjNF42RjbqbBl8nzh0
0DsPI0bgNpv3Km5Kxa7e9iJN7fLlbhjRSr7ozGltBW1IF3P3JpBbqNB1ua4sNpZYOUifrxsYXkyO
KPtT3yTEs1Nk2mWzX9FqMnrLBiI6IHT0B1fgA90Fcnq1j7SS8ob4PTxdBLgrdwmmclion6nzfLrF
hoJ1V+eB+iT+NFr4h3TLe20mGp1+98VJQrJWwDGdH87kdfPJ1TecUWXpiPDxR/zdD54LK+DExLiA
nVj316vrXy13WW0nBGPfubtYyjm/z1wqxUzuejhIBvzWoBSIMsmgzjU9V1w7tamL1a3ZHCp3JppY
PyZfMctWe5W7AKyz1WVRMCgIuOF/OWGRs6st0rsD3LMqABSPDHpmxHAA8ejGablsfZtuFJQloqBJ
0I8S7vqFQ3T73YHpmSQBT/iVJP/LGaomMQcWh13MUwT+SwZAmJkk64eAr8Tf173P/bdG1BXTTtId
Ra506kb4BK+p+jXENG9+o0WWa+5k9UDa9HsBgEyG5ZPpHyWmnfL6r4ESpLbrfkMSpyJLcvJ5v6ks
rRQImLxVVySKdFitPGiQbIFnRsjkbobgSlODgwlONvUvGkHk+DfBdlVnTXS4nEyHlwfleFxjhV4L
IB1BNWgjV/R+gXVFimeHKxQ1HNmRD98LQTjRC3f4v//HCWc1IJ3jNjCD9YPEEJY6nfj0PTLrdrmu
/Ymwm9BnzUzcG1jd+GjtXkqrameNiXYHN1NJExRQGKKtOhMJMm23ARx4y/CG0nQF47FiEi1/Sr/S
C/gWbZPCdNgl7YKpFlxPT1LOswy69xNWVTZclUiVR3gwIfy1MF/a0hOZfE4fPfuADqEgQjQVv94N
N4EgAK6YDgkl6mf2KfK+G6WLCLCa1W+WVOaNWDbL1qWYPhplXwLtAQ0uvRxS7fUtbY+xgG58YZwx
+J6TjvhbxvlYLku7jjEPKByI63orfmFHPhi6UuzH04GcowgNo3Lh07LI53c7/9m54N/OFgNDtAgE
u7t9Ob0qr93V6jr2pl07D0pQAuxC7cM+J5rhP5StQzkjSEBGpmSmnKiMErnluRCt6hFnZekozEb+
lGjF2Lll90TuunB0CtEoGa5ilxfGenz1RrZIH43/8D54m6V1rvhP0pL6TQkODRODKOYR4q7ShiLm
4foRN/lowUF2oNmlzKZ/8JDVCEka326JAlSL0Vk8PoplWXrH8vn4LUuF4iiEaAsmqmMHSMnG64fW
BWJh4zWKcPh+8XPDdjGNfVjjHadkqC278xJbt+lLFOJY1CFcchxDgpzXe6yxu4JXSPoGgbJ5bGvr
fVtVsSGR0mYjKXXfTqVbJbHK4aAj85gabW2tLUVuPsEZRlnV2atPiC7aEcdqDWLk7o8Fj66rNwqz
wbhuM0tN0PXnxzLvqsL2z50iNbSUsh+Iio+xK06wPflFE+kzM1jgtIc3ppX+ZwHo0xOypl3mK5as
9wYCYmr/kjjXo6ZnpMbjKAPFIaWqRRhGIbWLOu3jIKS7nPYG2jngxP085bzNC8PSL7FCOUgk1BLK
NIVOjVrhRdbPpxqofmf7mP5BN7Nm6+lfSXF4gIIXlHI6u0qKAqpGp5NRZeElu6vWQv8DEZHrUfTm
aDdfNtyZargYCFkhcLc0YCm3yOaKmEnO4cE4Ic8Hsvv2X5j1DATiFiRoW4Hlew97fMYySKHpAiP6
guW+6Qkt6O7IFQjZssPagatd+Qwj551F/fbGmOx6cUzZwaGFRSDJ7h7bpyuwGAic9WrL6wyu8f+v
QcCouCV/9GCg8K4f4C/HDB9u9JbL+fXCaKYX15m5fUeRFlqAImkzO+IXhAwfhZWeVf8cWY1NCFdC
28aQzDqKRYhdey0Ut8RMtK4dPp0lWTo7fiFQ5mkLwvvTC7YqDBLwouq4DOI/9ETgiMTjmH3YRjuL
Bu23GdSkW7LLgJYbaqFQUkq+kEO1Ipnn34zCCBwM7NdjYR44oaRFSAeEqVYoOZmUobQ3e1eo/fi/
KmJfFGhxiHWKYaKnq3KgnuZmi2I78sj0JmJeG0Zs0ee1KEfTyCc9+t4IAyIIH/x7/TKTGbw/tadH
VT9PTWlEJ9Ug6AaGPdOd0PEEOpNduMSXQNT7utQwGN12ps3X3jPzbVs2rzR+6fmzwvfgKQGfEoxF
DjQ43ARY7/m04oh3is6YbIIsjg2UkjhnSZW1Gn8WpOTe3sCuypn1H33Fx8b5WmOfXnkCG9jXToQm
QOOJYVKhYTIzvb8mXvJzh/IcupCsIyqwSVWfvzxMc8ejIeD/6m1p9G+vjH4pvPv1kp9aNyVh/b9L
pys7NN8HuciQqeXma6XV0GMbaxQmaSnOnyvYIlFUBF+XGlLHzh6erl4AdMfR2uOPdxFKKOUZZomv
G+ExBUhvYiQtcB3SDhDr4/MQozVHTc8QL+ovQZdbOQiuWlwA7QzG5AYpCCv9k4URZTFvvPhMj4zU
fJuwMJ9TRldAQiGhThp2IA80feiiqBuINQ3+S3OO3fJw7+YG0KRR2wMRxbASvzs7M5RFNaNIRh7l
27huEjvsfqn01P8P/QYqVptquDSQE6r6wFTXx6w4r6+YvZvz5wW847ct2NcJzt42gyqA7oSiIgXp
7btO7VCg3WYPpWj2kWIWfR0YmYwJvetuMfh0rQpwyykZmJLhtwBOjslc/T0XlJSZDQBShTmvsEvi
zKu3BnaUufFAM9INeUCELi+jZ9UDbutONmu0lDtcb71Iq0JKbdxJuGe11+mE49kBUrYYf1xm98lD
2jHz9vxDsOmAFx2ky4e3CaWKq4K/v0UhsrLVEEZNvFshMTIn2SzXsvRRE649ZFZZIwbhA1nat8RF
41r/D1erymMRS1FIaAyG21pNSpe94o6FDdcw4+qsobtkfRCXVmHpWPKf2QkEoPSm7PaD3SZqYgek
b2ZHO4d8QLfXtiWL3CKV8T55IKIqPJPt2mRAh/+DizEYkmUKAveM6Sz3r52WWbT+u3k6czVQWdLS
JwYIewkuTDkzMfdAte78haW/SbjzCnTf16uDln/l0+kOQl33Zacj4mWdg2GDpzadnj+ndB21HHvz
FtI70llp17xri+6h+irlw/YElU1Mn4naLO6hyPFV/5QwUGWu6d09OcLjwEdZoXzseewfjX/wlgwO
s9IfS/OhzKRQl0QzfM36gOXw7Ms7VVAtv8nyPrL3Xnq5lxmrGrBWG5ljw5trPeLA/Q6FizPMRucJ
wdVzLupMeddH4SMkjWAY58P3q8mn9wqBGTsYXza5q6ZF5mdge1t5bWr5Km2X0q9YKHwXWev3mj/U
R0yWlgoWbQIGvdjVW1LH82dAoDcg0t5yYDzKMPDXJPCVGJ+s5LcUQl1JCi1jarZiRKWbd0pWE9vT
XoiaGtoHdsJOnEBxXO0BJ8QPrfifR1MCbEflMiRBnvtXL7SqqNPpiIwonnSBvR9fQA3pms0G6GmM
mrASeCOktfagbbV4nKG07eF6/U0+q6gciUh7wkvJvj812hLS2wVjYDuC7KLZUWyPn8x9w0WWlAz4
2QjDphfPgccIDPGMHwVSFnfhI4nGZe8ro50sMpLEeqhX0DClMhnflj/NGnyGvYOSrpGmtsh3FqJu
BcFWDIFBLmuTxckOeHvCFCm6SwBgy83A6HltAWvS6NKQtnyG5v6mNNRyi1lCeM+WccZmOymdnFNe
1h92ye3s1kTFArhvdUTPEpFaYZRnN3pL7cMljI35lagtrP0H3qWQgCgU+ED5typM8xEZUFBifuRP
ibbTzREUwaA6No3k2690xSsgXO5owWyZhKP2m9kM3b0I4IufWNOHanL2hdOsapv0ZAo0SQ/p6g8T
VbuATH6F3eDhZfTAQ+g2vK0kx+O2rDVM3LEqlcegRh9+/oQiZlWBbecp9qvuNltLbC+YBEn/U3B0
yk6jY4qnF1Nhl2ojCouZwXy650ADacSGTA1BanwWDXyyct4gyFkxOXPKK2ws2cHA9GCbKBKlX6+7
sHmn45usOmFYdijCvkDUOoTgcuApDvMsxc0h3tOptRoeCC2mroxg+TuYiX5hOiDh/DicgRSbEA/Q
NEMjP+Q68F9Lk4dfaCKzZsk1NDl64/oI7mpa7eabbf3/v4JbEsnJfxyl6BGnsT3tnkLzAW4ILm5L
FhLzLgszIIetTQ2Y9fdfsXlhPaAxohZh0Mi9jMh6ZR6nHqjFeCg59oPunbNTxcIXyLSjNgvVLSXA
t7T6nNeM8xaMXvwl6LcFkyHidS9rGJ5qE9tWKYr9CsMxJepGiRdQ6lOWDbY8SoEEcUgksp/QfZlE
cHJH/FyYUAdMDQM8nPMh9XtAc6zbWVhE3xpJmOvEnCtPvAv//uyhb1NNea99TfJfA3r9WV9DSeyf
CynrH55vDDIGzrZfxu71QaTCpFGVqVy+H/ssDkoJOcjmc4YahZfnAUkHV9Q75c5ri1LOc8ujqEnQ
RAaiu/ufTHlXMmT3fCOgVbbd2baENC4JjuoNtwXrf5SzYZADrGRqA/E7L3IpmOhio5qxSQh+bF1w
dfP078OdbM/yeVp6fDR9t/fEKPhtRZ41oDNUn95HAYcLfTSeH90aR6G3zYtAEfC1Vanj540ZaPS5
13GZXsT+IsXoK/e1vsFxBFh3Cx/+S7U7yi2BwrZSvt1nmItAwmjeYKPlTxyv7rI8Vj9gS9PVEIYf
tMBbZyqP6y0w7rW63QFA0ytwpu8DHIeWDfVrs1J0eVpIjZNxHtVHE8bFif8EKUpgldVAQDCGvI33
Pdo4clJcq8qPxMdQCs2pWAA7Rkb9NisfOD95bObqQhrQdDVhJVQPEeZcWsWJCniYskT2QYJaB50D
eq+7aWPSAXFHNRV+fQ2kuaquTnMj5Qu/V3jFxpr9F6UyKTRyG2rG++VVt2TkMMW/a+VYDG6e0w33
167OLzvZ5IpHCAm+O3AIVX9xcYcoxoMZ/WJ/nVIyXH1vX93oUiICAyP7LzZsRsDfo7u4idcXlWCK
v/vDDeW3/UzyLHSEvYCXHcGINNUITW5ttrxEYreRpQTRZ7K0olV4/kF9/obQO94M+R5fcau+0N2T
SUKz2xjMFG3D5Fa4fmXSdJ/ndHvdjm+KHc2fqvqEq0IkCrzCq8VkSD7+rvWfxZ0rYyN+cb375sJx
Ea4zxKDzFTsB5wVHah8iL7tqXM2tGbhFVP35S5VF5lC+7canDivTM5mzlJNH8g4eKB/gsnWiSYgf
HOHqtWW8QTkUzEv5V4BxP8nbBqBtSlxhlBxTSHfGCrqiuA0tzc9AFH4kUeAVt7SL8h8EoEEOdddo
/s6Qk6oIL4/5/hf6HioUyhkNrfIfVUiyJiW5C7AUqMIggwQb76p3Kg6H2SGhT9XnOEZQzRXJRAQc
4Co5+dRGwSkv7RJj0dDymAq9Uhu5XF5NRoc0ouCboSSVqkUiLRRXvou0eG7xHFLuaUR2Y3U1G/5f
vLmdoh1euqW/dFNyer9+g+C1VhapeCpM48LsPEF+SRTFYk3TLDHBeci7L7b/UHundqBc4GnPKS+H
3U1IplJUfQl3xv4qd0K+3HWmkAovN6FhPgQqlhDrvcgowMrvLm7KQ1PpL3NNtbgahvX/9bTnVvLX
iNgw2v9KUIb92kgKg1TG/EpMAyQILVjiQyxgxhnjq8WSv8LMQIjI1YQZdhkZ0yYdyIUHJeepSjfa
9iDH9k4TtreCZIxWaGIIRAbYAnjHN86ADXWdQEyrTgWliO7Dp0rZqufYU/vBCMDdoZEYOSMMweiM
z1dtM4VlRdwixFfRLlM84qCw4ua3iDaY23R10NQ+uWpyc++8s9UrtX+fxTaeRp50l2/T4k8pEua5
Pf2vaLVkgQpaeSQnRRJzlCvZPdm3+XaUFRY/tkrW0OyE2PMyOXie1MsLsLubGFySXghBRXYHj5EZ
/ZbuiaGEffb28kj7LCKSTg9jzluHZNV4wVvPJ76cV7F/E26og+F4YgjH9gY4iHX+Za+1oA/Qazi8
MLV0QBYU4xoO/WOtAta31UThQmonXCfKlnyCGFgr7KJcSyX/nxGGOVbMmDdrAywhD1YrXhrQNj/a
hkK2H9k68McTqcSK6NlH3YWBcJr0qnZav1O6W+4wZ4eKVEL008WFa3Fix53HZ8uGBa5PEs+rfzvd
Bvv+glBUEZtFnPrVIK8E4VYPvU8OotWQY6tSyYYlTrfmoJ6aIk++uaU7JI/nkqC9yNfu8QwITdRV
ePISSNEWkj46OyTKBRatluP/N+EDjxqSAanPT0W73zHXFwmgcps9MV2E6mZtlghBELuarTHh4+Ql
0zUIguJJTHcTdCeCeaFm79zKo8jaC5bd3+PBWqxe5VDpkEfYB1ATddiO+RefxwfmqhPsZP36/cS5
j5BNWGAyoc5FzX/H3QInasN/u69n6Q/vJbM2bI5nsLCeeGId/eeXwi/gGOQ2YwTH3gniDAa4dOQp
uxg85VXU0MCKSy5S3W77ik5/uYtjosEjnFR6iQMckm3XDaP+7Covr7lGLp57bcuNRIGXtlkYdDf0
bBKNNxUZR49HCFYtDm1ANsSgbfbnmU1HhumMca9F2N6WUBFXJ5iy5jG69/vQiHTN18mqeQuP4uK3
5NIQHcOSz5vJnjDLrW+x/ez0B7jPFeOWPnhhNvLYn5BtqKNwBVfOJsusRzTMy4mipouiDxVzMvZb
QoQEIlL5S6dN2DyTfIerSsHqQ77bLtwNwQrLyS6o0aZDJKPZSMCNTn5DdoGY9TE5rydGA/gh2rzU
gXvRKKd08G4qa/D8bNUOWJ5QCU9TQ2dkyGL6OYBBLeFIYqJzV8zmcf7GZrvo97G8PamRuyJaX7de
NAzPJ0YUfQ8GnzrhMSQ5PEK21xIq8vFMVmvCsErIc8o1mBB0NSJxwFnUpU1KvcHZ+0qZDtn2R+dt
B3vIqcuHtEWmCEl1Wm/Tj+qQAyi/iDpwsYhEyPBt2qcRVBPLM+VIwv4Yfik5VRqCmjsHgEp/gApv
57jcuTVwRVUrqP5epCm6GxuHDq0RCZKzC3YjFVpjx6nS4BIj1wKN0rIQRd9VagcZMkThKXUaU87V
tfrnwvPbDwtkYaJRfSzRQvUq8Wv8Q76/AB0mRoMLwmK78ysRAXzugj5c8shVMY66CnkTDCLTShEe
5nb+1BGawKUf4mDDh98D867WOXLjHohaUkfgH6bbWal8q+/GolFjNUDHv9srWJ6PKQ+pqsLhDStN
eQ7NHir/CoRrmN99KsmwWgfn5+SfROsrHKPQOYoBfSn+hc10ch7hR2WfvFMWqr7a1JFlvMh6PewV
FcQIFKK5y6kK/2gRpfcpY/kZQzhBKTqIHV8zZqlBN5JHrutPBQQ2+GKzicM8bBneA2N6aaDnCl3a
r/nsqjrIX76kyV4mOcMVeFUYv+vxg7qRExI915JoxMdEiL6HQ2La8rSwuyEkm6nVrVsJ1H0dZHz1
u50Cj/RkPC7DvJy7cYwAeMfDSHX+gSw41JefV1jW0otz+qTVOfiRLKYs+JWLNsNjr7XmJ6+WKmp8
7OtNq+PGyxpsqzM7VZgtgYUD9q2wv61XcUIUkuSWK5220LS4/TF07PnT/iXrtE+DDNQGjJ8suDyO
aO5qprnp/Z9AFcXjCn+wn/nX1TKTvCrBpSsZQdria/diBugUZI5tbIkBcQk8O+YQgZeb87VzBzXV
5tf+zaQhRWMesIcfhl02BTB+zs3/Ka04Bp2FaiGLf12o0qc5CH2dTgDFOZUM6DBRApvXTDmvqsnt
iC8QTgXAwfJkhPw93SBa65lB7vnh3L+aObzl3AbFZC96aLxk5fwfttgIZ2BQ1KXmqlr0fss+QMJh
iHGFS9xxuYyku7PVJCpi78A/N/3O3e9MePORKAnGQa9KgDi/5irMubh8kvrdpamcQuK18dwCfECH
h/Bs2Fe9Ec/yPuOG+hFyHgz60SvrlcGKAtAPNu8NGektlPcYOUYCnq2KvBl3WvQ27WPXXUIBrm0B
dQfbHLJXQgTRi2uvbuhQc7vhxMFiQsCGGnq1ygLNkgw4SKhEfUfoXVRxSo56UqkrxkPGMafggCDY
9Oem7c/HsruUhb6uCYkm+MAsA2Ukt+/0KHyqYqXhVc9ZPAiMwXWvI4rTbrLfymubRr38Xy5V28PD
QQOLs8N6olywS1L+lT076/b1oI737AYi3zXV284iMuDgkY3WuEpwhERxUqMWmIVcJaU/QLoQAYJB
vpZc4HvLZ33MBofwNQ+LbrUwGjPjGn0nPfVNbaMgvDNB7Fryd/9mOwhf46LUm0WPqmAw8b+JylPa
CSJesF8upqu+L/+9q6VcJi/SWFwz5qSQHI16DwoyyWFOIqiuoiwzQWF0MT2WgaiyH/KVtL1dGY6/
vBLksoM4GARVAn+9trq0WyknRUL0r9kWeZ1HhnlpDhAi/+7cLommx1/mQPdTnypIEYhHjuPbrEml
q+QMxJpjA4qAe+YcgWTJtpJuvMYNEEQid+aGmo7i+iYqlvZ7ADdrCpXTyoBMdewWsj7k9xgVSltY
Tgh+6U8A0A9QnAM1pxtaKmLUWG+EcyFxczux5zohQyV05CGIVcNGuUasPJnq8WWy2afL4eiHQKEm
N295fFixcdd2GfvLRI7e9wGmO7imebK5J3ub1AR0Z8EoeHKuYjw3v1/OWLngBYTZ2ddZvg9f/2ho
69dIQSM9v9UfeOcvb6VfHQvi6jsdGpLSGfPBYcgs3bP6PjMhf7fDV11mL38k5jYDWyxo/HkLUm94
RfU8AteUv4PbPdKQGsW9hfs46H4cTj5Vt+pVLJD88Z1h6AoaFW1GwD3EG4mPmjLmZGWVVQI7t9Fn
f6x9TE99YVScykTM5M1iv9E31QH00Dsi0e48wK/yP2Aax9a6m/vFZShUocL1Tbid1uepDm273kLY
JCozpGO5YnMBlI2zryzQGY/wP+bMZLA7iasnFrAY8Ckobz7+WnDlD70332oli57sgKlcEVSa9cdT
Ywn68cKsngqBUlgrh2+f2BvUf8Rp8gsGKYoAncG4ggq+lCT/Q2kyVPn4unisEoLf5rxFxpk9jso/
oltYxAiia9OvYTSC/j3ezQf5QJqannazIf1i9GNLXnK/6IU202R2O6KGHyibCdVRt80pA9PFP3pI
DKrK/ldafY32Im2qXnEQ4omedkBldhr7sgrUvsX+D1e7+PzoMRRnPefj4P0EYlYS9dP/Da6PtY1r
GKlD8dbIo9h7Hh0Bmiws1pGs9tIvg2AoeFRq5//BwjuZS4D2snO/Vt12irTcyp79FmuZB1keRGoK
aB/ED4+QB46wRDmWCl3jqDvR3Wt0FcQl+iFEuPjembdZif7Eq8jUSyYbiC/ZndWS9dBhkLPVv+F8
0tV4iPBeIoMEabHqflGnrT9uMGYrYpGm7T4w24uRP1sVQfja9UzEnGdbld+qg+TW7wqNLo6YGFpo
D08YgGUKDnz8svtMbhLcbq8r3yNlf3D75kvpNBGcpVtoNuAyeXqgBkHnoTOMYe5hhjX+zqBVH49w
CE6gYfqFdr9VykSbos67QrNtIA+S7dS4+za59QrTjUV5b2YbhBVizlBlC5HljiFnEnMe0R2ALHGW
XzddgcZV1TK+UKUcsA7Zm2kKXw/75cS4BbAxWf/82U7/HSYTUoALCyXPNsIIL//4DEFG3pJit4GA
a9QL1n0KeC9L8BtRRg5onkLyyFmHCcND7Prh43Im42sI8uLOMWUoeVbJQ9h54Gz7O5zFHuasXK14
4QOw6WOVDGZ9d63/Fxzr/ZkGeMjfxivXEPAm+z4RPGRDol3aBk7rfdGlET4oLvGD0nVgoy+PjtMt
6wUNej1MlulUOxYlUMHlInGkgqq0rsrjLKgU1X0qIs9jhc0ZyxyCtIobPKCuY6yQKIc6z1jCHl+h
VMnDZP7QfzeImPRCvRsY6OwOnJa8uxPixUqEtHfJhi4LiL3jIXK2P0EPmfmKT6XtSpaylfs8qZ6P
NCPIdujZE2huAlyEabl2QBnUVzrcqjAJMJWmSMvEyHqR9IJt2lNZAJE5yjqOTOc71uik82/znunp
rWZt2/5BTh6WJct7iSYVESTrAU4qNNZs1llkh2Ec6tgn6ID/Ug8bB0AmSgu5mnmYiWhehaqQq2c3
cAWnRyx8bNgbqrHMlbhDpHCzy1CmBpxy538QEe3k2thE357nJXMz+KQ0RlrINP8s+8PXGxCBXE6U
epmBz8LSMlOVgp8pZkVHbo67+ZsRT5caGnUoQy6GIX2t5np7RlzL1CYBDRfPZUWQB+XcWZtkvVgj
8vKW6qIWJ2HsFqN350WaIe4RIcvsr1GEUhBiG+uJ75dS54HilSCkw/Xn7x72R3+XlTFhHyZTUUqf
N7Ou0/+eKtPEh9n9G3fRuQ5JDlVBfzq2zXEVtamFvHs0NlG/7jevmrhxYoj8u1sZkubjWR0zfnXQ
xTzpxKpCWb5zJZGeG0RNcY3hwDAkSeGKzU+P+5kXVxnLArmcoXnTO3DfOE97/HPKq8OaPDh1Zz7i
HVY18MDF4p56bgYlFH7LUmFJImy1RaOmsOaYSwyvteYL4IVaXuXpwwj+ouJ0z7kSzMHfz6TcOsCT
yO5XxlO2LXPkIwn5pYcNlRi6PCYNxtG+ePdTca5YhrAS2S7L6Z5HOr08y/Xwawc7273mPF6GyM01
rZ6oFkSRI6Sm6bgXOJrQpwuChe2+wWxJ9VGUtj0ApXpFhOb8M5FBp1M6azUU9vmSeZbexChYOzbn
UXejCpeWIBImDUFK76NBB9b2NebuHZU6z7Q37OQGXUMDnNTanOCscKdwCTEBi+nOkiHKGpKlN6Tk
+xyeDbfkf4D3X8bveXnY5vNubM8BxghJwnivgW7BO9KR1N+TWEx6znvR0Fchir6UXMOlJqYcpTeY
TozXfYw3zfmqQv3SkmW2jcXV8WgvVFYIqgnRj1HE+hX8vCMIEgOn7LMJya0K0jXLf7D06Nr79TO8
CEyLs+mbgNO2lW1sU4UEj14KYzgIHkioI1F2Mergp+AYZ5GEyIeMnA8pZqR2LHrH7RYFvN6ND4VJ
zSllj1oyWgHQGqSdce9MqPz62GYUOxBPcrF/RopE6KqDijYTUQn5wr+cz1XDmrKLm0YvnNwDLlBE
3Jbhm7csObcZu7PVWVt4lwdbxrNFmvu5kext2hN8OZuJu8CTjFDIQ1WflSD9VOtzrApaET5i/TIV
eEUYC44nt6HDiXxLwldidDYNByqUGvaoM/0CQ7nqChoe3y5xcW5APG8vVm7upCN8KbXkkT2Uv0P7
lVMXvdfq3vmjxsQnRVNOj8ijIcaQSDJVk5D85Wd64nFUVaI7Nd24Yj44Ons+bie6ccIUSoeEVgh2
E6SM28k5r3B/++eDT1eKnAOc2hSnWadfhLaWoTEfmMLG3AgOR/ed5B2LGkjfQhVmdAMCEAt99D6Z
9KaNPylG+XvR8SS+rw4A7BoJmwC+nkXwadIBaXU0+YNa+Qaq78cDTLvZRrnIYGc6LvQ47+ajxiBS
DAJ+adOMxUAWLTHFKDunWcB/2P8MGv3tyTLLV9BK/IpAtk2Ih3QQQCFuQdEKItDDbRyLUxHA3RBO
BUpoGk0QiZRuUoSVdVTaIlPBm1RLb6C2plXv57F2XNsL84Bpa9NgIarS41G7b2SNaeXR3Sb4bwXY
ypdAfxBkwqGcE/qI4JBv01N7uwfJyFK3kCPLGWUrN1NFe3xXC9eptWpY396kx56WFrWsgS++G2rX
G+UBS1oJc7JVkTCwFxjtMhPDl14WHefitI7Q0cEC9NIkMKDaWAH/MaUMw/b8tk2azeYlJBp34NsO
wZCQGQblecjZI2woPkkH6fYI73z6PhigTVb4cVfOR+gctkOOZPdy7k0FfqaI5E0dP7bD9eIj5jlN
zgqDWYzusjX4fAnCsI2HBPZJov57FCKmi5Nl3GFYMBeGm/244DgLq4x5P9Z6a30izgbJW8SZk7b2
nR0aFTexv9kB2PpnmZBjo9AM579qg14IGPyRDbtfGQrcwS4ds/fGsWph9+ziTd/caS6afKnfb1bc
hb9keF4p3cAEYUuz+lNX5MySwTCVeZnxmCa0MGlVQFI2c5CNNgM9NINXSiPjCg2atdgcrs4uGhio
BKPffe8TxCCAf9fWq/V/AgeKQ/HmcoqivKE03+gS4ms1WHVbHkuvwLNIPa0V2ayn6k3E1Ic573Vz
qpcIbZ4TB+PT5sH8G5fq/0U16r3O/p7TME1X4F9Ju78wfqgyOSlPbF+zdJYYxofdKA0xb3ubeyPh
uQTLg62bzVG2E+GXskuG+kngeak/pSmpe3BNZMIGozfIg0OjbZDD1sY6A97hUhm2S66EJFzkGyE9
diB8MA1CwTA9MU0J6tcAsEtJpDoQXYR1qI5lN9GwNF1UMRKGRceVoaPL4HICbyZFx99XgZfg5ayc
ePSBCZXvgQ+ArVxGQ05MWzz43dyenE5dZKjm934DFwK+1f1QnIeSksLW7UvdOWGU/uPo/cvYoZHu
bQb7lDlHNnNNS2hIORJYorV5vA+cQHDRBV1S/q4k3QokzADEEBoTWlGO2BcfLOpb/mphvOxPLjWo
Wkykh4gMw982+jXUPi04/8Jx+QLJSiKKEhAu2h5YdPV7L7do+QMiUeulzzDQiVXF08XixQfIx9VN
aYBGJg5iVcl4KjQl5XW4TeNT/EfmWv+OQ/7ovKJVCYzZhVgUpWnGjLvpwr3P7R/cDty9+ADoWJXS
Je+K85bZ8APEm1LEfqlgfLwwbDQKVphTc29GEzyfvy7yK8Es0YI1JXKTDwc3OulcwNcq15MWtQZk
ElVLL7cbmwv67iGw+/0xti7gTvKGR2Hde1V2HgSQ6dgK96PT4CpzClNOpjRW8JWj/42Jxa+Y8QeX
aDMshOCa7726QIanPQO5NUoLtMvdipcXVYkFpSviixrDhDvbBh1FxjDG0CYP3PtUktKOBM0LUswW
QML8d59nOg+RmRFVOJ2h8FQSHLjXwdqqRrx8H4b3GntunmQlId1Nvfpa4TykzhtQqW2i0fN+eWg/
XzybK4z4tYhsqMRZLllwrMjZZCdimglnuJQPRVUGoNzFXrawFCjKF+r4o7ZOc5UL+/zky6NrPUrC
w038HUMjKLBbi4090KGj2T82T2k7DHJdhx/EB/C3WNvcq9zlH6gkts8iB9CBxrWt8jXIngBBmU57
GORfCaRXzJrdDEGrN3KRWZlRyADZ3B77HT1PVJA3761MAcX0UbIbyASILQbGO42/NjrrMVi7wSwL
uTIG1w0xfKyQS900+M57SAv5EUYjLMsa0UvMxQkHxmakYC1aPQyIEkalMr6lag5KHQ8DBS/bg70Z
KCMpXoUiIqw7YX4ugB1BGXO1sKmOrtoc+fc5dXVwHBPfehvCk/u1SbSY+bDqo77GfOCe1jBTEcFf
mT8SbAF8cO2T8P/aD4FtbmX+Ld47sZRaNWBksU6U5OPLJaswXcgSWP4+IoJDKMfE8+bUNoQP+KtU
cpSSF67tQmzNyUdOZXpSlMNpqLFsVqGJn051F3u1Qg3JSV370W5ssqpiJVd0FMj3XF7yM63nJxj+
O+sBxMH5VL9PFetNrDlYC0X3kCeckNwa4AoQ2HMedt2jUd3Ksc5fbcw4jZxW1+UfyOYSQUVq738i
N4LKcazQcz3cOlN8NLScjwzi2Oar440uaabpB5l6SaVBOLfqMHpmKavkfkkTwuL+QLkqvXVpE/u4
bo//Z+hH7U1jBN/vd9fFP3IPzhKMFZFDjr0kfoC3+0lUOYNcmdMck8KmK2DH0GS/x7AKB1PicmUy
HBtPoa2HD6bfK51Tp2JY3X2jynCIT6GjX6ean6q+OVDPOyu6lVPghxTm8oRoFjvLu+KhePVpjkhK
8q85+G9ydzIH2Fw4tyx5kqV/U60t58mlaVcUnuuWx3y4Ivg89WW7Fj5p3p5yVwHMq+Tv5Gk89woD
5YhsCPU8buwihZCIWJlPKl/jisjReOktgXNBY8+aw+wXI6s8OzObVQ2im0scYqEPghKENhPwq8LF
0fzwyRKDSj/Y4Z3yWXo+dYfTVYLSMZyl5JwwI7iNN3wSswwPPCXhIpjAl2WjFf+Jm4vCBvTmXwer
W/kI2xOWaDyq1Y5dWZ+4PFmSaLPvycy2LBR272vLixkz5qpbVeoKKC8/n3eIHheXFUnvqKvhSy2m
CceqIl+I8OYQtMlDfV/b5vmR4DT2rb4pzJrshqry9okrZ0Xt1lRcGwyBSA9d+3KCE8+86NuZl80Y
Kju3zA4oFZQz4uxF3/kxVIjWhbBt1p8dZ6JtWFeN4tns0ZiwVghnNKK4MzX/+FV9p16EaaCF844/
H1OZKI+U5ukQhOyFFqRY0zvlnJUw4bwDUt1bnDrbdz0qTi886XOzX6GSPNuAn8pPSSpgoRpw0OwY
ExhWFyZYSuhnnx92UIipiO9c6kOzcH3uzMWOVxf7MvobMPC2QZ34Au92DL98+pI7X1eJeD02wny8
nw6I7CRRbz8QzHr/FebHLQLuGayMkEqGPYBlZt1cgQxsLO/l4aomRjF1k/j4spHenxT2BB/F97N4
Gc/bCPWnCMBAnZpFLC4Z8V2NU6b5CwGO1FKtuzsm8b2xhz8rWeacmMP2W16IvkSlq+wiagFtCXkX
C7M4Nh5E5uU6HHAE7mVMqVtm2tF6taoAlU3gGBhDe6uNYmXto2RO9ApGoApVH8i2lT8j/8DXPNxd
EUV/onBYx5iTALJ8UBojkI+Ka4HJRgFnx4FKWqkWI1YEqVTixTOpRO1uOZH6LzaXZS1DHmwMs+vd
/SmIZ4NWCzMz4PI9584Oj6jzWtov785WfUfCEpW7j06PIj2wy39HYe85CM9nlALJysEcP/7tY2Om
w2iZwswPmmV7KUCBYlt/GGqx4E6E6LG+m5ouzp4+nSmKVetrLD1FKLpjZDhhCIzDGaJ2+y18fiRi
8gK00lU85DNvhGGZwtqB6bKcvb/ZjX2TR/wLQiaGY5WfMipwMJi+7lyizKBz6QxzH4YFTGndcEyK
agWB74Vv/+pZ7VMtvrxs1G8n7rM3qOF09gkB2UfBMAJnrQnMraXpfVpIQuC60TLUU8jIQn7EOCj0
tzNpY54B1EZgAH3h0gRNOTU+iP4ndqi4Iig7ugT5sPAd1mDKc3XP2SN444MyrwFc1iqiJt50n0HE
Z+SNIXkGc3saNfjTcAjkt/PeOlUp+TjKCW/A+6Bxc32hOvZGix3E9/QyHCMmLGuM/Cvs4ZJsswww
P+L9kBn0dN+UkO1jnLwTmhWsqHMKW9VpxLMZ+oZv7pAfXRVJEPNo++39jDsckMAwvSxvhVXlPEHc
4EARBW83afQ82jMUJTChf5pyYpHqybtyvUHZ37SNehUHMeMlqyi/27l3v7i68hlP+Qzu0ueD6jtc
BUDU0kMQDLo9WJdNLiChrk6XlrwWLKHDHtcU3RXLAtP4Kb7QvwUApsXsSRMx3MKrldq+smDaa/QM
sPQLjGTdOJ5om8QTEPrwFtNWw4OqPHXDaH9xwyW23yPJP2cgo+gspkFFp8NjPg4rRRRwpoan6jkk
tvpnpgqfdajx2Ojexe5OMkVQJfa86aq6CmUu2KBeOC5GcrijrLBRYP2DCT59j5IKgQJXKHHfz4OJ
n7dZpmA0U9mCDvx4nOVPwYOzrGRUZJGSOcykzIRM//5PDcjgL1hbQI5CBs9g++qKcOc0PjER0Yzh
NwN+7uOSz+Ni4LlCujqpy/UyNjfgl7fc4BwwthP+ggTqxmPPhsp4157Z63QYSpn2qfjOeiaxCnJK
gjBg1/G9CGlxXG2fcnGNun1gHJhasP2oo9CjHBUJ2PlNu6MMEbvc2+zRanvdIspzytlooAmoEIzI
2cgteJpq33S1etHeVAFFe28BZF+t+uQCwz/YqtTCo02OVqAKg4in8Ne3NTZ4qVU+wCjeWAtvJP2t
8qmqSKq7eNfoYwp3t62iKAKZRbKtJPOqdesPS7r6g+eYcPiVo7K6sAYYNY2Aw8kmVCU03Vo18NpP
2GildLrA2Qivx93b1XNKahu6jzx78on2JC23LYqkmRA0p8ssJzA66SE5BUWmDfH78Y7x8uOaO6cg
HI2Xtant+gxz7zu1QJNh/odpAvBuA6V9HzvqvNK7HdUzgZn3eYe7HTM4OVTo7DzHd8d1c1Bv78YW
jzXuiNhwI06tD8/gLt3NiPXvuM/agnN3psCQBBdrIiZJHbpxEL8jtfaYo/406EOBFAu0fFCRXy6J
Lmp8xNMl/0es+6ojYl7xuwk5EX06ZK88pZNk45UoAlNl+kHysnBGXRdg1TpxMEh/wEO9KJ3grblE
8JZfgPRT9DVeALoTCWS8ga7aaca8MyYjx/ToRNue5JefrqQAJpuLcG7ffSf/B4yEvJ3DTb4CQ5Nb
wqg6J6EDt+tSjPsUBK4GCaDXLnvbWsEjP+oG7BJsL/1xUfPwjX4f9EqZKNJ+evMt6qtolgFni+R9
2m/ebEaGov5HbPxhn4NuEk5rf8BTtm3ftM97ZjQdZ/+vznMIIFCu2p2JKci+IHKN8obJs6pqrect
GZ8UTHHQBP1qLif8j+63V8waZrW3IKDeg9X0FuUG/S/BXibZ7IhW4nNrDfzBgPWku9TsJlLs5gBE
cOqL9eHBRL+fXk9KdRdkJ7dpeeGfWs9ZyHK1KfYNoN+MYovjwz1rC+EPobCWTgTwehsCCGBksEMx
Dz8oIEE3RNbBHIOMN63Z034ZPywmROUExDjobN5vNvgpTLyXvk6cjI7lnSq0PN1i5QV82Q0BoFDP
cA3BU+kbr3Nu8Wsgv812VxTRqltYQiC2GLiqNSUm8kGqsFWtlgdKJPTvwihgoilJHJ2L0OAAWIVj
0GY5+mfKkst7dsTTzMtuBkqOvDn4Fs8RHwwdf9ns9U8vHS7OJDD3XCJGvOpJxZ6ONu8HAm0IxLeS
k3FzivxUVf2YCXX44vM+GSnudTgoBbSO+MHlwkj8mdfuXWzHPiAB7nKKjmiJis5vaM3+l3fMEEdw
YTZZv/jKuMa1Vg+MtWyET8mSZs8CvvyBl0LBNAPA202XZ7I7xhY1NLqwzWBKso7LU7/zbhe4Vwh2
4uAXjtrguqpr3V3aPwIU/1EYpgHTlS2pLYU1o62PBhjhjQvRM7dmFLSKVbPMTv7489Qx71H3ItF/
Hm+0o4Mp1JJRI4ZVPNmgbprHsB2fJFhxh+3EK6KDzxf1scRrwMHUN1zAwTMDzHB4qjBTfZ8vHAiA
meU6TLfGx8q6gqyhtAiB0f8vrR7rnkuuRPD5NgOunPzqFyFWNdmFkwS3AdqDBPyp26T5pIXaUNDX
JNR0emyg4utOg9nN0qVO3DhBwQfFP59blmcJXRBcj/XMSP7KWSJvGkWCSnOPC6d8hwj+10KC1a3s
aDAOty5Itjn0mzVeBaJIO7+LHS5MvIFYFuT61dXXzd9uk08J/+GB59g/4qom/I4fQ2flvuOKaYma
jyILKDAjreboBk0mpusqpJOAYT1EKFJ5zNLbVhrtmxJnbGZo1RBZ++nQS4jJivWVXRYcv9gXocjP
kSRxjNnYDRuevQrATgd5iVA5SBb/Xx7TAEavcyIpjQ7LCDO6TJoZCPrPC86QVMs7X1VhN/iBbQMv
VAvUr/d3JhPedRr6jPv2z0CraMaqDUgKVLQbbqSj/NXDVByTFRv56Ew5xx0MGDPXPP100kj2SXBz
c56bTfrPCiP7dkHSXn++ndyOFi3RRjPBnT+xaZKQ9QbNk2D9ne8/BVIFZHtB9HjR0k2rus2O5TS0
CCm1WfYHwqPhkJ2wxKl4dC44UoCRD/shMxgKA9izW5A7gj5fu6ocAbtRF+ecB9T7/7HOKoC1YPF+
BJr+0Avmee7tT9Z9hzeh8mLEroSazAuE07DAwGCucYVw5g7zuy+cK9aYs4hy8pnRzM2wF8EGsLeU
Gn0j5TZKZYnCENPt0FwCPMpbU+FJRfXOgxyS0BuCx4uVdbVevheAi51CJocfVD7w/W98GjNGwGQ+
3FNRnCIaR26nS64twctOegBKnc7a0hZ/xNlowCrzXFgD1JsbNKu8OLB7qeVaC9Vso/SAP82FB741
jFR3j5i2XUra/JkmREtnY9KmAgP0YbVHs1yTUF0P2XEakAE6OQh4cYsWhVFA6ARFCy2wTCckDRBm
w0/HvO825ZDZrSDnd7pvr/Em/rQcAF64T8HjpINybsXjyZvjB6+nejUxPn4/PdnBQSmWThKobT6i
pWquo6f3zXaYuJCPZ4xAzTWi8B1hTh3FnmgfzUqXQMjKXSo3i5wOSk8HKhSQI0S+GgQXTYGOUO94
VDizSDofmQc3X2ywjdJGZJ3NoSNeWesyU9aOtShj+bf0IrtR6/g5cuzgac4HK0H4eVHmS81YNtxu
edE4G1EA0Zesy04CfJaWrZMyJThJ6sBw6NDTsKNfOM1W0J/naKwEo/TGcfbTzOa8hrZbFOSF9WHC
hJOv+GUDRxll9OuUfQEYhRs4FnR9snQDVLt4tuC8Wwb1mILd5U8bBLzt/tDFBFL+V4PqCOC33LAu
xvT7mikag5odyvdRM919RoCfVccVkZCjx6O4G2dcrjzdZh+maark9fdWwQY/zgxvlwGomxBDCYHV
4DZVXQwVc1L4XYuMVicQuD8whpu3lcoe4fSnKI/vBCTtlYBouVUF8A0gleRDZYMQg5Vtp9gWt8dE
BVodX20FofLw64DevaNXOJJrcKa2/XwKKlsN4KOkg5cPPhfktulKgeuVhH9FEyzCBjWY75rvmR2R
aUeOSh4eBgI6ZaTHiIXHUaxz3VRmdexWdqrQa+61e75IloSWQIQLYKVv2EIJ4dyKP2KDS22WOQJS
fkvpdhi2VpY98q88varxCsA1CGqY/TJPqSKohsh06Xq8S4wjodb8KswHGTPrjBx+VCH3G3VAYNsa
lubHkq6dZrHbCtHCo6nvZpl08hAjHfinR0XdWpSCz17zFi5xDWMUBbQwIKAubL2vvQIWukNtz/29
ynliu1PCWfsqM1QbpM7Sa5kScoo41NzvemYRbHFr5aNqJZczaC42Z3EivAwdwfztNaxGDnbxVFmh
0Ay8GCAJATcylMxINtwVevQMJKhFX0ur+5Wk4/7Dwbs2dOzw3R+NY3PrW9sgNQmhLC4s80PGebHi
zfENMN2UZ/m7JydhXlNkfmoz8shA+VFgDVh5aWkK8ySFl5oE4ypSZf2aQdTA8m0D6x2fHzBnf0Dd
Aeh184UIWVAJD1m7e7cJHZ5kQQXfOGuHtI44j9StoOZo0lwygTvFwSg9C+jPK9yDeu4Q/vkVvvaH
lbldCPX81xiB45nf46gB9mMfSxMZVIHuJZr+pS3xx/WywMdZycyDtUeznxhO0hrQgZlsFiV0ktLj
LDWuvUnmSp6QiM5+BFG0B3iDvhX/1xnwdU0Xnz6lQbXvTT4Olb1hJgnR25HP6fnFbnDosOxgBNL7
Zs/sj++fb2oOnffrUxkewBimGIvGnPpLW2kzwzl2n9P93MZOqj6x4LdC4I3xKNzCh82AZHT2SyN7
kx3jDXz+HmCco2qm+Y1Y6AjmD5VicGWPBhTdLqHjtTAy40w1S028mY8/DEkyzVp/WQ6zeE/WPY/L
tcMghjIIefG664/d4TxK1FEjd66e8o+NZlL888EjlK87ArmXZD6hNY0UbN1Q3tGjTBbTrkXvDmrB
on0vKPeIMSm//XxHYDOsdq/80gQF9TcMy+Itq/RV0WJ2fxMCq01He/LipcJ8hs20bg1nxahBMBSe
9cssyashiGfdyYtfoAcZzM+5P4nZNenZ9vBseAFehYtCGnEVaDGO9mG/7sm5OgPOEwY9KhMRUUI8
UH+czq4Lz/QLPlxp4tk8pqu2asKyfpeovR/Pl1Vkrb0Eqk6lMlbot6bcpDFrGdovKqGa/7fEEWV/
cyhCkUY0Ns2xA2UrBYwZOSIBrehBXksXx34ctlOQ+abwoeHm46Locz1u73OZfKefFJQKOb0hTe7n
3pt+ofd0stxm3xEbT9qy0/Mmc+nOCtNLEYqO+YtgWC0s4AcNOPiBohDG790TixosemFnkpG0K2VD
NVnxmWVaHwJvNvTxbRSh9u5em70rk8KAj3QZlWdZV0hc0Aq7yB99S78GtaZtwvYvRZbqFzoV4Fd5
/mYRxZLLqdncnX7oUjw0PYzDx8hZn/QL5qgayLtTnT7Ihwmhzi3XEVUldiOyWlyx5c0TLZMu7yDh
lhPqKJ4x73STVtTq2pRTwOXqC6yfTKW5qpXrkjG5NTbTvSjkdrDTz3UXMylOx45Uj/p3eWQ1o+zo
U9gHRRtWoQm+Ijr5XpDwfjY6Cim6CNUAzrz+4p6DRlEpuEeJvm8BETgbtyAcADiXZ+H7OZGuEvUH
LFqxQnNZvJftv1yaLHiHxl9c82nS6qnVraWHLbfr7eM9A455p0DFz9ARjOFWFOA6g5pcRN/V3UKx
W4biYYki6Mn6rxpHVfxdwnhzNh+yOPjAkKbgXC5oTJZGpMJfSnCmJl2EiAL5l8sp7wjEdf6MZvpa
ugj68HLE6cKd90mMMc1VskBeq4yBp6BiZ2hI1JCqn/fC4F8xMgQ0mjkbQos0XdgJIXcX17KbLTx3
PRTpRD75X2g86IBTux5xz0JEasgs8i/Plfnm+4ipjZQ47zWY8i2lYbeV9hY67413uLMvp6lygYaL
NqprfRmU40hHNuRDIUF2H1CnB2goKojIH9meVR45mVDz/S6MJyM5ekFFhQy5ONRCKxdtY+ZSPSpg
VqcwJfNPhUztTXH3I0FW5x+1zBriqJjCRbh4msMBn8NKg6UcPzZEUAJsQ+yHQNA0Xp2cCQJ/8fKu
86qFih1iA7K0yzVZyNPvrBDzOa/gsM7VACwWD2ymXEKO5UXLLhe4EI1pBx5WLewB2h+u2/lOXlIK
Pt8oS5LzwCNfNV52xP6JnjHX8nMHTyoTVNDMHwXGje/iVV8NDsj0dE85M30Ba1vw7QxlS7chHuqE
iVy6KAR/Jmwuk50k81X5V5OFLwyIxwfrE/r3LqkhsWLSMWj/xGcgM7vUnDt9RoaDGaXnmg1Qc/69
m0qYnRZuR48cfCcorvoqoj4ZResK1I6GSk512BrXwgWbaXcFh0B86MupKyGVXVD2mESgBK7I1dBS
JK0EPXMevzrihRN0OjILICFdqUGfVURKSx+k4zq/0wGVs75bKZkbVyo9uaS09okppxz37T5UmB8+
AEvzHnGezrheCnDNlU+9R/f3GccqPuYlVVfaf0uU5TdzPRY1Mo4ScW468GTpnW33ea/y6HDiO3J9
iaouNdhLnpsHbbMJTQXJks24D6Q5JoP4Ku8VqbQ+ivdIgvs33RWKdRzdSyMbNUCGT+t2kM963nz7
2r+sAoB+W1G1jzY8wiksP9IBvkwTkObyfkxeJJ26ZLpqDsWi76PW/UXihWOgwDQefA+L9LRirczD
cxkbG9yYWeBR0zs3TWeJ51+1HaZTlj6eY3fNH2cdYBZMGiJxmNYoiWDhi4KjLv4j883DZzXyc1jj
2KbIPafLlOlY4ojnx2FLk9cUKat3IVV87kkRjLhV0Zdyp4xP+aoY8hWeMusYWEp5lHs8KOHzPFuQ
cPzYYZKZF2Cc0qPi1x0CTXX7Ejl8hIWaaxGxub0PTt+FRfZs1pGpVwFvp9ijfiwcPBCagwLrGyBT
8Ffsbgx0vC2PdeKGjNBdAh3qZi5pQgaNRJbb95Y86ggxuTs4a2lrsdMxLll9W1dyHwd+4eDVGRRH
QAdv8XsXHKGVJoqQC5QUotr1rCJKfh5slB+PvRSdF8Wn7uUkyzAi/BGUq52+8ntPIctqtQHXjBNN
VjK/hKYGFgUUTd12u+tamANQq06h8u1QZ/gm9Xr3HvxvBL3/PoQqblPFJmuoN5dWMYfnlt6OV2xM
8NBtB8HwVJqUMsTFDBNwzpcqTO4t9NgNVl0tgfTJIYq4OPkI2yvDCyAl0K1RF9OkuGLZT+9yiWZD
TFvhfM91bDgcQftvEIYTkmVYlztbk+tP/Js67Wv2g8UKFWqsf/Yk7rZ8Ch1xluiQpszctzjqOh9y
5sCghMS9JrnynoKQfZCzdaP+b93DD79O3D3NWyGg+bYUegKR0KhF0TZOG/TlSlipZ9eVNrTlcpQH
Nxu2fA0ZND5jvFVr3NseOWV0NCemqvqMLJo3iaSHgPwSrLCKStBcVS/2TU6uo1mWS4xdIyd3GlrA
qvI4REDH34OaSCQz5k7UMuU0Fjsp5fsM6taIcb8thUCFfKnzzOkBazlOorEaTrnxSBPEPKcWvarT
2noKqbURY1koxeQfq5mDpj9hauyyospESdPRVryt14rkr73QKP1r84GknDBoV6LeBZC5xFG3TYNA
Nq+XSRSKPcUAGJZyv1gQGRMEpTj0K3lQI+0CsSiJl74W2b6/s0BQKaF5g8m+v5SiDNd5Za9Od98h
4zQqD4UoBqJmAW1OuQvj+m+RHoAnpjH9oKUiHGR2lkOH6nqOMvYDZrHIyMIqY7lZqhWjAUW5Puso
UsvvAZnr33TvejnZqvk6Yv4v7ggqKMJGzkUpHoLIDZYNdbGCYSlbCfFCpqivXMRQnG6aQ54OZ4KX
W/KB/yFwniy/cwcZo2P+xRLL6DMi9esR2vgdObTqpwxXPkjruyCsaK7NlyA5iBkXrpC6xIRJRyw6
H5M/akMQ+bX9ukPdfDGmXDmfF374CVFLE6VDL6SIbbg3dBRpsEjkLUbNVYErbZbsLdoMX8+Vp3oG
V+S/GpGoDAhlLwBv0DFR9PV0HHKuN5iGmb4ME4j6iF7qcvteAlVRFllEnWEVqwYuxN9hC6o0V0go
b20VBmZl4kGywyjxAgkGaVdo9sIpOLjZI3f14H0Swfv10XsTbWUaDWJqiEk69aE9bVWdZpp6ucSW
T99E2jby5lk9y1kJqSa642+xsiw9AHCYXuori2zFGrG1fX4hy7rKv1ithci4vqgMIz20m/wyNtr6
7me7hGdOlP11LnptFzpULpVkGQEE6zXTGI0EOc+wJHSEpmRp/ygjO+O+Dv7TXZe+iFwzD2SKKtaB
CjzEys6OnM0WMS+m+5+X/tIBxqYVDC3u+Atw+rWAB+/pFnM4fqOWFTHRyvYl9F1AJr56uOPYkDwP
2oI9XkUgzHg1fGLn10tBGfbq2LSOF0yHYd+g2v9dXmxwQ1gADdUr85bu4DblVcyCh2n3wbvywrdZ
aXoIxyTmPc/5hZPd21QnqnuBR39EOp3h9zAqzhyUv8jgkKReFcBkcRm3w/I1zVlHEiCpcP7JJw81
UR7m2nkPpOwthLwz0W4WN9XC798equ9O87kqo7ARL39uRAdH7p4BUpBS3wmvZgCLdnn+va9ibpVD
hK224AdezFrud5arAyYLR0T7PAEkY3tal9zTni5aavGiZzTDTMcBltVET2IedhwvDV2UBQn2jXPL
tGBbzWHB0SR2wTsf4Yl+RPyQDWywwYbDZXjkOqdAjJJxtOJrmgMPkUboCzG+qOmoVxxgbz0PW0l6
1iHt8RzDhOARsLOYAvTp6K0C18UbYebK+5DJwLOjQp87F1dTqbe73ujc0m3CygrJnSqyPhOg6ywF
O7qZuaJ5tYkxHZ3R3AkdGpwMurWjy3sm5VzSbf1ZmL4ZvsPIHGdN57DCkLIRQbsrEa+PbcdTNYzf
9Tmh3xahhVAIQtUz9jEKhOO6y9iBRkuiL8AkAgRNi+AtSZBiu1lwL7cOjGgOFakedYtfl4KrjhE3
jgnaGGN9hG/+vL48vFuLrWScpI1aVj9Hga+6UEI+JiK+nUNnnYT12zTJOJRccxMUcX5ckqdl5dcN
7vn0lk3XxkITxLoV6CTEPYc/wMu2F5GzBG+537zd9sSQDGiQd/eC59c1+kghdgWyNfcwHJWzljzo
Jbd/bFV0GfgaMISwvAiRuPOMrSpyDxl0g6gdHcf5L1bW5XIS5tIKHV0EI7ZysFsZOeZn/GT0rirn
T2hOgJLGMezdBrmJ7tY6RKm/TRZBlxbcKmMiDL9g1j7cFT5Gk0zzuamLf+gn5eq6nNKGd1VaoSUY
fxw10jx21kRXq8pTHG64ERWqeU7Z9d4EmQ5yzRYsuhmjQvRFouf9l6QzkFLaCpNqmj8vbr1eAkBB
nd0hCLLtLedU35joy9YTr4IIUGpEdprpp707vmUcNvsVgYXmMbhxlVhyPPHLfGI75RUHKViUkLzB
yF7xsyHlpUT7To1p5av7kF0wyQWkExg/geR/4uLCtYh2vYvDj/WDWadwQVib5CB55el3JbKKFCDl
5YXcPuq9qJM6v8AMFcJ6fWMATXtfUjUWJpSmZOuOzxLa6BUU0Y8iYeuU91AtxjouSrdrks1nq4A8
ymaGx4jNzt7yzpnDt0/Cw8g7NRUu/8z5XctaoOA47/FRHGyfPYyqnxsSIVf8aDEP1zR0RSwOOR3C
VIY0kCPPQWdzp8CwqDbv4QI8FB9q0rtK45CySrmL/7Sbv/AD49SeyUoH3p9gy0aEyWc9U9ae7YTT
mPLt8E0KD6vfrm/wpD2JELeL06wweTTAF6LzxoO8dgfVXF39PKzILrqXcWOZc2BfrkIoKzPYjie3
+3rhQn+hR8bmx02KPLWO1+zcWLwxTyX74EoO7PEKMRPE4+FN564jscQpvx7SsaZjE/fJE0AglaKa
0K5/68Rjv4+d5E8cMbtR5xZ1vxO5a+b4SulGvUwupIrM3XQ2NHyzeOTHZjwGiLAiN+VX7prWx5l0
4kiFILcZrVT8+Fvi+xNYfTJpdQXA8LNUKgjDKwLTqwzoiiPXcNxERJQM/XradkIQcYiizb/8bnBr
1pyB1p1aSnxl+5Xz+mMVIYP+b/GSRgsEEyROMsBNPlLYLZmEDbEHVn4cK2qSDFdEM8gOH3V6J3NA
uT6rm16KwXqnVdukwx9m9BJteBSn4ev7Hvrss6bSgFnjODnRmh+1NyIfgPlPyAFd8Xl6Fctg3lnu
x7UnKDENLna/Laws5UQnwDYiFfeCK4haeNPDybC1TvcXetSqJ2cFHJVDrUtJWR0nk/FZ3EyWesH0
NEaKaOeSVoroNX8lm0IYMOHepVpNl0U6W5XdMc43iM1REoiQacWib5FoIpUUNfbMxk1V9Beka6tD
RvdGxDLLONqR6iNbBsxWoff0FfgZ9wlTVtUUiGMKphKrKySTEp6g87NPM+LjmwtNvqDKn5UIiJEd
c+ThPfZyKMeAwcgcxHUJoGGU58Q6BgSojSStC9kBc+w4qIUCurCgYzpfESe5mxnaGmm27iOQSzjw
fS1/rub9amYoJ5BhAwuw6pHUJQZoxm2mlL1Gd6M2RedmvSuKjTa1s+VaW7x2PrAvEREUnfdY2w/m
NHJkNmEAzjG0rqrB3XKkaqvnJoC5cdFrENHYpDpgq1SWlFNxU5nOxsJJPQlxhjGJrIQxeX4tPEuB
ppudsWGMp00VIMxeosfP2Pdz/poAPw4DPJcsjcCqSOw8zbf+77P95IqBZWXzTAYtma/li4Gg9+1m
o5d2L5Nfr0brHg5Edu81OYAA4shZU07Uz57ox51qF12la5hz6erhpHgDzf8bqPx+dIU3U/GMMvHl
iPC/zA2+Srf4xZhuK8ZiWbON68J3aFMhrKhkUAomxf6p9//2CUxwwoFNm0PhWCjXweGp3RF54+x6
+D/1xdpuFp9QIUoQGivD1NBSWY2OVyWH6937ZzPQ3BBw6WXOqhQ/3jD3Y7bJ3yAdRaH7jIVhm+O8
tCWJd1s9B0k4dh/kThPbzFU1nUFhVgXlgsLSyPlyv3FdQumPQrFnZ29rAa39acX9ke6A78XM4VmI
4oqwv6ykmMpFODSgelJ4IsxKKIlsq50EBroDXceTNhaPvB33W8VP1puJXDU3p2w/nYvR6FBClqnK
0cItx5oSM7Cc0t04o9+v41pfpx/Fr3xVXOwsGFIOZjzSFqLqAaw7vx0LNU85w3ogeeVR5jNPf+tt
tiuE7pjpgnNmwD+s2+yrS0YpEpCBMItlzhqyYjWGNxnj6aQskW1rKTwlsrYwwzvYgkJDVr5oSaYX
vCAGnfQXvxe2uTPItB3PbyA/dnAW3qtw/JVT4ExXy0cJzIvZ84MP78wdm3c0Vp6vITl3MC+M2kGq
hvlPtAHXz9D6ZW/QzSwlXoNhIqwkcEOGmgj2TW9FeJKgrQqDvLTG+5h8pIRthrjlYoI215GSv828
/DZr7ErBtdWaJp12lJ78Kk1vILIrYKTrGGqxVhIhYWXNAYIJ+xokJCA1uacS/MoUtArStLHNdQjg
+GWoECZ6Z7b0GNXYNC9Dk5TTups4Sca0l1A3CX7acJK2U4Q+BWUnMnLvwfOpcA85PzpkR51T7JoN
aJLSm/TQAxFXTIjSKPhehWREpNPP2z049tMc3CGsSjGa4Vc22Gl1/oALg1oG5p7FskSP/pu1CL7B
dDV/eaKtiXbea/BiaymYsK17qWnHBREj4cd52JIMPGHchVQbGnWkJUTWzJB1RC03diK39jHGntYw
LKW0P24VetKeqQ6gy8A4bVzhv2i9Yr+iiRqQ+xJiN5PHEoIJxxXE7gmBvIMIvnLAGlovMt37/gy1
8Faemcd0dUcofyBmIPpl8sWX5NFEHc1qz+pPVRs3II7kGszNCoKiK0Zj+ANEuDhvwRQsXwzRZiCC
Io/P93W9a4TZxfOwbhv/cpavBKAdBAarKvP3ZcyxWohPP6f/pX7NGsOsjiu96edEBeNGeV9YVsOK
rlRTQox6XBIZ32gg3L8Ihg0t9IJRypnuEloiT9CsAblVwsYSXKupFjTSn/R0upjsZ0Bt6py/+KKq
7gY8Em4K18hj+zFPfqL5/EGNvyoPnUoeimKwVi0ETIFVWCD7zPyw2ued1VlXDkbWWMFS7DOaBFlZ
/+ytRpJThyYbHDTbhGI/xiHzN4pGDAQqpPTi9TNjsPwOfV1NU0vaBm0+aKLK4Kcr0IwAUPu6pHMi
owGtoAGwhxzRAtviy1LCpb0oxg/lmFzEJrLS42rGSNpchjegXdQuutJuDQ7FXY6jVHBK+2RdZMsQ
WFq+Ct5bmDN81vbmA9fbG4p2lLBNk09yueBWQtAPh6WGFqh9kQce3SI6WafryKc01zBn3+wxwwow
gT5sFMzjlLzjyC03IogqNyKcEWhvlEHcohvMvot5QKVZ1SJ95XwBzHh7qikspcZvXljSN1HDbMux
HJQEfb58tId0N0iqojU1II2fJhBjW3YXE2Z8XZ3p7qqjUKEt53Hiymw++GD3NSU3tONrfDPz46aI
rxLChKWfzOofrsiuOLvGe7dwbcFnfpZemrGr9BC0BGMMyOIwWW0UyxijAW8A1Ba/V9F8JtOqGXgN
lHejhkj8s8D/tco+urYU2lOFRZJ+JcbmNEqvkMOWpfF1xssSdUMsaf5rI8WWRs8w1hZpUWiRdqCA
m4+7iOMu+43xYzglCzfVFgkEpw0Y3tdJw087tVRWnBrgmHaUzLwU9TZIHUUsh9LvGd3lwtYgIDJB
xEae9DWvbdlcT18XcILnaLa8WCEmG9MkEx5P/WIJyfyjlIsRTRDv45w+1FZiDmRotsainPLPKRRL
TZhn6S7FEenOwAAY0EjB4CsPeI34kmaILeVSxXaaNwFiO9ru0wfLpKhePZKb8PyTTK9u2IL21UnH
7WNJuf4E9sgrmzNZsT0Gbyvbyq7Q0iJ/l14NCajDp+mVRXKOhzROLh2AFIDZyiVZ+T6pPqrgx7ty
M7yxzsTpkdxZ50ScljbaSf2F0C6uSR0QBNKKwXs6UO6jXRQhWd4xtG+GCRQdA53YdUBBlqU1uiE7
V9HAoYY84nC7LBI2myaF5jpuf7gV2YAAcUR8n/TA1bmO6/WhDE18Tv1tRQtI1AFiyqO7UMLISuyE
5/EBRYFcdXP/7wEwmsSA5jsCjPh5tMmBs7L/l6dReguftuo9gcWikCNSehnwhY2ScL3LXgKN7Sk/
/F0R1ruOz924H4seZhFz/iAcWOq0gQx5wzz5WeDKPcRl6R/Z8NeCY5xv8PdTRDl5VoeC4Cp3QOeZ
UvHVlU3lsGnl/aDedV3fDiiAVMmH2d9TpjZUwG0UY/CzC3df3/0ngVjqD4l2FiA/wSNrNQOnFetZ
sEAqx2DOO/9M8dC9mx8rvbmb9dRELppJ8Ov+i72LWdERKsQKlRH4by4TZQwcK/TvG2Pg4fS078xC
monmxz2fEEqFsBFBVUOoeZSdH18tyLfx4SyrU/7YLpaeKAnuAY4lpwbIRaCCY5oXmco3C0mWvkUL
or01ieEA3QM7C5vizMO3WwbN8104u/xNTde1Yb+MG9lUtfFwdwr8doPsOSWKMY7SFMCsAnGonMR9
qUhvpM+Joj0W2s+F0uDIudJsGS/Ca450QBNfTmP+dYLaT5nh0X1NA8qkb5djnypg2abJywYZwBde
zY97bbAKRLp02ATzHnPuAiC/sDFtz24fdS+sTaXzKpfM2txVWBWxwt9QIBB7JrDMsaohwNpYkx/P
GXD8spMMdY+6swH56P2IVpgPIqu6589EiWGNp8Nzb6uFUNN+4bB7dPWOw+qewnTtlVgdfoRQXPY8
RyGh1MupOZ8BRBOe0/w0whtAqoWz5jKuerJWK16ralurl5nqaxSChXW0HNebRW7o6WmuJMeJkHcM
uypWLBfVKtC5dov+np03BWBAr+gvwx6F8we1K6o4tfNm8JySFn760ufXVGI+wBAp+t/sMfaeRdsV
aLSMYJijZIb3oTY4OUdVxtH8G12KyVimjujAhneQag2Qa00FJ12m9wuFxtaq3FNtXQyGm+sdvOWw
/jcuVUpjy7ckmOlDemKmpZcez9bJSphmhotzk1F5RhdUQ2vlAX7kumbB/Aw7PjdUUTPVBQgxaYJV
ks61t3B7KV2o/YokoEKBWBzxRFpkbJAskFV4OXAOHWqqPisLZB5SnGhdffwyHeWYit3NRbnAtcfj
4RxGQbzLoB7b1L4YJVooP4emGI7XZp1D9wWKYwVoz0jRr2hTfxYyS4jwe+KBdVo/MUCWX0ziPToW
Ea7+ZI5ewsUvnagkXxwkiFUDeeWO0DS1bH6NuhHrXSfWDcMTdBwd5bc5Dia9HIPpAnw+7/Of52LF
IEpSOzlyORwkfGz9ThpXNE3WRar0znLOwK/yamGnunANpZMWgQoqkC3x+N0dIWMtXW+U13HB5e1a
sT0ioEUkAFCH8ijbJNosBfvMC/mVSE9c8aNImstckM9CMs1j44wAQd75j/LTlR4jZ7a4R/nHjpJN
UgLtdhGDXAqR4+Ljj0fVoQR5rabBQN5tyDohnAmRJNk2YjkIg/VOhh9HZAOyKlXvrarX1SZN576O
hu+4TzBvI8pab+ZYS3IYFNyrVqOmRqm+Rwq6nAsWTDezIfHSJdg7IjSLCFlE/YMooL1D6tODGJ7H
t2+SH2bMNLXHtFj3G+rOxRIU6TKMJc841m84z9Ekmu+JD9XyfB7HFLoy8Hh6J3ztfvsB1YiYgP3U
JkVbS1oFO8xh5f8YphV1cEXPwDdLpa4xZYg7O2cJu90cHsNwZsyIheTViwnc6mVj5+DGuFbyzB8X
U0WvYKl/RrEc4NbDso2Lu6r+Ubq4/bUW9uB+tz5WqgSjS5QT4y4SmO/r02MNDhWT7489eCweFt5o
FXzAL9hKfujLQ6NpbEfb0b6HSpe73eVVyCfRSyknWU9GGOoDKB58L5niCmEVGGirgfM6eQ3pIU5L
NbhPMhB9deLjmR4U4/uo59BHzUnTAcN49vHduft287XOl5FxYyyWGrl3DGfQot9nTO6MFStQr81p
pwcois/HQ8REAbg8E6hJI4D7d4V0gq226RyA9EYL3L1ecwP7Xwm3NSZZnENoFxRs4AYX1jRRY7N+
aT83t9bocutgFHRk6qLlRkSmifwWrACG20uRqw4t32XwTOJp8alPKcKwfod7QWzPfY9BnwgEko1q
WLzcAnPZT7YEXk9q1dK6/yw8sDE4jcE5nPHicyPkRclF7oMO+J2EKBD1yEIQSv19+k8hvoqocONC
hNIjlIXZ/bcEU2YUUIU+R4HClxYtb/mO1JYobh4GSCWaziS8oy5kSRdLds+uRY+/o9b4AQRph/UT
ejoxbqmgvn/YgOB6oIyc5pjGg+hXYjJv8UYo/jqjlrnr8z3C2VVOd3YV6Q51Gk5Y1AdQKVjaaQQU
GoO6j82tsGPVZ8BK5mnC3FrNLt5mgXZb5lf8Ux9i6Njv8KnVefmhjRgcEkuhyhfkNMK8OeAykVPL
K6aWOnP2KR7ARy0kxyS8DV/wNUkgF3ND0oSA/GwWBa74eW4I8nfsQMMSrcQq6lQe33FZ+mGezkX0
qD8FTU7utNhyQdcDogOYugRgTsCG3RqrSaiItFYkYmonxhldQWzslNrChxJ3+BPw7Ait9yHPgWPY
FL/GDf5a8cKeTHYQ2F0FXJiT+wZo1J2EC6rCU5ZjUKOT9NRyq5xM5i0W0JyECvBf3zyiKQnOuwst
zTjzii16g1QF3c7k2aubQxiis3CvQ32tXgZjMLk4dgcHQfauNIYYQE+PniJvXCkC8UOFlY/CKw4Z
HgVEbM95k8exOBj7R4wl48rXx89Ux3gtrVOM86K4T3CtFoBlnlYOe4Jod8+GevTOJarmOP9BVaVJ
C9btyJg35QrPLYUVnmowfPzMz7ikAo7ZFXUSj70kT12R5b0dqvVfRmIP+gcgvdXmTXaR7cHxJErL
Op+fthb8s67lH8ZgZUpUOTIEifC1TKCQDMY80uI/rIWrRMEgkEVHoCCznIzGwYSQVcDWTUGqNRH3
EFFEYOuVEbJ4RvQQAyRj7mfMbAW9KAVpCcBpHMy3vSkqcUETHb53RJ9OrM2arHXuIPv9eQfpnVO/
Jd4t1gTvytqGXC6YxEuHuWUo7tRUw+wt/ouNJkgFaEAP2gP6MCKkZdKwmAJTpbd1mFdwEZNBzIN6
Fn36kJ2X/4gl2QuUTFxlN5GUGZrRzRp6U/hv1Y0qeeqgScQBDRLhn4xFUBKvqGZuF2G7HkQvHgaL
DaoH3268LNBrfK2kwjJeXKcRnJj9DDLuSvgLczIBOel11Dmg+A+JdkTfTGqPZ3q2K4VHqcZcFeIC
tbxOWilkWmaHtbv5vriifI7RXimdkPRqrv0FuoGzdmDdpojhXIVcbwKEWZDLjiJbPbEdNNQzRCQJ
qLgT2dV3DPgh2i8zfLmhTByGJKk1bVewr143JMSCitZJFBErTI87kkW7Vn3fmwV0sqTLzvK0K2LP
WbOMwQ4uUwH+we9BpaQ3m9s1Uy9slZ8BdaO2dZbOWKT8bpOMhLX3xv+6kE8EGanGGslvYF6wPfNO
PvpmVJhoFR+6we/0Ge0F+0kdnTUrm3pIg/71Hq/LXxBjZ9JKzDYwgdIlih/RRkuFFZkPw5D1I8nM
iqMEcNIMn8bowRlKYlalr3UDtrAJhdmxOXMKR520G78ht3SZCEGRjcnqIsEAI33WAO/TDAmSl+yT
ct+Y5tLBTbIRfHVyruRKdmb0H/xJtzWaEig2qtWM5fHNe4LV3/6UUMFeC6vZ8j1NDbGez5i0ZxMW
ysmKG0bUToKPsfk6KnChAo46uVBs8CpWqzx+GvWkb+EAvdOl4ei1gxxc3mBAQcKRQp8p3UxbBp9F
fdeMA5TAbTuYgkzBFt+5uH5YKnqgF78eJfXV7kUj3KfWuTBoRqrMRsKKDEuCzBBEtyH14OzUGNfp
AC+VUIqJpBWn8ztl+W/X5oLlzFrmlG63vKD0Ss9rMmHXYqK5i2kLaUFgOA8FZiagIzqLNbqIFUm8
wQzdHdEGVCv9V91Fi6YVNnuG9ZDBN57K5OhLaojPPQbpPHtJtd/VohrShdp3wCu7Vqzjrb/bXuAj
hB4iA1/OfOnK8raLdW0Hk+Q04bVeENbtDJQpfAx00VJeR1M1kEigewnm9Y9A9Vuj/qo4nvuY4Use
q1Qj/AIIgxfTi2QKOQTmg7ytWQsAFWShq9hj97/Inl1dlrfEqAd9fAIk0U4IQiPh2FyjwtieHj5R
dC0Gg59TLUvtXX+qrgwgsLSUrOi905mGIeT3G5R5jPOkLF3bhQSjaNQqcwpUBIxjib6mhwDN+sgj
BgVF9A1fl3rZt/6iFBKvxYN6XbuAdq4X9bf2GsSflfWdWHaEclPOvQ9kPhzRxkLBKB3JwdhbFulV
HMFSmh8vCVlTv4ayFcdvgn+wiFlnFjEDYJ4ICWJfmdGL4QALjdDJuaPBG4YXaiBrOqdU6aEr7XLN
zHD7f98FnWcv9PRarfkPPq8lVWu05S4W+p/AnwzHOBxiBgp40frwic5HiR67SQPZ9OLQccIg+TMY
C0lmLTmzcm34xs5FkNm+3ZHxOFyI/E4zj3PAiyTO/kzNhtG5qxRMu5hLRd3+wigPU0R1YkB5CPL4
WmzI1Dg6vICFSIyVy27wO+LyllzsYgJSeeaP6yvcPUb3g12TmDSNhif94kXpwby8PZTqTt4eMen5
erkMnO9QI7OLAqlZTNDVW1hYxBtc3RYDicu24KDfSQ0LZBt1vkwsMv3R19plxc7DL9MqquaAZX4q
8Po2qixYoPT/5uNxtF7Fa60A2nHwyp5XnmNZKpV2GF/H5cWnG4bu0Yb6ULDYckaXb5dh15ok5uOj
z0yhBvNezjp/amAITme6qrbj2JluHgTVxDUj0YuT0cPOsNjI3V6HdbpuPsLlXD4CBAOSQxV+J2/v
MYNgZnYOhW0dj7IPNTD2hOqL+A0x7VcJzoGPDzJaKZOKshz1y7+rdBiDAlocx5QuYdLvAoVnMmWM
seh8nU+4608EZjWly6y4gCs0sITVERUbXeB6Q8xrWcS2RlkZ3QKbrlL7B5gvmggNrOgp+FBcZSG8
ZAjI9PXMlitazfTR0gaJAJc7HRJEsG+KR9YrGx3zFpoPFCHryx2h0r3XjKKQWsw7CVY3OtLwfVUn
I72WkbatOpOddSWTegscxv4V+60nwTrQLZxQhDhS/4WoxfV0vBCjNHB78kl6ZZ8BxvijRbeyiMAV
qEngxQDbv3pvrqoAjFqZfwAt4mQon5/P+1VZOq4dWLx0Epedw4KWbyCF5QIU+sTCSx6j7COMz1wt
FatEMugUVBKa9RH9bqcBV+GvSKCL3hePQyuHKSjvIx83CSh24XU1BMSGT61b55nPNXNEmU4nwvKM
8iMbhWJGyIEapYrxjK94ruzs7fXXGlGlbQUpXF/DiG0YDDxpYU4+zzQzITrrG17z6NyfIiQYOSje
45nB2H+aK4DP7KkfcgZBsVbJ2UnzcT8n2RLmIas9pzuI0mhw+aNZUzHXiXrnVfrIveLeMXZCr1sS
9qQnEtRGhh/+wytENZRz+i8NEuM3V8uiomwKJYR4eLEzp27UqqvhjrqeAuuJRtrrHxhzpuPwMHvO
3kBN8Bis4NC4oZ4v9K/bcZMI2dWY1Fnv84IfDQzwMc113jzxx42t+xF+7gFKdvm6gidMZGZzq/cS
34G/kRkHr9qzJwKxKzxNYd46bb28ZguV//A5rSKykRojWi0pXyrSTXKt0pb0Vomh4euvNhH+sQC6
tNEgGHLJG+6IrXFZsBy26Qmeim1H/VGYgrE3Ngq3qjjC2ebjblBtNLHrCBmZRaeK1VG6JfiwGt+j
6yUkl2ulUWXIjGE0g1xWOi/swL1lrfusXcWo/O3LIc60OdjKyGfBrRHTZWeWgaHcRC5+q/d+RU61
J55teHqMtEcEjFuv504h6hMPzeYJiB/pk7Bm/suAPHYwDbbdx+q/BW5GDpOQ3wY0ey3nnRqthiU9
+AUa9zSKmkB59KCcyNM8FjTBlPDrjyxAy+lxuYbs/t+hU1ib6Hc7FJX5gFi1bIz2N6eQnoktn9FH
+GwSiYsk1SQxqZc4xeuqv7ydF+5lOYuphIE26h2/NVZgJmlmDbJJ0+M13MD6uE4qihwRcqrq2XdV
TTa2kFaS8ZMzGcfP8rAYkdSZYwDZUTv2VTszO/I1y05RqnHc8FS3jPYvYm2Lg7wvALAl8TJyJC1J
D9LpbHc0+TuBil002YeYuOS+52DJFaKtmY4PWNwlgGgFsCeXHjdb9UA/RiNiQYb3HIIBJdz08c8F
DTMEoELN1YsC4GiGamqSRA4GPYRFG/4nTCb5TPqVFqK0pv8dZG0GzLtQevHK9dy1p5RMBl1dbUXv
nHF5gW9ECXyihmT2Kv64vN33RIvekUefJwCpCvU8Tu/0OauRuRTHRJiGm2NHYrCjULnFzpW4yAtz
IdTeknQ4HWjq0HK4VbdrQqSiNPiyyKBp4inScOG/YOx5hf/Hu63Du0/wrn5QiPg3Si6UP04CpHPr
kbFb+w0inKjuDm0Wk3vRvgYfH1KVrIDpCfR1iRcwE2sq21TSLiWs8o/oOR5gIm6pGmP9bUeoI2JG
rx2JtvdmR54qEUGPnIg6C7apBkyaD8ajiEbFje4DbY6o83y6H9xLdeLxrvLb18ERZHcfdjz6Z40h
DaN2nlG3Q4TjgLLFvXBHZ/Z4IcrTj8jLlZLHVBOAgulQPIoPSgZ6iGCEmPs5fDErp0pA+NoO8m2s
TuXvmKJqjjLssTrI29cEtLBv/nBe/n+n54Mco00R0cHJJBacRqTJgXP0BepgYcmY78/j6VXRhRl7
mvytaEW1Q5KdR2PcfHenOQ66s3lcKCTA3Z3xZyMvTVGDIjBIv4PM4RwBaQ3M5NXQyBGR3QkxZk9Q
BDFOiuIpynfJsiole0PUCNZ7dHrRUrxCdwe5RSxeP6FLFPzEnDBSEurgJSQLUOpVpzo85d/i1EMh
fCsHAmUfLpymABiAyKhbJwIk5sErFIVBCYpH0PaOBPP16GXD9ISMCZey5rukNJhWUuiqMWZGwXEN
0D9AX3RUGp5phVfKvS0Mx/NYYCnHzkhDxgZp2i7+umF0m/2pX8PbHSfNxANBFapKkfKzplzook+a
frU7eDpg9FSAInRtqntrloEgi6mjviMmmLzKKblUS3eLnoqE+slq1xpmibtjhnwOpJylu484hsBh
4gmf+S97UIH588B9oZRK4YkzD7Q4uCU5AnaNgTWL68CCO0cXh9PhB+KXk0W1jdq4YZIs72trIWW4
VK9cug3qXef0kcZ+T9sAwBPcJZafMy0lhpwa9888t9IJ4EIwfsJbEFqqzE9jS21pziNclyZJ5oWN
DO3DHrKgbQImSBrIEPW9AKawa1n6Y4iBJgElEGXlVaA3zU2A02grg1fJGx1e5OtwFrFP9cz8weon
DTsYveGXq8DdZulOKp6NvlSsuHVwr9CW3fdENn4nmEuIsH5LoCK5dtRQsyP/6QK0tvHxBZNzBygI
+1kXlI90ES3J+2GdaFsBUJqI6d63Yepva4Cl7tujlevJlkAtziibokRfIo1/Q+uA8+DwjWDJad0W
UvcegHXTbELVhBCmXc34dSsoMUKenaW23kHsjn0Rloizy9AsfdJOkryQSeTfER5lQsTM2RHKE7sJ
2qL5gVXuitwVPHktuH5/MOdiw5TYygIlL7xdRNMUndrwjzEasP6rI1EIqh6Us86ZGb65ZKFFh6h+
aHZ+FOvnzmzqH4CLgpyuCpdkaRRrNoMWMQq7qWpNUg1QOR9WYIL5qxfRG15Z7fAHRvbsy1YgVmOR
KBjftTJ1BptCS5JEx1iUx20Pv47KURm6SrBXP686gPo0yijkw5gvEWvNXt5pv08C1IvFtuuQ7pBZ
kW8c23NXBd+WKZe0TIl9eEI8VunhBFTvfDUIin62AT1qVmSMXbDIRXlJYJga0KLE6QDz6G/audXJ
QHe227LAQa31RpeO5hnJVqWn8OHmC2O4joSAu0X87Zj4samZQ1GnJSI/6qR4lifBOxe/43T9rQSa
mIm95IAxXbs5d8DN4v9Zw9wywwHwKA2zTkcHDj721MumRhW6iset9AlMc1iixLzAF1uCSn13ukXT
+rT+ELd0qma+HJLI17R0z9VKcRXSZNwUgZ3E5YhmztlBAwO81+6BaEhXsYu7KgP0jZ/GnvZMwN7a
TQvBON7cl3IGgj5ulBo4aPkVNLlI2tbwKMWM86AhNd4xQBjBKfAL36ys38ZiAVr+Lte45rr2InCR
2s/xg8HSjN3v89HnhljZqP85ksUScRBmrvecYvFsvdBu9fpuH/METLwP1l3tPiWxCHv5C84iVnRa
Tf95y2QQnpo3RaQSkD1lFNriv7FwKuDyYFB71tCV9fNaJnpZSPt+UNbzhlg2UHA5/6sqnxyqfwGe
KE7Kn8iCFSiaqnh2prq5Q8GkEmcrfOu31PwV6ZEoNGPDzP1zfHW7scjk4X5g4sQbrGQr5I20DsRZ
jp/BP6u39P7kTCGK5XE/qVBWJkVQqW4URmpwtLBbh8adqeEQ+ReAb/JKqTV/4CTyMuo82XGeb34A
UIm5tKONxwSFzAHfHIypyNlN+VcnxPpeM2voU35BAtsqs2398wkikDDJovmtTgQe05KtCssQCw1k
J3J0lVn0VpwQ1wNlkKg9Jh5YcUd7oF/7FwhSCrInAsn4opVhUPiXbROGx5wnuJXOy7ZW6CwNYHtG
8P9psHgkZGomxSvZGiT0KnhdcHZ4BqdfU5EFIZs0GWROR2nqjx13B3pK/jbQkgR4ry4qg0ctN7vg
YvxfRwfDhmdJ79zvMfrGFq8tq9hrn+DHAnT8cwEvGSNBp6vrOLLUmfHrpFlS5ndP8VBpXzsFtju/
24Ud5TJt4dCqFBpxGVwRdQFABMegYNSZdydtM1o4tq8hjmklUZNO+7+sKyOOBXl/uXhrMO7QPrhn
VnmzulOYKm8HFecqrpe/ELxCMkXjxzSc8LfV6XShJv22pNjIB8WUOGIVRrLvkKkstutGVScpXh2F
cCHf4zWBc/goMhW3K3LopY60ufqFHq8dlwGsOIZchwqMjqhneTfHMeTdZdyFTL2IXNTLAKEjslac
7FuPV8Xcw0DIk0yzj06zzqg0qyaLLZbP82yBfn8MS25kX0W79+WtjAU8K8lGu4ymOAEGhZdJOxwl
iKPljaHijc19RbOMlBhxR5bxdq0wqGNsJuE/rQMFu2kygQY5mplnoEns0cbJ66xPqNvGB07xy4Ed
yt3ON4YX3PFMHU0qO5PaC5Yi3r9qH+OJtGRHkc1hzr9cmRijBiIQEYktotQie09+H5THTwcy2eFc
TIXHl6cP5xJUDgLK2PlLjKDnJ5P71/vRFiNTnaTQprq1Ij8F5/3YiO9RCNyjRnZfvZRUwZx7ARM9
2JmQHn+ZKTPp8WZmZKOiWMgb8h2DJTInj+90BlRMqKc/OTJlQ6D3H/4oGfpdHKIYg3wz83M9v/07
hHELTnZMaiztBpvTlt2u3NELtDeHs6AFQnY3WM2wmt55d0KTytd2XH9zQWpxrmGCq2fgwbDQNha7
GyirG++hFpWId+cBxhlZoXgLTL/f92m3qDzBTRuKZtBzzXLygMJguXaADeAiWEWDXFxE7c1GkLSL
YReB3Js38cLj0Yr+1ZwR6duV+NazGD07hERogjq8X/70AU6cf1+ods5Df9JfSaLxBxiS62qVu7Zu
xuc2IyUETsYmy9JrIqxlcrwTBHWd+A/QtC1BWWxR03ANTn7RUgrL/ieAGVz6y5+tMoQOOARm/wJA
7CdfuhdNTtDr2q75WZUSlnsy6DkVyMMe9D/S/B6E44aZF5KJyNLSDpjzvNE+6nwLXi63w7PBHh1r
hu12mKgLx7Nv3mMGhuu9AyQJ63L2f3uRLg6ntiFlxA4HJHTN2KWSzCDT+SKW846fvTVxe0Qtxa7x
RWb8w5A5ztgV6v0ZmZiV0ZFP2TityAx3ftHOUy/Qb3phcXeuP5+dyB0v5mqHsQ+Djjzwm4zmSakv
bMV6zVG0DPGHpbKud/dnujPJ0oaC8svNi7eYSWCVgT2ctdp1ZmdCmfAarQy7K6LcCzcOCZN13JU6
8ttW693P2G6QDuYilFtLWHUhV7B8ApbgLVX6SjMkPZLWY1xh1JiLqPAxRhjyzu4A6eIS5ZJKJkXa
BKDXCfzZ/fdxJ+vvjZQDYPR6pxGUG2Z1Piok7YWWnHgJEbQTCuWigkVry2aSgmtON+KaelTx5cBD
NGXdikBBfEWQqu0r22cQotNHIn0370bvCnJmuwBSH4f5jQisxrH6DXSiykAc0sephqeMzbRI2LY7
dnf4UJyig2EKjGtuAWAgvcJ0gg7eRUS0tNZK1VqtAQEacwW0+85Zowna0Zg5wchknpva2GslT2YR
SH51jHXdx43+g+uhDQzj5TLudSo+nuBguWquGEDkHnkTuajEeJ6hZNFGU9RaaLbzc5AYvq0T9woT
dVk87kakaycndm2iKojV1u8Oy2ktJUioWc4OdzN3hdRdPLJwtoBQybfjtTta/MGdAv20kr/ISsAx
e2B9FZHDGdXJPGGZAo6V23ppr6zyu1zr3YYTOw/AEXYEhedZlGpmOVv5JDD9btykpS3menktsbHg
hch26LCXSvrDB6jn04OomRdilo7QIAPz88jC29ZXPd5TWXSw/R46c4HqXZZ9I6ibw3GC0YKq+TU3
HOyW4wScUv1aGZ7r641fFtdD5NWHdnSDt8+9etXiurlhQ0zjct2+mMGxqIHNafNdnnee3GkYOO4m
6WDGcBFn+jLWAPCHrGUChpa3MSftimtea1zfAuKMmxWylvzQIukCm3zPTZCgLsfilEtYlLudJAcV
6+NpOznJVcxl6plH3w99tqHo76tagQbGfshImyXE69YYYAiFVmDXvizWa80C4mHW6D0RrUVcWVBj
N9uUpTo4uLgeuhRXyVSYI/Rdi+WkjSREPoUw780hFxya+nFzDJvb7RnWlEXNZBi7KNUd4nXXH50z
bsUe70+o7/rf4mjksR/rslz1LTwtRkA1/kZ+qiqBbbFBS/CjAwaJhvWmG9ZAU8V5EPKPVVnA1hs0
9KrSbwNRtqWYsLTmVVz0Fqh9QxsjQUiNnH4qoCQr+UI4r7f38SPAvAEjam1pTb6srg2xw7qoEeCB
hJXE4QEtcM5uQZblxQJDkSN6w4r3OOld7vqlvN94SuXe5fA4ChTW6zQdjoTFqThby96y3lBJXmmL
lF9/JvHguig/VOoBrn9YgBJ0Hp8hldQazzTbxSGbYleKrxHCF5T98FhkpmPCFQhvYJHNBlgtOI8W
45D00NxT/DYwUeQJYODf6EQlQnIvVVcGjaLp0DWfirpGmEg5xAdV9vsfsNU8V6lh3RL5+fXCzHni
6DhwROq5TEWa3C1cDQrkxVsyq/d/Cy0iO2o9fnuCAUdlVZ+KuDSm/p8vZoZ9oRbG0izMOZ9H4i3g
mMRQg9OVph/wLDmlf6G1ecQiWuJN+EzpiZwcDpuxY2OIkVeXpSMJxe7hMlpYub5ilQ5tbcXU2xMy
CljS992+8xOooBZgy128dtPw/luQPoZMYI7PCi3T17MFXkhGJSAx6QjnEkxNVHf0UXZHBuqT0A3S
BuiwccSCSsNP9ynMjQVEE8XsJuxfm/JYCIQuTUy9lOzuie5vB5nFPbdB/BwFbbczsInlwwp9zc4V
3Fp6DNkNV+JxmM7tgY5U5ru1dau2q8+lrzfcFmMcp9CjhXMxffmCso1PDwrj4HvjwgmXmIwDIczW
FsYMu5hET2WDWAA4xFgdxTkSuAF6Bb4D164GXFl4A0jLTQWmdMCpiOND1qTFR5Bb6ncL/wMbiVbt
GXQehxyX2t0de7ZRC5q9AN9QB/Sz5K1PKntDZLeVTPeGLUBrUMJxTXaDxh1dDiVp6Vy0h7RbCJZl
COpBqIkHMh5NQhouoi8HGNYt1KpeQMsIByAC2+LPCvzrJye4Zf2+oMub2SoYuzi00BBo3TesDSfB
yJJG1qJu6hbfEHCAetlLVUw6HmIZIQc/lezES+9BCIoWrIXLDews5jwBrWXbcr+vloSaMDvsJtAr
SkAZjWHAQcbS7lVDb6aeQXM96MRRnljs3TgG/r9rLSHreZ6FMtcZHNhhVejwKqF1uRsesZf0aKnR
ctGeVeN0LN3y8vNQebCI0fkjG8A4rJOxurZcj9cnUQ3u/nV0Kw5Kw9Z5GhMhIBMsBtEf86d3xL3N
4KqyS0Q1RzAuvm2U+pUVv/AQtLMjftX2lIEKRx7Zg+VE1NCHm92nzOKpU3MuGFkoEpWHIDhhEltW
4+WtRAIHec4lsfZtPk0WHuyBrAU1tZlNLAEU9no8k0soTpL1l1hNUOQVgOt6nU1ZvXMFEINBcP4U
aDGT0qaFpqA/Rby4ZfBD9T8ujt1lueqHN3ugjv/f4uw5JdC8G3lR/ckaLjMdAdxmmAG+Rs6hwOpz
iMbT4PEutYXj+ET7gpySBWkhgUsWKbn+Pwnvce4G5hjQDUyQcY+dSUwT2OaWB6aLvn1rNMxtsuNB
gUN0dZ/Fr4hwTuu+II50QPAXGNGatydVTLfdHJQ1REvA1WPZFCS95lrL7HLjv/l24QxMb35s3Y+F
9pwlAFy7ffWxDhOirxNZDG184A3LGADp/+XL0v5AVqrg/zX3g3U4BLzoHGDTN13oqev1aGsq7ObX
XGYB7Dxzn79/57V84f71fwcpMWAMQUNoVg+FoPEBV2CWyCA8/hEjEmLfsN1WFiTrAq+Ts3kvcx/D
WKW1w4D4WH2gtiFJhJqrLB0yTzaP/itcWtmf0hDjFagCEg/k9rhFvW734/LoNbcFGVP/RetzGT8a
W2bk2lMeKncIOllmueoDN6lVZ6O+G/F+P+TxIVhd9mAYFVYupb2/wycghib3q6D910ZBw6tlDqvx
jeB4nMyev4NMrPI23tvf2hGcehmp3bxjjXNLkjH3jA9HIRwKiLgv+vOWV1ZzVB4gA4p61jcUOZKM
2PiFbw/S0kbgDhXS7cjIK8F0U7EyMBylS4AvzIMXL+vYABFhXpt+xNLTbMwZPpVjXIcSKUfkrfDe
iFJm+Cy6sVqaOHsi3owvmQHNLGTpDe6v1uf6J0wNRjjIA/RxZTFaF37RCjzW1h3fIWtZsZlXZAEI
OgIVrF6+TnNXGh7NaHQkkIldsDDvt5nC+TB5BpZKO3v1Yp0GqKE2o1K1aiyCiAl6iimRbacdrT3B
+DzrOq/yAUP+AA5cSbknD36SSk/tJX4o89QJj6tDTxlqOT911Lsg2nuHL3dzPxre0GJEsZzrqDpb
+FfUfCWSxQCB3Sal/kIByuzcVNHCtY2GUeqpn9avaKWkPzHmaUxaCKzuNFrbIvJQ6x6ds4dbB9+d
a6ZbQECIb0Pe57IaUDAuybLihE+yx3fHckTgbohacLlxNke4jnDdCCXM24ynmAHmRINClb0feLqL
U3P7uoydY9wX6Xx82bfGm2DJS+ylstAAVWQ3bLjG019fANs3u718uqJi1pYHxH4iL6+tNqJmf0oO
WzXYQ/sd2JiSXc7BI0+FX2b9u1PH8+BDt6xeiVYBi4Ij5/hMx30eRA87QdREpRqP3/N4a9u703oV
e5Q1mA/OcPpi2EZ7aK4l3D2jJI2WfKFGZeIhcLe0e3j64nydqip20VTiUqtu/uTElJnuiRprEJ65
F8gXiZFGWLA2k7egDZPhWfSxahIasQM79ZSzje57Z+JtSQDEEs1wZs7M7HwbangEgmsFuPmkqqwA
6uFK30PATadyvVeEIzlHkEO2iSM9QXH22s1INXaJUmw2yXweRd26AoNsFm29tnH10PlPeUnV/f+u
PH/aV3AX5cV0SpXl0n4pGs2UZinwmaRydyjtwvRJQgk7HHmyqwQntD+r3wcvuh1lfGcrLibG3dwD
4Gz9TrWsehZYQM1TiQ+7ECa2ps2nIkkbgGvG00wKzqrKX+VEAe2eeymVfIE14yccvD5zweXLtFDY
su9lMj0Qq8depi1gVgecy61qby/hIckMQEyNh/ZnT703cFD9N4m/NAz6x09mz7c4XzMgndux39ZX
7lYsBmhTWTkX8TgZ0eOQ5m1eNTuuMTM8H+esqrDUNi38rc+ea31yqxa/bLp/z47uYDoWeGLJnJpq
0yzL9GA+XfrXvBWjaeyyzSQvdqpDcnio4yfVxEl2Sbw2AQSNl+a9X2onrRtWrs6x06OMsRupDCw+
TcR5lHGUI8JX32ohT1bvMlWgNUt5a+3Q2AaIYhaEjKZycjGoTvp84bUtw0H/MKjR7agpchnhVOaf
oK3tJr3kCIujrloCahIoign/l9UTkXxwHDsijUitDlXG0sR5jpUFVH5pPvmMeG/wznZ+f9xFhdmz
UL/2YzECKqLo19vvsEWGObpZj/XukVDrkHo1jnS3hy8+NXtF29A82Wz/OISkJxR7pImJjSnc5Dq8
LtqYgv6gRggL5MBfFkHJfHTZ9uoKxE9KclCjJ8B7gDqum1/8T/pzvp2UDwjEVv3uol2owFM3k+LS
8uZ9frZe8QXABMXFnY4lNE4SdDOFquCwql7jNyt/6FkNr1cNU2Cj6Kjede5uzXxBA9clM0Bs+kvk
2JDVqylJKHtGn7Ikbe5U2WSm/pUXxQ9RwRe0oBAUR1hMmU3iz4A0PHzKVIFbcUq7I/XFwnAaIf4v
f/6qFBkpEqlzazUX1mEbPnxUCV/N+CfMZ7qBsdBTNwjpiGwvVZjOWMyZxZBx1mpXM+mwwx/JnI4w
Aq7x4bJCTAyQV1v06SvUuGKxFuSrOqpEKJM7uijvDKE2v468+Da9v3txxemL38fYvmiE6jSU1dNW
4oWwiYmXZr/ifa2Qwwre44uYh+6rF43LW9QesNMtMuXWZqkPUIaYCdXfURSQs1EKN7ODQoD+rmF4
IgBnM1sfqOptbeunhMrrxlNx9K9dA7Bpp/yYRQl7GdKPyq68VCAEIzlC7AKtNqDcs4/psIAdl1YI
aUjKUwMESwXVFAvbcGX+6vm4sgkrDCCuY+zzlkYdGYAojp+L9I7Z3MRRxD4wa30L7W/NurkJ2DV3
BNWsi1OYkXdxXrmNXghsdNZjDEYmC2kFxpPs7uJJPScBagOwiuJi0UilYGmtVXUBSdZLO3aa0Qif
8nwl6ZamY7Wy1rfswAr96Ze9p+1Z5bQzDO755/1tBiY4NltsdnCZiK5k2IYWV81JD52c2UTdOA05
mkKmXSehD/PP5NzZ/Q6u07DjD7N/FWpCk///pdjifRiwdvQmMjy92zjB6ALtRzmimklEealrnjpg
WpRfZqbrlOBwL/1ySp98Di29BzZKt373eDxJ1hwBrov2Pq44G+b1mrNFrc/z+wRJ8Hv7F2MzxHzj
W6uIGMMFK/JIoTcKpqjbXKhb9dkz0jAUpF167LtKcO09LzC4ELHOvISFcx9/M+L3sDNlpKrysnHD
VcxIi98hLUC26wec2muzSC8dn9VQapKnUqMkJYG+o04nBeXdoBvjHEArz/tmaiUqj2o6IhwiaJ3w
k4Pz81+zDnQ0b6AzCmqGwb87zDXi21CwhCXwkJB6pfx3VAw/t13925qzjWU8Zb82XPOj1oNH3C8i
u6Fy9uXmtxUMqSc74f8u9s4KrCaMMNmlgLIt86akK6+Gy8O0m301pFauUckEicM/TyGxxNtb+KJK
cUHn0b+cT1WgaJmWJ+JWxJdsGFgO/ZuvvIFf2xJAQl5t+k/Bvf9mkxh27/AUFRVk1xScEtr3kWgk
XA9J2CLJToiIZJaInbArel7VUXgrWdexygZzbi0njnDS6pDBqdcClyYCUNdh9ip7HuTvFTrT4/sG
Cc3PMGRRQ/B7hdTeZR4pu/mNUQIxx/Z2Np2U0p2ubUNcAs41q1wReqCeigzKjKcqZr0gjVGoaJa4
5C+WqYr8kSjTb7YfaAqXikksUa1K1wW3oWyRHMeRmJdJHHZQ0KUFMv21ibESVdts68nYlDgu/Scq
VR6cyf2594G71H70SBpATS/0nz+vsFyIOdW3Det8yKZTJDhzYOkWvLgS9DPg8r6mmlcp2Gxf3Faz
yetXRsx/OJafmppFM7TraVHu+lXJ9N41sqYQvXDLeSPnBUkREfGkuclxcPkhJH68IMCH73S1hQ1o
M/yoIdixCg8owru2yyL7zM/yhy66Y7qkOGZB+5woHaQchUB8PH0Q/Q04OdHpWjf3XL9uR26TYdV6
EoHzOkWygB7+F+1QRJGFma7pdXZQ/DQ25gdzqBrqgOi3u3nfwiZAuZ2T1LJHi2W2AgkH8FscpU3o
8UjsoLEcwy99Sd1GxToM0ABkxjafie8JZ5n4+sd3twdxwEwA3iTAVRI+aBF1MDZ1sK8bQYIwZjnw
1ZZy+sMQo1jAgPoECog5QSO+avj5bsdUMrLmBJ/lnfELOqUxpJYEOBh7R1QVHmD0xnM27rUBlneZ
ILDRe8RKvpRiblPHm7EijBqw7bHGe1B6jflX4gYTD9ee7mWljZLJ6/Zx9/MViYe/MvQgRj0n8iGn
quSyn4qb5SAXSyc8cuxzkN4oRHa8fDiHQtK9eEywPk1MXts2uwfZOHLm5XCCwYQPexFCV9x7qTE/
88GZYMASqJgLl60uLyWU95303ncIBC2utNg9rKOBYNof2SG/csfG1acpbzwycD7sFq20csDK0jZL
1twc7mmFkkvc4eGFtxjPvcqI3WH2SxL7fDONojxk5V8p7hETXN8cwZTj2xSEnmXYg33WGfu/QM+M
nDRKxPKFIvh9ijCRRzbw58mwhjEjHv+tD9esjmftCjN9W7Kg0ucCtplz8C6+aK2blj/BOIZABFCr
9lJjLs+3uMNhI+i51oL/hn8en6/AYheU+QGRPJcUVDzY70nmig66vUbJV3H47FvTFOCEyfqDdymP
YM6J/rvv66cQC1/uaY/ugcNmOXVO7Q4Vut78MKhGFu5J7VPa7OogDbSHdaS8760r/aR+AiiJSxgv
TfASydvQv2l0ASUAk421N8eu+NrrdPBxbikKtXBuUxumgm07N6CRyZXNhTLndWRDeFW+ng28jAwE
XG3qrD2+ytYskS08ZDBIuDm0H2nGHBig6EvAgmfA+inNgQ96eZf+Kd3J9372lU3VNNp/2NH5c/lk
snvcsemAsdA321xkowv6v95Ebd4VwPwiYkge3w3J41ZOmk+/teysoWx5GjxX49j7lt3N+qxV5z+0
WwSumnZkTap1KXdvnBJP9AJWApVGAeF+NTLqu+KbbAt/vmEug3RwKYqa9mA0LmUgTlaady05FYfx
+Pd7JF2GqDErWCGPUJth4OhktFlms1bWrOVvbUFOJfjehwuSP2MFJ+37u5Kqj+to54UwNGQqacTQ
QMXYF1hMDC+e/XdnuWl6PKT11wO/wh4eRoAa48OdpYus33pzvSawgRMlrycx4oO9S6LdJ1o2loe9
nAlI4I8IVoMdrLKFKuiZPLe+oPQg1w6KdD1YF/BwmxuTX0GFZhpL9nWmfUoGwITmcIcdyqumO1ix
c5Cf3pUnpTUnnmNAAQcHFbTPe8h0xcK2FnPuPq9iASSAnNhNeXOImFQMbf8+UB4QF4xf+Qh6G2WY
fXQ+iKpd0LVtOP/BG3nO6ciBau7aw/SZdU6j/2r85SpKMxzKZ5bU8B2mwILPji/3p4/iQyn9TKNU
ugwEC6PPkUQxIsxQCVt5YRvcPQ8uWxNIC8wsW1K5Poh91iOS8ol5fvZTI3YFs9QxYBjxaRLpOF8q
EKVmlfo65AxhLg6uTjMb19I8F5jUX1zyot7vVDq+2YR0ZeILcH74ISxa727fyR5m1nuarrg4ccq5
3frmknBOe82yZJDvYK1XQr5VjFzvCeFMofo7Uc3KkQDqOHaif4JiX1AbAqrURENRTGABYOvGnS7S
TrFDGg8JiFuuawGooU23nGNNzL6JHg0c/Xbe13hToMIhJMNGCILhmZACQF9fn5VXfoMid/brR6CN
LPqFy9/25RQ+xuDdhiDxynmBHL496ZQ2Uztu9Nqabmk+akMVNtKS0+5rNglbrKnA1YIRZg63dtf8
wu35kh6DO+/E4nRkVtJgiO49YA9rIpju0j0GVsW7HlNnm7N/+rS+iuwR54/qts7baFp+prTlcYTV
LBb84khcNIX2PXNfVHMVW32tITKPoqJANT+D52ar2cdwEC5C2AQ3vl6O8DTLFNQDkU2QP89gni3F
qS8btkNiLqYj3pFakmx5bv1Lm6WCJzQtCaIg04UXY4NCp+3MWYVsT952W9ukfdUez9Sc7UPN4p0o
yuP/BkM3nvFYEC0KFtyYsRcLxpEGJqpJSb+wmHlDpXg+Q+sIEsZ97HpdtKhm1ldZwlMUdpe6kTeK
EkEhk/sE/Qwi/6aOqmfz4Jq9/j9dSk0R29OqPaK/JASjMWuITG2jJfMCNuZFn53UBIyPlq7u3N2E
AK3hh44HFor3QL1O8eEwGRrE1fET299cSgYzaFuTotslBq4mFbMfhv2Z0yfVAN38jzfP8w/Vc3Uz
XnJ2OAyUh0Krel5iJ2cHbWVn9WuNMaEa3A4KB1kZ89MFPCMqzHMtKdxqxufA124+FESvdad3jgkY
qkRF2qDUd32OSZb12NS2wKXHqTUyHbU7r6N+JjueU+nqQaNUEla+qM7W7t8XdTmdS2mn6iUbRYAR
QkIRE2C2hY+NLh6csODbMQ1EVhlzBDTckaCt+M1AQHmvgswMeUoeF83gazf/Pe4ZTIyzb+ByitiB
a3SMIn57MvB8iPTE1X4IT36lqxNwvtQENl4DHfEm8SGcwpdv6M8vx5RfjkN9iYCaJrroMLoRIJKb
0vSFYnEovVUCPDOSLM1QuKlIRgIMITbQCa7faXphv191IybZtLm1C8bamI8zuBAJheG1Qq9YK3zH
Rgfse8D6cTVxDintg7Tb2qPPlul2l1qay/rQwMGKD1L1xY3L2jwDxfbc4Xvxv3E43cPep+6X3xez
0Sz9zAQvQko5oZrosmCpN26mTwpkwRNFfLOfGrq6sP+OA+n75A8EvqxBPBgUFiLPPOIGR66MzGXD
fFqz7MG3RZ689JmTxjU7lsUHmFQich9IWXf+UFj4ZeHJC6gYE8oeh3cT6EoovbV358hB0PfDRt35
jsmBfuNDxGahATbP6rXTBkC/ppRKg4S++7+6yQKkBDJrGDhjBKj3UGmoXYxpHXjQlob1vkauEA72
GgpVkY15F+qtdiUbtyK8M2MS47Nqia7hQME5a2agM/NpLv65lWONQTBXTcJXjWKNR8bammo+3dUI
T/ZC3f+Moooy3Q+KmMXsBVf/o65WyLOMsFkWyRMI5s1QVeRTcNDyfEd+MvPT5Fz6DIg9Ie5wKQeB
bLXfoybEo2ppW4Z4ttt+ERsn1ntW0LJws4vWmdh5IOTjh5cXSWaaKjTPnmeUVPSp/OESPuhBpdrO
7U4K/EvhAmPyX80inatOHXFmNM5wweJysqKcGWSTh2WrVYjIKWAcOY0nZ1ekFveggo9RTPlwr3aS
qHV8fNBzm5pFC7teTEoaA2qFOJaYAgzNRXkx6O+0rvdUfPbauyfAq66+CYb31ilwU3OLufYRvWIn
rO2FfVhxOAUDS11EcB7AQ2im/f7wpEfKPDZtMbAQ/7PGanpuiSQZFkrVYuktFItwamevyjpqVuAJ
qNxSj02dgYls/q7lUf1j6mpyJB0vAklCvf996eiZ+p4hzrxsxQHnNgsek/GTesjL7pxG+4DWrZQ7
viF62tVZHd7JhvS3brjy0/IkpLC2JlXExnuDw5SgaFu3IMQom7f/5GKVJL8n3vZ0dsDNAC4qQ7xA
aiG4QCpHIm61/aPNMSucJQ+0bC3xyrieiE/KWcZUyc6fu7s5g2fJ+UK2v2ItuUudNua+hIDlAQrs
bHaR8ZOo5hwNazXi8tN5L2QJjg7juRFCOYWv5eYrclNWifiQUvYIH551EL3/cBOuIgnbxo68ef7O
dxb/g+zEm2beQY1+I8fSyNQ8U+aSTPRhy3vVsp7fsMJVZHsXGsfRg+F6FqXTPYd0S9nsjDIVbPBN
bdM7AeeiAtN3F+vUgiQTMIw/UAr2amRm+OGag89U6NTIDEZEqMwdTwYeR2/xKyOjBkwr/I6CINxz
cw0jjltWQSpo1vVk21MSd7h5ZxNJaPU1oYRWJqKv6hZZZOexN1t+01qA9C0UGK1QQ2uantF3+Ck/
PQ2Mr2fPBCKAww0OUZgjV9E3U0Ct7DR0TTv1n1tlkBA2ns+6kItqUfK5JPy3NBSJpyDC3Aj3VVBK
33HzcK1K7DpPGlr6RUc9MGTjHK12mi6ky5tZVdXhCx4TX8ARPKDbpjjc8dSH2hXEj30TFinrVLHB
jkEYdIndvXTuG8JFvTlDK5utL5glJAf+RXUa+wapnWwbxtA/y66DjoJe+OTrKuqbxwfQEdfmg/8b
1W0nZnqBkPd7V89G0tisj4eXYG/gEIivtJ46yKE/JERcOME7QoYAsMUuFsobqGghbot4hGGJGSYn
md8YWLzgTRmfe/v6F4wyl/3v3TdBIRh92bommIBbfp7CY5fFQg93j7f6Ch22tLO8ih7YTx12nrfZ
5l+1NI3DkTC6grbN8HIeYL/AiEi/aI0FZwa9ZMoHIJPLLdhfeEVWNPWp9vr8OEJY1FE5rKLUlqqc
BK7vTbbbLMH1ma+0f+WBc6x7d8Eh/dxQR79K2wWam0lnETQR1eRyGFKjWZFqarIXl4At29rwB0Ru
q+WkrgR04D+I5SRgyhFHJl81MigqSHz4CeirZDkHCd/vv7PqhcilDjEecNQX6mQSU2Ayv2QNeUJv
o4vXn16N6hHBwbvekYwAY8bBlPjkXwpHTYNgShRyM4Gy9rFFzyR+PujkCw83ArRe/XUw+p1fjBPL
+Vt2JTPR+BYx4ESZNpWlK1FcPVwhvAAt7LXrHesTTfOJGcoB5qHGh/UWlYXWpGZEeUUALzifLfKm
Ip9f5pvxvD1oOt/N0ZTAjBvO8BmAT5ZFTvITqBKPrEFbp20DI0FJAYfNTc0JNamf7vrTE/YtCgdh
mZ6Ml9t2ix589PFObZFSC90gh1qrHMi5U4KB+HAR9pb8HemUOgkrWWyTP59Q2SOi4j7Rq+B6xXyj
mHisBfJzP5KB+FqLWQ8e7ply8KEwQy4357pqczYhcQTJiyClrwlM1PlKHrz6P9/hnu/2FvwIjW9C
NBI9JS/WUoTXUOvJaJnJozRFqF7yunLQmwbS/4iK4Rk7vdRZx0xqD3b3+R0RnrDzwsku2EFMp7ff
1qP4MYY9Dyyh2nIzfVrtG/0cFceWAgRnwFpG0SVyPIfAPUfzhIdNQ6H4X2A0vLU2BQUzk4NeREVz
8Kl5eTi0q0DkgtPYq4fsJYufjkspsxlsJu5NKlWz9KMp5EQ6m2xXNXCCCwI5uYPsJj1o/VnnKqzc
gW4bkXzduj8RiFxriwIVzCSVa4dq6ASKekodLDL/AOIyXkMlgU+w6w/FZSfQoxr1aHcWn1Bg5EV5
e8jTwb9uzPbAYO4AeTP/SyTkouawxAkq2kec0sGrDCdIxYcUt+YvItSPVVmdkzlxtbCbOXr5kQs6
fwOUCu/G6QfsapMPg18LwYqryQuN/4+S42Wpo6Ag7r+iw8+EsxbIAQz2CPcBhSSOm4VDPK3b3hyq
mLD5N3R21utEmAPAoGbZD4F18YZcMYsDDjBW6buZj8/v+GOD5l2PNW+UevioUyU2PbBUsgaQ5sSG
CYoqsDOsLV69Ga71u4Uht7YJBVyqwk/b8dHJ2h16zm1+N323yRfQ11Z+eqZioqhPnHoc06pcrHdP
dkXKk0NWQb0VBPPo0cEVNsKQozOm8y4xoV1DQ4Ysw7yrzyqJfKUNcPmd6XDOeOwluqpuUdvhSGzQ
MFadxWXvoO5Cz0xbLHcc6iD8kQEyN3vSZHD5Jx769DJihlTRu/63QvfeelixZgUwiXKnY3b0/2mv
M9ZN3Jez+fQSQ0KxtJAf4Ev/gBcaD0jcrQ5vr0MJ3l8K3LrP74t2X/l3X+CZQ/ZcbduL/zVCzLdX
NrqGEO+6jlzEHgGfVZ+XjeZeLHNiCsROKxKIISJ668qMyLzevKaNkLfqa86m6JcsGYeF34iFFgcg
KrEOd59amQxeccrP3/quqc6O1Qt3uIlPvGWd2iYCYPOzs8qlbn+eYoZEnL1Mnaqwf/dIiacJcYJG
03tmpmtQietPsWn0gkhb70JDASz2qdOVOSVw0Z+0aSy21S2sXc4j1VcoBqUs1dSoadN4C0g8H/Xi
BKDvDtOrndBVTJE6RZZo1aZ1/PUVCVypcj7v5oZjRF2uA0zuwXGSugzvt9A1tuqkhSRXm06wnj15
4Xny7G0jY0lmxpdAnRaW9WiNZ3JgKgp1JNdF4t3A+1O5/9PYyd+7IeX6NFrWaEXUt6dzAtKIHAwa
16w6RQBvYYqAt4gC4otPoC/4Q20iJ/po4/PsR3OTpELdGaT2Gr67hutAlL5ED7wg6HV0lhz0Q6EU
5L+E6GmNlMSwkIdypT4WUjMIYwKaHPZ8KcPK75Nc94l/GpHaI0g1J2iSElexeeVhh9aUU9QhOWuv
S2Jji1aohjDdwEanq2Fu2XcE0uncEiEBRSwFEnJOsjAKr8Jp2Pd5yjmsRIu4JhNPMsN8Nzbp2T8x
vHt7LcCPlX32kLKFTqGWESYHp+v5OPb9FqnNM7jkOHot/2SKvnzipbKwPixM83doW4YhsZ0VXio9
gtqI07pZhFOQFY3uii29Y7kwHOfkU6K1xP+Tv09bw5lpH8kZx4oIReXeEryywK/d7ZOXRIhetiEQ
BAXj6TRytaOwAO93bfy6W659PdZl+YoCyn7RWmgVEyASjJLz0mfmx78dtcFwpQIc2BcLpMnHDbzG
rKYK8aj2XXI31VK+rvhB2hnLshGn00/DRRpq5ZyuARHoVHUyLe12tQ2+0AyMqDZJIvIk9/FcIqeF
7yHz9dKupqAPk9P/cOXlD84/Pk7LeEbuBxaB6eqFWxRxlmsDCjbW7V50hZeOYkYs20pPGPqmach2
bBOj87zw6zRwkPPD7qvwMWNmslKTFYZVbNc8C/z32Z/+RjSwK3Qpt/WJlZjmI9F2nffNDRxzoUjO
eP8wlPnCIKRH5MYgQzD2AreCVhNAW0Hjq31z3dtxbGBiGgnQqAzQWOqlg7iH8QE2yfPochVhOD8G
LszrAjsX7C8X2ngoULHphVYYgwQL1Jt5GEdNkpj6zJ53cQkU7Og7R/K5NEBt3Eii0HHXXfU/tcZL
Q7nkIV99NS7C2B6GMbwSLHKAnt9Kij+FI/SYujl0M5bpmpQGlk9zyAMHbmRPlNz6a3B8Br7MxT6h
7lOg4GcVq7rDwXbeWPGcfaivRWnJzEmA/7Wu+hINCLhwTgotZjA02QFaTJoy9s4L75GQK3HE0/Eq
zo5Ux4GVZRvsYp0gcZcFbhlB4sdHrBv0qv8Z6L9Hvdmg/cpng8nkEWWOyUMC+pyI3roiKh3aZQMI
pJjAcoT2cMgiSv/K/AfqYTdIKj6SvykwDZ3esf8MxV2BJzlAnZ7Jc7FdoUCwV1TbtmeZW9eEO1nJ
psBcQhcAFRxf29D+tEow8ihmjhiWElg6W1yXOcpuatKDS/L0ZWq0qJmy09LXdJJqLb2z4ioB1SUP
AwdXTM4epONeWohlOEue2ioVxhb9ECaT6OJYT2sUmcNvVhO1rgG2gJUMfnk5buLqPJMmhsM3jOfA
cB3RqvD17PAvjGxNvWV9rp69jwvBsDr8SvuwFV/NgAXjT70jl7wOSKj11U1E/bMEcV+OFpvEJjZu
Se33eycj5h7lZvXBz5ifTI2x9P8baTmD01sxAc/abv41rw/rfPtR6YWl8ChT7ITmfsvFjVKdC73r
lKdoXXRpI0bhdjAOXXx+e0cy0Kmsa4fUvz1s8aBfSnb7lnVVTmXSQuUkEVgd6G5vRZioGZZ1Vpn4
722olHHLBke2tBr1pQfH6f6TxzqoRRG58fDrd5mB49KRmdwKJv4p8ITH9PqyX9tIMUahOazbZWyR
Oh4+PRlcd7/FOeNb9FDG7z+NcP9IF7QKUudO/2qzXKOupcvp73gasVG6gQhOobsFegZJbqNuv/k3
Owjrh5sTjhkz/o7RG6lNx1TLf5KZyQxGtTJLVpkjdSZbCK4WAg2csrtSxoqunCCdb2oboam8dMwE
K7lbXl4FpQ/g4azQXD8FalM2KCZtg+L9FTGLd1xvV5QuxGtGm0iKy6hy6yRYeW798FjhSqdwWbC8
mKL6rMZI0aLHNX8Jwb3BxDorrLR86pk7EiyQBk2yLyYhexSp/ZA5uFQOPFC3+2hir3rYGPLt7uiE
bgF+ZAAtGjk4NZs6NdPbAcUKNbQBGo8rPhWZpGC3h9lVw6h9h8bfVsOJJkIGowdzfc5DEc0iqwD+
kuzsq4XR69A5nsNFTT+F82BiZR/ieHAbL6YB0KlBrft9X7a9736e6vybtqMr/XZFBjKyuziVWR1p
M/7ths8fN0KtpBPI+yzw/oZisDSHYwJVFZn/MOtdlPbcKGJBKSb5Nu3E48MwIUhIHNNzlO9Xvc73
4Cx0W00axajhxVcC09ciEcsd8/U4rRwrzk7+9mt2q60iX8kKf41CVg/xmTA3S1QIRL/0sAJ2JUJA
xfj7yrDq0+GnCPMC8hDthtnb/ocFg/1JCjs56YPZSQa8r1FiULCiBscvmWqX5+s66kYOwVZ7soSK
PhynAjdtC0cGNBsXMH2GDn2ZUn6n+HtSmisLQzkc64JUWcMfgTloK3Ekihc+GqShJnyJODorYxDy
AgqsijfNa8Xlc3JSEnfAbiOByBCcWGT0iQNgl5qSjL+bSU40dkZ/Bvgh+deHTqJ0Uhn4DNHA/8gn
0AUHyxrbQIUCMeB7UQBdEa29UyaX7kHtzgwD/YmCN8EnP58rtTS4W9TUm1+5b1BtCtGu1Y0O70nl
TisxQUR4e9QRd4qTWMe6bNMXcBYeius1Bf1I+492Ch3tn6ql9PaqGGl4OvvsIjTOXEY3KM1i7mRg
EsA/75NlrKXAVEN2oRr4ibcmkUUH2AiNJ/gCd18h2SzSNYAPXCnDvEs/BaarA51oBlSDtYUImOSd
dKNn6nDKAEUnfj/F1qAcVIZpveabXI3QqD8VMSQ0d/NZUyoVmxcu9CXJvZGSxSu/28LyFOQMh2mi
2LMRncYVzQFrHzPWe74G51/ksNntNwfq51i7qZ4w7wS79MDcRE4pJpphoSyZefSxOsZ7f2q4xwf7
Hs805l+dPp82HYCBkgJCX/bW9J/hSYU1x3tZqXca2n5rfKw/SVak93gObB2LGeyxb/VRFWArdmDS
rGeyWlWbSWWjznPXCfu7yTWCr5DaoPMh9YMZ/TiGH23Ynmqyc97JgpxvE5Q2bQvoa77+telKluqS
w+5I+0CVSo22LUCAw041UtRbB++jcbSApWytNSrlrZQaCSP72AUAkpATwviiRi5MnPws/TRHIUo6
wTT3VoE84qbtSEmxawBju7l9UB9v5DUZAlw9/mCeb48BxeMq38kzgjHQhiXqeg9YFtqISW1PMtEW
PrmMa4Y3MtI8QZ6G0rPA9yjLhq6xLHHMVi4Gsp6CZznetGpVDbu6syOf0ZesmggdjLepqC6g0AvS
NEr9l2oUNFt+Js2yrLh8yEH30BE2XEMO2MmUE6wF0otsxM4txPUoCdclJQpUDAKAvOseshWp737L
eJPxCDVvsHO0bzlOg/gwk7O1AYZ6/TGnO5jF+ijRCDUIzWU4tiPutKkjiFUaUvtU6hDXah3RdxQS
iEg0QvRKlzpi3TOpkW+Jp9YAQEQc31sQ72hVOeCE3x+UaX3Kp4+jh7VZEW9N/wSbn/HWX512q7E0
DRopyxxby9FcQ4274+r3EANcVm9374KsAvBIUHM13vnegLXNqDMXSjZpEizI4uy2QnyesOvpquqh
XI8v3X+g6mcc9QCZhVovWdWB4iAsykS/VNBeSeQnB/cxpIhd66IQepP4y8gTj8LKAAu/OX1e+m+K
4rXGqh+O4QwAOXyO7sAdldUUDx3oHhuyXaXIp8Wt9Bo2gMI8v2OqA4QaQ5JsAAygFV1rGNczmM22
yuA47Evrwsvxws3kTg5El1vVtDD/PCR62WVlExZ3uyNAHTIjwA1r2zCkjTyi/N1ejh+mI4P5MJIg
kNq5ZmEZVPCLFl8oqW4N/y8JCfr6Mc/k3WNwTbeqKMvjxEMUNrDQGe1jnR7E3aEhoT1wch4cItZY
w8vpLpPuSw3hUzCb/89lm8sfaPWs+HdBXVi86km51gZo4PsErXWmWxaytWh1kxeOyeuSM6ER+7Wf
EOQ/dxwnL6GalWFwQzy5Hc/sXGmNlr6fYd25SjCpfVkt5Qiw5SePKxADknzLzq1lu5IZszgavKrT
0MkAl+TaGRvBJo4pjdCy6xBGDyMVx3h+4O4kXLT+j8xoYcLWC5O5rS3Olc0Yb+dvZbPJc2a1dk+l
sgN43qzExbmeOhzO/CcVKLS7bB7WaXMqH4aKQ2sUg7Br87EbB4dKdDNqa4UkCF24pnUpNDvvqqjC
fMtba6ai2Og4P4SS5wdZxkOMF2L+zsQGfvqVrDo4Kd/tKAR6mHFptee/4RZJyGrfgHwn6AVc2H0W
wmOBWDjGhTknNXnqenJrwC0a7dSNZzhntUwL5kNWolcMhZrtJhPCtGbiZ2n15sOsXkBCC4q7fYZa
Q8FGUIPya5Esp+2LpehNkBLAxx+ZF6bTZlpXkmRVkUFO00PzAF/59q8MsQ6LG2vbYLuZowKu6qw3
u+B7f5Dby9N3UzbhavCWmTu1kejjCfbisM+zF+lpNvzr+iP2CjmaeQTgPQ6P2yQW0CktuVc+I8H7
bbs2pW9nh/FsAw0ZILHAc3GsnfCDcEKb1+YleFKbXQNA7NexVHPKnXPrEVE/wIGcAcv7tu27Jbt6
JfqbwluSGiQAdjH0l5+rj/ZAxUFyNQwj6n3yjfATgoVUYzzavUTLd5AgTHvceQwdy9DN+HVRd31V
g1RYx8P6ELSE5n8D84yGbLw3nmeNqWSWivy7HAgbLl1DyIEg0Y/N0Pehmar8g60NM5h6b6PKMaRW
ZSkxtXZo09ruHIU6U0mnX07Q17VPqPabDaW1rujj1m9ffC78OMOesJ8xQsSAEYl7yx4/HE6FAcF4
0pORN46sJV7nm8zz4+loRytS8+G0V+Vmc3Fz8SkF+HL7zySIxdvcJN9PxIA8jrmxKq9vlTprEOwT
nSSu3eMkrC8pTeUiTYOOdRNaEhpeG6D7MxmreuAoIH6V66tDzAEvxmeQNvNWbPUavj/rKuIudJbJ
QCbdDZU2DBHROIh/PftfLPRhOIk5+GuD3spQVtFRzsBIs/GptQOTCHa4MNyKmdZIoD1s+Tlum9N4
UOLtzWtsMXUtVkQNKGIW/KLr86yxhg/0A77OFASfcTnqSQt7C616mATiDmjM+HzOitnWoNinCOPV
vr7+4AOpCBu2skpcag8S1zRBrEyECJ8T2/nKDOpLB5jhkF3mtOxd3hAYl8qnWUA97SNEOcxU+7DV
aJ6aUsDMPs8AR3JxIGWIUUmkVXkVt4Y87krAads0ge6HBo4BWhfxigbS3mQPQWYB+exMEw6Q6Xer
iVsrii94J4RUbSgpEqivlimZ3ablHwFJ2mg+7ifJ/dFEskwdEWlyH4QA0DhXTff+ey0tqdmAAPGF
Pe1quCQGKy5gD0UYt4PZuaBs462IUs0+2huqy5GnR2KZkBAQDFK2Q/3L8cR8dFjjeBqx2tLSMLFA
PRJeHiGJEkTwXj20ZHKjRXDTUCkBWtKZ2XYmfce3XekOIBp8KU3m96WK9/0Jb+SnQg5kelGnb+cF
AP2irL2uGAxv4H1mLcrty1w3+d0eQDnigNU4cflIo7l4j5QZ0gK3AKSa1Ks19nmHsFpWQdJOWLqB
EpTi473p6HMB6WoiLJV4a1flxpLNYU+JE3619j2Qzld58y9n2dNRD36TD+KN0LvDWjCdcy/7DAVL
+3wEcSs8r+VJ6JfpOzw8XZsXBHMaonEp6RVeJJrvHjG0FiI6FNY1Ts31sLULiSkkaltmsJzxKEob
567K80cGV/jDlCU/CCJ9B+XV66OD1hsd+nNo/FBVWMhjI5irlUWfgl++Z+EqX6EsyMeMZmsK0KDz
TqQJFwuOBIGNh4H33UclVSXOYwQ66YFRu2fGbSXxvMnsWcscDPFPAy0pAZBCBgDbWqXlb10duyXz
HIMjL9iPhUNiBjgLEJn1ci60hO6uVZhEXYTuRJGckavh9LNhHDn511mQ65eO434qRxZ8Bkvmr/p+
ak2dJ1HcyiErDpPy6lcw7NkohaLs68G1krozAefM7L3PjK/pbdJJG1l1/T08Vg32fHL+t327qINo
CmKZrh9mfl30s9Y7fQ9fbrNYIRp+hn6AYa4zNQ9uOngExzpBOJLx8wWrehrrp9OeFt0nd3reIT2N
8TgQAjCZUzb0NzFb8H+FHrd5PcZT5ouREfPKnBlqqTVQnGSkVvc1CnI7aJRToJZoVrjePlpUBQuW
eCzfr59vqJeIjQX3VgYsC8J2SrpPj3tD+pFN0EgO2Y1dTqg91vI/3CDKf2kjvDluJosNHR/dVpG1
Whwh4Ylv50YBc9tKSNqQVVpJvIx/POKuXQhG/yQcaQvsMCkxWWRawtKSzZ0Cqpoe1x/XxvErIdoc
Kt7btYngAeOd9jqbwHOLpCDsq7P9WCBZ0Vv2xXNMUgIOy28D/fHQvbJbwYghJocjIUwqwpa28/OD
23JF5iytswBv16JWXr50qv6t0MnlkpgjfjZg1dEn7H6xsLgKQdSsYh05ix0NTSjbrS9gonSAC6+Q
lY8wVyKF0SAN94gt6tnc1k23bnNlIohIwG9+eTmEAZQjBXTdnoXzXsbyUu+bWIseL5427l0mCYgo
vjqD3QaGvA7jDJVgpPppZB6Z4poe/oq/E80ZIQ++O+DTKwfUaUL9/u6//+cc5eSAkf18ConNfEC/
YzCmNaoA/vt3JO0fWjP6UnyhlPIsyYS0u+4FhZmpq7AskJQbn77k6aujsT7G1iOqe7C3ucBYjFA6
Os/1NxFPp7dvZwYt4TnpIcanl6lAeA74XtjXX9CgiZk5nknShuz4w76BRSYh+pXF9hpelZUJgsGh
+K9p/5GIIgruZQieSekntxa7M9t+zUO09U2qD5De7hKpZH9ZbHXHPrS72hYzt+Zc7q3D2WQDBXCe
sGoTVPMl7qDZXu4HmI+c2hfyN60Eke1GfMlBn5LH3frYBf2m6JTnTAvRyLo5On1JFfsSYC/4FxjQ
y2rrF4KXrGPgH/h9lQDCNAhU5CnEO4KYRxMiFlkO/RHqLR4abOPk7q+1NgROw+QjaeTuUdTULESb
pYq2usoggdNmseSyrZJBabXz3dYpAdkEyB1Z2sOqu8LMq7MB3n8p2q09oz5+QvZLiLX6D9RNAOwc
/7/Ai9Xp7/deXRQsE9hUVUyz0ChyD4CCdnfBanCyku0PKGyYA/U+OspnwDwfN2Bayth5rDO9NiET
ulL09n8mHjWv4H4Fdb6OtgLkD82yh0DkEqaBfYc99Udg1a92XJBbiEWYShNDum7JHivTNb2TIAOR
RhNHuL2gezUHkNK475QcQyyssfDThbfG1bMwVx0aYPvgJZn0ILOdNCXv9zZKnJvIXY9hnodqV8gy
2oAXJ3iWJMVc41u32CoI0YoWGZz9z6KXDZ9IXYX/RIUMRecw1ODQR8zkwe0YWZB96N2gKVn2ClDJ
08T2XojpmX6tH7Io8DVY4zwYG4DreujXG5XbXBwZhYdMad8uzgFZPtau0GcezfTECU+d7MviNRYb
9PwlWx5oeLGRM2zr2wa8j6Ua5IBj5F77h9vlPqsR1gJO+PFZQWAXjqyBUgAR7jMZ1jrmAifBMe4v
nUGnRJ4IXDvzvXRsmj3BOiA2hRQ08ueTObbItWhzY4NvUTA6+IyhWzHiOsrtNvY3bf5hjRnd/rAQ
1tJjcUglhPyD05/vqw/kUKESxs0SzJWbLcjIkRZHfzmNAS4J3Pi637avfiDBEwKf4fZG7cfsLQT8
zwxstoipyPS8rpkOwSfD6pF2E9tkPnN9GpQcKU6A34blky2X81XfHhpIVRvu5M8xfjORa7Zn+/mL
FKUo0yNacpCAm2zbqOtrKBhxlbq1TUoCr1ThK5pFT4udxxuFvPtirtCimVzblZuPuzxXfjeeSNRj
fclWzNbOJFjIR0k5NxEpkk73K24LizJJHPamLD9DjPdSGoUeG+D36/XNzngcoftx+iGOnY4/DihF
wP+qlg6SAOdbb6kAPUiR1KpeEz4PCyCF6WhTmErEv9Rd5I8zNzcrVKD+k60zKndW4YXYNZ7HFcI0
In8MA+Zz5XGlNnsvRXbBni9mFuxrOOGMUa4RCGmwK5W4ZqdkecIrTbkFbG6Je3mbEAlKl7d1SuRr
l81so7h5/VWsbBbP9s3OT4BV5jwjF/tFYKug2T6DrC1jU3PpfJJCr4U6+2GjiQkPqIfDm/QWax/x
idOW+3YenADce/F794Wyen9G6bosXUrcoTAcadY+mt9QeUBQVWR71Sf6Y7hAm/bRf8O9rRtCgNR6
YaVMkaspJVWxPVvM9htkvoI5rfm4MhYxxBnsxrGpZ+USlXoR8ajSJZHw5QTKVRFsqz+IGWBTfzwX
BgAXeBGunsv7nLXMqq32oGrEMKBg6mhdGxp8bUd1j2AbrHmR4CnD9vrN49UuZdadhOCCTrqwgyDp
msU4rt2TY0j7SWxPYxqsrpHrYCyrpwX1vKdaPF4Y+hg3PSVhWlA5sgiWXEmELkBql5pVEl2rB8RU
zTc3kTZtoUjBf5hPstTAWlFkB9zKBb2CBGkD6bpXWihOCgFTTSaxJbGwBFWuNFZvXZb7CYLG4lxq
BrlKyr74zaxVbTfAuM77bP5J0EOKafpybtM09cLVEAOrEaIf/ZeH+1aC1cQgicR+CVJWPC3PHPu8
Z0/vkw/mkmKbHxXn5GV1vTvdWgsUk0hzBtyiHhoQwEibKx4s0h5uGlxJH9e6SaLW0xcwzS83Scm2
FO0DuCRPKU643PLumcRnZTXz5Ol9bjZ6YJGBKDq3SKOsRYPjJzpUFzomnm06XNEvNJwobJkMkNIb
wJ1OgfPjoAVt14aS26Og3vYSjsFfClLt+/ACDzFYrD9Exz3+WMLzsLO92esrByJ1sEaVYfaLPyPE
Ks4a8bUhUWLDWO9P9cbEWyrYz+FY9cD5V+XcCsm8AG2kpaY3K6pFiE4E8DtvW5e9xv6oTXxHP+nF
dS1Pfm39SHLauCF/PKNmBljnkILwMVswaEDG6yrttbuSZxd7Fcy0LrG2/CsqnhXoHGk2V7f76K9X
DJgtjqM9DKnk+V8TGcbZ9WM4S2pBHl4MZxhjs6hJ9B1eiKiSght2xhNqZIwxxosrIDnxATnq1ZEc
4uN78jdroad5MkiTpYu3dkiI49d60//kuEqfibFaHBvWRzy/P2sSkAi1jI7bJJc49jRtEA344GDP
shrpNocLV/kzmvK+T6vNmuxIx+17xLCLHTj/Kx08DAGUUZgyu4Y4ML92AezCeVF7LGUX2eGClHHf
56/JhQDYMzb3opEUQSm8AzpLVF8yU2jyPehgwytJXKBvdzPcpUSX04wsWU+F6Bh7lN5m5G7bpXLt
oT0GV2gMGMOCo7ngkiQaY/lL2kdGE0YuDWaEgkm+xKXe9C7vJLWV/RC5ZylQ09HCxhinkUHbSO1g
gMDU9cFiBS2ylOQIxyh2RfHfZqDu4v62c0uHU+JCMC79GozLeDYGsZBoSNu+o4MkexbR4GqHku2S
bqChEIzODls8ZiGSxfb/C6yOzsKfcVHm1LhgsQieNoYH+gqXuz0a6EjPy3Xcn7/KruwrFNhQI96K
UC19i09UDXM81VErhlJWvEdqCjHh8bUksNTBhxQXulZnwaQdl9mqHX4OGjkKcuFEthxvoLkTTQYk
CxLMuTR8e72jehJboF311oz1Ow5NCT+1QmXfQlYdWPmvdlpvJhcVR4vJu+3fhjz2+w1Tr465Z/hb
V8hJVwd9pTLI4u2MpppSfBOfu8LvSyiLOpd3Mzc3PCQbMoMNK/sPDOynvIQxTP4QiqRkS9EbdL2A
817NUAUCEF4MZbhFxb/cs0GWUlMD+Cf4iK6B1iVx1+s0Iwx7QvdwjdIuPIJyoQKDbcsrrNAcbtKI
eLEPZHbMVEw55DkfzAgSpQY69/02Ck9CJ4bFVNCoiJpbPbfKg+0C/ZBqNAoJqsp86J4y3KLdVeGC
roZCCk4c2tkGfhUFU/XWR9x+TQj/ZHOE/hFHCSN2uqOqM4mieHEOul+3fcYT2abDSa81ItyfRrNo
yFW10BwwEJ0aRG3HcLaLWr65d4BFPZeD96nA5ACJaUIa4FF91j4yzRfPlW5cKTWJGVLumwy8cEoL
VPb4+lDG40k8ozLSQU5g1Zby3o7/LrOSmNv36Hk+6yYnpaHP450VX5vwXmKi45Hi5Gm/KVNs5VY9
XuNTNfg2/RYHjzc91ZEUAOHsf8wMyg+LrHMfpNMBVZbKzFFwsqtk6BYXSGYXJqtaIuGiyMNYO2HD
Ionx3jHsmETEsQMgT1zeF1a1Wox8NrQQUKN4Ulz9E7oSCdzOtE0mlqfTeFrHbam784R2wPf++GE5
9F8wLnkrLKqFSCtJioFm0ftO24iqeN3+imCd+cS9WnuUAGJtXf4P/SFnH0qEtG6xAmxYRwOegwcr
7o38gi646BXrass8reTTrtQVIWWETwLp0VMSI2cgXwr0aoZak5yuqrOk7GNaEBIRwe1dkWo77xxN
cPpEWzE56193BLnHhf/piDxDhilXNaE5uFIee384GgHhHet2RkQLkNqdZ/ujNwvjrl/1WFohpfA0
nId3sey3+V686aVIzNVAfQVbSbHmEbVy8o+ULmOooLTEg2CqCPl+nrRqu+hGjJI7LwOKPjwkzAEM
OCWZZBr+OOvccXM0Qc+L8ex5hxVFLDyhKgfbrgXEMGswBj/9Ph1+nIimxJx9ABI6D1W0XRxmLLZV
SsDATbagMUvj/2aouSPC7beZx1oqSNuQKT0UKX/15EnJQpRF2GyvyVcXLQl6zZid9htL1SpDJmsc
OP0Q+83BkdXEcg6fKYcXBSZ7HpRQgnkH3vYWSW1rS9phbuQDV9FhTwsSyQAeLtpq7gTYDo68D+U2
bm0GridU1CKtXMoSVxmN6zteY4xj3IPRAJUyt7PG4RhTDpklavY9LoizgQifEKxOg4bGavwAtRrm
tBIlu2k3kqvEuc49nVT60pozzlakiaOB/XrkclLzXzsBTw1pqzHftXem2mEDuuBsqhrfLiMuUl9Y
R5X3ko3CzYdS60iZt/CYQWyEqEXVm/0XlRYwYyiKMuWDK1JSMgKO3BU4zB7hSPWmotRCWgqCt9hN
5byROblX3zsRk/fDX6SRo0PTYE0Ecg6iTuy7UR2Xy9pRFnxvkJffqhxd3EV0ri/zBdaiQvX5JHrW
7/3XZZT/adaGeOblarf58ySREkW/yg73s+VMKlIE+aQwD2Q21SzhXGYdJb7mkAX1sG5XDhHxvC25
xkOOcAdeNB3I/os8LvAYqUKV+4AI0/2lY2muLyKtrWxDmHU/WElM0hRNv4HB+GqdhVslfe2AYtw2
tQxfD4gPhG5+U5/Bg9fjN7u+hw5XaUX55rpz5YcGZAH2BeHZof7TcNKaHUfNbjDo7kQRsIMLin7H
yypuU50HL4O/rJCtnkJfqzcWnegK/JJhF4D9VSbJbbnPBiacJ0DEpWrh9EYmtw14lSVK3jZUJRAc
6mEAxlGyWGsTBhnzDx4+1NudWvRwzO7Lxb60UnpOkW56WwVAKpgsW7D0RGTh3QSS29rVChKg9GhY
Cjp5akyY8dMDjSEPmZ8Ul1dCcnnf7p6uIP69VaI94wDKLvgXrg96NcygvqcHj+JztIlTspCr3hq6
XUVhGZiFarLrGdThmJCF7Sp+grLtPXdQpZg3FMrX4/IwwXttuR9YwP/yKHFTuegh3RxvVSUy/9yn
tzuXC6GVxCKD76ubuTyLsZhJdGr1LMT6kJHVwGx5v4V8oRazwpkTh6t+ivRvQDSHPdFydQg+3rea
FuiFZfmrWfzJ2lLY3HoWGG3ZC0A6WSTLnMElGyOkeZaMJcnL6wgKSSeZQFgC9w7TO8w/h+Oi6ASG
xvQsgz+M14E4cf8rlVV+p8nciHcoKwJqGcnRH944QelHjmuNt7nYaUkt5c7fBCCPHqaCTsxEB4BG
4R6VSeFpYpe88/4Hy7L6NAd6wmMcR5ofoZ/w97jzFjvXjFqc8NE4oDz3HKF3/4dHkQY4D+2XJiLi
wLjhkEE8s471gSi89ClzM+S3plhcmcGAzgvzaU+dX907mWtsqOCSs9TNeVDw9E4b2zhu0m3uvQvF
sVB4A4eLNlx5VOuKQQ3SY/YEFsr/11qRn2CECv4f5yORo4sqKK3STuXfO2IuxSzEzTtyJn0d3P/m
BVYIym2pLMgaiLjm14muX02zx5CIwwhUup2r9xdKDBvWLglio8JbgIyAwVEbCDbyb7+d4YwQiITg
SzXafSkoV4hXHnNkopxscO+tR1pJ9Zz1qY6Gsc8yVK7k56XsLcrQw5dfEriKt+RdezgKHY5e0aKQ
ZBFDGN3EWy9GHvT4cStg+HHgrZ3CuPLzwoipfoD+of2eJ83Ag2S+guKD+V5dahXdpJB2Xk2jH/RY
EDdB6vuXM0WcR6pRey/nZf/pG5RMU41sODLiiFo0A9+YyW1Wmb057HfDNPYrty019Fk8dYhIxx5y
bR9/ERlgWZ3PQ6/4M3TWm/9esFL3fMRZGcEVPsdQhUbs9wLmaGRDnXuYu/lQuRkLBIImpEOxsTNq
aNXKkogk3vuaFWSIFOhHIdLN4agnn9l1vRH44ehTlwXB44OwvNgznIJTtSm3tqZDlNFM7y6nSy4R
FEMY53xnyUPranvAH7wDVrOQ4DTL1btPWxrSM1bHrsUQY0ziZJYxVH7k+I0CYycVTXnRAy8bMiK1
VQAhkNPdxWAmKKYfgS+Dv2e5doxXIleWbVZrEfCaa5fWKgb+HG2jZ3y/oXwkq9Uh+jrxiR4EgIyu
3qcvAkUI9bsPSv8cvToZ3giHjKla8fEigVMPyVbumw14rvgQnPTAlg9LbPJcaKRQ3nI9SQg0OdwI
TLvrG11ymcnpPjDzgTpIcPOBC06jC2svAx70/g+WzPFYj+MueJ8cgFlB0NnZ9FBv48NNXxlOxPUb
CO60A4SdMhN81VvQSLauJis3S45RZZYGkB9i3IwA0qsZyEGeRXcfJYAzHjvsTcfLT+Zhq/p8gcSx
lyLp6F0T7u4+oNI2f9fOrG2JDo1GKPKcXUE0BzORKgVE0LqSBuv/A5OgSaabLhIdDzKZ5E0Jb/76
fp4RBHNNRh8wuVWIDSNrVIdsdeKa/2VS88Q6eaH687rmYTyPTRkpxVkKs2VG4JfJ8p1I6fnem+iF
mGXmErsJeH1TmrBgHAXoyVFLKYyk+3yPbp8UHgGWFUwic4mN+slTvJcwDDKOuBzhUwPOJ4j3XnSd
5oRoQAA5emtbNTrRkcs87Avavr6Yp6DjJbnPw6EhvNhGHm+F3GXATmLfawlM1KWUq1SfnAaQ28gY
pMtUVBnAV9aEqrlvpwDmUS70WExchgfJoTTj7zHS7VwVbCPLfEBODJ7nM4RXVamBU7tqnLN6EocD
ONDU7ix8XsGZk5ec8q6hpcqmPWIo9PsTIMEUUSj7RoXdzo0uuGjjN2fq6UxFmjNWbe0ne5I/ut+f
UWgkKcKThpFk54O/FqlINvmIe2fibTy7yntCQI1nnfaEnUvoCovzUMHgKXdlJtvRZy+HvLG1wc4e
FACnNSVaUTeoTAhTGJOPVfD2vl0nRtlRtSMgogXaDMoOLBGzBeofy2Ok/GSiR8cXKLnPadpBx1x/
czP+vpxhh6eyXVhwbbiGd7BS+vp70g6FsBo/j4Fk5rBdcI0p5XPqnbPdyDvOGop8fX7py5ttqTFc
L2R5eZQL4WwysthbtswwOCtVNqdc3x/NXLgLmlbKo5rFe/tYa/At9yXfbf5ZYb3xC6G9BsHlnMVt
Lt3k5fV8Dl5EHFulNEk0W+iZBSwgthRMAl6y00mgKxEUOGTjxWGFKrlQO4XUlZMzZDnHQvLtPJlf
IjPkjwBN9AlkE5+wqo9+KSid+bhjtuItVGn3zziHU7QBZdiTWs8L3cVoV6iYhgdokL+5aYVP/Lm8
rMMSecD7dJIN3v3+ozFhUbadxFQ7nE6/udKydPyDJq9wI59noMaNoqFjPsHk3sm21S0kcbWS4t4U
+tYbM2edDosQiLF+JneY90IO0jWSoRWzEq9CQATU2NPe7gbABWtI3npplTSYPwL+l2yJWY9qcjyK
vuzZdTO7L6N8BV7gr+na4kXMMIwpmP1NTcjNY3G6Y5F3vL2X5YESjaJpgUwbmtMcrrzze0Yid/kK
j/zeRw6lHE47yC38rUPUaXl1+Edq9OkyY/9uyZO7rFyOwIYvz9eoDAOO0urXT73HleLyWsT4dLMh
e5N6A3eTIu29lsoUxKJyiHGkFAaS5RjOPB95tnajK/OL61vMz/RrIxccnfR752/C6BViR/iY1OA+
XUCVRs2VXHYAs7qCYkg1g1QvNSOa5RF/Uo1fbtDuuzvPAQdB1YgeUeO93lCDEIq0QBNf1vFJWUac
a07KjurDjjUQEKLxRKqM4qFY32TMGTO2mKxIBD7SVlE9IBy4iSwxegT6Q2kypcVQqpYh4aDrmVPi
PPXpNpJ+wobZXeaaFKo5kcZY6u3AKuSXfqtfzFyABFigoHv7JkvMK/hMLzkiVzPCYxx2RvUZEfs7
u/UWFLikrfsGK9IAhiAOW4eHdZDmuxaIpnNi0zlNgY+Y+9Ew7B4fYhoSJgSMLwV+j8eRvKrFLpnB
T/KQf3TqpozQ016AMuKZYjJ5deJrmeOc/RHM8+21nAfxwOggQuzGckW+Z7/c2NdcoIO0D/fo1v56
UeU0CUuFYbJR/rTWPhxys1cxV2T7B1/eRs4ZY3Z8DZdwJzkYLQVCBwv7iODSicvh0aNhoPEbe4l8
vzRZwUq0VjOquKS9uDpJ7k604ygR128TmiPG78Ph/pYHTBNkVd4dRp5ZhExrTRRn7xg8aGOl9ARb
WbmBAOYtoIWvI+wAYaGWR8BQRbOmR4rIIh5vNB/t6EKu6gLNGeY30iv6SAi3t2Ez7+SSoGRAgVsl
4oXdCcvLxJs0Znt13ssbE1/Mv4n4fw1AS2YdGBO/IvmLnp54btIwD0cExKwcX11dkZ3FL4PcP2ZG
49hEu4l+EhMdg5AAzCLBSIzARP2BtV4ehk00giEAxo6pXvNBDgKok+6Ubz/mFZ0yY0DMhsC1R5hH
DdTAt99vFD7FiivGanUucpu4NksnYE9cmo/wgnTsIv0M93Q2kZVTQx5ZRmEijgxy4q57GBTkCdLC
tA/Min1mhooMlFSo46NxTTS8v+uA2n1TdbGbo3tCKrs6ajFi2kHZbZNDJM1bic8WABvtsM/OOLZo
m+GyBxsB581PF0lQs/gz805FmVuA9zFXOncAlNgO7UAqFEgJpgb+fOkWNMGxmFpjF4k4FsG8wabG
d6xcGSHK7flPRJGpQkph7rOBvl71Nik63/0P3/9/iWGc+SCrO8jisJyY1675Fmpzk5KfwBz+nQRU
i+3ccFs8o7iYlZpnBuBbX9IjI11t9jUEFTovwsh2zMM42+3ebWRWlr6LW4lv5gvTMS7k/cjl8p/E
RxZVmGWndviyFJqQVkugH6AvGnkOlC1yh04rEsdWitxtJJDlL/3FXCGFE+kCR0tuCoMdNdy9P87m
+TU/FAW4SnfxwW8JDZoQ8aVK3vPFbfRwvpXTE6upgUMgElRYp0eaY8mphoVLbimfPzxRUSu5ik9P
UgYn4Rp+v8D/3NUPF+DR4QoGacmaKU8KwhW1A6QUAa2K3QRShz0ZWoyLLyYoYSsnwmdnJmCqA4In
F1d8zBbF4K7AxdQvY+t44gRVQBZ0fdMjo5/0Y4VkQ1sMNh0XAATySKTcRn1BbZtFyJlCkABRuNj2
72OjB5SMUejluGfNK0e9Oj6XYAaO7e5LNC6eTfRGG5CYsw2jXpyEtSdOErVXFdwx1pnlWwWUiRXm
EzUU8pRydKWXyQrHSVcwv6drgyv8sAYThvZsP0IdeKF6+NSTA5Sxs2NGl15GUum3suS0mBx38hsV
qFrEiQ9DmDkDYjyJyHrvsZzesFmemGw89o3Xfyon0SD0JDM4y8hdMZaDF8pOX79B1kRFDstxl9er
6+1oFRGYi8/sBVL+4iA9h4uus1Q85P/iJ19p0CtckXmjK49C0aR7i3vMdswjK3QcYhI6+yc/I7Uv
OOssnFEjsTPUHmsMLmIrTkN1oUIE2EbXAJYU0Y9P4xiBLoqJi1DdhGFO+cfOGEeYI9pCWIFpPVsV
i1grY5LBG2q7LlFkhkvHZBL46vw0mLPhd0sTuv+60NF2FUyqYcYuNgI5hgN5sAszyIwVMdtyMOgj
ExHpEdJCXEkGSw3ywvSEylP/M6z+zbB9/652hE1DcumvATpgffOPEUBD6YCKYR2ahJSv8PwOBj13
AIuvHbxXsykWBXsol4CDM5zwseS5erNjLQUhfoRFwcLPc9QR4UksvgpjuSW1nO3lULYX9lD/nprn
9SizBDPWZK0AaYmgBoa1jM9BCYLd1p9XbLLTfJ9Q9AnmaAj34KvNWE+4YildHxIPMZBdFcWONMuq
B9riDPZ900qDBxjYSIHY0LsxHYo33eKT2bFwSF2UYqaLa1xpCkp+m3StRChhg5LCGZqA2OyiTCCT
MZpagUPVqo9RYtcCkaGpBvQjuP/7NtvWlJlTDiGGLUVGR0jdY1b6eIbUkh+FtTVQhQajcEfIedaJ
Pak7INVkdQnuaLf6vPnHSE7Yr85SkRTg/kE+55SplT9jMi7lbDSDg+CfcIu+Gm+8pXNQqe7HxDoj
quLqMyV+JiNqMuLODMAu+zjc3/7C21UBoGjxks+jlpqBZMUnXLSva9fmlj98eZYthvo4ggONvRbO
1k+OPmIlL7RLWYs6vci3RU7Z89e/Thy5wkbQ8Yw5yUBlqy6INXXoDhxlHqCm40KjDWsDZPuixzzJ
iUri7ySLLsCNj42IADlksLIAa1Yp0pNYErgArYJ+znU/3usP656k/GONeImvmPLGWWhhdImf3435
olK4M4+kZTaq1PalwXxz+A/TkXE0FOqoa9inVjIrbiOXLeHFYhydqWp1h3k24sf/UjsPiGNR8whc
UqhGOv15EHgiXQQYvvA2krK0vL/1SpDWG66ViaJ85yYTQqrhWcHwLNNFRk+I4ejvhPs0+uf2DA8G
h4j9I5HPdt5vvlyp1BuLIn+qw55leI4liFxYPPPiNukdtS0F5zFrYREQyAMs7BCnv34mG0Vr9nu8
ooFBPWqB4Jpf/4lowD2Eq8e9tq7cl0aN2rz+j5E7mLihGUNrNystlTGcUMR4arPwLmUkw3IEBwZ/
HuwPuYvrzrbU3vJSn/2uplPEazqUK6jZCWXK4rj+NC6OsEJDDowyq6zhwx1ZQ9L+tlZvrlDoc0XZ
Ne2qSK6tDTwMpIjQwCbULO7aOCW2315n6bhndJdvtnVrg3PjMEOIXN0Uj6Oyt+X87mTFGdQ5qOUC
JC11Z98Sd6N0m8LstcXo5KgWoPv7UmV/7enZwdEYlFflQ2HG5/PdcWPItDoftNNa4sNoPaxhm1Na
OQihBqQSB33yfqQjCXhikPJflDo3UFQkIwXia1hMSqouS4WrXoCt3EFnoP9QtlO8pPS+5k64buVD
gs/xkH/VaCtDhPEmX/GT2TRjBvnGjxygtdVfhUWYv0kFro3mvLXXq9d7p1iVgS9tdHVcC7ijJbNH
ckq8X81egsBRI/fSQRtf45pV6XvymLw6iM5L9D0pYt4h/9hY5uRTj/7ZqAXE4bU5uw96chot+D2s
oCLVN68hTkwv5FZnisAXsnYMaIsSp2hmUNuyIKnya4fM+5nt4104rnlQFp0X4yJnOsbfaI0MPm+h
V3nCnsHoFlo7+FQtPDR6dpek3ut/ZwIVQCkTKSrFusRO1BdzmSzOdvmSShV/5MbXBxolMJ3I+BSH
onXNRnpF4tE48GWCelkpvc4FJkwWE93SIh76tvZbBVM98lUHKjgzGKBTpwFePRA/krl8aGLhEsfl
dGcnJiAYdxR8r1rpjJskryssJGRWI7qhtokSpo/z/bJMmeImtWmy3hJwCAFTzNQPcdtKpFUF5duU
g/w3+ENbc8ilflH1oLAp9jUMVuK7CS+Q7Lk0wVkN1VB97JUWZIUkntRBCQSgSUSegu6rht/x1bCj
fOfCQ2LUFV+/24G2gdKEfwuWX9tSP5+I+HCgCCEt2/7nmz5NlyCN4YlPQ8yUQ5pTVzRmLc8Nu8y6
p2N4YpBZ2iPQb783ksKodbQujUjnuilfmYWIUQS+sUYD3qtWanGBDpVmy2xRM69eVkJf0BtJLesE
Xkukfp2F9QXCcKoJzpqfc+IE3TWq60VPM9Q/700vq0O1mX7TfsEddE0URL1W578hLRjp0HVXgDl3
SdZpmhUuKUAJsZLKiwLTVrFFDSJFxg7Mz6trWCcEqeYc7KoovsbXDVbNnEt63694Xw9vxpRuWmal
s/PXdjVPE53cTT9V7VTjD5iqdBtE3Oy79OVV1TsruRk+Ml4X6kRPfNncQO6brbi/Wa7UJ/fJYZXT
YJT92blDqQ81AgvN+DoPAe6T06opomo/RLnYICAnOf4TV3duTCSYc9LQHrHWmIF/qU9fs8uRSQdO
pv0Cy82Ad2RMXYyBDR6+pAX+g8rwq1d7Axln5yHBkHHsKwbPex1YTZKH9SlW0pmYMGkGuQAheroL
/6rJaQCigBAxqL76FzutKqco8sxnGkJey6tT8+kk6A+qIUssSBXMQm6WBoLcNOKEV+ZYo+GfhAjR
Vq0KRH35UeEcX4R/FHNHhigmvkjiUrOTQ8frMK6FBSmtxhmavYmghHJPd1N7r5RXDIantCzjMxpZ
pbGclvBnsQftOIjjIGz4GYE5YuFqEsK19kN8YZoaqFTxlcwYLkill8AKVCW1vbl0UN8bp+ZOCJZp
NE53GL39Srv0As/fVHnCz/NIox5/2RTygDlsDqu4mFTToVc6s5zjdBo5Yby8b/2O7b0HopFuXgbb
WsgntJgQ4uRiKp0w2+ZA9Ot+ArZQC9TU/qXQZxSyoMsNFkldtWq+rtBDeB+1G63UvbiODcAv3wiE
nm86RfW7pC65Un56uUAZizA2zjtl0uhF+Pq37/WlnCyfFPYgZi6PDPAaatmPkqCzbEjRqtvctYcH
ylnAKQPX4CRrWDIG2DTpJxYRbhi7rHu7zd2o+KY0AxH05pOyDQD5fkFPsY212YgE1NmHLIKRRScK
pe9C1a4cIAPy5D4xalXVvXTnzW1s0SZV+l4S2EXrWJ38MyVawEfrzQ4oIogX1r97xPJlrdYF1oqx
GOi5MEl4rZhLmLDHli4GWpV91YPF00MEwxv11U1aLPMLcglEyuCGKqf5V+M2N4T5aw7pi5bMENrq
D8tau2t5h0018FcwCzS2Lj9diUWYGH3kdxQM6TlWcEKwq70z/W/ZD2cPkJKcSodExZhydENrCo+C
+0dArHhbH12lWVxkdiNacgzB+RPklIhQkfnoxyj1o/SPbzgTFguoMlD6PHMLjuw2T1Z7P4eLxnfJ
pZciq2EvejYdGhK3tu6lOXcdp/PWppZJLOOja5aafcWaOh33M2gsr1VkpHkQeBut9GWB+ei5sDpb
jVlG0tUFIT2SMk6tiqf86FjVTIJ8zVFnB+wX8QpoBdvb5zvrMUNBJEUSkN5y/RTvwz9tnG9JWGMo
GzCx5wcUBjsZ5sRmxvVjJQvcXSOwDkJgyKXGVnq1qijV80VnSE/4qB6+2weiqtKRuTMFnH8HRUVV
UHGaQOFXyrgKU0/mVkNrilp9gnbxqjrOhQ0v6ox+21P91Pvw2tXpf9NfrFdUAF2LdmrKPgEq9LoT
GqnAbZNyMHJmEy+9VmbPDjOEyA1UtipbetQEMDZWoXXM4Ewm6Fjn0roT+wGfK9DZkc9l0YLhhpKw
B4/+qWDUhMLq1CUw86ckIe+bgQ9LTLT+RZe1I1wM/G/1AMmgxvaRPOKjxnBMdsz+7wWbYQVRTwgP
8qbeLyj0G0eBzSBJ7IOOhXzkTIk5oQoD8RGtFXfETP2XQz81aoAFkexJKcW9PJXWRa2f9hHk7gYc
TOzhS2NxsXZDHerXloaOgMiNNmxE7RjxFnKTmDNLWOqrzcOzaLQ2pc1oCNS1px6Xksz9hxJxsErW
W8nezTmdwj0gHxjsE4IU0nVr7O2Ik28Lqg2aWcHNUcjmGXbEMv7L8lve4dN8uetfdcEx97quqsSA
MVHUYD/TwDYrPAAlMDgx4ezb4IXByCw4NwJ7Hn54EMC6JNb53hd0tHG7LPbdNtYQh4+ZfYcw0try
b6iXGWti30XfD0eAyyBYfPvdkL9aEIVHaxKs4243Z15bRAO1j7ec5GayOhGYDD/iEQXkCXj806gx
7JqxCv1cOUquJWWwVFwJPHUeIvWFCyuLg75BXFjMcFIdq8DnLKusRp3PjW6HZ4fh0hhK7qtQBy1p
A0uLffHtfqstpqT0rTWUpPcNbODo1MaeTqNydlDtzXhAeKw4QD/RybJp1gVLqDFn5RHb06A/XO/b
zzWF3Lvs/DligeLMgxcO/bCWH1UfP1oLMrtt5rFlElQABQRHYB6hLx/eQCGLHKqkA5FWacuwYyGq
L3X1Nou/8sivDN7/TmITK5Io6GSkOF8aenoP5yhfZXIPtCjI18fVfqTWmK27cWFWKFyRCUMxkOdQ
zN5uFAC0g/uiCXgWgjhf/D2dtLgMi41t+xt+O4FoB/9auXr0tt/g96zwIeiSQdG249wG6JGEdIuU
Z0LImKVxbd1k8dPOKikC7fmDPQPB02Mo62kAbmWnZBrNsgpYgsN/Tz6LuTPepxU/6vIT/jRrp7Xl
MqA1JbgIk0Tkb4z8MXT5qzTFGg0IH/YvA+ErCAcpRKS0LJs9cYJrXqX2Hl/AB3USXCMFSfXRBEU0
B0dcJdCX4GKPZZStp2xCtqIkGOk2UJtSAVrct4CBiw1abGe2SqBbkzOMxufVl24coa0kMMmzimmK
6yAJ1Ajfw8rFaiTAg5U6loHSVsYv7nDsTItYQR8c+0/a9vX5+QD653oD0k6d1LgmE4YWo5WpryHs
edFb6/qhWJceHvv48VWWOTsDPT1bcxbPexm53/VoEJ7VSnUdRb1Ji7WxjKWWGzkEZykOcOGQUpLm
s3qBeRmBzO21HB1dvaj8BugZvsv/x5V3gmed2GfceAsVODiEN1cMXhT1Oib55qWSsUHHmxzoRqk5
tgff8dvWlSGXqRHDUnkkVxb/zKs6+LAG1wvLWz/YE5+WD/nUuCDkmv2CrhmvDwL/2t0JgCfYeFj4
cfUUaX/psqVdFJzwNDvm6wbfdEXyLNuEB+7jDr+KBc+wcjh0/fJvEiDFw/fO/nFQuAUrJEpaMN/K
BEl2MSj3H0pQPs2u4saGxzk2STh7M+rkxC+wVG79CUx3XPa1lv8FaoBtJNFXsABjpErtmmSk5p/m
DAoJRXPmFHKKsbyzkZmZZa2ezxAYyiXQkqTl4duTrosFKsUMK01SqCDk0w1eFAJvmLkcXVEAQ2zi
8BramxR8gnrnE6w5dv6tbgjMaw9A9cr2GVVd1LjyKBwQf+z1jPQnuog3Fs906ZLpU0+5JQ00w6T2
pLkaxIeleRAjcJQetS0B3WeYIDZSYIdLPC0VDOqTfhfUgI8toZtsomSuWbcYrjuZYBfqW50MGpUV
GWyy/VxGyPlr7+79Qe88QysIpgTTogE4rWhCa7HuKszt1gVfYUuguj584oDN8CbZxaexMY314X1q
HVE7MsLHxb85gQhGca95km0qSkMvsVpeD0qXA+H68A2RWNZZUuUcWxqC9Eh/rdCwqhFhz3NO6Q7M
PyoA8acVsP2kNHWrrGUMpi3pJHxXw4aAUjpSsalbVFSYG/lo7gVocZ4XPTj588umJWkWsdc9nEUu
3Enzr4Kr3LWw9hZQyxWyHn9nd5j0vHKMmqkjQodAzCAWjlKIsN2IFi5j+u4CWP+Hdlkl1usecxMm
f/qkKYwicqwIe3q+ORwvHW2Mh8nReyOCs5rfAw3VWG2tC8jzX27+K2whQbMEwHjU7mvWr+IybAq6
GWceVakZtHfkGe6GaELdHMfmUwPBk+sheaE6Jyi+JtetbNKziPN+fKqkTIPPN3d2nolVq7bgbDrK
wItJ/oeLRB4KMO7iqiQaTRqXPTOzUjlkXAIQcMQ0QpJvIkseKED5RGM+4ExDZ3rndhtz+D+Q52uD
++36JYoAdSLjFQrS4cyn2rMxOOxpVZ6pXZPtUKEKu9ynVPbtS2wlmwaJRc9BialJuYUf6C9NqwGc
G61pulhJGHErfH3KATd/YITaBbwB9I8Lzn6boAiZaUdPMe8xtsL0W05RbdQy2YqqmBqK7/vgy8hu
56X0/lYUmStQNu/E6ZQGs8LICW74L2QmMd1GgfkhlKYZEbE3KDZKsF5pIlcCy1rgCZ+eKpNe7X9m
mKYFXT+khEIwy7DhmrzEXJH59g81kmK2uZUzCrpfx8geU4OjygqVy69tHOFuG0jw0/a6wi5v+oY3
+dUs+u0JxATUxhHbU3hXJZCjcpJf3T4JXEWM/tTALHlC0j3PFpvDIBRmW4Z/rdJD2a8vlvGkOXtg
VIzG8DzM3Sd6yIIBuJkbPO8C6/dvMWOrWvoCWwgH81DSAHMbRyk5sg9NQABnaQl3ejxxtWTnjHbb
qB7t9a1vwlep3HvHBWEPUBgN2BJTAeCQWMzyWAIADkLO+irPFaEkWEGDE0qQi0RUA+KYP8SC4Cj7
yuqE5hkOj6uJVvXqLxVRgO+l6YfM4yegirjBc9rVuPGZRm98mtr6DspMqSnZTvG3IiVHyEjLSeuh
n05EINmDSPTEIdh0atz8VMTBGge4gOjhAMZLTZnZA+SnCdpF6ewmW3Q9RkTvQRz3PWo3P7QGIb4r
KWYW3Dm4t1YhcF/iC/Cb9pqHdEN5MAjGQjrG9Er/yNQ7fQm5h2Aksn/op903zbkQsCtQXv5KDENx
ZY0oeomgFskIick0pWBcELhHvxOi361sHhvCZBMgMzMRH6cKx7DnhZ1BB48ImvpP7i0ghO6X5Y+Q
yV5qR9elmHoRykjy9OcwzaZK+dqcOuNzSsg+0qy7hCmkbqfC9WxBpP3UKFXmGC6jhumxb6G+Uqmt
rz4mSg++aQsTGJau9bJd4YK5fktkIB0kbzwgJV1mbi67nKJGyS6qx0zrQDXuOu4UHx+iun5vK9/R
+C8msX8ioAwEGzcPDG6Gb12PHUqkYYkttmknV5TCBqwHHQhPFoAQzTAHZ0EKdNtenbFcpiIEhoaN
Nz8IObJsNxWm0LUZNUOMEEdco9AXmaYfKDa7mUWFikTjjkotCg3vnlWPfWhemA5zCaLnk3Gry94t
hVzVGQhAMRioaJOVxsvGB/zp24vOfTSrMfo/qzOS0JLu7VSmsE28ZdA8Vbq4XS72fuMNQuaCc8WW
8AH1d5ZvRLWWYz/Fo3fNMBW8U8Sfzu8yiRUdQkx53xLE8tGrHp3uwFtAp3/ztyL5c+Q7HMN19oga
ZCUpHMzDwY8eaKMm+ZYc3flF8Ixr7Zr0fp7JD5/praCllEsDTNugY4+JYKyp6M5enuTB5Rfk7qnj
DAgyTLIpaWfuJ/8mKwU5UMPbtyPS+vfIUM3rR/l8/Y2NJrOITB3ZRT9CCKYHnnSh1+UD0LTGzXmO
EvnsCYLEpgA6HEclBQcQXERxIo8g8cduOBuuGe0ouu/WHCbyckHdUpANS3BvsikP5gLR2YkQU4FD
lWTE4FWwaGD9CLEUQJ1F1k67+IIyfA//LDbH0IdGe1lECc3mbFOJd8HnOYwthkOQoAxqCsmeAJYK
dWGi6jelYJC+3at2EBLC8ctYpgZCJYS7HOHzFJYob/5bTsgdYRMyuc1VvVYtQef+aljZbkfa465h
gCd4Z+MrY23h4MsR8SjDbV993qdJqYuPCSc8AYy0KvpXGeImHBpfp0Ry6kJ6HBgDCpI+QzeRdmNr
9AeIGy/RqLndYuhxxThgilHFdtcdpMYn8S1PsVIasfb4BHcHxkrj0ymanOvPDJHWxISebPl4PDkn
9LTEMH7cZLXvwhfs+0rPsSIkQ4KRBSeBRYwlWyFpSD4tmFdO2jjL75N24Oyg3bZGCuVCxVEYfxiR
cwrIkuNHetMYmACjKWiapyhBoBsyiM8UaiQ0gR5PYQxuHA0dFdFSGoVcgwaD29e1MQBbjApOrs7r
4QaQ8dz6/gVbNtTQhrR6nE8UnCK1IaolbsyY7Z/Lm47XvWa5lLPP3k8rhqAr95K1r7wOPE2GEloU
gUqnOlkYiEq4P7E2hKemyBhGBsGzQIyGZ6jgoq8unLD74M+v0NFy6CyDRmrTKgiXJMJg0CLms1Y3
9SJw+6ksqFipUUiP4MP7h7+Kg22KZF/reSam+3U2j1TG3pzAXSHjkznL5Xa4kBhGDShpCXwQfaOu
Id/S6hh5y8JXTVE13er58Sq3TcyXrAWtVf5qTqomavS8ODTjbttSg6wkAfV4QX2T0n+TqxaBCaUK
N/w0iPzuh+Gci/I1baHoz7rft/y3dYpBh5J6BQ3CNGE/q9ajyaKmnVv9PdyiS/3aR4QAM9hG+ED8
TeKBWmmVfx+ky3IdPwk09uAGjI8uq3hDwjQ4FbU4FJcXF8Yycbr/5Sy7q2Q/fNDgjNp2eGVL6+7q
8O8RJBL4ZuzwadLObtVamU6yZAyCEeTKkuHUeHK/IfkMzQsBFYlsH/yFyeaNlIcOxa8PAjp+QLLu
QwIEUY4fDyvxDmqEIy6SCaU2cvJvpzTiWxnG2tM0pJdS8yJJjgG3ZKWt4VvcYQUSjD2SBpUbrt59
uCZ1P6dvuCgSr4IDNZrpO/uehroJLoLqxpYiWg7lwXMVw2sbjA5OZlLNfJFZ8ZHOT0/JbSOqjdCg
HLGZHLaM1L9nAmU0w9/AcNIi9zx47E+oG6Y7CrK+m6Ofq5SpJ3dtQd0/hcdfM4+izdb5EMQBoKUF
wGMVqU5yAlV4LM9FI7VcVVqmUUsIPDmKfmP8VdY+0OZ5mHqE8aP/ufmQXrNt+FEXLKQaerVcKdJ9
I2tP8e8/1+Hj+iF+51+VAxaK0NUOzK7xzzExQcvmB5fV8IGmCl+Vd9AKa2rAHNipPH8Zy9SzWn+g
7V1/him4k7UaRPMtGkZ42S09GpXuDFYTzbqsTYUnogqO5Ted9PZoSh0liGk9ILmejKYJgc2DEPPs
T0iFE3QPM9FR31ivEzvHX8latIsKVEi9o7qTgoxoju4YGGGYlJggvSqbPkqe/F8eE8V0a8AMN0Vm
gbnzviviqbwhXDCXtDRFgVNKcUulZI3qyoZ8aLMWnys14Rt1qFZEElH0MNTSGFk2bpDQN3vb5E6Y
U1vNgTkrPbwl3Ek+9E1C+ytU9ynSEa9Ra2+LIcM6ah/czR8kgg9rlH4PQhn0mqguPpP1InMXkjGa
NJo4QZob8AjcZ5BKlDOE00WxYT0+hC0O+Qj5wImAif6yflnzD+L4qXM5AOCogByJmx1Ddd4W1GIs
AIe9nng4wa+EKEBOB1dxb5bfVkYaQ+le4I8kFeT01NJYKfAOeSoq8fjrde+RyVBif5ylVCYXseiD
s5h9gjknlBYeZyvbeCUwhviRlgZ28L/4udVwfw6s8dOwB56Xd/ashRUC2/oC3iGTMzI9jIi1i9Zv
6je3dBRqa242ij+wykjg9nKKKySime6eBbaOnwOXF3QubCZfGQPI+Zjvk0mbVme3ystqS4JThlKC
h6FB3c5Uk0fe4TnRPZzGpj8codqMY7Jzh3xSDMN5neFcOnLxNiHIzx8zVEAwQ5VCI2iutbe5Oasj
IQB/a1n2dFWt5o9/dzGP2OMNXcnl62yZ7xxdmiLe3NuWXODOsfQAzKAYH6gwkpX/tOO4YmuV22SD
4v7hPlo2aJ48N5snJ9JH+Nc/lAN+7PrxUsYKxaCH/0utRSLqnZJJdrgk++eytIbb0TAj2PL0TxrL
BgbdQLTvywDlm7fK3Gz4UI7JJpTeWjhKA5Cw9vvtZ7JEr7qTTBeIYQjNdfcgBM77pwarlD8As18Q
BvcipK8Jsq8QESaWnvdn/6KZxEivFaMfyCyPpXlhlkfXm8wisoehMYIT6flJXiTFLkXmoyZcF5yn
cXoCAta+ij6OK5TLgsAhfbDWDZQn318Hnu0waZ+bbBCSclkv+rGKNfulFkmn24C8w++PrpcjWq58
p7NCP0offKuGgXl6r7MMi0Pbh0H6+DNr/xF3m20kc+3pCMf+jChy0CFgkkLr42k0JzMu2EkOZ9SC
2Dw4dDpJQF8wSFW8JVnvMy2SDPN6LTFg5lL5k/rzqzOupG5sE5DJgCS+zQspgS3cOUt85wxX5jcC
Epe/9oQ6C4T8fjCfnO/mSC8aWCI5OnztYzgzuoYDSNSY8G0WiknRX04DVqqxsAbXsBe31mS74Tdp
01+Dq5XziSm5CXcfEjM1inmUdSQk7kgwOrX+eLgcf8BsCHfgeHyzsdZO7pQyo9S6LfrxLbv/N+Kv
UYdGHEAZYISRfcvRhwYNoWI1hUIMLijlh5LCvV/ZyJijaHvOewuLKhL5Aqs50V6X5nIlewoXvWu2
MSL90xoRFAJSmVVMhDQlWDiWce/iPso+wMwCo9nxs/7URjNgf/IcIMV6g+mTWl5iPbboylp9/JeJ
leHAEUYu7EmbCjxMWk+Rjv1W/4dvCZbk6/14Se9owSF9OBjlJc6nC3NFlEKi4G9mS0SvfRbx9t08
x1URhk/Bbe5S7k9leA+0sYMhA1L53/LcDNpXXWl32p4+7/dAfqGIBYs4WV+643ldDNgJvqJEwNur
u/4wx7OvflBpgu+mXhgjECdWSfEvpGXb3vhoz5bmrJYb/AlQPDLaWLqOVtCBApUM1/NfBFWZyr+R
QFhK/dLhC65z5j4trfho/T0BIDIYXAxnGTiRMJR3/ASP1535FcF3L0LfSkByAir6g3WcdkFQ59mm
QJ1dRa/1AMvK8+SDo93mklA3mTL3jMIjJA3KYtf4VHN+mgq43oeauxgVylOEvcYo6nfoBgp2+h9S
fu6rtKQ5roQOrVxQmKLoN7E/OjL8+SZG64L3m2rGctRJihEXJbFHdLq0LsHnHcOb/SB1oRH0/cVM
7PDaoaF3ITBvoe+gJbzPqlsifPeAK/CxLW0h9PUDwoB1RuADFswzNT/DGFHPYuTJVIYD9N6tA0fZ
xKchda8lfcFcDSO05dcohIIRqNCFa6//FXkMLqPJS4bCqldqeHB7iXJiQRnEV4B9hdwxcDz9a+nH
ri1I2V9PqWzjObrF+72Gqn0QztKaAqO6fIUqTwOIqSBvkENyfRWIkeYkX9KbXSqDmKvpkQof+e7d
Tft2S9baohY8OEWDCC8davisReWseB3ULnvFub6+Fbf2hmdqq84NF6z5edZqaAS5nuMSLumtcn1c
U9UaD1JUDSpOZ3kLEpIrJocO7TmSCEfilsmWiP4doeTycC02RKMVQ1Twi+/ugN6RazUkvGEj7BIw
+MZD9pPA+4yfO+FOEyWcURMecJDmoWr4W0AIoZHgdrX62Oa0P+Nokk8AihAbmuU6qnBFR9g6dt/5
v8OwKUNZBFz6I3p1gmVcFDMfb9Q35eWje3PjFoUJbMx//6i2bZmdZZswLj6qMd6p7DKv/kdAh8vj
lnwnXpsMRzpJAAJVOwo2HxCYfKZJoqES0dySeC91aQdx1Jw8hPXEJti/ChgP9X1LHV6xG+1iWt0F
dTAnuY8ckURFulY5Soc0cbl/PRSaozx9CgHUGVxXFfVm406YbX4+SbO1fXPjKYfAcbnCleQyUAw0
TyDDzzzh+HMeP+Wyy7uR1egz3Reve0DcN3KInZufb+NAy6HZ4JrBgVLskyZlEEgEffAcl021msYE
fNjQHLIcEYOTi16/CQqaslhsJbOhihYiYOBQV4rRtKpbByTA8II5kG9HB8hkBYS/YU4REQTpvl8k
0rizj66AzoG3RhXD+i4OZpVoodwZWfbRZ8bMw6psRmRwd3eGHr4HawwF4LZ3+thXZ7kANE4lMwAx
JmjNOfAauesT6jWTD0cw4QNRPmalTcnANDn6AGP8oVyYjaSpByuOWpMbOzPTJzG0XGfhMBxIS+Ez
OzBfi+be+bfZwZID35dPOiSnEjDg3mj7f7o3B5Vlt/vgGOMTDmZWjCXxMYWOOdJQLCV074f9h1LB
NKDOrIkO6GrQEzMMsXfW432d97oZUsUPgePQIIc0PwmBHtoqWC78vWHcMQ9uAy63Ehy9OyuDK4sf
Hs39NB8TvHSKzJLqIxmwvB7w0LFU0sF6yMc9wdHBZGTzUl4HomRuhDz2hWSXeltBBRvRHXwpXSNq
c9ObiP02qqRP0jWnEydwmA0SvcAfsTzE8f9c7K8Fd67b5mqD3l+2VBTefa7MwAjCK8QVPCNmDiz2
8BQ7DUyPGqzobhKdvI507pMnZyXTFyAqJ3X6thuaguP589nE5v+AoMlog+eBUdBr5hvNEWw7kcaD
H8iuxVVaGJROSISHRcrhyFghe4jt0q/bUvpHrNx6f6GehPTQNibTlSesBM3gc1nW7RbRxxIUuJOl
qllgo3aYzto+JOuLkQ8uvlDpilDrrpFYSDrmJqh52k+lxSylX11m4PpnrKw7FbSYxADfIZ/SYsKh
+U1B/ueCuzrwnc9GXv7SGhalb81+Qzrp6rm0Gy8vMR4YczezCn2FwJwV5PksVMq3n9fP8TRWQQdl
IvHUQGPtxMhILrTkIcwM2fI4RflUksxm3GxP9+DBkn08AiRMlMmdQnlsyNxbVD/6/T4pEJacB6gj
nDgfltqek45J9iJV2RJI/yQB91Rc1vb94fudNvsOHhDRyFlTxMROz56H8u+rpSMBpk/aszoxKZFi
qh/fCGDSgYpVdefvuOyH0pG+HYjrZlnDcEQ3Vc4T2sexCm52ws8K9LDSjKJ+Bg97I9iBNfvcR32X
XC5MAhAm+49wKSdZPjtBI7pC8OvPZcEmJ/VXgBGImSqKiiidXopYFZ8GFMHINZUNhinyAyrEgVIj
FFoxmaYybF38bDX/5geg5qlRbl2VNr6eU3aShpQRjplKiFVcTha+3lWo22GA8J1Eg3byQ0qABIEt
+vTQ8++XNLTpHXCdqLpYeZUhNxX2tlTEZ1edoF/ePzJ+iZkdCw8aCVjotl0tFaqRAKVKfoFQMRr7
h3Ikbo0LSIb2gjhZBjZQHrTcGwmUj+Zixr6P6v54Y6azCVdbginb3w1skovEZBzJc8Zxyr3SjC2p
3CtqchaaWWB7A0CBbbkvLS7fHo+5B6g7HhJXbSLU2g6TqFxlwaTa6Z8rw8BPGK3VNgSTebRwno6p
Fh1LU6TF4y2TRLV06/zLPITz2O9yLGDN+dDypoc74px7NojeGYYERsK8wvRyFhZct6KOs8C8viul
JqdZd2txtbRcXxEnW0BkzwE0GvY6U+EHYUb3HWQClK6IAmCHDZC5jVkf7aMA9+z1ECMvH1nvzFt1
JX3PNZefZLT+LTkzlcPTG7OJRzO52pZ32TTKv92gpNM5kCBFXpRKmLAjJVG0XtUE07MPYHk3H2DI
TTtXxXf34nqn0PW6c33zLDtL+/tQWaHWtxDB7xCA4hoCtsvIhpXEmTvZorfLKPwSdnnwtyMEUxsZ
7LJT5GwXFdNuJmvCgkCmNIEi2aPwWx+nAJUgfeZ/DfcZvwC9WGsSMA3MC0qBnRP1H6pB/3asMnqe
t0LS3LxMI6C7xnuayWGBHP/dudNJeV9Jq0Qjp1KP8HvRHXpiTkegd8s44nNbp1Aiwo/xl7D9TjAS
S9f94x8DBaziDgBIus41O8HIrTq9Hu9U0spL6pZ/SZAP5qdOKh6x/TeyXZodAXQhMRAwMYCAQEsF
dnXizf2sL7eKLiH/CoDyUtQFQhotaUM/7+Ij7rzM3xtbty1lIkNSepX0cGv8XoiJGalMrly3tUyd
qzJjFFud8mK9N+KfNVDiAMKgVOBjtqMh0CRmM5M84MzitAQdh4OnM0thTulJv3yVYxJr149O+/Gu
tttLlwahoxSwdDeJd01kRM5FyO0p3Y56u2j7wV5HR7iweEG/D2lXSBYzwkfgsYNkIKCm4qEGuKHV
iWMZ38AqCZkGmrlHI6MU5fX20FYgDn5tGqaFdnxxmE6uOm/EJpvSLHVSpjo4Ixq9VkZ8oT/prx6J
ZHqs+QwQj7tr5cZt2PC2ukzaD2ku/AfUQUzHkZdIXXNlYGNKpMIoc/BsvEKMye5cl+J/Nt4EzGcB
11zrlErqvwyTK8dqOpkQ8TdtCeWS/XBAYPaMpfznEqUiehoxldBqhJCKkBPXWBLrv8MAjiCtEini
iVKrNPVfCcjtywXnvUPfRFgpMgWFmfEtajsBkgauVHeqCnkJQ4hWGelGSY7j1vE2kNWk8Vb20xBu
bOQdW4iC9flpnEoS20SG8uzEHe42ywylBgRjWmz6Ws4UwqcYaTfiQ0x3vdIchTRqR5/w++0YI0oY
oTOtso+uVAgFh9S21PMcHAjuCDXBHJjlpz0hrbZ52QaBHVqvF045r+hRA0Dnax7nPx2geoOYdxoL
BM1fv9P1UfKn1hreraOVz49uftj6BNW6F02zjVpVVMsR0vdFpO4IsVNtyL0Tg9cN91fhNg7eVp5/
RIT9CFPnOmdx1mHHZVcRBBwOQ0Nj20SDskKpsC1v7+N/S8IiY1oBUCBPlM2hrXGkbIuIWvDJ7HSN
XoEao5y3ijB3g4CfmT/U+2x70ekTs7YBxnln2BeSGhPQQy5lKKXXAPYuiCo7D7TIABuGJqLwinTO
0o7UwDuidLbCKvg5dFyBO8/2zcU2Sb0p67Wb5Fjd789PFZvIVFwwv45WyRDlcYCzS70wYNEd3OsN
R9beISw2CaoiU7pNeO+OqgpZEBjhb6Blxq5knyDQJoaPPw2HwL6xiaGej3TQD458sRT1x6yKbPTB
Dpz6GC0DQeKJR7sqV6sCoUHESJpKCEyv/IitIoIsU/i+wNveEJw2kh2uG+VCzZt0IIvsD/yUe5cX
7eysR5plfUuX6mZDVKJqPY+99W9gW5bKbc2rw9J3GJO8UTAx7IJMEcnmk/XfMNJn7ExWUAqPBBQ4
KSvG/NZpEiRPnPiBr3jdvZRUXoi6oPx92H1c6i9ztMPCqO1y7jb842STD1Q9ObBdSei7KHNEd9ey
cnSbbcJqbjyMQ/hxQJwSRkrk/C5K1M4xqvCVOtDySVCHQPtKnVdaY3coUKX1xKkQFEO5MSdG07dx
2/BauwNz4jLGLkAJyzzHRih8iIweuhfFagXR3sLd49qcvmNduKviQn/1YgTsfrPDE6ZXyQquzGDk
Dzm/9RtdSxR1IsqDXRcACFKgTfy7ZnUYUxS20kI1RWzB93ex540Mkf73UD6VtZ6iSOR4uB5yx1ka
leK70q6WGcqCVTmgf6kpP9HevbEw28pS9I+xrwYIL07YOHabc+uxeeeoxFdHF9IHXZEyq/DX0jWq
Ci72ekNwaeDm/8gylut0cStu/wK2idw+h+SjClU/HqNV2C48qj37GV3bL8hplrg/PI6y763aQfy/
agcNlt9S39Zas30YMtsLgMqLCH1IDWo1dkAdsykzOn7ls9q+4yBHkXT41f9wYqm8OoNxGRZmAyY1
Bdkt4e0cVMLaMDY/R5xZ6dFjPXy3PxXLXZia2lJAN8g66wwaMi0QnatqRh8l0HbE3Uz3GAozWU0o
g2YVbBR3yy+z90XiwBaKpzuXrgILIqLwMwVo3++Jroa0sdD6E5jZ/2uL0tikLS9CqgBSC/drYUzU
cqLCXl3ixd1scVBcU7v/Jcs/hXkDI7BRXS9RplzE7Tet65PdKWOaLWRsw5Y7kGtbv0OkOv7xUP7G
zHjV28z8AE1NjQ96NHpLuQlHk9lMMo8fsX8a4mpOSG2fLbieAAThOaQoosYJnAWxrU5TrFP6SF3m
fhe/zIVGfTlvTjVcZAfl7WKpfnZwGY89+I8wM+wSfUjS4kpxhyMG81RUbeW6wPgg2ETQnorN/oEn
lr8bUcj2y4XqHFgFciWO9wiOVltpTUQ4LgzTEhr/SlELn6v9bUU3cPI0kGB5bRjsx+ckschgML4j
51w2s4u67hX4C1o2QOe/JbYNiPGYsnJcwdlkCZMzj59GidPaYkx6a4N4J7NveEiBlZold1YJMqjC
bikwIizOnOEs0KuBYR2DqbgBrew3mBRHbroZSCA9EBL9wJOuJLAue5hzBm7qf9c9rYvvLrUlALSM
S6f1C/gxbtE2RC6fhJlFJMM5rDMTF7nCwwuVvSWHEC/SG/1y0WqlW7OKnc4BnfoMr80IKORU3GXc
BW4dKEO9c1U/pE7+nQoRPeT1g7/HUd6xXU3Xa7Hb9+RJvrMrim4N8kRZb/oQA0AScpWX9tHgHzV5
vFYDkSxB4fbU0wAWBqeudj/Sv+wU1mB8jkDhjLSSGfpkzCjJpRvIBrINjUqsfYmmc8jMZl6wpIHU
PY8IFzDXvMvfF2jDkzZaAx77781zc3yQ9kryyTWyoYheEKojcb9Fpdc2grp9+ZJYHscdQJ4gJFfA
UBX5SaWNG06BywKsNx84WAKk5I91qAqzhmXb0mpknT+ENE6UU5i1fzxAdKDuL9QNBdcAg1Vnmn0f
qy6E1eoHyo/vFQKrEJU9uIyW4eS2Uef1CKSn84hplWCp9LinaGn06BHa5cEhL/GtKu31X/DqI7Ez
WV9LxTMjU/fYyzEd/J8FCwPx+aXegp47Yv9faAKKPHsewwoJ8m7GT0FYSCDroVa02JYANJDGVJdO
Q325MwN8F0wctcz1/kIa1UZrRu70DPXwVCAgwAs9R2UOg/qBgd4Oqk+VcsHwNJXTGKUomSE9Mg/e
/CO/Lzx8X/GHif2H5TqDdHewWwhnNG+723IBOe4fq0gbfJHLwAIWc1vCJfRbQsAhnYmIWC61vG/K
eMStQVlY5fANmlEE7N285TvQ4u2c6B3yu2IUMCqKKJ+/i1LCWzZzPCBJML4a+guSOm1Q/jE1X3Y6
EfAPp0Zhz/XmITSA989XhbXOTp0KVV1ENIOiAakB9UiB9GxLyneUNiPtxfSt/yReGaZvB+hIcfrN
7219Of3Xvr+tkXqBos06W86KPN9zOanyAquCdCbN1wHDjaUIMVxhq1TeQ9XyQvNP8MafPlOwnNVv
f112HCgSjYprm+NnhNl5jWDU6z7WrekT6kTTQqpGV5arO47k2h4I3AlQscguhQjyi7pJPqh41ATt
4YpM+5U0ZRnpPpgipwH+cmIvvgDa86o/j3xiOUpLu8Yf1J26kUM1+Loh5FF/35DyR7e+KLhHDBUM
voq0ZvdN7IjntsueLbsQVhmL/p40+nUYYJsl8l2sTEpUTuu688L5cQzf0fZWdzcil3+Tz5Zt6+kD
JfZ1ZZASptnkUnPQO3s89DP90b0FnWFxIjjsjKh38FlRuTu/IOj77hccF8M7L7ji8ADIMx7hQR7T
CNG2mhn61F8A+NAO8G2jXFtwzo3EeaMneJ4+/LBgzXmxpT/YdmPuDUQTSzV1azUv3R5V+tfVz6Cg
NgFzG6C6wlQ4+Oo40vGCUUnC2mx1CdVuau92AeoA6BKbggG3pODkppcUL2vOg8CWlEM/URS8tF7D
y8l03Xpg9pijTlpF0itWEIpnhHDRsHeR8lW1EHLhK0wx/94NVYAxLdQjxYu5XZRARgvCB2eTy+eq
2Sz0rl7CwhOHS1a8ByczfOKbHaDS+k6lpOuwzVF9zhfvNRpeVF4FuUleYRROZT/sEPe3eBiSbP1b
XHNRZpk8c8iJ5l/nITqwk7kfPS+j29ASMs/3vWqvZwC6DUVfulroFCX5L/9pDpbdTcGpNer2SkL+
eDMDNcTcz6Avtc2zvzliAiZrA8UQdCOPY+8m79vCor6A6N5dKINMe/lVovKQh+qvVBskP/+FoVqE
9pwYrjZMLqRZOChm+upH3xiErP7g7NGw3kw4f0jUlwwXIRrzJrYmdBK/J8cOY+H1AR93r60YrQtC
q9e+FlWKiF2s5F5KtrUp8/CdXDIicZMR6DjtAYZsmjl61S/5qVyU3K4BAEXaY9RXC0TQEfM36KvV
1N1LbhzPmJGQQIVDsy2xaz+gt7+XJ/fzqBwaNwBpfZx4C5d8XhY+jSP8yjbQaFsLn5D4SZL5IjGs
ExdK2eo9quL/ymGwWhaRCSDc9wnVON/UyHM76ZTW4iYdznoEvVzzkgR/vwC1Mc7i1etumAxD9Y/r
wnNAnOcLmAz9kxEpi0QTWbGZsHHzb0T8AdJoLrcDMlNl/gS7fNpgaSYpnTAg3t2x5240VZFIkWkZ
V9rbrIVPr31xAJ12yfvDQZBYIND5uiwn118V+vmig8xM+KJiyqrLttM1vklT6s+Sixs8kcdp0jAu
OAHTCk9ifKh8kmwY4eMAL+viz01z9mTNssnkMbqHoLZwspR0gB9ykdT3HtPl3E6+iiNZhKnNHX3j
NSTiP6yRG3b5+RqZVHGwJcE34QpNSUi6HyIjSMmRCUJXspPpBxvPdQ2TjHS1/qz40elpbB5S+wmR
U9g+MY5ylIC5cQ2Ux1NkOZ+GBegWM6vTPSNneVpp6X65+N5Lv9czTrUpTTsZhcMy1plc6xPVmNqo
jxXwgfqy1cqQFagcxdSWDAxMgsvan32XH2zFRWhqEBHp0cgLWn70IcqH6geFsDqCCNL8RdAYRqSZ
hQc20jLWGRlrqeIsstX98fBpoj5PxaFdQkNwP7AeTLU5NAqMlGcJ/6czjNMyv3+8fpe68I/3Dscb
egrcohYsygwURAUqMmOhFJlBnxm6xoBmB+NMaf6qXppA26UI9ePUDUBjBPA6lMuD6c8EwzGIm31w
J1omOBUhjhM11F7UAyAaPDSsz50twvK3nwNW8NNbpIcF9a6z+maWWmQsRM9nQASdOvc92K8qn8Dd
siUyYIAXlGIMkcfZZtJ9CCt1tv7xepdCz9un09K5rf2so35bLkBfq9s9cFyXCsl9XtUkgmtntDzH
Klu/axAMQ+0J0xFTJwTwaNgU0EsEPVPHR3CdKIv9Mlg6rzwdM2gghIV0eSBVZwXEmNwY2mDF2QK8
Tzk1nvaS4ANLuerzsbPCDkiUBsZtuaitt9XOJ1a06XjppgWmIhuG7RV661yU4IJ4GK2M/Udc4HZd
eU5hSsSu/Cv28kUQrjBmuXR9vk+LvaBsAlLwlrwTkGx2abwZTDptxnT5ApE2kYo6k87QnqdkXneE
9gWovJMxch2Of2D7k0YuGyuPeM4j8+KSCys0O6f0HOhR9K/I0XONWsfP1aX+/3MjnvWHLVRn4TZN
FkZ5Ht498HCtzybzBnbr7iSjyYKjyqTt7xoyYqtGjpdM3vl8UAyl/Fw4osUcTH/H2lwg3V4a1k/Y
WjnsyIi3j6m9xYtOtnT8OXybbODsrFjKaY503TLQVm2ZtQkBoclJE/lgfFfzkgHpjjoHvIpC4U/u
O4yXOXD4slvnyDoW8l5X+aydG+xMRGEz57Ns//6elx0Rqk/AczxlZPwfT67RXtNOK9PxSpYBvbZX
yxioG1hyhik+OGVZGnqBRCPs3LwLR9Na0CQ05QJndLCuYK7LRr2ims17VwtWkDtnOLTeKypN7RSg
4kNdKfvJbpPFJKMDJBMhMWG8YBkJa3SFZIbAQSMxaX2qjCFtL57La4RuBDKz8c0GTDJX2MNAC8I3
27QU8gFxA5CqGj+kcfkA2rc1xQVFsTAnL04fsGs5CtSmD0+JJekQsU0ci8CKWEh7kGLGIx2YDm7I
i22Vdj1oKGWpBqzryXD7anfdobG8pQeerG5cQQJ2ZQWNvC5pVIbRzQTsPX00n0X02AY0qwBgZEQc
GzQqhJLk28hqpUtKp7E5YyVGb63pnvYtQbutTtzcdiwUIuFl503PZpE68/1xCCOWPy/pdQ5d2FzZ
/489BOo4OiRa7hkruVPEkuN/Yzwk0a9894ZHjwuhLsrvGXYPZPdpvrvjw4XEqfbXI/rvjQuVFzUS
q0KdMuJyDzWOeB6CWInM7njSpJnYvxrTUWpnZucQ0/Q/uQXe51H2Cz5PTXm5xPQbLTS5s5pRLBHk
ZW4i2+u8nzjFiIO4flW3BxmborM9nfDKWLIPD14katAzD6zhDq8f6QwhK1piVwln58TMpyyTjQIa
idVNWtYTd96b08OI29RAAwASBLI+QGzfcaaEt9I2FF6+vlFt8Dtj5RVxYRTHMIfKz7AxNcRizgln
ePh7xw/Edhjfc/0YSwN3IHUDCX4lsiCvgiFuCY1dwp4OvTAmmiiR4r0aqUtrIB/plZDcOQ9E+lPn
BHWiLeLqt/SqBJV9BUctL/8dUVmx7M/XMQ9+LMupop4UvKhjQ68apTD4Df3PPQpZjhUihLiCBrqs
QfT7V69zEPyJrC9vxZEM0RJGQte+YB8/Ti/sMSh3m5fhwU60laTwNBfPZTMGFbynevDnTz7rsyRN
PE3yibZptGL6RzVoG4YjgA8lwWQBESPuNiUz4SFhQlY0W7VooZb1PoKTGvVe+AVLjFVqACdci7R8
p1eFNjjRmbcNxx4uqLFqCTaLNxKV+eGZOzBzgCPMzo/BAk+GlP8v2PsCDALDM2dxMIifePZuu9ZM
2p3H8qXl1x7OkTGSrT1OfJ1mZ6ILjGPmYmJYOn5rmsDIxWxgxAYIc4DAiHkTJsnCIvfFj3OqmoO/
mohFWtR1sViCZA47byEET/UQ6NRgDCXHjAz6SAqSm4B8b03VEurouGKrEQcVIbQ5IOfCSx2vpQs4
bcxihyv/7rmT3xBfgMimop6ysoY6EMNCvc+vscAU9JiuGC2RrtykgCmAs1Bzf/Sc5+ZbiAx+VGze
0v58nc0BEUi2VptOrv7cGGscm3FBJcfUxexnc6+vUTodT10GhkdxaZDrbdD7uYmBZlqOKVnN+3fB
HMya5xsSstxGJAyV28mFd5d+MKqhWeg4seu/yANLceBZ01564Uq70ciMnm6h3gEu0d8/ogAnbZJn
Qn3xYqxhHE6nR8qjKq3ho/ttvnPimOcsWExaLy143cfMw6tOPPCVugbdjtAtIEP75Y+U+uplEQZN
gL9/QzT6YhCpIlZmwCd4cxek5a3R5B6qsavbKWN5XsxsgOQBtsYxEAbgoTFpPVP+qzuDT6WBL9XN
KzSK2BOfweRnZAjGFdsc5tKzNdWeFjeBoDUTi5QFPeLreVvzWpnhrgiJTLOOpOeALoLy6N10iBoq
logjfvY8Np/6rjwUgirt2Qh6Z5G4plqwNhnW1uzU9rn/gm3lynvhZgvhb8XU1TEvW8q5BfL5wXd6
CPQa4Is8tqXs/EoHb1eNO2N5yZFKir3sH3JdHdukf7ZLT2xr/fJeDVzhFs0v82K2IVFvxYkNiH3Z
YDflCceaCb3A2rbg6HjAMe/K7RdFxtGheKR4rn2P2wqnm2IetYfBXlDogYxhcAn/XVW7do6Amv10
cn9/x+C4+wPdRVMZz9GBqcADiOAKWaQcy/5sGCW+LdM4Y2Kll29LYD0Zuz6n/3TVbWPnJq3n+nQy
IFY+WGuSC+kh3FX1SwoM5b0RrxJ/VvRFawtxmuOVuZ4sM8nhY5cBPbc6XEIze5tROOrYRGskatkH
iVUT74+RWZ0qrvmRWFaCJkNfO9ywVlwbmADctJRINQzQZUsaUyoRYO9CCakIlysl0dFU17StzvLD
YNl93HTZ7PohkJ5RV7cbmzJi+/Y/vY42b0zPqZnV5sdhUCXxvr0ip4pizSyMgjblPja4eYmjLOcb
oH1zFvHuQWsqUfXDqnveg9AJyjO5ihKezXN10GHJdEpu5bbW9cSJ4tHZr8L1RXBjgqM6L8esp5ns
RAbvzjR5kZzqOyJKcUxDfDPM+Cy0dPKEO2pBc837tY6/qkO7ATv0Fbm4zMbJ3kgYtvnr1ATm+cS8
JUx8xnkiLjTHm02rKVFSKCa5qulzMj8DT7hW0+Rjn2Wqk9LC3L8oR6pJFizLW02hDP9UGabjitQ9
RLMq2qXi7jK0bcIU1rQ8A2Gh8A/mukdKenI08BTkF8NQWVLt0hlDXfgV7FpwJ5eUlAMJbBb2gga6
5MnPFTZmK6H786ulyTCy+KgTGbHsc6aczkzQS088+3yfWMGwMtJjYWC2WFoBQnp637QkT/3UCDFR
GRAunJqmtGJ5fOYpySN8/DPmRdfmBCgZNdFD0ylvuWsMz85o3Rk1u8s04F+IS+V5SKpOrXCLlJ1N
CsXMiuMeE767vCQqG96XVu1pRBRpdT1iwgfxZVdNgvV9NOw2lY2Z2JGKrBqr7J2jHgVdIEZY96FB
IiUfw52susIhuo8Jvoec0BS31WVKtIL/m0sA6Ll+baopyRmfdjofPtIbpfauys4kSxw3tWZddCAB
H3tD8yLT11EFXJFDEEQEkyIXURD9bQN3IaFx6lov8T1sO8xqRQ94EI3IUCb5ruyttJmL6Ue0ne3i
/hCvZtt2N6sOsGWN3VzqAYN26nMMm9xqP7Xo7PHqvx7IbDAfAsGGIE0ryY26714YYctnTh9yXZM6
TZ6ovivDn0aVoRNcAUXLIN+mnYRZJWaRrSRRAiLeQbZj3YlZOLFqzQrvz7ubE/1GIR+QctE4f3lo
IA1DB2AdOg8JKyzo64IrO96BDV9yfM5uR1+ja3RZo1cNhhRq9UtIlTWXvzvJzXBdzkWJ59xnFOBs
jHjolmfSjdFab3V5IB8q2qPXwQCF0uqlsvgR5aMW0CyiMh+ZK3HxzoJ/ImmNEreELynDeTOB1IfZ
fD2SE2xKLaF2D69SHk9FRJmmOvcdheHT/poFD9gz5nPiWGggjxRa2cPAWj7423R/7fVmgImluhQT
PkxLSKhpT2uX5b/tCCuOooayivDB06MDOhVKcZzum3pHcY023SXcL9omnDZTttrRcdgYoALpKr+x
gNM7MO36W+KnvWC0C5/3zyG2sxuInk5bI6FUbCKBZTugcXQJHwPfsXK6qRQ5eW+eYBab97dGQFPh
jJF/0hyax7fEew+T1igoCH+db+sfghQmcHNTED3zCsb4WtrN2XFwZkV5GPt/h4I6SzM5t4RyCi8C
LjteyF+qAqGAOtaTWaH130q+jTqViCKjlHXohwtxPUByfHoDHFGd4ILlhpeos7hWE2XYNrFDOQib
Il7/g/WfdtvjGnUxUrogd2l9FcXabxd45faMrOuhFgeHttfLt+CLtjNcI5CPf2IDwpJ2VNBc/7+c
2sa96MGmoEqxlpeDss93o82/jdhGARfXGxBczzA+NZvc6wG/SKbAv7qgVwzCqFnwUiEErrlP5bu1
xXl3WiVh1GdW8YREwX7NvlJIAX9I23IioYcKXdPCpKQuG9qwInHUQXNpA69rX7FD+Tk03495R1v/
pq+URB3F4cmQnL9FocEvN/uqrgpenhO7ab65ha2DYKjA0a8jEE2wGq5+9zcuxE4c5mb9jmzF7jTf
tmiwUlDfXsnMFHsJoV+WkWsSoFyqZ7vgpQU0NdcwQwkXuK+nskWnNPMRRYOrdOdFlrDCrmLRhFto
pb38OKB5ju6gr8PBmDhVtTXvFPjSoF/3xY0NFX6PcEJyHOcCR+j5PrSn0EqeyOOMtsMRNJj6lvhm
bgwteqk86xhBF/JbVVdyOINSBscC1hkKBlSkSudpEpfILYTr3NI8I/kV/Itn7K6nkQCtCrW7XkfF
Dc6mNldvnSXh6AkeRVR6PlfpTQ/VzJVLJ0NHzgzQdBftf9jmmlmbfR5ehHu8K1daKC6wfPL6yEod
TD+ac4LnBCldeGGKzi1Ynl5GzryDO37KHhjlbbt70B2bYz5/CMNiNfUH6m3kJXwJMkt6bky6YkfY
vcl4BB037RAC59HmROhca1vOukCfBAz0xkrK21zRQpKoRcPrz+p2IyR2mmnVAWl7QpDXtGEYd9E4
Ox8Gwt/+LuaQ0MI8GPFGTL8fBbH6Sv4SLh5K933wzWR5SsMOmXr/RRFaep9jhZPbtXNOagVirt8M
wu1FBNnACrH+OiK6mw3R73j8lh9jVb7CR8+eepIlvjcDCyRcDaHipbjiDgYa27rb78TotUW8WhIf
RcpVIZRj8OYeBvUhe4Nf0fIebDaDag3VFnKDXjjSHuuSMKLnWLhjkCDpc5boHk30miZoctO4GgFd
4t8rGUbfGYu5MFYSozqVfosGQ37Tf+d0wRpPUt+iLkpWLVCqcVV53mQwePjaxte9LgTv7TWqaEED
tLKZb5dG4jdUPHCujh4E7yMBDFTKVqKeRAwPsTA3xgtRUf06LVGARbwZg4gmlmkWI8YDcosy7e/x
L95rXai0/bFBcPG5bnp7an2mlSs6pab97EGryKWJGgMpLq83FQkZxnz9hX/tb41Bj9CMvvrErNXD
8zLQ1I6O6juopPixcLQ4fWKLEAjGFIMco1Qj9hniNr2RAf7H4AynDxI63OxabvhEiI2FgUCMLLjc
Hjsj0+3qX7yUxqSF72MLvRD/TIY61/5A09JddcTImKxLJRRjUWo6qYVnfO+H7VwRwYpJLSFgh0HI
/S1kFq/u5ISNInjiE4nnxpQF3kp9QhpNefS0AqEafXZw1h+0aki3DwRml0xlqrjYyE/1xS5qAk9q
cu6Gdj8ZFA7N8SuuuOof0kYSUBRgQ8+g3wf4y6AjWORPdUaQvneUG3Iz4Sj826Qqyvp/EsfMO61x
dUJfMjVI2Q2YZ0NrpQacc8UenhAIbAX0QIanfPr3CmaeAovdqonu4X4lCS2J2jEyipG92mHaqS3r
9rZ6HUgnAju/VGeqRQoiXgMSSn6YzDnFtPw+UE9B4qBXgVu9Dy3wWhECzu/zWL2Olcw9up62oFaB
RLcInr5NrQCEp7qFypwuLZ5D4OIxunXzfN4hpEc44kVFJB1BmwfKeSun7uoT7YsGiUbwpef6TTvf
xA8JDiFGDOQrrkpJIRYYY97VRrGWU+oaheon0A9TYTeIPbSeD7c0hlAVp+LWvW/U4L4Dv2m8+TsN
J4vxyqgziLeQn0tOCNzVSyYtbY7S5DHLA7BBCvBeWiY1wK75/8hR+R7tO3IeoFWNzSpe0mQCKXsB
TCk1F/U8oLUaR+friguaVzSCsc1ZziPvvM9+KD5xW5O8zJaQhIN03869hH/yZT/Cqlz6cjcjY/9O
K9zQIjGPbcwuIsHM98e9LIEM0AffTY3VoqpmUPCH3oYKTx4vkKjdbNWHt6+q3MpszH23JGLfdGMG
BDdTnYgDTu03b5ZyDjR36pypM+6GUh7IzN+LGl/YTvYER9lgKuIwLbg9iDvl6v+OMvhfxf1xNzRy
XjEPFDbKxI6m78FnbhAcSjWC6oKYMb/rpaJ8Od1aVQMj+1WnPT1e0vIZzlExJNVapTnnbNAMDDIq
/9RwmZ8NcCQwJaQnZFmNvBX/GkMjiw3uWs9pP1/mEOsrOxS07Hlv1oKKq3kuU+JdSmk7WwRbnfrC
7d/IlGJhciKJQDJrLtbRc6PHteXXl7mGSoox5gN0nKp9mJ22y7oeH30TVzOu/I3kanXAx1hqp+IY
wi4PPHEypcDhTltldNxPZ3SJztLIBeO8JCG+vZjGyj4QVuoOVMRzcQwnKqrXTvutsW1yQewPyquR
WD6vIy76NlPJiDDIwga+1SR/DWIy70hTQwBJxvkL4OajH8fD5EQOuaeYfWfURYvhq5r6sx/L0ERS
0FYxtJcVvta4ssoUJnrktPA/PTiUdMZZuSpgESNR/HHFDSvzymyosIxbbg2MvcOGZ+mChS/wDUX5
8Lf31UI5Xqowcse/bMzXHmhGQVj4B9PrzF6cfjM/NWbB2jcw7oTNiJHOt6yJn5PXB0t2BXGI7dSP
garbGc6zr895nTNt3LCPmqRpqkZFZisM9kpzHY2rfIu+1aM+kAqP6PKzUpWN3z6G0F8ze/jNoRG5
JFh3Qco1z6QA/37JQ9mIleJqT5s8RKaggu1ALoKpQennsZulZyQ/trWs4hwrZ9SEXuDXev4PMmnr
i3EgtzGSoMdyiAZW0s4C63G0uvXiOcTB+pa14wkbcIxUVTAzukKLNVAQSyItx2G+1iv+wduk5oG5
ME02yklWdTWXRMp/IMSPSCeGVbKi6f9z8SsQW02Q/hFydD2VSZaZuS/hX/4zIez2rVQenROf8RV5
A/9kW206gyaJXSoIPiVAxx4uuXoGv1tkJ1YPnaOUo0fpcLQkxPbnzuN3JS/RP8qoBbAMwhzgwtWm
hgXcyYVfHzKp8XlSnpdL6Lag8kdtj01JqIxhizsbIuwbYsn8i522/JG18ytOB3hvcqItk+PKGUrk
NcDrfKnx10KJeernNSBYjEpYkvbTEkoMiKuPtNGFq2bqqwJrvTOSPOHYW30YGHfB4IWJMO45vnUI
ZYRz68MmsLbNQhA3ghwj9qKGPYEq5D98etN8iwcYq4b4m75MEqZkCIDBaTqYz5DNOIUjgOxFLriE
vQYO12wmzdU5NuaddiFyCIZEXKtBYwrFr7UDtRh0M+SB2hvlB8EeD4HI0LSjrJRA8RGI5BAcC/qG
+71VSHjHixMCXL/SDayknr+ykkyyIHQUGkm1pzjvsDxpsR2LSImPVDCuK/O9tFGkBZaktM0sJFR1
ZLsV9x+H3kXRcYGZxBSRyUFaCPlraYI/kx8duZeOhJ6BKCBt8GjMNIH1asG876yIheeXWt+5tbhK
8bawM9hGSwJ48cdCFd6mNlg8AM+HyukMFVGGcM67IywbgigXasNHnMXbeUtWfFWS2dGfVfkd+/3q
2lNRBn/DkxQuLqSFh64zDUIkXK13/hcq9ToDdmTcR+Ji1c9OreAjIZgeuvLUiqPbDC18I0XLQdzc
m/d7KrUG/qc6RcmjPT7ASS7AETrRaT8curiPOi7AlBZuX7IChSvaXogJyKa2QWV8i3rvP3UQy8Tc
mbuQwFmQKmhlWYNlV3Gjq4VVH4qZjfpIcKAupHIRCwTtELqFnSeRajMzHIT4tgdDsDn3lAM/d47n
EhctTUbBpZ9QYjyVWbeg4O7e5qUi0URMSwEOW3G5OSsPRjakpl14jvRqbqqfvnbBwFaVg6tPtutB
oKkqnMIO+4LKQ2VnaxrvzUjxztm+CIuC3hhn8iPPbd2vqXZOy405x1AYPSqNZWokceItEl7mbXXg
ryAuayzxq2EAlFelDZZNnHYKu9lTeSgO2jmbQ2uVIrkHJEAjKJgxHOby6Ibc32MG9WHJu2yKSbPz
zcx+bOz7bomWVr/s46G4BLj0BpTc4Eu+ErQ1ST6JHvX8GgqeNcpcxdl1eN4r20ghrXfUkzX+4I3P
M2Jcu09OZKWqkGyZQPWGujKSfT1p2YstKSSVm0mQnkA64+MLnX55M1ojjgAZ3D1PY3hK9b8F6oJm
uD5rxyNMXQwWQ8ehv3+WOu7YHoiSkTY0hI9BBqR/WPBxn0eN9cNZJtjbqsUVippxXztozQAmYE03
g0DuJjRRSNAm85JhJkKhzwsR4XTwEWMAgr9jHYwkgWXMbWHmLUadvlYIO4mEOdNxAdUwP5YF95Rz
B7KvmdZGDCQu6sZtqWDgodmxQsQY7LOmlnLuj0NXavSQ2aP5uBMlmFJKQw6nc+AjFcf6r/3UeLcT
h30HM88G3C0emsX/oXtysO1Fy7bEl24l6RrDiZyqR+roIXmsMK/p7Qh3p62FthC0O2SUEGxP8YB2
5Y9Ecu3MQZ5Xz3glva4pO1YuQflNiZCd0A523yeN3tf1XXOKHNKnqGJ/m+chCoMeTkestZrrt+pi
FS/nbr80njq2902dMPI/hl+WQzhaA/GU4O1jtp4VNqH22QdOh3iG+T3g9PTwI/DJ4uZSVZyxpIy7
DVJXA+i0JSMn1Z4dum4FQyoWXOu4v6oV91wsIMOSFyORfm3/jRTU/CyhVMFjo7xsP95WC/JLB45g
JG/KF/8ZNXYyxoDHXcyZ0zys29UAGPpvs7+R0xPE0qXZikxVPz3O6TsDQMVuBfcW7cr97PPZkOwt
idJdpE/xxII84DyRz8e4t4zaWhrlfbI4z9FTVc11DexNkAtXpsb2iQ/uWN2sw3VHNNoI6Q8DPrxP
j8jyRMwlXYObZSdJmM0wP/uOraNk1wpxZ4AQL+E4SFgWlDNIyV0aH2O7whtVcMDz2ElfiyExzQtL
veUdE9fQH2wA9WPheh9JBH0+FI1GpABwK99kRrKZAzw+QcRpplDfIkZocgJd9rzKxG6zdn4tSHMn
r2vzrDQ7vKPBUg7CJIEjeorQnkgNlgNJv5mq6ih5G2I2yrIpLw8n/785tIpdW0A3XchxyA+sxbnX
kJ2uysvLP6mImkGPehY3NEHGzsWKKtKTJ0TQ5D5erIKwDdqZBp964qxZzqhD5hnkvLlZ2Q4VmahM
Yzvd0vhdTW5FZ9YQKpe8h7GG/HJR4gC95Iv/v/qmeDBCqnlQ9mUGuMuIGFEV0pD9wzAwexftyA7c
SDuvARCXgyyNk+QNmszeWAccL2BB7hNsXDOPv7Y0RMXITJCvmPTvnOYj+BLBAUBxG77FEqXGuAaM
rEyj8DT5ATGLlkO+ctalzweQPBY3HEU73eAP9zcj4A9iSZVm0ChOwnhhLattTkNF/zTrY8PuO3Pe
yf1koykz/DU+NWQAzVwefwI02Y/H7IhhFhrbhYRjrXTpXPk5i5YziNMFvthHcMq/eWApkf68h86a
hzLFt13T1+RM4+c0aYLVkw/jOO+qanUTjzu4n96glIIwh83kmOeQiSx/ppZR29SHA3IWQLOXMm1n
tS3Zpca8jgf+XBzrYQW4Zul4yGjtWiWaS3tBjBJeJ4KmDNAvqbBr7Gp2SDokfbhL4QfszJgukOWk
v2vEU36gnC/HKL6aLNa2Kta0Cwy5cYHqKj/IrZkXZn7aq5GS9hS7I95qUD26WV4kLyM6W4Bh5o3N
j4F/CEqjmGABOchDIB6hCV0UhhixY8fyuDGr+956sS25cCmhtP3BURR0XaarFbTCIZ7RsbpTGcUt
AgVpqRquvmdoeRy72NtDA3cqsc4OJRj/8QXjjFHpoEtylj+q00P0xsL/iBkXkqNbiZRW5tPMCTOQ
ySIT+mxlSiAejM+KfQrfy6SLwLxXBBAYurTQPZ+xMHU1DIEIf3KtoBoQZs7N2E2ANa+FzGJ93rFW
nKgBWSOAPDkE+wtz7iJoBdLhVktkZYeMPUQDXlagYFlLJPltxgiDbJ+F+UyYYV+OSIeqzRxsTl/5
7lQYe1ZJAET4mtfwywiqHTrfjX/RJO0FHnxKFemVlC6cu7lwV96hQo51tHaLuTwJEe1rJhWG6qDV
OtepoB0UZRvN27qB/jTBaKx8qnnAysKpzLx5O+GrKQ5wmhUPkYe3twM1Hs6HILva50jckt0LiPz5
WlLqa8PhPH/cC5237nIJYT/QjRhEjxlfjemxc0yycJf8Wtvf9FIysbz0Pv6p8OMw775+HWcDFthn
J8GNW6XtD+KrYVM4WpfJB2YBD3xRyLqJyRZZRtTLiZG8jFBrYmWePDPI4IyawsW3bHq/4gEjeJvU
+u8En56m+tfgT41f6JcW/QJcycTCtS9hs5fef9uimGvABve055qaKUfME3BegZjrU1UMOBfM3F5k
963UvqqDEF4yuJf6RLIE1p9+dUewXfWhv5E7wijGKMKSunx6C2Gat6MCXVp+aWqBLfTRCgAjIdYa
fKFZ8VF1TtqN4pNNRF6g5DYTdJllI6eO6aJqiYrdfw2gO9PwggkVppD2Co5zcljYJyeB42P5Bvfo
0brGGbi2oQYQUFjd3q2/Z8hgghIkpqNiY1wra1WuKb9O3y9HCd4iStv4pHuRZInY+cppcZi+dVCa
1fkDC/XvLwEF8giq424+qTqQIaZGNs4W9k8C0rYuI/goe3XBMcfrKcFCYAvtQZ4csBGz4/XfogZP
yUWipryQbLiUzDZdTNK+KhGVmwvbXwy2nZZwT8z6eiJ8a6MFR2u1tUeiF809LGWe0IlOYIu1r1gg
gQ2A33zeCLixE//f5T4YXIihEK6qPYdAu3dGL9nQkd1IFuZZ8qNsDKseCbI1IQra75TPa7KV4KQS
sk/kkM+XUQRr1vyh1usYnbNh115aFHDX8+mh+NX4amGp39m+bxQ05wSHD4VjYAdho5GbSDJlgXjS
g1bCfTv3fnHT3/VQuWlR5cGMTALXQjsgXYKN/Q+8lvd11B0T+tFzfrt15ZfuxWCcpEkUXnuMQDhy
ljqMaLPYJT6qUVr2R6zD+PE8R24TfZRTAX9B64k+dixkLUjZ1C9eJYioobrpyAcXzRmoUap46db9
2xnIbveyP0xy6nv92i9crUQ6IrQRBaX2vBFLKitRw6uRcQMW6PjU0CvSdF9k6hrZiN6iWrYsdX2b
ykIgVYuP3dfE93QeolDHL2qGBf7XZ2PiidfIqXg7x/rrr6vi4u2xMniHEpHXxRW5DSeWG38WRvxL
mWVMO+6NpW9YIUstbFwjtmQLsBrjmGhmxeBA2NC+TucOPdcutiA8FXr/qrxnbY17AXeF2hglPe0v
4/Sh1FYMIVZOkMokrf13Vd1X8FXlC9v2vFQ++xl+sf6z3kflTReEAR3N8YYuov9UmSS88DHIkP82
IgBGQn1zpZwUOTFfmKrK93lvTQkYXVymMWBMWJLsYFYDaGP2Ef3WeEdlq/lqVnUGcH3ZcHnbGWgm
/Ik67Eldem042zTwCT4FBHEMyp+j7onTT8rG36qI6CwrlLw7GrSiq7cR+GW9pFfQOa5Go4jP//6f
Gm7wR+DBI3bnhWynyrOJZrlexK2zNXcm6ESttiq7BMjpL8fCn7wdc4d7ouwlVS0dK7S73ik0WFBB
lUnk6pB0TmnqY8KlUkAN9/LpDq3TzYp3ZQ/3uzOrPEu5yWK3nAipgQWocCACaRbjVG/5LfZbqVTQ
A47K88ZtAguMZqmIu+BrrqjoMh7gM3LWtlemfwmwcD8NU/hel5AVWvyODAfcv3GSi95hHxsEBQsm
+XRp5Ofw7sanmPcAlI7UTGSCZDOSXJj1wr3N+HuNjUpyZbtrBHux3K6whr19iykAetCgDCTtROiJ
d1+uTntkdhrOZpbMJ/gviiWdzAKWqbwdG5YwrfP2dIR0vQDdVm1T8bW0F4rlJU9koDdFlvmkx+lA
amWSdIkwR30STHW6jdL1V8ru+mkFJ6P2GRAOmLcpiPSGorecTos15MyV+Ea08c5PMTjpZXJDm7g7
yPcVlj8rqLwvC90fvLKCpscW7qSazDsRcL10m1vjVy4M6P7JUB+EMEAs2tUh968UpBixpNfBUUkA
rqniTQZi6dsbywYUn7lw4jQgYiTsapdHfnT5VS2d1+AOkDa/w4aGMJ0QgAjfIaq2YPky3aetcZPf
mJER4DaTtDoFyimG4wjK9SJIidaTIM4BUDdvSrLNG5xKLGD9WnnAjzMAW8edkBzuJ/YvPeaZbBuy
9NJ6c2B1KeHi3gp6yjjJKzWRH3J3w0ykCffnmczTMIBB4d2lCD/KN2QIxy5mIsTgOVJlwcNMwZj+
l0ZNxOkMH2yQiT51sb+wAfXwD4yJzL6fZEA7YOXzm+5wrvzzsg4mikxfjbzP5ZdCRQVPu6pSYHi9
f0sEqWGPgTPgNG/XEoNf28BwAc78D9GX0n/UmRPH6h+Cfn0YkR+WN8KF2jq1H32KL2oupDTcTZiG
l2ip1oVOcfQG4SAebA+Ix4rJNZMZcXvmPb7LJ0pxZDv+vZ+gTUy3xfaqCgPqqIs+cQX7NXDmw7jk
8ynoQP7QWo+za7PXKlxsyN1MvOExYMNc0UV6s1448Cx6+IXfV1V4pOm1KIjgS1D1c3WygwgLGpgj
SWGngSinySGnEQH9KoNPk8/5kfIw0I04UAD6frYFm0GQc8l5oSdEWuhW27uyp+8WyUGivQhGTWBk
Itb0ZH/rBS51I34SRJW0B7VKMz/gtGLHthn4EAvgNmSDS9OQf/oXxpaKFHhwPHBKtqAdIchCOd2L
OzLhNqLFIfCEs2E0RfCqi77tZek4dHQ4PKktc+3LlIju48COLGWFFflCNduIOvOo1+eknLvdRhMY
lxqNM2cqfZ2V3qu15okEdGlB4wbRJuZrmyiYDgA6Qbzc4+u94dqjbtpZ7WPkP/HFPtnqe9hG9Ysl
CtiK3ghZDdIxQC9Fc/DIMYlL6ErHBV4gTthBz8vLSJw5c897inh6ZWMs+PDO6+BEiobZM+74ZfAm
a0IGtyY+qmDVuisHOPF7S10VBtyr7dZihEWO4N35bUjWDLVVtUBYx/G8kzTre3wym2XrS+1QRsvk
Lkee1Hr2Gjk+w7oBpHPDGhSMHXeAau1OBvPD7/HQsnMvBRDL9FbnEk2IZrM4w2MUkm0sNDiN2Tkb
Ca7jtPqIdXtdaJPZpOiSFtNK5stQlXiiGkl69ZIx8wlUIq8zxifiLisuM3YUILHx86vfJWYjg8ca
2TffIRGRjKZqGLiXwey6995im9wFtgFXt3jmE+ogKuAZlywHWTcTXPJLlnkIp6pYLgMc8DBa58sk
VXAKuYsarrJLCC7AjIivzlox/U47T0y0fOmi6zfXpG9qisn82u0tIYusbXppPBVFG+p+w7B/dzUg
9EGiCCruXF2ELtVNp1mXS0NVHN7/N0Qvuy7oLbyLeyg2xZLKeNqN+crZ4563ODMVh8IQvgGidziW
YWyYr3/YQyYfUdz13uujMIYe6Y8m/tyPoW3Wr3RURuHW7wf34w0CB2x7ilC8IgSerdbX5wAhoFPG
PymrU2x5unSWn5R4eqWC36wvS6Zr+GAmWVY2CSDjebMKKMAoixgN61z18qNFHOf5vVe10FkdpagZ
/T1n95tX3kAzH3c8YOj+xt925uUKQRCWwCMqdq6q+ca2KV0z7ufWh1IHNQSi6BaBpQyU9KnQmq/D
bMg+sDSVxCwKN3auPYCUUssBbZK93GppwMV+MDpdEcpfZaH1sKMCfWOjG7T1Wk3PTSd6LXSOitrV
03WEOgXYF4aZ4E+jmcIVDhcLL7wFwk2BEv6sLaQJtEUDf8AtwHdb2dxVqCfc9zr2MMOOUbgxw6mF
w+r8iJ0AqxBYZXogQjYG08wrsngD5Gy/FEGXUrswp1ayQuvSt/oKVWJXqVVPrpttEq8bVyfdmIB7
cMbWrNuXpJ+eGq+AUxGtS6iosydgPZMA3P6T+jAZ2YYGntKt1xrIbZ4Mu91Ns9gM/PhcdEGnATZL
9TYIcxBYhfDsQpFUgkQkOFTmFFnAzlC8sI+vrK8rnkinyshTBqYTJB1rs8YUqLPDXOdZd3infs8V
qGXJKBXkXrNdYTt2R67Csh198n/oLMa1S68i1F9QlXscW53KR3sco2RQ/SY4DT265LYgVx8RIpvK
m9HWwel1s2G+3FEFVFE2Epj1oVMnsWTLfm6C3zr8a3DTy7LMplrTpVb64Wyr05eIPELp5ZUpTsAY
P0SZVG/+lbUVavu8PBMcPtFIs2UPoxSBRBOKnpsS3Lpo6/NUXa4QikkTd6d/5RSTATcUvX55oVTP
QGgbR04rgG2p6ICiAuuhqXTNOO/KKvE3Tu2qAxg3RHYIZ6utqlCP27ptjDb4N2P+oQGXXHAgTrLU
fkpV6oIMeKnd90x637Q9ItiSg05080opQxJhVL/RKedpiuunTzwxXv7bzPTjaIRSnNXaADcAwI04
G62d/4Ul3Ul7fo+NKt+nF/XqbjE+FzUhO5+Z+Gclt1IwBqgaPa5lAvMZabAqRX6MmPslCPCw/ZtJ
jdAy+RdeMztc1d4u+Q7K0RoWbOjMd8YXXtl7N8NKHFAHisrhpVV01+nXDPwTwrNedXq/go82xGvj
LUjj6Y80j25zaiZ7Uzzffw238QPJPRkMvpfrYl3NV9na1g3fmfmkp88JB9ErOObd/CticzZxoW3D
Jo1weLwYB7rNHta4Ij6GGo9xKOxAs+tVt+pH8NCqc4eMdFfwzBpJ0CqF3DVV4EJhmA8jA2JlhKsz
POcyl6JdtI9m9qywO5sbnS/sSyQddus4NRb638rimsgAWFjhogGNiQtMsDpffQyxSSNpo4aPQgX0
bPLS/KY/AX6VwWLSee3xb5Qo9qHY28fZkVGn+1hKE/M409bpRtuVCX/qgyPWzZHwMJCZo4AXoy36
J4lSKdVboZcziadWllyVJCcqJY5t0o+83lqPgT92Ktzcs+RNLJV82oq/sWIoTJiuKuwUlDg4/Mt8
zVdWayb8N/yZlDPmIMyh4RfgFp3yq5brB22WGBP+ryLM60X87n6h69Na6Omyh7CLt25LFmDWfOB5
D+gXoct5bVZPcg0aY59O+x0amaE35hBl4QHAsykCl6fF9qlpI79tb8nHIhdLJaAuChvvATcJ0Zmz
McS0iKYvAStto571LEsmNNfdtjIoPywqktiQoidtU/0HUPU0ne+Au5X7vuTjxkvEyabfobpn82j9
xA8nGG6xxQtx8CrIux7eMMalws+KvszWpKui3LBLAlcWno18NllruOyYmblS8yhcFjVw2CKYupC8
QGSlgveI+uf3BgY0RA8/093VB3ZtByajYfFMJgaaZvv4VT/xUA72dXahxU4yN/l/ZtmTcul2MHDw
/aQctAbotn5MKdExYd75atrjtsXnij4OiIsOabdIPRI4PeL72YsXuiLogRRGylfYHH0MfiheaGDn
CisxNam37IWv3hSX9fKRlGragn9CLMLkqj5FeXYtxz4DCWBUaW9HqxyzupqHM3FJ1AKbGe2q15Uk
1Cf8RFoRCdxsA7JZ+elRJzGvuBuS+DI/JCNM/m/CPNd7p8dBv5P7oGnRfO6eHT99Mhg7tkKtlsKO
N11ydfNP4isVnghmmgH9a2olAPj33PSUwbarHVjKP4fzNtWrqy5tZ8YDhU4nuN2nM1zv3XzsP6CJ
jHIh7hY76uNSaCTsvy7rE6HnZ2jP3nkx0DaDIKzp3K44a3X7gi2VaEFPBrn7OhN5SHpFD8G+c+UF
mkc2srl2lcVNcW41MG4uCs6wO3xT0qhWDVZU2AVFG375n7VRxddj2dyLGtjAoiTvB/WSuDvreL8H
+Z5kpjAgGk7QOMZ/Ntl2b37cmIne2jAj/DCvlzooc8YIFXfYgfn6xeR70/E2mZExbPX8OLAKa9O/
8LLsQDVtuXSFtnpzdnOWvIR3NOWkIuFkxuSndo9emhXpQV1v+yM3jsncd+6Sw/yrJV82d9iIdCL1
+uEXrEFXNrvU2pQ3pe+oDDFyAtXaiOt6wkERDvOGLBFIEiwxIOuhJqUXT6t4PYRmUBwE97/XNA3x
MyqVqj2sIEH9BlK1v+M3v5sAjupZ2aCuU6QXrSK+1f36NV33kC0lxKrpEoC8OFOjmlAkiuzoMGGO
QB4pm0GfZI1ay8OpDiiSSUo24wQKmmtQlc4dQaAv35kEuH7mhDtb4soyUAIskBufv8H9N838FEJr
mWMeDuUv9FAB+phoK8tnJtZX7bF3CTDFpmkuWv8sC2Xv+CoUp8e+w1jK5rrx80ax5T5/jxQLR/Cb
3Jv2tY6JqdSg15qaxpIqASGE7htuEMMDebs9GdJJ5ZpXM7KBV46iXREHnPENu2fKNZ3f6VHTzw+v
P1qlv3TPJffelHF0Is6Mmk/ZCUC3rZTZ4O2yCGtfEZx0XggNpWXBuiIxPVvQpCK6jvDoNiHVk8fA
awfxbSzf75qko3Ta6JbXMFOmHqsI2r/dPud7zTemcQnGBSCtp6kqEBhJfavSmzrnk805qo7PkEPS
9JhC7iN/yfgZwSVUSb27lXhOilFvukpNLAnKpXDikvUnSe8utKVRCGTmNUstubG4DjY2p77VEbab
U2Fmr9WRQ+l9Kpm2Yb5lFiYYGbIzxVlRafmcPvACRtLKeKVfbbOmRm7kH81vyOSjM1IesUp9J4vc
qZPLXPpjfqdrxb6cwh92bvplXWTJdKywMz4XPrv5Ihhnjb1TIF/QgAZXVd1wqVd3WMy3eCGlo0m9
OkcPfJqKy6CWTh5E5Bar71632l6azH3f9Sgh2dMIE/WoOtBPM0NNFGOu5fO1vK5RQt2KUz/A5QIL
Db69W7BuMXQMNMKUoqTKNsES+z4WYGD8xGbdRwe+Ocb0yO+fdHXL8I9qF5aSYg/ZZf1TJi5mz8lt
BcMlcIc1Xx4aKeh4ojCEQs/tZ1VAY8SvoDp4jRuo11x0IKkcvISJk/eoVv9yZKXmCTzrDH6Ab898
ujv3tpWF4fHHw5KeY2g3I2StOCib678P/6jPNSALd23kdXYt5BfLYsyA74nXX1LGKTo9BcsU4/r2
f6VfXP6ohLvLU4j/9GeCeUPNQ8/yeOBpJDrcxp8YkMVpsqZS3H6d7m+9w9ljtWK9veGusivL7Eoq
zbGOILen+XcmyGt/EyiLT4ipESgSeu7U8eaNfjV1g/U9gJCNEycag4ymD0yUSoTK0hFmvpBrYTTd
SQiNpJYegF6Hts2Y6K0mQKUByhbl1qqHPXmCFq/vMjQPuY4M+OXCwoDdRvE0lDLU9u+JQ8/LNj0n
QYweLff28vC15I1SS3xTNHMvzmYkyL3woC7bIkMGb8/4RZ6pBVyDyJl8R6WUl2HWxrPREzs8DLz3
d95HP3WhNC2PKEE1vG+J5Ri9DLMKpTnK0ZQalUxlFwErG+i5e1CilUx1rjSGQBBap7LZ9FLfdqbj
2oEkZZqrKTnuwSjfYYHmPZ50JuoU9yRdt3PcQ+u5gpL6tcl4isaOEbKpukfvaLv92MCz/0Up02IL
YiY44Rjs34CX1N88Nx43DHE9pyQFi1lQl6NCt9DEtz8rHTOcLywN9TGSrwIf5sBvYsOcz654vodo
cZ0IB0Xxt9DiCKiY5pvtsTzpcgqvh7qLqcD+Re5dbxpcIjF1iVplqFBxnu8U0KQHG0/wzQdt6NXi
L+BXqR5t/yV6RL/Pn+iQZaIH4nJdfxLZYrdW4oIbdHx9oo8vUjnTOquAeZPEZ/dGDZLioueecMCy
22l+VUg5AMYFAHD8mbxlAagn61cJGKGdJtrFSrk1DY5Fb5nt+LYs3CVlk+jqyzA8uNckGb5v0uq6
qTpszfb8jQ+4hg53vawJBCu7bEOYv9WJoOEb17xXoP+jiHmSE3ilkHiTnQPnk9/voyGutwolc3nF
SX3ThfIdSHLgmNKhpGHUSRRE7E6dyjQ48tjXV+zOPGig91QLYl3BmkhSgK2gD+Llr9s2bMCAOGdt
LHpuqBwFs2Cas7koYRFRBsFpS9nutP/wxJZZerypfvGtzaNbYG+mwTcj4rwKgcbqX+Fk8LvAdsGF
fIFeOM57/SQxK5sd6Ni1nlUsc0jqj6jA4Si8jIG1D4ATOp06i9PnpJAypMh6QHk7QkKppAayQ35Y
LhKeWnva41f6bhRCS1XRN6RUIxLUrxFnTGSTc9DCVO49eITi5WgnChYr4GNzwDd4CQjcB5c2/qep
6DTYuqcZ1sXl8BuOuDCBVxEffqaGYRUu27AvPdVQOsetPlfil6r3Mi3r4zuvfZpcuQwqg5aWKw61
JkQY/nsVWyhJbjl9OhA1jhvrdnZt+9NO0IIdek7uLmmMxia5oIEiAWx+QiDbs8PHASXOV3Rx0bA/
KvN80fhHpVrXhEhWY9rWnGag3YIuNqUCWqBoEIy9Qw2do4C3ex31ieZ5R5bP6Kn1FPXGQ5vE4J1V
g9n6XBEgN0L12lwOsA5je4WV+Ff1H7k8G6j+8v/PZT0lCH9ZmiSixcyK1Od8/4QTLpfPSQ0LM9kT
AcxezhBRqx2CmyETfKEvGb3coWpxlfAJTcOK5aRLLo1kLNA6XVLa3rybClPVfzpLvpGkOobWNm0C
n07bj/GRzNMqHRBiUoKXaIe94lgVuLlKSJzgL/SpsGHf2YogOmWAp4K6EBmG9OPBhOlbwisrZfJu
9TwocTUzhWnfojL+nwu6xb62tUNmFJSGaARdKb5NZ6/f0uo058lsw9oMSW2Y9nk1h04nB8oTtH+e
WGyhb6qViU9eMLt/wTWvtrR099Zke8DA2IsebVj3hbganfPJjqYnpT6zqU8XwA6YLAkWkJaxANTT
aJ8TPmZBALzzzKERto4h9gSfjcpfqTFM5BV69SWilgRJvjWaq5MvmAw+8D+u0EPPYYjtFfB4QRUy
jZRfNl3J47cYyabtR/Hinfs0Rqq1WAwyEAEusUG/hSIw9RKpmFdpYmLVEH3UKxzdSxvb6JqDvHv5
VQvheZmHpGA419nIVtH1LUfTpOs89XuxDFs+N8QM5i6erzlG2iMAQPYcFL267dPLxZonVsgEGI7E
682r9nJsXZ/ZZU8Na+54+GYBe3NveaD+Il5bNI4S2yzJlL1KPrXGXjDgBCFfwRkikg7G7P/D9Bxz
NufsL31FgAARw29lHUF8GKivI4cCMqp62oelm8YwV7jBnu82t1YiYRRRHYjEq97wDuJOEz5/GnXE
U5TxB4LiDVpYW57EgPO6YqAyBibQ+2s/EMjrYuyR0hyJF8JkfO4Yt+tKx9HKzmvBFU1qD8TJgTZe
pB+qJqD3CgeNRyiKS3Ktr9vpInO7dVcbocn3X0xPfOl8czcc9x/SJwVHDoleJn7vWAnY5xTVEoMG
Ku8EbuColfZvsD47ONHIS1/zjiDs8f6vtQXSGjB3cVJffse/75lZ76PINiaXC5VTjZ5XBYw52xSo
jeTYujzw3ucQfZBPmZ7F9Nlkic1PrAkowqaJNfsI356txalLk1cR37fBgWVKsppPwgiD3JG6r4t4
S54uXkrZmapiE/99M7zgkHp8jvf33oXYEPB0FelxtOauWztCpN0ljaiLAV87fLK8NB/b7h52YzBU
mgAPIKdzTCEsIikGDfxtnE0OnpzmgQJ5rujyWKBnuBI/sLrMoaDbbLeDPtye9BnVKhkrH9kwVFrR
Zc81AZfbgHG9GohHyIo3GcO3msxuw4zEZKRdsG83BFSmVSsS/VxJvhClLPsc/BvXzNUMVgOpwH7+
mdK8tO75kxvDrLnoi6G85NDbTipm9kOvRsv994JNvF6MMbDzC5NA3MGTeHdmq4PkViU9bJpzc4S6
+VpnImJwlbxp1yBnMb14adAtytlWSmz2uV18NekxwRWrX3JF5ZWjopLCaMEP7Nn+uUZEbT7Bwr1K
6mRxhavrc8rUIFJYXsB1WmBULVX+wqtpVub3yTZm13Algkyb53nPU0OyYu8fM+WUoUgjWXfZn5vI
uDsj37pwiJhDR/Hi73yDHCK9Lb9R36nOJYWKvC4S0YKRs896Wtc8lETzObVJxjl/wnselyAxRv+m
buYo+QgH77n8K6ssOzbMJMCca4SJp2f7sKfoL/DcbH+EOzzxKv1E79tuDtHHG7F13v4/NqhKTR6U
OEsv3Hu23TMKcfp1D4rO/v0RySjliQau5KhI7ykOe/Z1fGQNoiQ29F2V5gBTsGzrZC+wul+yFq8o
AJWzvljNi9HjtsxGxVwKsy9kTMdfvGlyNMHHC1T8YUtaZLxRSmDQrCJO6DUrXJXkdLCHAsRj/KnJ
vUefoBaw2aoIYLy7rBgX/YiCx/EYLNPAl7+/U9UkGlEopzFuqLujBstpu1fPfAwclScb+AiPQCPY
RokjFS4mg1yaO8B14iM+L0/Csi4YjEJq/8Wvd0//dv/0x3Iy/zYeuA6F0lUB+1ka95E3IpllEm7T
Xs0UBzFyjGwQkDqbGOAUuws4sgK08YxHW0yQzD78lJwHl2bfmYmKcJZ7TiMzL/Gzg7OPZ3yg5oIr
BR02bEgv+hQ9SECccuVfN1xKLMUvOl7K+9NAEq+rBKJO/QaQs8JO2ljEb1Ecle9lYxu6OcQeKGMw
CdIEoTHGPWjKFm5542fk5f184oyaZdU1HvRC7IAiquTsxqZxft8/jrZK3xtiQ7szh3iKczxULC1v
Yx1SiY14gdUFYnV9ob4Uza8pUvKKpWRi3D9z2jZ8co9XnF/6APC3dMMPQucKUaYlf4sEmqMGwk+5
aCoJoqAFy3y39UUKYBtUdaIrvRzC+Id7xfuIeke/+LHsgYhuxzLghDbEm/lb/8Kr3ZT5j8aeXOVc
gT+KFhUt721Pn0ostCDjypHoxdaiHbE/p2L4AKUkEtYCJhwvKHAkRYTNmC5mtc7WMB0YtaxP/RVI
fNg4AwNC5T3c8x2vdRLEf/NXedwuuPDeVbpnVuezKpOjyE/fPETKvHrlcgUfP8V82vRE+8GE3Qvm
/+eBUgYggk7u16y/rzIK0mDCoeV9WJmNpRlQN1J/JujxpfGbpOBSzG8/Cvo8KLXYu9PhHaOW5KFT
92tUXH7yO6uKEoGBsTraJR13bJtSlGTN5pEiIxkgJ0r0Tv5d4302l+1bmS5bAcVyxGVzzKaG7X32
ujXfLMtVCH2DE+PP5wj1lLS2NNofQarnyBFCBnSpV42Ac4joOsKJAsBsVH+bdX+G4Xx5ksDKJdzJ
XfzYxYWvEv2qwacROk1c+KfKF6H3AcgQr6lZt+IE/B25PQ205mLBLtRLOHXWwk6MNADECdTIdEGe
LBPsSekySefQL/rN4cPXV8IIjqEXQEHXH1Qw5jMpNoEsxPNf9MlZsX4bkx5IOhX8qzoLJQp7spTD
Zui2mYNpdiHeGcQ8n9g9eOD7HLR9zOmfLOTFjHFpgRjeyVEeBq+zbGaKevOMx+NhBjneS80+QkBr
FK86H7H2LabiXMfSi+2wInyVTt6HdZBrcryrALpBLjf0yqV6kKHhc8teOj/4R7P6+RsDAYvR6LW1
pPTHEB6SCpEbZRB8HdIaKc5Utc4NrEyKHPrE4Jya0Ia632tS9AcdzavSW3GX6PQ1CC6PKjGpvKLR
j19kjD7bmOuTHT8d/Z/ZOa9I+3SmS58psHqA8HzbzFa/JaPwPxVBN7K5uOZXZ383v1IYd+91EEhR
z4dxe4uobYGEOL4RoVLd/KEiIcbyTZdkSJbToweqg3AGVkVlWJsZ96e/1K1/vvNc9pQbgjRgJREf
rrV8cikLY7icGja0SqJrcnY2evlGcwNZiEp554XZqYgwHOMudwIvaRFY9MBQ2ac8cAywheEKdLmP
YsWh31+fmCm7h+eZjNEt0yPa4LTk+Xq6ycacF6fMKRFNBTRnTEJg/4RbVgyzRjfgM06OuEyUoNFB
Y6fQzk0ym4T4LuEOIbrU9dlUhcIpufyEG2FXGababJC3qYqQUfG7K1LrXQ8U/reUpU14yCpqcS55
STlcXtB0E3gWxd+fPzbg437dwA5hgEGI9fYp4cwXh94fg5Vi3xYCHMum0Q7/SAYs+CDERKg5qwsy
NN9efKm+D37vKFRCeeZru5vlv8UIh0FzHLwct9NzpysqYtxMkzhS/Pg8j13bwp9HvdET4u/FKNFt
eCIBAOIf9rZPiL8rp4N023WDckHjuNj/GnqJoQ18uqsGgUBcMVWbxj2FMrFPZgvokSAPuiIvMALR
6kTRBjWeGvmPpfDQQhrBpaA2eRlm51A5Wlddtbcon/sajkjbw4dMuoli8jH64D81UDMRi71nGkiP
JDQPlrjjpLLEIkXJI3TScovmuXCF8UCSU791j4LBI4okYXuQT+MIPud5N1n1bzoS8S48Bp9yfFdm
UVbXjZgYtvB/MMBALBKgzFP+jpSbLR2ZvFj4mNPOic5hzOf+MUbv7rKyiEZoophR40sqLnPp7gxY
wvUJZkCQ4zW7zi8VQMgYco5/ww9UVxrCKQ3myFImwEL0CpYJ0Kh/K/lH94uyd8bX4fasj66nsoeX
9BFQkUEXq/anZ0goCwXxkLkRIbVGde6n5aSH2JxJC6iRp3I4escKRyoyoLD6VBt9mt1AlonWm6fV
vlYu9YG95EEe95Mw5vEOi1+Yu3KZQKFlFh4vIWkYQoskcAmQRQ+BKi924G7Yt+MsOb7U1wTQtpVT
4Fx8O6C+2AKJfjzERjYULXg7lMTU3PyR2hAT+vT/H7n5ZiWJ60jzuJf847AV4N42C+f7cgyOp4o/
mxLrpbB4O1klZEPKDwv/2V+mKqwP6OYyCwxsi8BymuHs5UiT6DpdXs5UneguNVfBuyMwp3axYM+W
5K1FjfDxk8Q5B3PsIZ15B47HMH+7az7t51foG1Nf7CUzLu99KVOJVxN+mFpdoJ+C/Zd2i88RpSWD
ZHLa/ShIvlYdYe5HnBbOaiNegVQKo12qFVwXtptBROijwK6fEJJ+fXDuSHsnivtDDjpC+k4kBFOg
ARqJo8/tOv3Tt4gn0q5/gSzCJCeP7SLBgPWTNfpmet8TdUOinn2izTNDqJpin3Xbaz5RJT9BlEeN
n4DE8ZNvmSWsaIzn37T6e3b+Vvrby0EcgrLYyCgLK3RMC/uewupIP6YkGrTYrivcpBEmvB/oDlum
8SQ/lHKW3YqvAGKZilpUp2qiLYP82CLfLq2DcyMkmI9Yv34+gSR1K0H17n0xWpL7La3JIiziH36G
W4yJihpIRUJOsK1le5AIgUlLed41GzaaZwQBMc711Qm+mkljyiAfHQ8oq0Rk4JfrpGKeat3FjX4N
iDu4Ll8amHATXMlsdogYo/gMlVeDYjdsYjTNjYCjlVkkH7cabnhDrkVJHTsqdGJu7eZ28+hsYiXK
EdRy0n5Olr3gmJOg91ODB3FcGlBuEbsNQct10RTUQc/5X0Q0Yba+sEkRfGG9vJy9vB7fKW3lMx1m
la3omXn9fzsXla5drF6ePe+8oZlaA9esDAkvAJF0VBr5MiTqY9fCrKvl1SXARl4CzIlFKqBFuRRa
qXE3rrdvohxx4Sd+FA4snDp6FXaCEFqEJ1LBrU62V18lMbTbsDINoXsmWFQjEOq5VM77vMxEg1NN
7qOdQOoq6OGhY5htWN2jRhV7J+7jkheZ01u+Ob9tIwm2LP6GMGaGwpiLOutTlcS2GArLkYXq94hZ
XHq3kCwuZ6glMOKC/eX2ryYveZFbOhgnezz0zt7vYkAC8LNsYlCpVwBkqbrBnIG2FCR/WienP9lY
I53bpCdSiWHkReHh7DBRILryE5+YZ0csFCNuK0fyRPxQyLtE17jO1sV4ptL1NS3dqc4iMgILXkHx
MOKwg4q86P1rN+7Sz5x7VutWwz6G3WyscWPawj9yQsfLjGDrZKs/gH8bAjgni6rZWluaBpG2UrlQ
m4VFN8Imd9zzTVtifGCOJWPiUQlWGMulDOF/j6YzF/bL7D5GC+6IHp80khanodPBhMx/Bldm6WD8
JfDkIOMRbUZDmAdsb7NHwSlFP6kxIhoEUkQd6mgX1iiJis4n1alb/MkBUeY8dANbSsgg1InsrjGn
GDQI8YyJ9wT6gk4HJKblBwarTquPXDpHFcGHWX1fYI3QBI+e0nSIvIm0mpVRzAdGRRy4GoO0WMOq
5QFTp30gN4Caz1it3zt1NUWUlhjVLsaZ53ZZLcmhQCm9pMpndfVCiUHKx6k6olAlE/YgUHX9Mg/W
Ah+cs/UVhB5lg617FlOBlPoVvaUIDJPoyqHm7yi4a87rGZgMlZ9QRYTs/46btDHNHIK3DUdmtc06
inix7IX0MN+Jd00ZOo8aBGGYOWAZ4tHcw0fFl2MRj1UtjTXpTOXg1x28+6s7CDtUE5getAvNuujx
6oCyBEK2ZqLQDJhCL8/3vrkYTFXGISx+AAPHdZ1MeR4sxOSfuUimYBI48a2WllHog5dx9o9AAXs/
UGGZJ0rjDgo2q4L9oa04YZI2mO1Xw7FYjxDVq5e0hq4eOJgT06hB7ra64+wx3I+7J22WTIdmaoJO
TToorB+aLcVITT+gj1xvXrQSrzs6TCWdK2M10jgfydgBF9E/H5oqD8kZVc3+AKFPaAqod3bVMZEp
RR1AmrHvwpR447X/VchXeE2HXLBuYSUFmHgpxrQ5n5Z0SiXprrjzKOqMnksdATl0zHkW2OyqI86f
wlAN9+UKVJUjmrLegORY4XkS+/hRo4H5xQrpLbjVeaDxl4fvwXBeiJMlYE92ghN+rwRKxVu9WORR
iZY7cbpd8fdDzmLA6BmKp5vOhsfV7Owimtypo6fH6bAI8SUSETRjqVzbSNF2PzyrVNlM5Ei7kujW
bOaEWSF3hqbOnnVlZ2PXgcliQQp0//xa0Dxvy7Zrm5zJYOp03e52Q4BwyBh1HNlFr+rTj2zZjm6q
aN93ZVCS9ZOH0AQSk950ngl3ow8QhqgIUNbOCEzwUsHScXP0T/+Hnc58uZgMBSqycaO3Hoh3GGaZ
PgbkWmweOPzPelkeBZfLL5zbRy3hwYx/KRFcp2RWaEE8XQHx1cHPaHNcneO1Ay4rm1eBhkVe3Nsu
rbmBZZ0Q9FZ21dv4Hw2pUG6D+kGnETc8fcp7IY/X7ZqXOrSoWH7eHkAjbjBQ6XJ/ck5qNJTtJO8p
4GoJWXBBaLs19IsR0asbbIhZNWHzqzJOs6QuP+ATsLb9qA4BXfMgMEJGOxEhT4Uh8Ue/t/pcZlcy
e/gdntraq1A0a1bSNv4bgdPeflmJ2ioBAJoG8Tgmod3fBeIpYKfQMZn5b6ytJ1s8iFsGTIiCzEtk
m3zj4EGAWpKXChsqLAOUujeJSdRZEZbfsJT6f8teM/YavC0fJXDGkQZneclXJZobp7AN4fP6CMSs
lWcvMsyoleNmbj3UGwSBeNoInayk2fSW0Dbpy5og6KUG8SJviuFW36OeSltnHCTzN7cs/UwB1oQ7
shP9V0lcBoROYuBHYvKz+pkzMlzyqjpSR9GxBDWu0Dcr7o32P+FCwMrcP7Ca1NX0UyquiHU81K8Q
YEA9uiEWxYvucHcw/9SOGBRJas5waz+w2WZhTL/jqoBt5SqEuSD54q7EXfhK1pZhMzAJDVCnjtwq
diEFZ4qmb4w/dWlZMewQwSgSAWkZqrDhpCynq+0W8zGI+ivOjgIYn4b+wF/L4hpUwLWCy6EWIF0f
2X97XPWfP4Gxva834QyWenfdwehLRZzzAziUo5TKHH/UUDSuqfHFlAzc2U9bqHXuIoR/ADgQ63nF
PfDAaeMtfVNtyRpdrNqJs0U+CM3jpz+qoHNJ07Ky7UGKZ75MmzxtjaC7yJi7C+HKvbgQxWyz9hHS
sYmUGdbjxmp27j8/VAnrBRtJUzQ4EJ7Wt2D+sPxcRkzvzyTfx91EiyTkg26KIkL4oUCNtzRZgsFj
BjqA+sMe5gBXeDZyWBnHEaYg27AmUqet2ypou9p5ltbX0AEkQeU24nP3hAXOl4iDp8kTeflZfa5f
wxZA3EQqQMSYkyKP36OLsoPgiMeheV5Sg/B+jvG3B9vaGdxL7TS0YitZGH/kra7qpqXk8r3RNPmI
jrS3a2TTzV4JmtpZDGBvExsqh5uk8+PHVY6fOr15pt/Osju2aP5xwR8immd+3I/OOm9rIgiH/WZM
JcVTFuMIOM1M6VoxPFdF7NIpcVTeqBMcViPCkHYfqwXk59kkNuuXwv4wJplerme2z34U/agCsnjA
AYH6Gls1H8MFJTNiMYS2EssyCs6BR4S5xMSY+Gydtn2G53G9as9cXnFw0pLhR4Wt++u1wuIZMxaZ
O+tjGhmzh/AyApPG+HUJGMvHH/tyyam0ci7Rag3A2ty1vv9PRe44lg7lMlM3d0LXRwar3s+VQcGg
5FO2KGqsTKP1qqa4zILoXMXk58FFkCfafpLETNjq/ND36y6tP50Rb6A0FSjjdvvjVNM8wkSpkkLY
mn672EIYTud+fWhppKOmVgfpDn9Kn6c2K695WPFJgUF6pQrn2VBA+mNNjH2MSEFeDbIPCWRpUzbu
IYkv8UM8mKQrLLTSNPNeGHU3i48IaNGbO+/4vGs0qPIB1bkbvZGd87Lv5SRt6r5N3ZpbR1aseA0C
ghSQOEgDjJhualdrdV9pzwPVWme+F6VgafoNvxAimWxLk4eUBuyBjK3TbZ7eG79zl3mJRBFBFrGr
Lndu3EBkHjT5wTpVDlKyyqeW7SwKgBCBY9uXA03HvaxD3S346N6ItBO8XW/1qxRiCjXtugnF4yvt
jHCKDFKjrEbwD7zrBtFx+m7JBYB69NXe/JKxwn3eePSQcjn8G9E/fS3bKosJePZSgOHDnTCsESOc
2wUHAMus4SrZv+qMBNhEco971HonwXQ0J/Hz9pOKX3yHFmEfhwGLetUav1YlngCZobHr+2OTYRlX
G1TLVMsyq+I/fSUZ40Ygap9w86kNQqyG5rNGQkaSWJRjSSiORDbm4nF8+1fnydsFDXpTpEiE9nrM
UaiDrbwgqlX92bd3FuUR9BvrztJF5oSPuldpDlegjwcVHGHZLgWr4rDGT4Xj4I3aB8mM0LJ3RwSL
KySPuoEI+lpchLdKiiWmm1Tp5nJzt6yZ2A4jsgJtIgx5I5wSLn4KqUSjnaU1Ip9CfUIa/39LiWbv
KWQ5wC7HzsQwuSh4hHYCeWj9Agf2jpDvPewe/HkrgJ4UJD9AfnaHCoZ8jogFQ0Ic/mDHfvg2CJRV
kB+mug18NHou60CgdBXUKVJ74DmjvyOee14AHAQEV2o1Qpo8dmLtTKlw9tAXkkoMqif/Ajvypxqj
/20IoFdc9wUraz9ZcLIMqCvQ7p0DFPuooTJ/dPQgrl/CI925P9wzJX3TYySZHMn0KvxyaFY9WNLF
Lavdcb3zpNtk71x+U0INQ3B0FWbUwevR6wf8U/mB2auCxeIgHmgsk+odHWWgv85Lwl7lW2nZhXBX
vN3YEljaTTVWVsHtnD+UyR5M93zt5p5OC3ZF/uiHOCtWJTYQ3suGNoZwF6z6R+PQuONzCezIhi2K
m/4bqKgh6bmfy2+kTXui8ycqqtb0cRCiI/CtnqqHNLhqJd8IBF3udotYU0XH9jn7XIhBY5RZ2z2c
fJ+74MmmTude6CYXbgOybwSq+RxBqE+gQZR885ewlcDbaMQPkBuc/IsN99g+FNkN/+N+LR+x2yCM
lzXMrTUwg4XX4Ogx7sFd86U0sIrQuWcDpSpA+na2d8M8jJe4fNah6Rz3UUjwGTRmLgox1vCTz4s0
3HMQYoF2YmkeH/j8vYJY5tOYsh6/Zt4nx0RbawfYlxIYPKSgCIQ3DT+y8hSd+MNGhgf7UFzQpxtb
OgadhKUF/1jfBsH/mJzA1KkR1w2/7Pt4yK36ZUjw4keSKi/zXaf3i68xwj+Ia5wpEgSHMYUo9fXn
/vvElVB2bYQniAhfwUlXAvnofaZJvxvypsQ7yA9ivl6lwCBDkNvUmYzfbKCGdVsttnkPohr5laNW
7qyQDDZsVXEV/llpuBUwwH2wkoYuDtl+9+L4Dhg4RQ0kDYN+Y87xeRV0GGSynZfJKJX+iGUjd7E2
IQM5jq8kLt/Kqb+iOepyaCqU8k38wdCtk6AKAq0g4f8vEfvU14rX6i3WTLGjG/g3qXfzJhNbj5JL
7FXqCGgidxNfuDFHpKu+k/zjlhK1x15QteEz9NGo0K0j5Dkcrf5+UE0c845IaJUB8kLW6lA3Tvx4
iQ8ZnDx65fexm23gfp+lkNs41VdkTdYaEZ753OUrlkt+vj2ZyF1hs6fkpwnRvNwX0bcdpScG0O2K
yp+c7sKiVPkL+CLCXNq+mPDTxXf3AAVT9rKcJNsuhnAqXF1026om6v7zKgNloV3KGelLXJ8V8o8r
K9aJ+X2Atv2iuQHuStmHfmcq81O0XtBjuSEVxQx/cxtsZ30wkuqU+32Q81KwBSlC7jLmaMuECicT
Mu7Xz+K1eHlsihCuNNseX6OJ9MTjbRjfFrKZXgUdUFVmq1rJuGgRYUojtayItYLNCBaMJhF/lVeZ
zwxepISNXpV7TAjtoXQDxi/I9dgRAwV1DVGmkZNENxEsJgpA5FVANbl9esRIfQmXl0VazUS+ObUe
mrsM7HVmVaBw+irc/c2SQWFr0b/pe9Alndj6J5pSkusai4db4fa1mX5BM/QU+2xjiwTlV2Z5p2W7
hfpe34Y/kztPB1JsXQWQSeImi6TRi315+3KByfwQVR1Zx2bJEzvZ+htCnItbsriwLnK0wRVrWyp0
CP9TBOuneZ1mbJM3BRp7IYd7/Eqljnhc2WySYQLh4WIzfT5BcdBvyehLdWSxMEXHyoGFVkE3/pxg
94GEtZb2dqbmYIQX0Z9LqGEIIEKE8S/dYKCqb+TTbc7lKqUiJDgAKSjdGpixjhVMXIz+otrCrLYp
tcJBtDRHRVNXU4iUQnZ+QWbTj76Ut01zS5jgyfQ2L04AZ4LIL2zxchInbHF318DrPB5B60DML/PM
LqFabDoB6TE/jT69smEzRnnWGcVMZd3cq/ZgGmgdn3SXX5Y0+QSrbD3yIwlgqfSa40ECYeFc/h6X
9WlfKM/wXnoLXnyPWRNIwksP8ImTmR9oGntGNW3FWoBAJjXEOVX6DqT1G8fE7FQknCBtcLpcen9Z
SpCk1mbkVLC0hCsoeeJZ4evVWlDZKdd/553UnAQQ+chsXCdyhHTvEmRkWfGAUboGVG/KQB5/h8LM
uZOYNS811ym0tslh/y3gnixyQ/ssTbUMQYhdiI4FLm6ZPsQ4i+lVY8LZCgdQRffCaDv6jQqkM4tm
21TcvcdPzlj79pkXs6z71EHO1sEd9zFSHctR7+uF6fdvNlR+KP4GCSpZIH/n9cOszDtwKFZXlCT2
9fPecTFUZKJ2i0XQjCOmKAqKemSAm4KWyE6rpu93V6E8uAJVj22oxR7RFhebRtG/2GJ2kQT6iGoo
6dYaM9B/9gqAfh8/6l8mC2uPq0um89hOl8SFFirn93TZRvbnhC+C9DqRtZrRfXQWfp2H8SFQA5K/
G4SvH+ESs7CbK+0f1U6Kzt0vHlTQUhBSTZ/76O8usiMULrz7MtH69afFoEBQpt3DuyvR75okzh/o
S9H3I0jClUfUssXLJEMSIG7VgMo9bfGbTYU2qNLwKX2XJWiBCXRp9BJfMSBUSCx6j2W0Lfke+6nF
HgeJwndCdYOJyhMGlxa2fmkDABChwt1kwJWf5J7i0wIOr0fn7MJ90Xh2Eid3rcfAFJo+ZpY/o/1O
UlgtAUQZ75gvWAyJY/olUbhTWoMlIvWMKefp++Yi+VVPvwR/fY777eojwhIwSZ+z//sdcmgMqpgK
Sps+xXj+RzJb8o6hqjQjVYq3R1R6AJiVB5H9CaplOgWJ4cvApyD+c7uN+8VY6Y4SnYCjq64FNWsY
r4vzLP9QflhWFdFj7DQZRlzuZISNbdQtH+g2Gr0Pj0ZxCk7O3lnfDLw5VlZyngZQI/VnB4lDOwrN
DlREmG2qKJ0lWnflJAwA45WFAB92kzC8ZNwNlmfAW6qAcByj1juuNmggMnIDlBfSaa25NZ16dm7c
BfTznHDr3DhqdEWGk47qzYFHARCDJvjDT4Rpo99d8S88Lf8af0mCSfdbmcjcgjOypD1Qq2zpOACE
E2LITpcjm97uT2+ZN9uhsjUF6QUsjJfHpnxztJIiXhQb2d72OX7f/Kfaz0E7f2DAcfbnz8z/Epl4
RMGWStm0MhGu9f7kPx+rVTsfD/cAFc8+al9NR1XksweDAHA4c1r+sdc+TzBQqOV7Hv6b+YyOGNLL
CCHwtOePNIhZsWM6XLhcttXqvjNbLIoriPNoZRR58da1B26f0XmFESQGTOZra9Lqnzw4m5yjsk1h
xD4ab5sWQ9wnp9VLZyToLCep4Nj8ZmlAepRzCWiMiJS+FSm448gw+21tC4vv0akL00/OZ+2RyjBQ
uRcvnWcW9Os64l3HzIjc6oBH1wSzUdgroD22n85PEMKbFlxA/ao0qgyhfbg7zO32bMW/IWFKA+z4
qDYcEiND12hLjX5b0sDJDj9PuKCyo86aNX4NB7KhWcvza/AQMqodJVnRuKQ4pNDWM1/hUnu+na0t
b1leqzB31He5rg+I+cR8WXtrjJngybrrzH+G9hXIcltmkPo/uEn3lhbDW89uFm3HyvqNmlTCl/zC
ei4xaP1iG86UyjKo729iiHov2dzne9Is30FNcubQIN5MJ/tEzebO/Fyc32yHCfY/TP0fWun1Q3pA
u1MA5zDxqBl3IdxtmD94p8ruVtUgewQpTWlmlXaluy4kKzMzlVmLC73DoUoDwLo42l7Vu9nxlj7N
jrB0K36f9ZwUK1dWCeULCoFEAPUCVlJ/lh0mL6e11asBRyY9+rkaRFTnOC3MxHMgTt4WofOKryuo
W8YZmQrsQLtzEydFi7TGTInGCDUKuH52NrPUBqRydSbHhYQn5r27/eLkHZ2Eo2VWDQFozR+Ej7aE
UE2LS6QAPmM02uFIly/OipeQiXpPRCLmS4OF1hD6J/Z7xHKZAltn0ulgoS6I7ZEm6xv6XGqCQmq3
2qDsHLaRQIDQeQHfLV9sac5qs52x6M10OhAPMprWs+DyT1E+XpmBSQzsMfVFXOENBP8L/+9w7zlb
2kxe1WapvuSNQ80v3ASLvYll3D1O47/BOy1U2f1hpo0jdice2vsoZk5evxR9LL+lsC8erXMlPNA0
A61VawUj/7HG9S/wQwNoRwsoejypB+kU4xmHAIZxtyxoko1QiB1azpRDPVSM8ETJyx5Wc9AutHZm
MtVy84W+KaUETMmk50PN0wR94mkUdTYpQ0ra5yCweRmIjpPYFxV4MEe6ejoxBKQex2fYDFQOxLYw
FA/sxljJCjYFj+mxoJkMxZWZfn9g0t3I5QDOBtxMOJgWMzScPm26rUJOMaD9vt1CSktDOn0X8TT2
5qyH7gqiW/pCjuQQ8b3jkhdYHIkYFQ5NkC74xZWaZ2z+vXidGhIy6frwkhaEJN7w0ukYrp+DfOJd
ZU6vApE8hpkwU1J7FQh8d9dNoliBi8FFTsuSLRrBSE+VDucHJdBXK7M6ERtu2fZYu8M1s7z32vdF
h5axOZxxJ1BThtuSCK0mcft38TbYo/ywmZIGvmRyMGuIp3EcgoijZPrwWvT4sCWhKAAxo55DwkLP
iIc0KmihY9i6wyZhlpAaedMdGk2FYZLe2WzV0Adb/ubjRtEZbL1Vgn8tPG+5hAg5EvwH12jjixFU
cvOyiwkpR0W74iocqqGPoUbYlyaysRY4vZ5zjJoH2mwxd2HtPiFlO+qyM9dDQq4OP1NurO6cJqJV
8zkwqqWQ+sSCXKQ8/NW84TFpcPN6YXSBcBzJ+SPlnvkF7K8MJQwjH8FBz49SkiEVala1drh2LpdA
5DwnJksKDV6VBByxJ1kRVa9sWm0y7YpaCzbiRaVv+ddgNjv4MJokF1MlhYEVfsHB+UI1TCIfZr2O
l6+X85pvVK44jPrqYZAuCCJQ83o9gP/m31oTCNS5qjuhd3/k4Tbr9zD7OAtxHkcNO+SorgyEhfDm
7q5v5qZ+T+co0KGfdFZvGCELzZTB4jp5J5EuEAKrCgjXpyBQp3MVEFIK28/duOGzIjd8u+J3aJpD
qOiOWDC7pMTkNFLjvQWQIy/EpxJlhharU6eTQWgGt40scgRSc/xi+4hih0yLF7vrOgQz/qdv20NG
sHsCTCYYDYQVI0D6RM6Pq9J5I/o4VDeFECITtej9PIIWr2xFcekNqdJYF7awqPkOzhlTHUpVUPv0
63Gf3XeSLpGzhyekOnQ7IbbzP3oIEJGa5l43LrhDT2Lxi4WPz8CJ9G0t2lJW8iChgnGIIlHF9oKN
1ziD3WvKkuaAN9rw3OYN9d8xlDzJU0ekTFqkamVuGR+Q2VqA103/YkId6KZo5d0nkR0XCqwr+IBe
smcNAUDPiXhh4R5dF/C601B7HLH4zieMvx4D/qO7nvXKRcBvgwl6lcoEM4Fx3yvEkulH6jx13kVL
WV7HP4OJpKyAh+SkItwppz7rojTKBYTZxnbyEl4EB8jX0sQLCZhp4U8aLkg4LUsem0qPVzzzZedp
iB40CQi2OCXxVm/PCDJUcCejBqNg0YrnzUZXX/JodlkbtMQW9Tv22W/FJvreYxFzlgKMC2y7xow/
G6rxCy3ucgESPDNzXxIgN32fCXNA6A8TmBgJ3vG2x++6tNgSIefa6H1lSfujiLEiARpHBg1Ta9/P
pe8/CtSmwVVj5CRuxidR6Ymm2MObPSAziU4cWyqN6Is7Ud/QRqXD2MFu0aZ5QytIsgiqtzZ071gA
CCkiCbc/yQ9e1bPraxiVrBcqaqvrcG5zV96QZAxz3EqSDkS6dnmA5wReCvBuSz5bhX8zZv85bsfm
WonhKkxawrEqSZ2GOv1UkRB56b8654J0oUCb+QnvzCwJWoPObh6HGrISEF8C7kMxBpzbPYUQp3ow
jUVJzaLamB3NyE/TGjePIz6D2qoDeXeN2WVY2qvUbvCjJ4O8BUqs1yU4MNG5PjTXz+4y6O7B/bZW
/T0tvFfGyWLnn4wOyJj71R758PjQQ0JqBGAKjLXcVtqc7EcbtsT/jpXr1PSZ7vV6MUViUV1yDDtl
KU/dWooNzTM0C9QMRfYHs/y2kaO4K6a8gQri7b1Ea/0G3U2E/oLEm19mC6l8XkYwYMAW8moFty7R
UfOBD/xG0lSOMB+nb5IKnubUNqokbH9DNK55WjEDm6R/q54EpZ6CTV2EET1yak55HGXKryhR5fo9
k7mUyQKsfr8l9gFk4PfA9od+rl4IrX+CMJK2yYQWT2W5R2hqeKmthaYHqBG0RklTGQVNbBlm+feB
9z2a9F+4SUgs7qqJuluXoTZ8GAy75a4HSFFm4qQ0YPDtfbkMZYlwbkjT5u0XqIpNd/949vvgwTmK
HLRICdkHl8Vsku8IA5b5mB9s/PlpGrGsqBWGwnZO8tmK9eIP3YxLmKkbiPIyHHsIC/5TjtjisYhC
etGEYn6vuFTMrTxQO7OcEd0fuIpUaTa6YQ+t1bU+P/5ZCjX/qOWaPiWJjxePW+f0tRrzv/8/Rqey
Gim7PENSVYmPDFHwFgJHlNljbReq/MOgrEi0eArhBSbDWq5vocidjW5F0iG+ji4UjsHRbf5FiKQQ
8elyTng71UuhS5gmyvImMECIoVjAnxmm4zWZGKT4mB556K7YBNNq/NkkEjkSBdC0WSUb5K3U1QN6
TdvjtxGzDHIDbkBus/Lseh36zvzqg5e/RN9PNnjzLyl7zlWtF5zBvURerPiRhdcyFG6gSLMmkfjA
YeCMQh71Yrka4sPgoyEJkWJHmG+ayRPSw/haDEuOTFedca/4NEwDG1+FkGwhNGvcC4z6JJEuHxrX
gKYed5TNrvxVcKXW2PCi0ztSvq+u0DE7Idjwgoke6HELujjkox7fLkSbd0p4ZikUVXXvNQu3DWV6
DeejnlHfO0D1VX0xCRUdMwmCof5ZxsD06CmTPfhuBZ7uIfEK2taZbA5QHrHqN0OLs+jJQ3qow3Fz
mnrFw+5iVZmX7CPfNPoeQNHKyLmnm7JwZQGXFuQK6+WOM7zy47p2xSKavd0i4WOSdOxDWGNQjc6u
SNHl0uan50lnDaluNVfJv1UtNDayy8GOz/QCN9mwXqWKjYiIHWZaIaBE1ak7JRy7yOP5GURQPF+H
S138Hcw57Jdugbcl82e2q+g8NnPP7BAi7SP6KX6hKW1n/dWzTsHUrs/jmfTUG8IBdxZmwggVklvX
l1sCIicidMYqQnJW5SYjq+df3sPZz2mKTsVBk21S/991toPyEYtb/LpHVrO4rb3QU4x/ylC9m92e
IhbQjZb+uoKYtpXkEzl/SgxHZv63IZmFAC/K7AZG8jWmtMHfxDgFmOsKFMPu2vUbyNUSkpGmS6F/
iG/3y4Lxyg5bfZEbwa6uB2tpS1Kj5JD3phbgCqzMzpf4DHdYftEjFvDhiWOx36KlcN9VZoJjpEbd
+MKaY5VYm0WDkgzmn/tI7uHX6i5oPa+aY9K+ZH8PxbvV0oZR3kKSJR5Dl9wF1jE/rMWAdhtZHxbF
L9zYhUuYtcRL292c/udEWWGn2T5TTSj10cl+1NgIQdjdKlMZ8wHgatvJRgfPL6m8Z3kb2c3LdQ1z
/UjMTs/e9XobJXFCZB5vvI9W+L++x5CjBnt6GgvoG45vK+EbLs8Aihja/UCWevq63ELVqoC7KWzz
7Zf+uvBpWnpg7WUJioT6SarKatJWpthIn7nVp9VQU0LOuIg/8VscEBber48F6iv5xh4tE8de8srU
RpRqqNkB00mCpZVeQsNcVnTd6NSncTztE9A5sBa6JJp7hFqMFhF/IIEYcP8f2DNPT+O2oxNMOzkP
WUk1wdcwv9UDTp1gaiifgkZCcxx5ZREO/+Px8SSxE/sPmosH+iDXeQqOKnLbfsx2WXVULdXDWQmr
a0p89PNYNmgLs9U1BPTnJDgRkcNHyrGK9fsNe3sjASS5t9oPCz8a7h3pfTe10SXDRto/4ekQwSAT
jEH43GAmPYSKVUtkKBI3KdMXhG6950hUyvX7kxOyw0ts9f6EpDDXSRLMqs51zZq6amzOcM2GWWOg
MHnq1xVAvVulRb9/Y6rFCiT5q2lQ3VXgykSdAYPW0XF4CmwqsIyasdYqY2+9AECjm3WkKXbp0EsY
K0TQV41FaGSaXW45LiZPVWZQ+IMdSJwImCDNkzdGb92rFx+/HNB2u1Hn4B+98UWnKuNgjKDlvMoQ
GJ8+tZm5WPkfa+Ry+3iXFLcaEA4Vigmr7Gc3Ehi3042d7x+rBZ7J59ch8Itg+EYwMt05BuTgfHdu
R2JLJa3df9kXvcYYlfbJLID/AeiDSR9ZEmau49MxFutQg7n5+sQuvD9QbDuz+ra7HTx8c1qPJYO9
wt5OI1wzUU1vm8o1njAjESFXyqdJwUxCxVh79TIxfhzzkznGFeGiXdoiBoW68VE3Q9NN+Hj4Ofrp
iE2UXUpc0hupR4j0kPoCpSx7kqjnOl0Gdc327xdKLZVTnqJaju69AYNBv6RFcKnnJMdmYENX3onX
NVUgAIfB/0GxQpyNKrLOpw8pGDJ7ry2WEkuLoRSbN/rsdMkTQrHS+C1X/cWgXLrkxO/vcujIMP/G
clj0YRVOQN9BNUMwlFXS4alHVhZKRCt01ZVwtuv9zTmoWWV/dvx6k8DeJNzk8mlcBI1GkXNEM0ZU
0bS6MrMg2vuu1Fa1g7vY4fCuW/iwPXt+tcekTq04YtuEwnr2fbB75RuKuiPapdGTxEPMZlyHat3H
9YRVoQxXiWtVKawgXA1PthE1wSP//QlObE6jefrAVoXhFw5ooZdXrX/7FpKgn3EqVPJ26ZwpET4R
IALq/PvxKlgQSOOrwdPTl+mrF+JdOMdAb3nw7cbxE6b0RjEbSTdg82KV8FaYvUfL9lAvNObF9E+l
5bS8dbR6zLvq3hutNlSvJWFkGtFIn0/MqOC3tKxRu5Oo5Uxw+1UGcr42Ad72ajjy3mihioJVikFz
XMppvyPTORuvy/BoOLjLGHcLsxHL+IxjL78N+fBZ6LwuH9/GJ/H+bAGekFmMWlaIIzHa40t9SRzK
wCluRKwv699fSwUDEZTC/mv8W4xxxn+xufmGfnnzPCms3Bs1tT/dkH/wWQ1KKwypDuVrzZijoIE1
OvpkXUuC478L4f9NB37Oj2+QnAnV34J6G0FY4qZQStAyJ3aYsjCeSRsQL+fkjX6EfM5SoNsR8OQh
c9/OGXiwdewV1rZY1Fqzics+PNXTYdSP5E3pBZb8NKhrScuLm+GwcvBEEzSvwb3+w8FmC0UGVJaH
x483cQZxF+LYSsl7IxhFV3zk4eWWi5RgXHNMXw2trhucuUSB+1ZMYugv0LiZg+a3Xb6CcqK+Zbcd
186dJFlh3IslTpjgBcQA7X8dNfg2kwl4zNcLu0tnyVS/fQWa5KobF9p2XfHc1g65z+Es4Sv1cvVm
VlqXWZwrlI4OGyUVNsmnWT6M+YYkm1VTTf/QQUIcvLMMqKUVuKQfonKENbC09ZBCLSXhN0sqEAbl
zqQpuhN86OZDZ2F2DtjkZD+12ymEK1k6OKYvN+zmgYN5FaSY6ecuw3HdvKf40GLO/PbN0MDPQJwL
IFkxnPOLRaUZPJJT3QkFeSdUvLQA/DzIDmMIO36TnmeTxHpjy4pgkdgwGPWPC7fZI7BK3XpdF5v3
T4nmoI6Jfs2OVx7bFTq6QHR2IkOUKxUKdjQSQB4beWRqIlkp5Fwo1PDii3YMNX6kRxjG46b3V7fy
AfYnA4wCqYjSPb5+PjbzvXA5JPpBCZndsv8c4VrdGIJULrO3aS7Cpxzvfz/ziVRC7GsGDvkhp+0O
PlaBuJTYp/aXdzDMkop7B+hm2AzDg/wG0EfOxtEk+pU6delAenO1aqFuRJ163pDZtWCISegakLjs
WWrjMfXNIZo/yH5nw7Zx+M/uwHeARCaw0CrB+gbPM/fJRZ7AyqQj94J7ZZVkusqjRNJoTnIGyh+Z
VMMyct4ar0fdvzukRAlrvr+/K7vBtkvwHWNN+bJsac06MpJNFS5ffwxi16CRFqhjla7oDh78Wrst
R3z0c/uAIXh9kes9uVtdMlMbUrubLAhw3jGRkc2yOlLztdiPnwIUTnwwrRzZyPp5sbGsS+AxsYB6
Avf/L0GZWBZl76XqccLgPC2SB0omWlFVLu/I6ttsw3fLmp0+TdIomKMhtdzReNdINwdoAJq934YE
mxfCRuVPN5vNdEtbmTiSFJrQYvNKe15HGx7f7y8NKUk8t7OxSIcvOpGop0r3m68MR3Oz/wcjlU4t
L0y0k3Tr7XBCZZH2RsOKQC4GtMu0DqxDEvZJEgfJncoHD/q5a6llrrB93VxxoLU6GRc8lJYEe9La
CAy+9qwWHToeWfMzU2z+Q+0oKQKXCGE0LirLHJSNngUaPm7QpOvGSJyH0Tm7pmVuyxgKj+u7SB/V
s9M4npQnCKUg0WfJScTC5tSkvea9n2d4SQ+4Q/IcjyjPC/FL8lIeCjICa7satX73qhfacxlJtD2l
0i6+CaIPR1Fi33hu1DlBdAxipUYJdUScFKbmii/zCjOHtW9Fr/WVLwKL/af6VDk3XnND3FsMw7lH
5erADXoYikuQ/HVP2k/RhSr5jqcXyr5hLUFKniLbIdZf1y/iYaJm67wK/kScfzIInHaRZ4T8EIO1
rJyP+8dMz0VSegRZNK2/+0sfbSbBzZraiu/ELVjYxpSOj8jPul6aSzq6/TC73W2CJHytwoFre4VI
mt4hTtaYr7CpAsy7eNsQB+UHtgYWH4meTQYb5DF3Lu5qB3DzlnsikRY9fs/DU9+aggeJe0SQ0EVs
GLU+D9RPZ0J9eSZbVT7EXIi+G5QN8kmU8vi3whxaivEk7VEz0QHed1Xcv8NCCEwz4mOmbDt7qvFm
IOo+hc6rJgkrazsSAtjll7fimegxr12a+i1KBDViPqYuRJZGxg3vMQ4rTGtkAEUvXddjx4U7fqbW
6XIu0LBKuOU7m5lZoJFi3DIc4HWg+D2GxzOqzoIuJ9BarfCc2W5KAq6INpHJHUvenXwU2gA58fya
Ud1mBxRP2sV3jfMuhQV32CS+a4dLc2VjjAXnHPKTtZ3lYHJsj+xKXP3ZYHpKZ2vps992X9dQuHEN
5HM/hVZxEPSEKnfoWFev+XyPd9SxbtjhNNPv7D+NAvy2JFk8fziiZDDFZ6jkfRiPAvTJUc5B+GjG
7QgPCYsBmxah51DJhf/XJSOQejGbmmBc7OStNAHIETS36g7cuUsUhunXMWdCobo8R+bIJiOpllLH
/9UpQ4xMp5Ze1A8mIxWY47MCTQfxW48Ps9dJi3J/XWBNCvsBCu8/YmXHwKciIKC0Zr6yX4hUfJva
L43L8ojhYg6Yq+xxHCPl/0E9f30F39RiKGZxCKG+cVW1DQpDRYr0EQNYC9M+2+6/8eFRD9Kgl4id
SqTAndMSkLG0CDQh+DiFeM9UIoBhW3suIUvmnAMo8+9RJOlbW3pOX9uXJnTDeG8R0y32AtZgBLI6
Bbfwh92TEcj4+dcqhIBBVGlpYBXGPHdqI2TLnvwJYdLXTYEbP44ddBN84S7gZ0svth773sobR9A7
zGOeveSB1LZrrmLaR2YtxvYuLn2S7dvE9cLKGpinMQi35YFRo7h5yzCqsMpQWyUp2j9PrRSOjU1x
ESgDRU59EfDMtM4wiDaZoDru5pPjS7w4hCEzF728M/QfEnIcpqcRdXRpPn5DPkl0iuqi1r6s3Pfy
2QuKwlCd1A28n32NUUG/kZaZkuRXSJQOTdthUQMmR/Hf2pnHkgmNsDt+dsJPDxkGORtnHwmLtzuD
Z6ePVVVUe7ek2SWclmWyJ9l2qkg/S1MNcv1e49IJxJBuBE53/3kijuEDXIhcCrFtd/vhqMq6n+mp
SywwnTRGhY8zrbtR9e6FqhtOIzWdnBUCPBbSLLqS3yNRk+T0qKC0HHjEjWkdCoyIE0zKQm1lIiua
TmvKNabpgOiG4YQOPYBK/xyjwvBFE0wqhawmLsk1eXL8GxqHQDncJaytYdOMP0st5jkBPwpnSpEK
2ayZtbDsfHremrYeT11xfp68DwT9ceLg0ShGAoWCkQpzKCsJEJfehFHQHLnFziBPf1ygwyGaUDTa
ALLGjnir1H+RSBuphtS/BgcUD/HAFWCi4mSeRz4rN3bnXPhyd2Teom8qtAez1+eiOW6IOifM0lFX
Msi32Y2CC5GSrDnSgv3bS9L7qZbVMhUNvjJF5fVOEktscFJ8U5UIy7IyD5A55j7eAEcMingVrl5P
NtCGD1ZiSEtk09QdZZV5FZ84u9bO9K2IsSGjKZAEmn87BcZrxTQpmaBR3OEXMqFrN+RfPsMTkBQt
7TBccUZZP6RHnzs+geYJhFbsjcJAElhLUPkTxUfJmkXDVnhwG06nZV/1ak4uH5nrpuJA2j7Vu6ek
t0Dx2djEGmbbsXKdRj3lp6z3K+/6e4M7+yWRPDdaGxGlmicIpytKEcF155g5SOj32FGZMjEP3+aZ
0lC28y/O4k0v/O+WSDi5+bGfqLWqJ8CK3VO8p8eVIdiDGZ6cn96JTrZdCKwWC0zw7LxVme5kuB+x
o+DxeHGkBGaGa1NYO7dsnzOxNfgnsXEZwwFVAyO3wQo0gltbpKaEePEExpIdsmg1Pwi/O4QjTCEL
944Rpb8ElBUtHFuWoN3d87BeGJza+/n2/Fty80xEuoh2K1+VEEETKrtcUPxtiR+PyXyjGHk3O6pp
/ytcex+Rp52ya1Xtxd6mYvy5Ka5JSxEynCPg07mP02P+Ou2uwfa277cG3MI5BukN3wYIndSxfM7B
FFovrygbXKyl4DAEozGoSro79qYssYx24JXMaC1yJASQMxm+lvKSsCY1KdkVq12pyQ73wz3pCxAn
J1m1H9UXbkJhTavlO9RNe/9klb9P7QGwOmc+xWCUaggXXd74krpx+3muR/5Bo9C0cI0MIZjjFdIF
WlgFyolSWYBd+UnC5HAvTdm3T9hzTORUCHBJG1E1j6TJIhBu9Vc7NAFzgLu6UfApXik2G8VGuTwG
SC26+FWJFpud0MZT0xJKFyj7gQcHrQ0AyjK8FjjUei3emgOTOQnRTvcvZKu5pEbCGbkJ28PiOo8G
Jxy7X4/va1rSOX9YrsQ4LEqc0J9hxOccsXo7n07mYs8XZCjz98BiR69wgQHE7Zvx28MjSNkTXYFM
eNCWQIZt/irANA+m78N08lhpv8YgQhmPdIQw/ZDwvpHVso4o/DNTmMlaEDYcpdgzUcB8B/tIIJDF
H3bwCuNA8IpzbFdZqXKWs6gP18WW4AhLCAiVriVyhPsh9kiwRB1tbYtipX4syL2/vGAM/IttzzKz
knwbdNEY0vxVr4Db48tHxUZNaTfyc0wWBr+Mxw9Qoh5oPp9zJ/j2c9Yc4koHCZvY59SCX+1qb1nY
/y4TMiczxYxBKqFQF5V+NOq39ZBB5/+mXqlBEH/g+OFudMAk7taahxPXhy6ZX+cmTj+fgaeLj3SV
kfW3H0IQOKiLSAKO9GnbsT3cB/XD/aUlJdJQRXumk2cRA4zAJTwLiOZPQ/y+5cTY3+KI0ET5ETpo
AnzctxqXtJ+rlK0YDzO6O6n0Ceyk9uiltq5IbV/AaujiS1KDyapvO5DNcbZP8kkSUvbT/OMa0vmQ
DVRMKpYv4BuoTtmeaIYmZjQ7E7yHmX5Iw/ZlSU+5aLGTWb+c0SRi+kttyiMY7U2dtkzCobFoMAsB
hR7Fh0+L29E6rmbdEPXFeyA9+nYsOqvOt3zDKhkmZNcDQRUKrinA/YebpBxpb28/CGth4mSkWWXi
GqKREM4j/oyJ5mCd0vJ/pA0oQM1v1vZFPs+LD3DY3appUeVTKQe6TjuobN2kzjQNyHSTPOSbUHK4
4NT1gg2Xwr1LPijokzdxSIKtVB2QQ3vbqrZOaJFcEq2NAXbPfr1baifC1Js6aoKKPvDPZncQvfRu
NjbUjQDuPWINxz3DFqrmVHeaVOmXNwCFfoljYMnNIAVUFvwvaydHGLLoIfElIGYhaKzT35FtO/vJ
rI6t3iFM0CZKWPRCuTOrz/DtnFc4A+AeBVk2n/0TzL1LFql6WUNOwg8EgMHNk6WdsBzUZ90q/iBv
txO+7rtaEC7m8OLR9N2hjXPSXddy+9nAfij+OaTKrHkoENRctKYpE9mHhWQjeULq2VP+qAl7FRj8
oGcap4rDhbbCBoFSMSUjV8gIEEfIDIb9wLVwXUrXj44CtlkuR+MTJzVPseGNNeaQEtaLbYTzBPr0
lSjkVpTthBMrsG0AnH6NMDbNZRK26ic1ItGucaS5wU2IWcHDPBoMwj03yRrYBLL8cODKhZe94jIh
3j4ChyfqwXowvA/rJHyE8c6d4R/9b/wFdFnGtQZF4TqFwbzsiR29BVyjc7wUkCouRu2Ds2nc5HmU
ZfOJKvWJJtegANGBd7gu9x3oUmwqDOKQE9wJhi5Ii6dzu/dZx+o4zq2phWhim4XiSRK/QiSzdcRP
1JmTLcJ4IMoUGL7u6ZW9VRC1Z0dqGT01QDg5omOtWO86qXaEjEbbpd+ygBfqbNNP7XFntWRjInKW
SEyoxdD0EiFeeS34+uqpv6NFuI6jXucPb31bpEpSy+qOO07EAJ+sGeng4DIMopfjXUFhK1kziIZx
Q3Pf5zfi5bOzHGzgz341jQ2X9B9ZAt0xPIQEethRxlf7g4RQ6MF6mYvPtaxl3W2b1j4NYS8q0Epl
veormWTALqUfK23mS59P4vNJr8CsSkKFJD22tBIFQ5Ost8qRpkFDFykW2icvCTZukLKXyOrD+pmE
9A7ohlBsmsj9hQrRgjUxCRhWBHo1FpBPaKp/uDFMiKe4YIaWVIde+FIarybNLDFzj+AKrDNcBTGb
cDaR0Ek1iszmAqE/79VeCw2F1Aqx4vYPQMhL5zxm8YmtJdmxEm1ysOvBx6Yu6XWtBLtoNZ+D5qpx
tKgv2ipbSMgH1FkkPUsV36/B48EdB6Y/sTT494z/I4XlPMYlESulOqe7NigfegHhLl0b0pmYwXd4
VIL8RR+X2vCfD+nWHSt6PFjKb5OCWDY/VLnBK3Uq0/aAUaX7MSLBXeTfSdKR+3Mc/5PFoGlzr7iG
ChAJ8Wz7FOUmfec043Rv8baTI/+aly6ytH7tAjaIwKsbbUVyynbM+a3jb6NM8RBeLx+38ESGS5wA
nv4DiX8FPw7cDBlcmxRX0NqqDnEf5mapeSj0VreXU7t1Rn3hyUPeeYcaqa23iPwifYtJUVZ1038X
25KDFDtBScfBqYEweE6qBoJtU2PMLbRa9TPIlQactvm3E0f0PgwAAwjgZV6Ly2bIjj9Vbe6WrAug
B/RL9aK/BonStNQmy1/xZETByu5oN/hVBfu9YhywwBTKKQl0PKaWYQhvHU0qg1D5oJ06qE/NgYdz
iLeQeLLER1QvFq6Ge0YMiTpPJsOsDeIAQsLdhKn8ot3Xve4Ao4XSb4d7W+NDWsTAlMAOdgwpkbsM
0/HlV/yQjwrwe+uQ8a6cG+Nti0Q4CaES7pdwJ+lgenKw6YbetQfVBX0FZ9Bl/9QJPWM/oQtqDwh5
MyMgp00cTt6mx4Q5fDy9cNW26r95J/oeO+pceQr5Fr2FnJso9Q2MR5zGVn3mjAScS7CR0gdaRMBh
e0Hzhk97iG7XyC3awBARdladGEkd4dEEbIOHLqZq0Ahn9FRu1PPYBkDGge84jUkg7ulxyMd2ozfO
P81orxevRUspKQ0QdiLT0RWhdICqSuRqNpZ4hI6LZv27xJJp/f2K1Bt5RkcxWwHGgEunz2sEL4e2
2oBIiJyT/+s7EMYRkXURP4rnqI5fukA+ujLnYusyhpCBgx/ia4umh9G44RV+hSEtkAFT6xW1DuGO
DWbPCPeiXqdKMvquO7aLfLQR/pUBwFDUPKJbSrDN45eYFl+Hy+dXe6kZ6pCWlnIU/8ibizldvU3v
GHi8JZEoulNrEGUDtEx/83djxv3+lmnhfva6t1p66h87BOgpKbNO7lXSgIci0g4evCtj3WN4/Z43
ezc5j7v+EQZn9iFfA169ck4Hqm3ojkOCTUXj4My1Hj7piG8Mf8WGjoJUz7T2UbrdWU6eM+/e8Bfs
PFuMTss8B/SuOA1YgfcfjOLokp2boGXfIjRoParTQAxWtnYKXJm7CbkVpWwjHy2PgV32ii6yjNB8
r3fsFwokK4J/GaXaTKu4zbLkghWOB+/IRBtzXeMt2OJz8ocENbNk+fNycpKL7/mjwqYFuFrhbw01
GRmMD0gWX2lSR7OOHilT7d7PWrXWylhSMR7LtytX3YCKb71UNtWfPtpLysjdnoyT8k1xhXypKgWa
gDDsnEZrly5zBYJIRT889IH+Qwg/c8DOFiY9JdDpd1JW3vp5muKHX2aaOpkoN/Qn4DCFfljXEgL5
e/JN3+EA8UZ5oYvccElP4Dh/y52tToKyCD6bGMVSDdr9yDX91zzRVhZug7OcXwxqqNWuIewjlELh
J4y8PfCUTtW/U0+aZXA3/BRBGyNvE70VhSbfP8VACW7a013aMhbPSjOLEW8czIy3KXFQRUrk189o
JH6r+Rkczmgm4jLp5pexKctVN1Sa+7w+rzTje1AO2E0LYAq/f5Mz7FKbks1Shx6ZpXs7FUThHEwt
5QN/iFT46RC2LOmv5hlFZORD4MK8sBy9GNw21r7vJZ4SPwO+2GT/tXLQfsXhICiZMlAoVZdqChOj
JsztidTLMsUht0JG6qR0k69Z80EZn3nx5htFHUb0votYn1LSp+FCGXMrMNEiw1MglDGTzsaF22c5
zwwrmXL5Oo15OKJcXwoof5731ECT8x49HJNq8mvxZmk8Y387N3qBXGc5O42KAwoME76uNPsPeYYw
Z+Np+W6MgsnKrdSUocLplmsc5/l/sS+Xz9jAu0LM8irLMPN9wvyRh9a96X5SqwHUshLgnYzdjGn3
OWTwrj/1iSUrYSWf+1Z9kvSxSUJk1UblwVvujlwJP97fD8IrvuLo4Oa6ZnqQJO46k5+WZI99icLL
gf79UsIyLqG5JRr+gUSl+LnGcfTGMt3KB01N0dwgOWuy71pd3ofi14h/hMd419VCb6hbePU3Pts3
qquhQteoCsgUMnU81O0Yhnq5Fv3+3DYn8E7KQrXMV0uB8BGQP4BH0HqQdF8V/BwS/uIYN04wnEG5
OIr9dGtEoXpoZm6MVbWbwrcrO7krq4ZWbPqVG6K5mL3DG4bpv4LwSyEn+vyzG+rwde5MGuqiDpXD
IlsdEA6Qj1YUt1XDy1K679UN/7ibX3RbRyvcVzefZDrySdWNcCr0j1zgchBUGF1UZv/HCeKB0xHe
7YGMMOfSu5lZbP8NsDqf6xTOgqjaTvkgoOFjhS0n50XNycv8oy3uPgP1QGvilz1+jrsK0r7n/ZJn
OPKMpnTQrTie+WoSWHsxU7Wmr4QtfH72gVCwS01C5ub20EpwKNzYKxPStZHa2FQfCVl6NRl1KcOA
1cTdGfvaMfel6yoSkZEeHCMDxJ8c8+DCCkf8yEg5VujZG2OVcZBqScj6jDXn99AT7jfaz9p/7HMQ
DvnB7vMjQ0of5DEONr/D/1q6z5ZTy5DRJczPVGT0LvRMaGcbVx7xaOpiYqcVXAobPdNMnwco1qHY
yunSegfHdS1vc3+viqmjzsHGYtw9+UWtX61L/AwAYxJkaQ36UuOrGfllIekQeBMoAZBIxWWuyeH+
NNuR/0PRL2eGFEvTu2ksJa6ze7Q5Pg006m8o/Co4Bg+dy/9abPCqq54LpsL4de+H4YFSSqEG/TXf
Hlco9zZVavb72pWIbuh3NK8U+h8n4QJtgYbZfpmt1/ByRjVjjzIQspFpG620TQNj8GXfK2VKT4xr
UN9b1nSkKiFSsQYkLPJdycj3ST5Da8M/KmEs6ndM2ldjCzzW+muAzhNc5D47tGJpNRO5RgnuHBGt
ZIuhX2cKDSfZ7td5bAU/xRM9OUWlCrbwAVRTjL5PUOjjLJLPFaZHHcE6PokliojVChNdalGNKK7E
haXr4yjQR8C2q4kkqCjeuIFon+AF0D/GnIieImdhes0AGaa+hU4a5GMgI5SZ3LD+pg0N80lT6egk
dfNXy0XFvMqTXvclhN0Ugkz9NBuGEcLPwOl+0ujvLbQNSVZEugmvQzN3OJVLrW+bzT+vxDtid0c9
8fU1Ua52kUA3edt0ezjc6udutK7X5lKwXh4bgCwgArqQvhLQlzwDjHM9431CX/DZ/lOm/LyWbn9m
HUBfeqABV3v1nPUbx/oX5sHN5nj88n1XkxqsXUkZmm8oYC9wJ/gLQLwM0pOIlaGEbebuHKVpgYOd
l2ECk6ypXfyhXpMeQounrEbp8+0MU5DjBQo/chMnpoC2+4pQarnh0JX66BbswA2MbdTjBPeleA8x
usSikN9/vsTQORNPm7cjnLtxrVfWyLyT1vAmFfG8aKfgcrwtXgTlSmyxqBZqZfaFFrdCsgX7Qf3C
J44gdl8X7Zr6Sc4/IrkWAicBKfH7LrDDE7dOZmvtvF6bNHv1d8wNifrkJrtKoKIp+82yFIzH3oQc
UPHCuWzGlCutBJ5oBFfHApFFumbfo0hQbm6ONaAzaf8NQNZ4zUpQ6rSGToy6tC+pZcHSFZO1/PsT
J47A40mGWdHprBL4xq/BxphGENpXlCB0TIM20WAk5386v+CVp3JhomgSuL2taQUKdX6mARPqg6wB
wVc6rEb5wQfD0T5o2Me8l34OMaawFVOySAMgdyJO9CAX5pzYVVg8Knwoy/toaC/d6MPpOL9TILd9
Dtd7P4LP5xzbc77UHNP2tF/QDIOujbePd8ML02+u+V0OCUVAozjo0i0nr8X9+njAY/hnKzgdMPkD
v2ZsYV/jfuWSSfXKKQBmqqXIJxlbZB8neRwWzHcyl4hh7FlTx+i+sV+aQdSB9C3A+1qXBPxtC2/8
ST7JHosg7lmifDQ6YRkSeahsqS/zJpvbq5QvqOJNGOOh6oAG1Z23woABfHOCNkb9U0ANudAx7mmW
lDbc3yWfpkofOjM4Qb2KPZaBnCwOqqdGJ5jbzb8NjhBuMxtDwnjnKrT+Clr6DMRpLzSMyxwh6Qb1
C6mnGCOwWGqt66Q3OaU5WHwbbxGPfoCDNv1D5Xot1XVzHAbvPnbOiiozTYuQTZf7HJZpOUexlUut
eQqY/qdZ17SQfv9+BsWkc54Tj3OoXwpG3njxXKJBU4ytN5zYzG5mRuWSTgQVZU65feNCOGBQyfFn
KnloCRQ32dOUX5vrYG0Cs6bP2DV4CuAH/bDB/d1kT08Yg3XAZR38SWlqOXREHGljyM+/wQeRdwTO
F3fai8NOdg/q03ofq/xNEO5eFUwoRl3M6jbWEGn9462ElmJ2qmUGahkOgINrcROIF/efgn4qwPyQ
uF0VCMVhoCFE3AGXmV2jr62AjM9jI+ptnjR3WdNbwf2V0m56M5faKcAZ8NDFG6Qvi96lCS/K7UCy
UGaDOi1nRxZSZHsnm5h9RGg4xwaZRl7/FxoOkRc3BXy1EqPcDsrhKNHMV2xtqq7sx92izep4dvT8
U1ln5DKfy1sW+3hkqYLCxEiDKdAy2vTSzBOwEM4Ds+NdGzFSy2g2VjvFajj+PgPF9MIk1wvRnlX3
6u7vdsvk1s9qsd6qvXK2fOkI8wKajEg9mlLwg6ZdbrGMv3YycL3OVMGGoGkIUQlPI8WJL7whT3aA
/CRTS5nON6ekRN88YMCNjy/w5xq4/GS8t6bGmTrlN3TjqyikkzWXBtx7GxaDzMvpbuILNGDJ+9if
FA8SbnC8QtvvzZlKoN9nQqsUeHcxP2ygLP989XLMpb3625aO/uDX5i0+qE5giM9L1QVsluy/mHyt
7xjTYyvHRUNzKD7QrH3Z5bMb/dLiuXYI3B4BLB1ccOsIJ3+2dAkTTOmWNvEqrpnf7GM+csW9MvnW
xe9y+ZBsF60lHMNgCjMZWawQnB6trdfm2xvXR1I1lJj/Gbr7XV/M2jF93UMXEE6d8pR1fxUOhwW8
0zZNdqjqYvc5IEkEUhQOgOn9NfCswMBmBhk4sW3BhMbb11w2BX9OQsylRylRuzlhLbhS+jC6ymbp
0vO9Lc4EhBfmnmhiklyvbrbEQ/AeEg8z2ZpuyWlxq28sxHauy2hiMKtNV2y289v8QOt6ldF6mtRH
fa8dRMJh0RC4vqNVBybJBqeXrN+YVLtSrSTY/k1Q8VCfOPUVzJNvNXtOHkrZBVSqRRjDE9IGed4j
knFOrCzCUsjtkv6Ewz1Mys1mpgzFb4dNE9BmITvoGDfTiqzMPgHeC3svx/nEORFCSamrTi6Mj7Sv
ysVvFYsA0HzJhAlxjCoz8hcHCgA+NKtBhwRO+NPKSR4MSF557dLJDmLYqRfuDIwx/7AysyE3Spoq
KhNT0/BSdj6NgkqUstQoBSTTqM2E/0l+W1rotlzpkoziSh2iog1SEuRhyg7PQI/cD84JNtM+LzY1
oAcZEKQMLOxTWfkRhS3SdSuJjOxkxMulp1FdimAGTtORbgE4CHnPXNaz/RaLVSGcbhfkwXZLc9lo
UmZXKMJNpLRNAWzfcaDmwt3R9r4Uy4PKQgkHL4hrZBeq7K3GdbQ8AUL4AmE12kVQ6wTCtjg+y1fU
hbiPFP9nMNTgEW0s8WsaIJvfu7RC5bZEuCzgVYTmag/ik20scivClDpyi11pfgi6LunJvudP5J4S
qEkwS5E0/qRKG5NPMGi0e09RDGed9y/s3+YxnrswuSTrSL5PsRIE0M9ujOzw7T71veDBX0rEh4Ui
qzU9NHyNbR1xN+ZEVDtnhsvb9AS72l/Ina9W4U8aqkvPhjUJF5tYOk3t3CSGUsxXrvhw+AkJzBME
TvH+JFrCZf7pnPCz2v4uFMuFRoeRXpDJbKqONMlhTrXpwTqJ7goQV/JU69CgJZLO2ADzbY0p30e8
4vajSqeu8W3HZJrdQ1vEUAz5FlUJGck/w42jbKCmxDpOLRIlRAJPRwSb9IcF7A7Tr00mdFbSLAYQ
zJLhTCoucaFX+Nw9qcoHlv7ZKl/GUr0QgX8Eq7zrf2weMOXgHEcyBeE6tWnDrKyXImY/EugrV0aA
YxkRJRI0UOIqTfosSdiH7itYjEakkcXSSZ1pfln4ALhiQFj1rb7+0MXc6ql+VhTskixuKEGV79y5
LgeinBvDgY8YfdGwDyTjdVVga9QRScfCkrIsSpHxpuI93zeUZHPqh6HBSeplYQHN94FyQ7KeivJo
yY1w3274L2mjbZSBAAj9fpF+ns5gET1DcKWs3axiMcIeRMie5IPQZdHnafa+Y5SdzWIUbmifDdcq
O1k6zLceVba1k6IHl/AOBrXFdOWSv2v5G5yKLjkKyxmZj4gLWc/ZrqZXBnHNPELF6L+BD3zWsZSH
x432kz6foKhHiHg0wpNabWb8L7xYBVG49jGaWFbbQrnZRnWD4JMCB4U0GsxcY/cKqhAO7NUYjXBd
yfpbG/rAc0EEeWnRbVOG55C8SoEpOf+VCFTeYDHoxGHdnI8+SUisabOlMo5aYY3ECZ8LA2RbFcWQ
9qoRnDqSkCUX5NFjTE+vlUJZDKtnA/g2cAqDIVj4Ew6D60R/r89nqH1MYJqd+aKzEeV1XNGolCPX
6ihYGcp9VZhV9QqjKHiM2MiaoNZZYK+gsbgp6lCRP9oyXTWcx0oGGQm3s4Dr7c1OOnCKlK54PyCz
D6F0fNlnjIW67tRNw39cmynpVIkigqcEvWDLMwt7uznVH1hnwvJzrcf7oiIe3QSFKklL1QRiGOvM
uokkXtUZxN5Ul9l3gQHg+mSBfkSlZFctVV0ELuAAzVX9PoJqvlQ0A56ca7GQrEjmebZzrP7CgEKI
dzX8crQXIrjSbUGjLMRoiOVFgd6ET9qVrRe2niXpxLN7Vi2AkGutCPhEl2hjOJMx5MeJdLaf1FrE
Hwu+NPgsFQIuADMTWa+7H3lxQziPPEwfBeA03lCerGDASD9Pe3Ljm/AzKiGSQ85TrHyiTJKxbQdF
NR5+N4B0ISQj8tyqAUJl3rXzBVnjRXoWH7exqiT+vwnpKlOVvRC8W4RrQV0ivLVYmut6OpwaSBz3
OIciPKRXwolqRe7V4DXjUSvNy9ZWv8NJwRzr6SUp8LNfoQs5EUoSnX4VShlLVcNVhk/AITSoU7U3
JLdP7pgNDw7UJK0V+vMxfkHwBeLllcq7B8isN0S3DHDxNYFFH+czMYpakRKfrXcypjrRmVSdsf3Y
wGmKQJNnMRzlxa/phU9rCE/Tz3A2JNMj7V1Yup4tNwPkEBg9xBaNCq5l8D6fC47Bns9xUp5VDkJg
gNh++9nBo2FPBZP25QUIJgqqkXkuuvM7EuTp0lc+HwXgs8rEpov7jfwlKlc/OT6GUUqqAC4o3SKX
fVhR/GFof5yG9Q+8dYgZ64MOd5yPaAbE8GfWxnRNK73ZxhiHJgQxTiuzJUeICF0fOE9ec7dew/KL
7j+TurylWO1yHnyIxUWNp6vtTaDZ/8sJ6XlRC9Ds0D1O13/fh6UYpoxdkC/rC+fcKinRo98YotID
Ghy57nifjY/FSuPpdk3ROYtNgCC3iwvWoyzqVze+0hR+8xcX8xHhoPtIiZXV824AOg+vUxOy8jm2
qAkERtLyA0x/IRVrFM+9lSCE7c0u5qVDNSMnj7UyMaBYqeUW8rlgYSNe7Zpg3D4W4/3PwGVkMQ2I
1Hr19zLfeTyVfDWgftx/8BJj8Iug7B9g1QA4jVjpr4BfaQFdqI0Z/eiSOqNVOTDcsooRa+GvwZse
koiVX054s/0Wx6xjkahIET4t23YHw4MnXQrGzCtBdBF+ndJA24EnSs6HntFl6VDh8k534/I7o0bt
f/kFNEtHBvd3gtekDGeee2YMT/guBLpnB07bOTDNMS+9feAL1Tx2FG9naF3gStMcC5J4oP0t53FM
m/R9oXeHzGNQARBZz0AyqUQyWpEbkFPRI/Ft3S24i4TamrgZ7lCnjHEPSKb50RKIDHB97dDRZu9D
8IE4Sd7JesPcJTlxWGXjygiWPqZAozC7WMN15xSuobxj9L1jIujNECe3SdVK1ugr78BG0M8DBb6L
cE3feSiRTEi5/6MLJkt0GzKPdUaaYRFy58ghlDURLUjQtTxjyA+qWO0xyMWfNfQ6/bsAwFIipdYS
OAR8hX82DlAyavvEUblMLWVtd/0YbAzuKT/v+E7xcwwvsK/ikUnXpCh6BUU1UiiBNa2fNTz2KLoe
fFKgDm7ijqf50HjF2IleoWD5MTRaYGmgl50D97U75V+BQuPavwwe239pPopDa5gsyAmSCvg7Z3nZ
BYKKuQm8RhtotGyJSVFs98DnOYV6EyIfCQl4v1D0hsTiJazgYeWqpQGrgZP1rolfQsCo6x16IlpC
ChCUpt4eJcZtIKc+yZ9mRLYItwXSddln5Z01/OSUP12GeUQU51NuiBclYyViRS3xqwqRChih5UzD
DjL6jw1h3SkjaXZQdHQT1b+J09yrcuiRyN1uGFJ/xNrCZmG9ku2kYHZBbppVyxGD5P4sdnCbWkO8
wXRSrBh1/EYnPNi+SiXfWkh2BZaOKPmXsl1VQxJ1KFsHoBQzCKEv4JAgutlArxi6VVXCwXKqPEhg
16TQmoo1v8u5pb1yvjmPKv/owhdCATMLY9sNbxkBA0s7SAdKPL7CRl7Lm7HrEczfT/0TXlQr/WuI
M02kzNJmQBCe/86IZNqxPHzVZTgheqe8KBo+5NJyBzUp4ezMGQ7m4DjA+0pSoG5yadYWkNn7oM0L
jIlYaL3KMGfQ8lSrZI1dPXUXnvC6+zkm+CHAzMeeN+1I75EkXIBreEfM9gTCr/1DByF1O6E4s3Es
yzVAMlhJSaYn6gqoFoXzn5pAXnPzH1iQQRtXGhd4Y+mOCZXFchJWcPlQdqT1dx1mbblfbOEUIjG8
O10qrRSm3qFDBn+p3sz4Nm5NPcLGsQKrFyKz40ch23SmcGaWjQaWc62S4y6axwKDCtx4TFcOTl2+
PgUFPc+Y4zDqkZo0cfOpOSiLWiicfQIgHqgh1j2OglH6/1lh7E60niIikmYOwVQg2TpgEwwTb/U8
rhf9luQyBafFF8cN0KQU8N2AgBHcztlNKP5sVoOAuxRzHp7p1KAKXU8Wmb1GdxNQ2qlthIF+OCIe
2ce5nWpE06K3Q1DdEqhx35C17arjEFi+8JLG5xIVYyOmomYDV8bImx7OBqvTTfU+Ar/PzMkMqiEr
KL58qIRhE7O4rPa32Ns9o4kDAWQaJSClLPRmILBLZKP35GGCSrtYzc5CHqHfEGxhQTzdgSWqmqh6
sL7oI3zmZZ7WD+xShPezEWreq2mkebw2g+uvxcj3IYYOA93H72XKLn7iAf+hMD1J3gNI7vrFqlzF
pzMrNTkmC4FvFV6fDyBGbPh9Myb5o4OXVi4GCktgohfJg9kzf4Vo7NJQ7ZvFL5paZF32TWoQFXfd
robWwNcQaLEBmj2PRYkWEsBOkwniWHGyH70FMmGXOZtj05LFgNdcqDWR1SH7xj5/vXAdBIkj9Qm/
aPuddXMjIv3ZhE0CznE5IFNuAmR6c055VN4Uq5ySdqBcAuIiqLX4qDa2LbvmeAQDyLxfdhJrkE0g
n8RCOOI3prA3haEXmW91D35T7L9kSvYlD/tfJQJxlhqhyZKfxOM9rjYFSvXz1URKb1WUzldfaH45
kP1/EuCXEE4nrSR2tUhKUB1IiVJR8WSKbC9U45YsrhIBgQ4SPL3mJcMRf8sex+DnrizALCFsQmPR
YqvTShJdKv3TGgL/MNwBE+l3vdUyLjJUP56/g1nRApdmVgCaUUPlmYD/D0pJqHtXYk1MYwdKJSus
NdgFsB4aK6T1R6Gfkjk/Iy05yJ/flO9Z8/XRJleSA6Zgo8kMxjz1hRR7N/VkHSRH0pTQNyIeKgET
rxNmq4OIg7gzt7mTsXDzTg5T2qa8ZkiZnq37RPIX1USZJLa6IM1InmWu0n08SmRI+beJQB+GE1C1
YZWIxwCLnymC1inV6fzdZkAS2Wj5RxOEiGs1CCIT/IeJJ1zp7pdJQ8f/6n9FbNCUij2kHgKvpCMj
+A0r4D07vm/5oRn2WWdvMo7zHJrf1+qzh1L0MV/M95MxxCh6Xkk+ehA/OaGVo5O8IP1lFNRMshSC
ZsHAfyL5qRpmXLypBiMKtZVCQQBSlfVrrr5u0EEY5x5bBJ6cd2N7CnLjARFOvLkyY4mOePwEnbbK
ZQijdhDuxBtQbC9JOx9JL6AoPmD9vAJv+XTTmF1auSPA+jEnCeNg2nHzQtV6yaNPDWv342O0oxcN
93pqmhVCz19UIvq12qM2lzaTC71H2lZ3W3rOKiLUuZbgczocF3pM1CN9t0jY4XLDyW/UnU5rwt3S
lE8D0z8QCTexx4D8uWmq7VvtzM7dZbPaf1FbbsQ3l9UWAB2VgKbu9dRC9JVAFllK1FPIIYtPWgbt
qb5Bol7YSkkT5ZbGnZSJRoFxSuAbhk+xHuHTdS7JIRw8DbY/HCCFp1ORIRwlC/krs1cakmwY+QL2
MoazuRyICfYAO6nEKM/hDSMnRXD4FfwG+4VnRYZ8jWnnFVPVjB07XQQTyupjPXgrqHXCKxVfAU+9
EzxV93k444wKweGVRRhleWu16S5otzoRORoZYWfKEVgWVAt6+zSdW+R9GDK4GhRh1CL4Fo6Nyw6A
HhqNgIx3bjPkwHfI4Bp+lpFYrE3edhtOqBMWkuAabjMCjPCDXP/ZsTKh62thitVryZw2r8foHgfb
7do5ChnhkjdY8q3pvlc2aehTNqJIOEjz/KffQK/cKMxHMqgsE4xkoS/7njdusShOOefNXgEGKIg3
fX44Y/cfI2bIC5tvh/pQpH5n59ee4YcCbGzMSYpN/TTi7FQGylGVtKctjPhdrz+/4ToGwLTNpLYf
Rxfc0f75isGR71UukaCD2U6OhAgmnSLvy1AlaguMkOAK0gp7+C+X1D1gWeCUXAve9YmGwzQIM9Js
YyHnCO+rTPwD638jzV8T9xNtJwSH7ZM3n5C9XjpIMdvE2Mgof0W5h7FRuK28xgJCDpBVltIquZ+Y
QuvgRmlUV2CBgNg1Rna745spmI0f5CtOlV44zZoC01dUxBM6y0GUacGQAPGeukx5Eo0AKj47YlFt
pZHhwwtJd2E1M5iHzgUkSX91I7ozeLRsMoZP5ieYfHnAVi8KzwBcX7pPFuyhL9We60HvaASHfqB+
zVfsFYXpTKZFlUVmPOCKMUxeIQAooJPoQhJgz+qGkcCIoaI5DmODB8DuK0r/eTqEg24BiWt2tg3w
TUcmymGuiDd1CT0HIXcl+B0hywEOxMJgvbJAAgt8z1j7vlcT7Mt/VqlaNvHOdGMWXUog07ug6X4P
W126JQGrhpKD9yUhZTwstkr4R1nfv3koFn9AOoHs9V2/Vpdamb6VwBhCb7iys7XD4KAsXB8HWaDb
DNIjna4bO+dn929wPfanuLzQtvu1G0jxQFGKU7KhlpWLuyruDVBoq17VCytL2o2QcCk0IP8a0xdO
CfcXCkRMEhWFAL4Jcekim7qQZtAL8UHvKdUGJgijsJ4Ro18SW+sMGi0QQ41ovLK1CFtoGiFdmXSm
zWh+yhIrSFsQEhHO115zSCy2lVaPOHrJWx7wz6M0BDMAM7C/UKxOH5hZODrdrTgXHkruaUcVYZsP
SFNeOrdglSSLLktdKknOVbD1foPmhelQ2B1b3tf60sVPTgivi56lac1vE6dMZBwIaGleaIkF7J0y
iFQClJl3eqkDU9UNRLodjapMcULrNRxYrJdGlvY7HkhM6ZImmxA6yHyqH7XgFbs1iU4vJ9N1dYox
7YPcvSROtXNRVjLwNULbE7OSkScynf6mpkYwTjRdGQDIq8yUZ85ObDXmLdlQWNs1SevXYdLqbiVl
rUGoaZqESpauqCMYk+8xqh3Zcc7pY0/P3yR3G+TWMVNN2kNq7uHFdFmdm/G+DeepA/3Ctkwk0vBH
V12o7AseMD4UfN/TosI3Sl1TdPhywiIZoNH2wl13qD+ALvRPyKIrH7YboMBO/XsyTQcTQAWaIMO0
NTstkCuWAIcz4z4AwE6XgWVw5u+fHKS1mVEigIo1tGaxDCnLhER8UQ9YEQqYpH9sxAJrizOBbtGx
5Wv2atbU+4ySLF5E7Wq1y4xQbc7LDsuTGFApzk/NqsUJQGb+A/SS+BVisfSZwct/fj6O/qIKx0in
NYZdjwChsDw3JDE4UEYGfEvt4QpDKXKxdb490u2QerVaXrV3F6CxZW9vNopHF5wV/Qp1C7QhlmrX
7LOLaax0ywamPkFXuqiCeM+dihebJ7JQVuD1vjO10w8GeYGfxaUOuYXuQgUPdIdV/OzrXFIGE0/F
mGYIcowpuXBN/V66TX9CAIjW1PWi460wGMUZoVSqZu14L830AGkES32Ito/uqOtrWkleRebWoBJV
jjRdk6nWEH2OTzVgF1LUXHclZnWCwTiRZSacqvhsskj0zCHwqg2br4wV3VAjdOqaQx4Qd4w8e8PT
prv745fnKl4dfRKLC9Jlpl/0yY0p4FGsiQOeToJSe3y5BtOZ2AmzxeT9A5M0SSX1RXzFIcLhYx8r
Cbk1iqYAEmo0wHO8Rpw5CPNj4dHjagwrQmc9xxak6wDY/UXiXGv7pM3UzvEDGErBpn1Zs5Do1aLF
FKjq35Ioes0arlh0l0kSff+LWPBsU20cyNGWQNJaAnGyZ7qgIP94M+TYCKPy6Pch/83Uw3kQQ7eO
JDrP2AjwWrlHKF3vUtlIIQF/3LNTQLu9yogFyXa6DErzr95vk8xcMOwzx71KHg12GqsdR9acZqCI
0zZbeu4/blh8bJDsX4ufL10vneEZRT+kktTpdQPye4LiakvMbSOIg78c2o1NzvFVaFmLL+5erpOt
KIXm7KF8soqfeK1p1H3N1zgbdwlEOrtd63c68VfqVQVMG4T8MeFR8JOleCYelueDbSphLaWt54YM
vkjCyvha15C0Pf7UW3KerSbYHuLfiqFdTiM2khmVcIE04ucx2WNj5yoizIMTQ/WxUqX7dSRlTXMt
CEt4NKxDNmC19ViJmPzLgUmZdNjPyk8eluJ65HE3JDP9xJW16uiOW90rE4jF+L6etvGdQKygG+RE
ySKVnJMY93gQ5S99Glv8GUWOudONjl+b70xe5rRCWgggChZvn2iMJ387gTwIjJS3c+4j8JV4A/Mf
+xa4Nis1EQLOzcNVI8ZxDKOU6I8e3y/X5hWBKbOauab58W3n582O0JFLQtszlBLS6srUNqq9xuhv
PnbpfiwR2pipvcSTliEGxweTuZxV8/1Ip02cwXIxPeQDq6PnRVHdKKSj52pOTHDJCC6BEvcrnNil
lHIF1bx5NNbYvXBNMBBMU25e+iUhRhTWEI7RVkR92T5AI9m4HgtCW1IZQiyE3PpuGInWB5KV9gED
qAmz377AoGeQFWOTFF9N6RXawwL8V0VrPwetC4r83dIv41movkiXRB5TRyT0bhJMQ6g733pw7+BU
B0Y0iC9xN50Shm2TA4Z/rOxH/OtWi7oEDCyMp2DSHHz6SPDorgWGf8Wp7SKqcECWr1vhv2pBOTtm
LZdFmPaoOd0jpP/SWj3wFHaKtRJVUppwRrgUTwHJcYfXWLArYcGcqdDx9RG1UHvkKkKRXZhYfL7z
VWeGGgKtThTM0su9dUUurUoXzmXtfKFUshT6SJU8Y07iEFYptHqXBi/aQ7qAgrmBF+PLQB3Hl6qf
c13snbqT3YE1NUlcZwHW0tN+LYP49xynUv0cMC/LaYZ0SIo8W/Ro94/FEK6pssqgLiGcfIhSdkGG
Gt0Z8JSgbCCfPWHRm8PMTbRdB6EvDQ8BVicPcxN/Iyw2bi8j8LTDMfXLsCIR71WuaVyyoIzdl5v2
PWWtak7i7iuygADjizbtOBrtZC1kLblqDbXOGsP+ub1jjRI4OqgIvSxsY0iO6X+rsHlLTgqwSiEY
t4sJnCLPuNTNuMK05IG3vKmTrT+4msxef0jTVvVeJ9yjPBslCcSvNQQs8KLdjvGDJk24eA6+LGvT
9rqQSG6PsdU8/+Ei2shlbGcxlG4Qk7x+NODb8bmF5zEZVmtXyWd05X3wEvi0V6dRaGFl0R1lLpeg
Q38RmaRS6HfBY1TsD0YRAjpR/Q2HGTbBaSg4Ztw33ty7SGO0ZKDerePTHJ3MpZ6HSo3TpjwbC5oB
46J2/c36E8DHU4JMSGKdLkelmVZwODHz0S0lupjPIl7nWrKYdRiKPnFb2cQ3TIewk5kQUBa9U64a
V/U6pzEf69/1p4/KvLWAylbaRXjdV/grq+NTL6EMvvkuqz9qoaex0CzobUhdn3FRZfxmMqgH3ECd
DDPdfZFf0b8Y1WTFNkPCQV/W1jg/1NG278gTjwf/8jC+5aAE5ZsgRJlmIhI81TPvmdbiDGM7byH4
GxwVh/67n0qWBHe77dc1X83y7V65i2qASPt5vXfIDbvITK3WvJ4bl2TyooAjOqxx+CrvQWFEkTph
2rBHx5v3Nq0jKYA6JguYuT40kmkfkck1BDRsihIsrg7q5lcc078Fk/fW6odLbtdHIoi0mtBqvMHi
lfVrKO7LSadi/cSvPe7e6i5usUwQChU5VSXr73k2UIIDKK/gPu6Egq472ItTux4jgrLYM9EPJAnB
NgSulOiEFSYXklgRKIZ7vU1h2Hge2YXp5UDEgpfyEb5IMHQ6xVXpSB/RaNdjkthZMFK+wERgiuXI
eGjfzu+fzmIBxmEC/BXc6ehuygzCo3yKQSCmvs2JiKz+RDx8twGrS5FHLcKkrI7vxNjiX5CY9agq
4bWSLVUgUXtQBIcmqyh70ZyED0tLiHPurdOlkVaY2qYjjoQ8cuS1OEFF/vK0Cv0BXldscJrFfdUu
+pAMw1Y9N2MA1arzkbQwuns5tJDS1R0y9VMdSg//I96uiy2hKGDKcozEpRjh2T6R2dZt5g3HdYwH
/wGgUU3/rwjmvkzlPM563aAL49UcrCVk60jO3fnDdp3AWPyCdIbtrCqOLryfMR7hfNjAuA+PI/Zt
SdFkknD7gifGvnFCouE0k4EsKFau4dQcze5MdXocWya4684chn3KW8CtrT4qSnlJuMliPmc9IN32
0bLO77Ho7dmRmmuTuyfzZJAw6PCeROpj7WKy63uVQxfvbaBAdGXYpzXzgVZwHZpKqc6uuNGjo25r
QsKm+GzBk8Ji4JrKGO6/JS0CEhalQf0kbdGP3sOX5HH7gp/vPpxb4zvY2rIEDjC8gbU710oR0PNu
x0uER2NcjOrGMdpLNSCBHTpmNngWnGUmRlB5H/9jPrfYiY2V2Oi2aMo7nG8njMzYvFN/RtJb+p5B
g0UrJpzk6zkq5bchZHy+yYLY5nzqrvSeVNa+h8Jz3dC3dHmhoDzn4VJtIZHiMB98bTEmYQKInDrU
1GHq4U8ptsl6yDYGs/R1jBuFkSb5toFqOy5R77zBDJPID1Ba/poq4uqbpo6qAlqteduMKIi+GtEa
nnqwiB/peci6Z2Px0gXf1iNEjKRymviepCgUrki/bvycebFFEiWW5XlAwzaYNm4k474fQYXnd65B
DMKOw/nm0jMlQN76WvCpa6N4RUR8htlq2wL/0Wdg1AW5kBoeSBXAKpDavk9bsQl4BaZGXhPk9m86
s+yb2bdsvsmK3Bsfwf2wbvOUfa+MLcGihtliPRGI55JOaTY9Xv3JDtPhePNp0uV1KKTUyfHqwmkS
qJNgMCC/QDo/AdumVsxiqAJ+lwg4qnjtmWWl5C9m4wP5KkXHc1x/2MQCkAdAv3MfKkE+asJh9+TM
QHd+FStMUlc5P3cG7MM7GAmUx/ooaUnTDEoJ64juyA1Tmcf9NVZPmYbbol9yN+aGs4jZXb6rtQpc
3hEbQVqHR3HmXb7+Gta3t2KcD8zJtAi3odsB2HA28KU3hjoLf/dCbXbZZy2HFW8XMSnuveJ9Yo7p
4MhvcKLedOSNs+07U4KufrJKPI4KSDNPwGrTVMTiYh4JMtAqnEEz1n0a1fDPqzJz3u/uHEdF9r/c
4PmX5vbuXCgVqSyR9kNR1QbIMDmkRk0OlJrHSBNUiEiffOX7KeDYRXwjAz3jyp8xU7aIEQ5Li+fG
L9s94rdihRRzVT983XcgKa1XVujrSA2VHOocrnJNu4eol4d3YWhOZl21M0Yg0kCMAJJLTKoXFoVO
Vv03qFbbEg4GJu5zllcINwhgXIg16NTXlTSNeJaQ4v2mOUqdpBnNGqEHpvY6VXowdLHmnpGrPx9D
tiM2NlIWuN9jPWBAB8SLFEAxCWKBBqb7VsTgA0V5Z7ATBZlx2M/oDjdp4czcy6YsCpxAmyEDbQDY
Heap7djPQ/zzD1Vrvv/DtVIlBY79+QY9FD0MuYZ/Rz0re++qFEJZ+LWfDBYi2PELiFNFuF4ISnYi
1y5oRmG++S07QjweSLv0admrQgDC/YibbvbUnHpeCD5w0gb1gcSxTMjNQSFFjCK9jIqHFdzn0FWz
mRMquuKoCsIAdOnJyvaSEjUUDYOJ2H25Ajtw5MLfLCrH8aKEkFqyKVV8RgIdaLCVAuK9mj3J4fbq
nmjRXxW7F+RsOoq9zXbyrlIg6+LrVLPzz/vJMPf8V1WUAQFSlsBJcJDR8z7y1XS7iw7jvuqYkum4
K1FsyfcVacr6GKINhCb4/AgoocA6QghyWwkizlHUAJAdvGJxoNh2yqGSli6xOrK2s2frFcLl5FPh
Mw8lP3x/GD/uwA5Ait+6/eTl0iWErZWYDzU4w2pw9SJRJkFu/uYHcEqHLHTLun/i6JKCObnFrUAP
ePOcIMwUHX2yzTPF64QnTl4YPMz7+alSm1fLgRdK6YSytvAwR9CZVhB6xz8+1AccysSKRtCczrBC
pMjWRIudJsXCJwIHSeTBj61FnqeBNyi/nyyS7brQiTTqRfflLkjPWXYH/VDhtkRnAINbNGXN4gai
pMGELzpUfwyZK4kklm+7Rku5D5ArXcfSEAPx3U6WndP5AId8ADJQjs2cGlesqHjdaTGyUjs/ZJSr
QUY4ZJ25kONXqzmloUStUGBoLo9Nn8EPhDns6GPX2xa/Ba9FIqorbqVcQwMQrWrQhsbWgt1Xbw/u
OozRPru3Ou5LWZnPY7oAhOlwQoptaav6PEbzmxnitxD0iybb5j9Vr3yuPoIRytu/kjBqmeTXELcX
sElUAezxX6c86ABZD2CzELsBW3ug68g56CsC0UDDKRe34mIN0Wgkj4U3Mwkle7yt8e9lMYqDvCB9
VGd7Okv/5XFVJB4uZxj+d3lCPnRZuJ2RXSxsWLJccSIrz7yhBElWs+P8BrtMyYVQQlcmj+2eFl64
r8AfZc0gP4KSgsEBiVMXecjmdZyWvCjTcskiEFi/o60pwzvBVtMUyXQ4lW0QlfT7+5R8YkJBHeq2
9Trup9M2pJQ+2689cifII+L1PiFEg7jbBFYALd/mc/5s4PDbXMXjKRFBszMTxWSA9hH6jgqxZrEm
41wVPwym3KuHu76eCt1PwHThI1yx/cmXzDC/9Rql6+nPtrYaNF8T8p2b/nWT0blirEh3B/Z8Ykvh
/59x5YyE7NyhDWtJaG8vwvnUEvWbDQt8cthG+S39XbH3RRg2gpfgXrxHF2vaCVVsCHs0eKqp0iQ6
JPJ43ORwHLeJ2bZlng2ojx/VpO4LZ1W/oRWTS+D97uBBXS1VX3aCOx53ICypbfnzsCZan+RuoDNW
uJclZ3pyzMISFAq/vOAOow6Tr/XiCEo3Kqhw2Tk7/7cPxwcbvE6ZRK651BVu4dFOISoASVOYd+x7
ZWEvnCeRyKO2Extxe0Z5f9q04jxOMJjf8s71TFnrfqTIm/GvupRxQYggqANKVFa7pMu3u0rz0oNA
33617ElM49BpMC86038YUEqumnTY38CMSBtKOxrJN+od/+5yAvA7zlrCvTfqnniJ7TgMWiS9So4s
nIAEHiiAqBTTSMRp1FJE7+AcJxi1b0Cok0t7z5nThXZO1O03E+5EHzgRDRxFdVlZ5L4A7isU+02T
WHWSgY/i7+SFpKF7i9axK5xJwbNe6NYp7mIVtIjRENcq8v4BJyv8zSKV7YGeiF7hZ7BTizNrYy7z
wKq3wWztGlGswSuslSuWtVTaYStFI/19pD8m55fR6bUE8WXqJ8iigQs7llkF0/ewHPnCMWgSP6/H
BLbELgy6JjEJoJ+NOnp44ogxRq5cR46g4223C1zRH/RW0V1Bejo47KUMbWAqW8kfQV44CfU+mL8R
LWmeGp4AkANK9tf+bH5A7vE3Gdjak73ubzMhFyoNElqPzsgrcfd83YN2iYAg8CyoKcFGXaEaYJv1
y2RYocQhtnkMDG8eunu/okxDtRIpSVdPQTwwRVVGchL6yAE/5Y0qPOZ8u+obhq+H1bzfTcpiYf4u
J+8wx3GFYJmF4EO4qCAZvb+fiDsHC4cdktb+EPeBqOGakiUuzOgn69B0o9KAlVQxZcMpk4Tp3wgA
Q2t+3E/MTV6miEEN7KPu00DDyNc08Vo24Cp9Y71bnIwHpzLu9se8jI3ykKeZTB3QaoBTMPoQekMB
hnp5olT71azQ0rV8iC8/SRjn+Dh/m7DAhybcg9e5IodWNqQgq5fFbe3B8/o8zZe8ormgZ7JHtrAp
u6nVEB/2+n2wY/NAlgwXQJrr96Sm9m074/Iy5VLJ9p/GnV4XPRxHi+1Lt6fjr58RFOpVsBAgED2G
eWDym4LQdFBTlPV/hOiHwBgbFIbkTZstq+XMtZ0S6LlJf7Jwoi46sISEdRhyagY6lYb992NWHacQ
hdz851DSonoPRuyKCuc5KNpopg/3MY6nfRP+QIS91xWJup+c1EIeWmL67nkPHjR/sQ37VHaYoO2I
ehfJMJUmzVzVwPAkL3EGRZ+nvsIqODSB10UN8tz+Xit3L8/f/+O6oHONisDJ6I69JJ2AmUOAY/nu
rkMpyj1+Q2xo/wq0hxY3cDwD807IY294ohO4cw3qUeYmc8pwqnij2jIPAVBM82pNSDsFtiZ4WRxj
I6PIt6NwAU/JI7edvjNgxyZanr1Ou/grjkw8aDkFuIcZo6NaU0AJgNG+E9aSHsUriXxcYFuoviXT
S4yBmwsEth25EDaEsA4hae+NRwEq+hrwH5mwefzJAB34opn7WcixwFDIdgsmregCxUlKaYX4l43z
r2CXOqIQ7GSjO3sEEPAZOGkvFRWfga2L3/T5dYshdVZjkpmwzQhVqKX291mFyz0bxbiRRCyxHiSd
GtSPiND//GQdeYSBPePWKj7bY2birIP8U30p3TbpmZok92dwUAO0CsJnTlxd50fcszhLk5nZ+o58
UBZdLT0onHxEqcboQ3ad52H25RWpnk68uVJ/mOcnlKC2pjJcfIf8ui3b7twbUIhkZNzOKDNS4dXI
4GkFWU+TLKNM13nQHovYD1GcViiPHVRJH5QWJT4DIvc8Sqsd9gxzjHsovdwLbOFiM3YDqUl/VGs9
azNNkGkpFvTTozotFGjRVzfsXHhinN4NJm55ymqYTxg6CE5jwXXC3s1yJgg1HHCRkjsJKuxRoRaB
zxMAjF9GqXsiWZoE6H+G/beQ/bNZI9bokRRdOfl2h9B+TZORMJIEF48FmBljoHN2qpjteCTm5yPA
4XiTSxyBqFRgCc2MknjawiFl2q7esCnj95WeQJbo9tq0EDEpVqwLoFetAnzYhqKI5horYvvGkprN
G+SL+N3KAnafrfMz37/YXYVgmUV/OEI8NVbzLy1qfVElQVtfMDZlIj5j/5uN+PbeXlgBrvdmAH/i
fiw4vYdRgyW8qS/JwXmgVnODekT8/undUOxgftZ4iZtAJ29xC8jiQlx6jeFH7dIz0flMyl/bs84t
VCFl6PmyyjHuDCZ9mG4ay037j0GHpdprDZgNH47w9/ji5TBOlbnuJmxDQmf/D+/h6n2GbSKOXar5
8otVD0Vw5X2mJdIbXWPW0QAUaGPEMANhpWRjD3fEOMpKya7I5kmg29lRbL/s2Bv6gkloYJNemJ5b
VGoYdO/6yFulYuSBvclOyqL5obf5XDTOmlzt6AAjuNJFr9stxLlt3JEDq5L+odzztlHpoP+5fLKB
PbmKlQzv/IAfrJUt+jZIJQKDOIPWhoIPOzLNuLE/OkCM55Hg+CENkEMPCyvEdII3uGNaS+UZ+z2M
kpK0B1BUMAnrlUkmO2HbWdCDX1x5Lyvg9WaYo6gV8gzMnNDXtpb2igsOrB2NeAjgAK93a0Sx+F3E
YZX3sV4QowjOntzq5MtgZA0Kp4i/fsEO7wSZ6qk25+4geAS5I6RyVschsg+9F86Y4k2s9wPVL3+P
B0tC/xuFH1wBNz9hHf5X9M53zHTG4SNAca8vkfIBA7CwKGX2u8oa0PtiHrWkjxQFEbIG3G55P+3O
AkUNrPPE7olB7jAxi+3vWlmG8ld+zSk9Joxed5dOlbrLGIvunMOmsxhRlRIpezCVIpQ35nX4wgwU
BMbPJ3kL3Jihu5iWHTnSqG1VSfGUnOsFQN7EiP/FEBxx+2x+Wf6uOBCknZJ7ZXNm4RwiptFhn/XI
rMUvpZuiXxDkvsbIWSNbpyIU1yBBk1/3XfmkLc5H/88oFvYwV+En36x2AoUZ/KWir/EXu0wfX82A
am/OUirlx7Sg9GiQBWSIPGBRV+ZKzMPsWRrx2axt4fFhRjjTJjcoT2Ao3JgpR/puyybLw50XocBG
9yjSX5n5rk0qW+MYc9rK+QmHSfvxUMKw0fqKC44Jewh258DQHFMl0XpqQ2pKObRL+epwMtG8iKyo
N4xhIqHstUJu8dAKULpFon5wGGkvRFqXRctwFg3mU8VMEujS5Al2LVhObOZv3ZLC8m/2NH2gZMIz
Kh9elYXwLEt8zRMmHT78QLP7B7RYTKthwnxT4BSapSi2x5QbfNq7cAM5e570oNfeH6EEsr3pnxmx
e5gM652SBCgLJMdNzEqrFzgdnQNy5be2bz/fxPipeKYzb5Xr2Ki3tsBrSZfMwCkiI71O3wvAthhT
4bKKCWeIdnHDn/LalZ075kDkwyEvWZc4OnUQa1DkyVVS9rPdXvwHg0QZ+WapXqBsT1a77abBNA5r
ObZfmSK2YwNxKi02rrDY5ZvQHNisqRiBeORWtekGK+WW4k0WSWwXZAK+ciM/UlUQ4dZIwm19H0k3
itU10cQ5+OS5kMHwTAXS8XXA5M2j0F6dng8TP1Bun3BrEVNk+Sn42AB2FrBiRq7/Y4ZaQOJkPjc7
BIBqkje0c8itlpdu2SaMMdVjuwc5DPZx86zNFMinR7v8iWS4a8ZILKWfDI5eCbE01OPzSoLgWyug
kSV9dhj5Aneo2DOAI/vCkjBF/uENAzYrug/oLjkcBMr1YHwZS2E3s/SFpiNnbGaAWvcuyS1wYqF2
tr7vRNoBmCAMzaCrtvr8/vqGh3aUe90p2zjIfXvhAs0VTc52FVp6PxIaGswip8+uap/1ojUpA1fU
FDhcmSFfR2QKVWwZ+fNILMsHFJRMYjbYDO1Z+0pWkIZyfdmna46lbOWBu2od8ZGVlNjA7uMnT6fx
5UbZ8kHNstgmg0n6JkfTeP65DC8BvobXw4rtRZis+m0VNtGDh3qKl09Fgm0+nurTCHh41+wZZ3LQ
dk6B/BN9NVMvbK9gXenzAYG4nHVAPEObXkfQ562nL2XY1w/h+4ynJRAbtoPUYurQakAkDliKt2Kb
ccfWxYsw6mKn6rxZ3GF+wQ6q5SanuBUZeDBCjjhipxjkwvDCVMuWNM1UXUskdHqaLKs2vGN4h3F7
58xM43VDLhFe9VprhOteU4XROJRAU3rey6PhjXBpeqrA0P+RDXF8MiWZOgjwonA6+3xmAlqdejLn
j2SekO+HQ68UIqsodbFKHhHzqHX2deDIXDxb7/E5Pfl6wLUdS6Tm+976VhuOYYhDTn/75FTox0pT
VplmVWEY9GGAB7WGzrfB1wMSL/h1vfMc9FY9VND+G6Gvtw3kQPJ6M9/vqnP2uejtW+nmtsDtv7H9
2Xs+3NUo0Gds6aZokx7VyZpUh+Wx+u7ribFPoMCeMHt0XStxJdm/eqvcPy3d9QR5Yk6ZQwv0R3tp
0jlZEBfixcnv/Qd7bEVRT7y+25qNxiVpiZaZD3gcZU1o223uSdpuPczLAI3pl6h9zrOYNIxzAJwV
ZinqQLGy+b6LSeUNeILFPRzUJ6KR2iL0uQQ8LzNCTwLS+BQvh5gxBz0t/u9kmb6oxZwqTRWNbu2H
Pij6xjk1X3bFczTT+rNaIUpzQdbnvQTQ0N+mxFEXfFCLHH3Xt2ca6YU78uqeyMfbhr4MGYAHSyxz
nXh1zHqU+4N+VJM8E4fI7HOruxIcnGKfu1CLNEmLXak47EafLKt00ikPte8zDbvsPlfgrDFXMMIZ
KOgVrQFGFKVWkKC4sZmkWC174b3U6sIJ84x7mT34+nCw8ZLpTIi2QwjJDAK9EvUWQMY3Ix52seph
jPKZFOQSpXysxVNfgJeoJf/dMCmYcDt4rAqramDR8xkV66mE99fCIIe3/Kw3J7GLNQhnWB5I+wVT
72Uk6iewz4LRzRJNorapI0AOiYlCM691/W/4V/If2Ws7DYI2STo/tV5PDTSTTVBfLeqV9hIfwpUG
SW/Z5QSjOjPDRHYpELBhFHXsGTLT14TVOH39lTCKaimozWJV9/hsm6vb0Raqcti0MdW51mmYlgZY
kWFlkLFfuAhRuZQ1qU6Gp6aeK106HWK2dvHkqr3Qd89sg+YdNMe6aY40YlJhy75hGnmvqdBNejXu
avlrDmZ9sO/b+LnjgAZGhncnp2OK5pBhWxdoW1q2AuVDIgGsxhzkRJQSl2BiO2TQZrEJ0eNn5Ruk
8CtXvRA4Ji5vAFSlEzqvQ1+uoDsup2BV822bYenLPLkCr/Z1pl84VylZ6e6M0PshS4Wh6J0Oumkq
hr3Gvi9kDpOq4KdTPwJm9D+uhWsITxH9EU6debewuHrP4CWghNyl1gfoBKsnwgOEyAYskPjf7oJX
gntuaF/LK9ZL9Yt4XdfotQtxac7bR+hwqqdTNv5v6uBIH0Aya2uVL7CoDIjqRe1xDEeuT3eYBxcm
N7jvVvaxQcMaOVRUKEXjmTQBqgbAR3+MakAgWBOfg5DJ1MZQ9UiR+kfGtoakGTAXR/wubcVZOuRm
eUvu2m4oo1gpF3YPcrajiTJZaiQCwP+WcRBrD0pKjF0APH9riBkARjV4Sv0D44lBN8XrBJ/Wxdb0
gZxaffw699/9MrITcK9lKwSNHF7ZJgTJ56/uDMd7D/lGeY6Mo22/IO801RUxzRL838Bbft8Oegl0
rUhPG0flbeWzFIsUKHSbLRzrxLclgSovpBthQ6AKeJfEvdm6ITaGDH926woZmP0wQCoN7hCSTHr+
DpfmmT6aTDBrVMI8bk10U8WBS0JOupU+xBlf9ba/lCL1ycaFKA5Zj2MbcBzIpsBUqRVfB6aXLTUL
Ali6dhZfvPwAbtAP2573nl4UQq9rR/Ou/u+RGXxNfelZW0SUr6i6WPisJBJXxLAZWva8fXTJnzbB
je24M59AWo1KJ5AZGpeyJq9DzHKjhMFxwG66CYdofaiuJWvDtZ8WsShIzaP+ZZsdytRhffoe+CeE
6e3KhsgFy6IVcYURnJY71JeeIeeyngOBHFaKB6cGTmfkMJK0WDnqDBxillLO4XEJaHhiMC+BOQuh
hAG2JJOmEyisVf/clDVbrXQitKBNe7XEytpOWgk+uT4YpJhw5l2h9JDM5/oITFWSCbkpvE8n9UEr
fu2LKusSZMPYxtFz6Hs53yt7jIic/m7sacqBDaqziO+DlyDoVYVKQFXW+h0DQdhP+/IqEyfG0eU1
HRAXevBgByQ3Tleu+FWGb7SwJd/q3oCs1QZKRVm60uKlUdS3kCwErxFPtBxRo/swHFigB1u5IKYR
JMYkhKhINetG7mGF3gx5QH+nfIKe4hv74eEXWCgCwI0J0Al3CVtPva9XV8zIcp5cQUW0Gx6eHhQA
U96AePPz/cezIU9EM4D49/W2xq/4NmX3Wkfbq7UgOnId0T6VWvKOIlmW1zORDYa+l57moM4V9t9l
oPrEG2EVNrpgL3QbIs5ArGvUkGcgbPU/2ZMIK7zk7Q5apxCrR4c/UpXaz3GonkHa0MZsMwT/RLM+
wyXhoSc2NmPSnsFk6D9wOd384W9IwVLUqmafghxpmtzCf/BIU+k9pFa0fPL8j3UnujOxzM2Xpzif
cslBGM79qVPym0pzKTaDMYFYiHajfusMvLGihbl9+Z4CtM+FiGExrfbjs5rDWctNdMJ4gRfwjKhD
ihJ6VTSdV1hFsBfnMMlyKIX9t769RM5j1tw5m0HXb2kEPokYQJPapGlLenFFP3XZG/CEG3NN03rL
LRn/xbV2GNPRpbH7x4e2g3p5ZmSWfAXxmmj3hevLobUCUxVJ6/hDsOhUnek9AXvBh/dtdZ3qyApr
hTJBW4GRNoKXrOeHS6htyD7hNboB9mqjUWVXKLsqCSZBFlAe0ouqOuaGtW0awEfU4uKAgq8qjfSC
TBPRQaObWk3EkcwhfEvo/YM5/lLWgIN+2zfgJCLbvSZOF4xVsF8nrNSLlLyjxmd/itoWUtg0z08K
kJA4yJgCEkB2zexDEaMJ4yhXy9RrYd+PLqX5qlqh5ufB3xL9DpRNcbZqKSALxWMQLNW+tMSD6pIg
dZlKx8+0hzGx4xEHRVZAxp0T4dt0af2FvLxYpCamvkb4ge0AlI5AZU3bIvR1VmkFMmC5INh90dwe
QNfNJaYVIvNP8YD53bd5SXvXNZwKBhUSueCWFJK0MwEOWNcXVWD+Y3NYvMan/WNpvb/m7B2pvxw+
ICsh+mUsS20n9fShMHNeaeqqyIwqyoX0sNiTI6xZvhzJ6nbXHfTLaa/gO1i81024tVc+L0iG2ALm
rOiSxC29bMOaiX8RSuIgz5Ym7YIQRQMSC2RPHvCUaOQilPK9o5iDy+cK+rYTuO92KgSWlcAuGQuN
XwhwqScHkgODN+yIIeEt9bAVDo+LLF2uhDV7dwo4MdqMXJzbETDoN95Cpf5SBJhpOqpiXZYbTebH
xyURMM1+9aRJYGkpyE5004EOqkvmzfXDOp5UJ1WqvCviKKJZFZOJ4grkUv3RTC8J9F1POedF0YjY
c2fI4ELwG4Ad5y63VTrKcaEx/HgpKu9bZVzAnog2X0Gkk9l3zBf34ko4gpCjNiGKdCj9lh80ewyH
YWIsIo6oKSHBChBlRkbTLBTBmYHfvk/c2p/AHebv/XHJL0nOxcroZwUtYYbyktcBBLgJMX0C1LG9
fcyrpdoxdkcZNgLX3nDX5WstRaXmfcyGAy+OkwOKe9sqCAXNipcRZPDEEQG42PZRoWj2OdrnWG7B
/Z0mbUibTDn7pELQRrs/rPTLc9pGdRw7saXo/dFpaHbYc1ixiqcgaB862FuFeh6gAsx4COXFApSf
24DM5tLbCTN0d5APrsT2AnLcxbiHFinMjr/mQocXP/nA3LkhoRFjpmHWFeUN+oP6j5S6+U1ue+fv
l8L0tRuUvPdQqomM2nCxCDog0X17/fOD9YQsvv5auWedodwknzSVFR5llMkrajjL9gPhabjpsvNn
7vCdPDIUsiIZd5vSTWhu68CgGoThRUI7g0uzuDF8ZlxuTMp1jdMjk95T4Gb2JI+UFb+x3e8VLfTf
sqBzwThJ0gLc9qjKCNNskdYFs4dKm5BF9uql9AL9zm+hnx2eoMJOIK8cWznCsD0FKVdUWXGrr9fy
NXuS1ExccFkGDgdmCF2wLtNV4Xydk0eUL3RA8PWPZOcyoVQ6QRRSA8gB7R/EqKroinflFSj7ntJg
3QW6enwZG/SilH+8/mse7K1v0fStcA2rSTPd+cEn+Ky7qww6wc/dDBX27XvOog7BHXfcpEemABkU
M64Tcf+UOxJvUYnEBEf/tCFxYJe7B3LCMsHGfAog5ipM0LYklFmThoqQkiOPQ8Ypq1eq5dzxqfT5
Yv93UgcHvNC67I509iVZ/xdB6R72mfhcGWqIkNmi6KEHrY3d0DgKn49nEUVHhwleHV70YPQ8FfwG
XGbejGzRDpiF3ylPz+EV7F+q3oD0xOcrMXRHQ+GIGwyloUUDkUFdm1bbiQRKth99oTNIeY0NLOfL
SClKM8w1BWLt4SX7ob5zoDJwEytgPnrl/GUf4+APqFL05BdDOY1+jdrZsjEIdrYqGTli72ECAPvG
VQbzNKuTwV3Nw/f2BzKcZ43OfrgMvhSPt3ipdKZEtYdREH1Tilw8LALDe7/6zGbh+va8KjabcuwF
KyeKQVles7SYa23AepAsKrbo4Kvsst0sxLOZqK5stE/nPJAvm1DWd/db8N7SPHRZc2eI/yddyC5M
MFB/G8oBET60fvmV8dAJYfFRvxH0NnBkzlR3IBpZ4kosG8pj5BCxqT5KYQGKMQ/xLPOuckVBgJ8U
GYbj1LhgbqvEiC1NOpu332yZbIOJV8s+YYkIdHLogS9aIErhyCvs8wqVRt8ADpiJQG5Po/yvXoHk
ANTCTON9Sfh0OiNzBvaaJrBxugXutY0NVNVB7a9zSdXZ0dvSHeEpPdGjmtxrlm7qKACmRugoEUv9
l0Pd8GhERIWqQ6JHdSY6VgNInEtEFI9ZhJH6YYE8iNABhKZiKDcSS7PFdOcBW31qOiO2cQLvPTQm
IMyP912Xi9EwRPDFl5EqyaeHWHXIfLxNnkjupcdd4Kv47SNw7ZKPDxXptWIusPzwontYlZPsMcaM
n54VHRIEYo7+tJ0LGHBfLXqcYibIEqiOV+IygLMNky7Wbywst16JmFTfjQUDD83RGMa/7mYKDtEe
pWe7oIYrzNHyxnlgwurI8XNtSexOWx/UAvL+vYCAcys00sFbLsJOKzeofPI0LizopzV07E/wUvT4
vi486kTYBhocjgQ/gFZ9mGQc79ldNsXGgu5PmNrmK84m3AqAHJ6MQMcXh/BHJkGj/XacLPDhkPcf
v6ovex/6NxWbRtKbgiVq7FVUuDZ0eBdK+5cJbk0op7FJhfYFkLOsLuapZLs7ZumvI1Ccs6O8Oo2X
PRGcaBC7pjOgYnQuoTYLcWle3Duk6QOu7yBOz3vK3Gr8b7Gr0AxI9JE6vv35DEQo/uhVIhQiOZ/2
E7tJj5P6ef8R34fYXYlG/PryHB60FDCOZtxjQNQWtK5yhWPLB36PHfFYBFJfg62HFayOa/9YUhOk
0WcTJaiLNjUZd5s4GXvNEcyA7/5S/IPVPSILwd28dRDVH/UFd+KpBt15AnoS2wTq3HV2eW+wRZ+m
QFhY3W0IpE4VZXv9bj1k6CLFDdV27JB2DlmgaeMvYbTo9y9D7Urdh+9/xUI44H8nWLcoK7xCJuvL
sByc2447abqjhpTDk0nFBX6uDgFOmPgOazA5KDQx5uwV4ltHzzxH02qjabG4Bgt9LNAyHsJQSvD4
iWCaqURe8xnvdcM4zxhTgsORr2I7c5zZobZritCLAwgVqUaLuDDo6L6XxHEkWhTXaOudtoQjKmsJ
6/DC8bKdcYXY7Nmf5Qesa+13wunwDgARknOzzrNvTbN9C1RR/d8Nj8HXBzv9eA8FnT13FPm/M3YZ
DFnrnh9NN446vt+JdJ+/VyjDyu4Ru1jNVvz+B1NTat4SfLXN/PwsZpsqnJcJoQ7EN8C5sLXXVYXx
Oyni6UcaWfKtG4pedaTgmMyrCI/kvEFU29IVp/tNH51GlTcpRvapzjSZyeleDGrf92QzQBxgWGxp
HERuQ1h/DSsb2f+tQEEkp0b2/IVpeOhOHLqwGQ0i0yMGjHC4PfWcCuD0iIucctZKEw1D9+pcm3af
bzjKAsSzYaXD6oquz6DjWm6merPQI9Wo0HXPfCUAgdx6uK9KTJp57Jgitl8e1OWvTzU1e20CJan+
2Rwpr+SEwPGqdQdoy3i8WSt5XLNBoSspfdAk11yagEAqJDUBjunlCPO69wEHShR5CkQ7qBoTr5f1
ce6SeOcjXfrw2TLne6ILHMSZhgGKv+LsOReueaClI97bLUDrFs9IfyDbnCcJrIEVhlC/vteQi6K2
NPoM8yzxNh4QYdSes0UH9TuqQJyhz5i00KNhY4zTyzQqXJO/fC/wW9YWSvvbChdosPZr83fB6AZn
ELKX38E6VlL8ZJ/8zsYJXtHHPTc2QeMHqay1V5QYr5U2zRGg4YR/pKwEyn4wz6sPuZLPz4OYx73K
8F142kr1Sw6wtr39WbA4DkWT2KtDqvs4Zx0hAC06TruKGeNfYuGqm602rpMMSA+Y3zmf6+8Ka/2H
YN6+8ZJ+buyd7eEIRVQ0F2e+Bms+VUml8hLkIoRnNS9vXJkH1CzKr5RN1qKquwfrEx+NwjRYlWfv
sAvgmPtkvCqGSx8GkhNfCBT0p82tOR8PxZW171YywspizjS+0HvbWYTEFUMLpiPrv0z5jyaOZmGT
Lcu546xJvcnrrNh+UnQQOa4olemLg2cccIqF/MBosNPOYmamuX+cMHdaTJFQPz4to3gbn4jfCHXq
is1pMLf7HwW7BjCunFabyx7ac5aBFeCEo1OE1eTWg8gqPbJXO4UbI1sdqH54w4w5FhjMglFrv9qL
YGkSbtWq7yAP5mwQXs6xVtG9HVkobiGZUljJYvNYTJGgRzuJDf6Ta8Hv5IDxDfBHPiRENg4YVunX
Qnt5oyicYOrpRaoKQU+gxtXUIP2O0oYDfpcret8LVmYOj4VlghUtIkRtsSAWfr58J13ATB3/PIFI
7KFGmCBkz/DrKePzws5df9sAFFZ5ndYI5xlVBZ3wI8lR/oMUFq6tCb+4NU3MkvDII2Dfi6Cmiswm
WGyGgJ12kGFqAFV7grVfqyf6Id5CIQqcu/NJ8wiFFt241OXl0ha5kS2O122kdq0T08cToSMdNfTp
bBplN+QJWXRyYDPM+5RK+OkzlWV9ERAIGi8UOc1gxEMvLVNlHmTlGozS4H+CgHulOzmo+KtwHc1c
QEi3FkWjJlWmzDIzcpPBvF2cI857YRREWdyTHVo7Q2kvTRnRVsSJQqx9/brT/OAihcdEqTDMk0tr
3Pj3xleTMARw2eGEYdL+vi6rc0s1aIV3qNvVoLByha/+iGUWujPZKrD4V8iu3cBEEky6eRYjDrg8
XzFNS+Oi0uEoeFIzvnce5Ap6aEaS5ONLl/Brl+apzqzY+Dt5NAZu9L68EYq1F4WGNIJMp3azK0Qr
S9iAbefWNFPEF6uVlq3sveq7KNKWx85yhxCrtn0sXIZfat1On+wbsVzOtc+WIyYnKTUAthdZYlP6
YGs87whjWZjF5bIfYGp2oZDn83Aa8DoMaPlbr//W+7cPCYvHbIB22x979AavSvdsY3OUeS87vjVD
vlQ/6alEfJXUbe843k3WWrDqhV4ZAeMnLR5y8OwWIFFt5rsbC3VPTKPM9fp5NERU1Q4939ZQxjwd
EhXS5g/Rl0Lp4sC6oV4KM46iqr2L95tBs7z3QYgW8QOpwke7c2+RQ2HvKCO5cSt22568L6laWcZ+
ewwSDER7lXxNWwCoLDwB/glrkkf6zW5Kv+ner0tDPNYzkUjihhdCGBOwYJaKSQoO3Jo7D5PhRwkT
wy7bvQLu3DZzViu2mA2GMTKHjpD91wXKgmBln2v/LRHrYF0MDruZtDn/0DLgCB1H9259SsZLlodC
G+0iFF/zBj/djNjX7ubSlF7I46LTmi69+YiONomNIDAns0cQrPy4REr+Kt9nZQNfBaWtdnwN0D4r
M/MKn2UQEZOv50G9R//iw04gE+1RpMSqaiL+cdARvm6wTGWBRrrhxjmmlCHsLkSUBnyd+fGuXhaJ
fYQIz0CZwhT1tan/H2RJGg19xazbZYjQXPJaTFyFxVhu8cbWIPedpxonJer8qBE9453m5dG+kirl
xAyTtrm1ceCpiSa99bqfjvjzoUsk0XPxZHMORbymEqwT/ReUF56lzkEgy9gZ5kTYvnT9YtKHrDDc
Tyzhjez8mp6EN02puaCrRgspcs3+Po+2NLNpn9qtjDVaHw+miauECB9O4tudYwtAHg5kD05h6Aa6
n87XLORnRdBwc8HUdjuipcn4RgbxeeIq+2iUK+L4UaaJQ0uAz/MPXjxCuj9sC7XCkL4YLqICpwAM
gIyqVxStlLEszBP/A2iLhu8mp7ybPZwWVxYF5SpoVW/mnCW1UqFup6kHDRv0EkeClD4tNTWRUMDR
+Br9l7f8sFARP6j0q8FQezY+/+O6fhuE7kKW9ihpe+5ntWOYhPWG00aBAE+iCDplt9xClL3bcAhd
wnal1Z9NyTO9HPvbk1auvl2DnSAWAjxoYbTMXwbjJ/zNBIkghBSTS8xneCrCRC05h2V4xy5GQXHO
AeWm1Pivi1d8VIF6PkUvXRHYXATMTVYKOWwX5ZG3CDutzybzq6mqhSrOWuIM0QCx0G28gYVUpbSg
OADfmu+js7xPriS87TBHv03QIurwolnrchzSjktJv4boo8ltz/zlv+jenGZIR79cCh4++WI8/f/q
CQ+xCAlAXc2s5zzLU9FI3XcDvFp3XYkfQrXfWoxu1pqd/Kzt3skcg+ldabAzI3dFXsjLAprDEvFW
zfTyNbNwjUC59asKIsyln42eDglttNxHs9L2S0fVu6fgN/ZD97fs8Cf8KNayNuNPPICx/CovvqPC
O7BOU/x83SeFTbwOiP0J4p8ybMQ2/0GTLHh6UXdKRSdmAk6IkcyDop+2/4XzqTMPGgmHPejIgShc
YzCtc3yax3xfxw/BnqoURy7g203MgyWBF73ANtSzdHj2+PNDD+rEjvAj2UUPBqqDmhNYjlUhhe8T
URc7kF8BzsC03RqDOy5BNcagd3GNabij9pnLc3GbIw174nLtIcSEJwBzYnYN8DzgBT4E95owwgnG
nLPo6kj6TOc3tnb6L6JCoafJRJUyeRnJRDRJyRLaR0R2rjWu+Rg97pN8X4QKZuHhW34SA+sgj0sx
nPPwgANh8T0scthua2bB1HGpJb56Nw1doUwuQuN+sHXZvPGpSqDJTamWyLrDbm4HIOxLyGqpykr5
CzpJFnfLgx4p7g9Mi19gv42OHKlH069EfCaL6wnt+4kWFRSqOb10Mv7WzEqxXxiC1Gdnh4ga332p
Tc6x9GjALKNeoUPW1CWzaCHm3tMY2goC24fR6IQfq0u+73Srp1G3WAn7lkj87a8fRmYRM5yQY8nU
VNMGqlScMh54e7KGLNhsu2ZosFdhQObnpRQgaSsKWN4jPRpDlS66ozKKXzW0+0CTzqYgwcgp7n4D
eUxK0+ybt5zfgAbDn9f8fTIHqsIHiDIEwGMBU98TRkxrfpJSkGNjMxmlYchNqkGZnviRWtsWwpNy
hfnbl4iggKcFtT4J06yj8taRMNh0JYYHF2WsfwCL/v7+pI1WKvbgAUffjJXt8iP6GpqQMwO2uOwD
vQae/MyLSkofCSSgHMyQvdC/Y30mghlFIA7tVpmhr1yMl1LsrNmTCOei0/R0dFQX3+ajm1j4M9d1
x9dwiz2M+cEtT/4+1hAgKj0tq36MPdR6mu76eidrxH4rrS/Uu3IT2bYgpjDcbwx1tR/iPcKKWgz2
yB5nsCFlcts5F1U1KMi26MJmBRjUqmzxcrr12s48n98rVrFucHsiytv2/sBT+g2qnladAj0UwYFv
asSUipMstnqs90fuNyKKD2Jge4YLIaygIrW24mQ7SgxNYn/sQPFo3oHKPQjtjL+TYkayFJ1BXhIQ
4IYcO04T4zps3eTj4kdKIryMXmGc7FJgTE1Svu93TsHwNzt/9n4DpTyBgyItR2TRhRyUTp3HgYve
fZ//EVaf0/c5PFDMtsV/OwByTgOrNsU6r4lVbg0WImXwJESEYUWV1mtOUGViAq3/N7xFSzYbYv+w
8xAiWZQLvZb/khbBuWw6AmZhieZjKjesk0sJUOQcgb+INNcdyDAIZX31mOp6h2e8Ny8tmQ9+Fe0h
NDzET3HHy3p0NINQgkndhE/pTLLn9Zxs0z3zXtw5KJqzmv7VXuX+IzdhaYRLQ1w7LWmNi8jKKqbk
u0elUa53akag99VMja6a+kSoTIiQMTHIU05By4D4nqsj3zRF1WXe2QHYx4u9EQDxZ5XlkH7bdsRT
JitYqMea6o15I+E178eJTB55C7wrm8sP/PE6D+JHGsowjz91+AogDJlRlYrbN12yiif7KzdoLg5r
xEwokoBXFnRHAf8Cm7SGMNcSb0JwwN9ZhI6Y/PUXzA7wo4jAeGuWeWE1I/TapiddBAS6voUJ8f4c
NnqiXgxa8NS5zhl+L7AKryeL4NJl6n96kOcChnW5h/I+6nlGICGdW4fXHShWYvkcdrDPkjJQlGsT
DIfv7uCh0i2Ru6y8rGEk//MC/YYLDFfWtC1BSBWvsH1xYJQJjCoArkN2SgQG1Iw9Smw9+lvscpP4
CXb9SklLa8CZUUWbrloOm7RGDyBF9KpydjM18BElaSMu26OwzDsdDKkk3QIiNoXOt2ccHI9ft8O4
P16ES94M3DupFvymTH7POuwg5VoGmZApCBHb9OeJs1Ph1uzJAmL6x4NmKU0l+KiHbPPQrnbVV2Gz
2ccAjz2NAYy6eSwgtyZ5uU9mz6TUNHQB1INLQZSXTOU6J8DhRruk/cxytsr29RYjIsW9heTOnUdh
zXBW5b3Is9suWD8rLLnS3cWYNQskUea44Sfo1z7sMigl9P+dDj7l5Rm9i8gU9ZM9MYDu010e2o/J
y0iHoK3IucTXA7sotMW/sarLyJEuiqwh9tLcUwzguMXvvIB6TQgPOuIT2qTfkJsMscTVhXkSFWjn
+KVYjeFXAVrRCksV1tFPx4DsL1MbmCZMH84JWjB/NM81PSyS8Glx1lGUjpp5cj+TCKG4nyJMrAIR
xR8oErV+wkRH1x6GGjbbirXnjLzrAfKRB3zxeb6Ecn4+03AgncHyKKdCwOvgwRBrclr7y/KAAlNB
5JQbzzzSm7jwS4jkoF55ukXFWpcAFEQYMJNJEHkbLqeGc1osc06Cwt2uOOcYqjrzCawIh5/gJuiO
2WNAKV5GL/xxjpEj06iw0xKg0V48HLn99533bdYdO/aBW87rC3DkpScxTb01wcLoFRVG24XsXZgK
TqbD35sOJaTgAaCX+Jy5R4UXp3c4lUiFl6nIMUffZvCYCqi/sl26SX07r49LoK8uO2idXg6Hl5ad
Sg7Xv1p9tPM3M+yaz0PUEtx4W97OCDF05buWl6Vok2fY+ZWU1sr3MuH8lCO+3616dGWqc4M2WDvs
+L8/fwK5DbhmwXjvnWGlUgFqy1syeh+UgrXAveoZ0MRI9hMpIFpXKDVl4Hx26qyEny3LYzB/NQd9
YLqwywtXCsorWnns04zF44gnxKUsIDsnMxiGbtl4fhwuuuafg7Iq1oK9QlFI8nEEiBLllNBDAtZ6
q3o+oARy5HSs7U97cYO6BocL8mPPH2HbuOUUdtLPFu9wtz8j7hdtADWwhtVs6mjX+nMREFKixaFO
S2suWLreUHGlxuPw8l/3xEPvY7OgVQl/FrMVpV/Vu33XszA4whhwH7e2ZDSE7kkUTHKQBTfyYMQJ
LXaOgFPfrSFQzeRLHBzLRjlq+bjLJXSj5NQ2AU9NGsEBrOZ2h07X+KWWRlqANIR8lJyhtivYjsoB
uyPYEsxWkgdVoYxLCAHzETHsXNalZ9XVBbYy7YpO5SiG8kDUi9tqlVkRfvIp0/BKFmjDLx1Zl+Il
2YiDTGWdXtjcWksKvF79U60s/abpXGxmcdh7VwL50puj46ouDnSLNnIMG9lJqLoMXDfU3CjjI+h1
UssW3KQwbBdi1gxTu611uLD9hadxXlKsxZlWMUYovkQUuuY2g53rfWHjiL4A38BifjhqZXJ6o+XV
8t+S3XT7DtOkyQSljFnpYlDphMlypdDs0b1zF54gKXkkwIjW4XfHTdhYE+V2J9nWCRYlgLBQi9zs
R8nU+ATN5cfEnxGdU0loVB/jqNpvYt2anokRiyRduaaqM1rDFHFgPJGXLQd1/F1qzCYgTGHWZDk/
zQzv48/04LH/Nrlh1/kiNPAe8CuKaxPdLsnxphZvUQISqLAv8FtFDTyoyD1sWyOZEBRezN3nXMgD
tnRe1I7HxHaRxR3+oBWB+2pyvOQ4AKHHezelvwgTctr0TEDN/TIB5ejJNi8VZmO1djWDjffltQx7
rsp1Gvgi5RUZDZu32yFQZ57pil04S394rL3VKxZI3FVpEVgtrNae3/ocFiEOueZrkCtAN56jSjMD
sqFOuoq2McYGJwY0G7iXbj3RTIqGC9jb8N3tP/VQdkiW/Msg2SiDFYFsNoEJgWYy57pFCvleoKqC
cxlEU1ZIf1L3oPYqTjKgHlv11robvhe2EMQYGLB5yH7ybS155iPHaWi5MZC3v1mLy+YGQdII9QsS
3x1OJGiUoyrUZut9NYPAA6FIvSds38LPpoMO2icnh6JC6I6Vf1GTwdyWyuVtT8VYO8eLIDKPQi+7
RaTaOrN0RXFE2wpTGUP2FB8NvBUktXVon1vsT4VavSphFzDh0v1oVh4saFVwlzSgQ2LXXdjoDZJe
uvjih8BCwHa8IMRsjgVgZvgl/3mWzG8uBt4wioc+x2slyzlK7oaF3ejlkeSHKHvvhwWvYafl6Zhf
x+Ngt2+ooph1dZ9R7vhyZ4tSdQNJEZLsjMKdRXvGxjIK7Nd9bEHONy/CeSJeZ2ul0DZGSN4BNmtb
V6E0Dqi/g35S0FsN+TJxwI8Ry2HWcln0/aDOhdVuyZJflQv3XZoHvXD8svhtFhaGhAElG0hIBgHC
kdCcD8RkZipMOTLzAypkmyeDlSENXHgDQobSJQq7f8n4FU+WXQ1yYLc5zpaByE+6YknNc1QPeIqr
M4s7QqqqLssdmGcdhE7bmBFkKkevctFU8bNvkyKbcDQ10xFbvnRFQwpJ0HNodYBMJQUgToFv2Jt+
cSJdo6E7/Swrw1BEXJ6en6dwHBDV4Ef4xzw/9sLO2cwUTOYyOn6CCiKwoI5hVHXXRvGuy665ijOA
RJCVoW9GVQzsc+J1AmtDX0l2vzLXfwtJVhTZQRKFNCquU++8rKDuOP8O88LZCwRWJqPSsixCgN4c
/b/FtlowIR25SIaDoZcBZ5iVeEJzVy3kaLgqpG50qUJEMZaWaX16sXjJ7TDgLYYxdV3UR0v3okNv
f/hcxg8Bo3pphQbdGLifAXeI8DT2MOSo2DWIWaADuEU+ofi5SUzwk+ax/VEFBNm0jKFoH+PBCX8W
J1Skr3h27WnXTF+Sol7K5YR0pIIHbyNlwRxdElRSZsQojQyGTg3ibKgXHVz/hwWbWza/OdWF4pDb
YwRLXhMP6g7uSbd2/BHd2fPaIBih5IB0+8Fg3oFGacvmAgY/hPgfEybMiWvd/xe9ut70dlTm0+Tm
JFaiQvoK/1wMtfs2ZKyd6Tguca1MbNOSdtUJM8/jXFtUhtA5sEonH7TKHlJHZ93wfmI/ybCjI1lk
t6PWLw0g2G2yas5ubZhx5Z9zCL12pbiHn1Z9d7JNT76WIAG/xMm5wJkG08WY/CFn8HEsdj233GJ/
7bAUp3oX9t4F6q7+7i3iv3P92R2YBrO64A7fC94HTlBIkQhUU5iFNRv04T9+ItJvfWVliEgkpcwB
w9bQuRA2EHqqiayBDi/TUQdBOQI/BdMjptWLRcHwiVEZ0Qnr1p4VmaYBTuS/fyAvkjiEEIKmdHhN
Rufn0dzDAwr8l/neDhNs13MlODBMeIt9AuyEwmtl4gssA3+RbRIORG3t+g5G9VvzsHaW04ZfmNHC
9Ujq8WSKTrkM68oCojr5NqS4aHaDKSctoQgU4+npwqULxjrf8UJB/i3ukxi/CuDo6atzE1fNjxTp
DILZn2jSOo/I1u1HV7B7TtrKi4A1fCm8zcAl95/wXkFRWOt3U0RM9RMlGMNFdKCMsah/DfJHlypP
q+tap+S8efiISkypwtR3pWV8NxdWLbesIqxqaxb6lnH9bC3f18kO8bgCNiePERRRi4CPeQOTxTbJ
ZMHYzvvrgmXCnAuyrx1q5mUoXHYuX+2X54WCzJr0dc5fnY1Hh9kKYJacD1DZhGmIADjAIUbjdeX8
Nl6ydmkAcOB5T0E3GKVkdBizP8lzEQvE3zJ1srsvFpb4phqcF1TasZB2Ep4Tnxv92hhUqdt9MlST
faoqN0gV0Dp2D0SgqUHrdCkdx1jBPRKJyewETMzUYAwUeuyEJz4rwNQcqnMMDcZj+0l0iAFg3UFd
gxlSjdj2gEs+qouxy9r6KWk8agPjVdh/REtAQ+XoF3cbc994ylqnGbLqI2EViNV5Vga/Xr5Dbm1L
s1WQrsvdI4ZukRk87QDPxXGBYaaOKR09rp3NQApx3hLvmhVCZNojznYv9hyK2i5nQSY7YXQjuA+f
ly+wpjl6NGU+y3aNn80bqR5lf+Okyl9Q0CS07Q5I379kCn6+eC1xpmQVDbLiJuKG4FQT4p6+HXqs
jDs7uQpCa1WSulczpT/ejWur4kuPmKRqO6CpOGLeE7SX+4uJslEUXwopoCyVeFwJuj8HDB09X+OZ
BbBIlKhxt/nHnI6PKEYYHIm4wXyE24bRo1MTkb+IYN1W8UR9WRAE1rXt5EQhQGVaEZOHHYGeivwb
Da9dpzLMOTVHfdo+koZiyW6kIOk40rB+DgoaM+K+CgNG+KxqNQnMBy0gjXGc+EsdtgBNyvbEOzAM
rWTWuTY+mNgJakFDTvcGEiIcsfUpGhnOXNhy7ra90Ee2VEE+HUTEbLbwL5PWC8klE1ibn+kshpfk
VUes+u+vZlMrbmm4CdEcz5geH/2GFBWqaZJsCdJfFUDuYRDlpPOWtDkLsHKbZIhRWKGIuUI8dYUA
3sFnz6VVDVnunbcfnA+Wt3o+3uvIhMbyZrhRxaJEOSaelh5tP6ohxN5Tvcv9Q5MLhF8zBI2xeiCP
BumUsuH9BJEdDcemhHplz67/PzsuRrtQqVgWFGkHkQDZ7TAum2BBVcVLXjcQ9V+VtVOBPDqfVkTU
Rf/fU38NF+xijx2eMlyMlDQKfwzAZy4XH+oqCVg0/j8XLsKOZHGjtkQPV1e7Pqsp04IyaYuj+F2L
N+CL8r0jCOymb5nH23rZ81f1g7eRygm2RqsGvd5JjGkDBqoYbOImkffLLgMB7qE3uEhz5rTuBWwa
r7P7zDNuAsgsSXltVGC5B5MmNfIO/8bE8INNDaGp2OpcfkNRo5LaoC39YdNmzzRcxe6pQG1mFRIu
Y/woDe12EBAnXKqduxpH8048bhB7Qd1z9Vf3+ZOQoLiyi+7DZ1Bf15kuLRUwa6nPmPWZY6ab55EC
WVa9FC2qmXoPk+6GKX+sY36YiKGWdiN11MrMvqnRtJAKRCvV8pjtit4WjXn9iA6Jg5cpQ86Ccz4d
Fi/+b4OQSkD/gNPzj0AXX6OIhR8M8uxZNua4y0rnjARfax5LnlAAe7mW3jqjulLDTprcUVryk+wc
vscu5ES2x3IzWN8tRXFueG54lWhaOnzij73cUbv/S706FfRxinxj916h/a9CmtGnD6Qq2HEphUFP
Nzc/MLdGoDqaB7R1RZzSekvzQERR6IHgkwpvnL3qeOwhsDb8yQst1Rt8Qcs2Ab8I1t+klhYkjGvH
v/XJAY6qWW6GUeiCP3ECZGhj/mG/ErpOUm+TnZPLgCjnt9+FDD45RGSoKlIgAG3rbVOacpzQm1tp
+vK6BwzjE94LM1rM0PAe6ldFwP0NsYfsKm/2+9zIq6HOhhgCTgZqnrhfqRRi/3ldIJq48FjjTdUO
cl835A2SfSvWjR/DUaddYxJgQB1zuC1Nq8miOHEHCbMo3vTfVpsYppmKBVeruUSJeV2HwF29oHCX
sL+UZeAhY4ONxyNtVEyAARtS0uWySRHhoSTVdTGC46BR5Ozt7hK8eLN07Rgco5wh7gUWJ4S/ZtjE
+8k8QW0gtfh6CUnJ8Gh6asXD/IAkGBF98zc6ZoQtft4bIw2xBPSLgT0aTSvOsv8dNuVDuS23T2DM
SOuQ9J6eYKJRyB2gY9/46DWiiHGM4fnGYqVUJ5m0jLo9uIm4BgwT23b4xg0s9bDAe2J0lYGFsLGB
HqjUwc0sVTbThttcq6NvoMGsSwhOp2aFvchcdpOZqv/HBvWu6+J7KGkexRGFTPuI4yrjzsmQG5rF
11d+Gb2ygeScZmdpT6dcxsMyTX+pkiYnYozhrxdNk8eBygbiQlhziVpXr1EuqQy9EYR8VdzrZAty
3gM69QViFbqPIZXqmb/IUWWl0bmzkysWDFm2bTgTKPJHotUktt08xt+zzMjv5L06Bo/wfvW9PyZU
VsFSTdDaMB9XDjRfRkp3VQXC6cjounaxb9iBGG92zRGZ9LvyfaSRU5Ms6wXCaBcXP772zm36WNhz
YTpI3W2n73CFrg4D7G368phqTbIeL9+rt4nX6/OIDLBv2k3RNE08MTQFRJM0CGa4SfvF+1tsBfD6
pEK9yb/krE9WbEbt6xNVhmOlqCvL+XX8H6y3bzTce0faakWajE4lJa/7KXl0Ehi9NokvyKyZzG6m
5umEGV9TIinxyEp8ZovKlXXIsJ6kzFkZ3vSiRQ09KFkydjM6DO3is1IPXAMfKVkT3iDlYU2pALmD
u5furRdkVo9Av4/CKw1aqH34zZ0mTdWk/RL+4JAvrDRLK76XbLCNx/DUea+yrLnnKdyJ5EilO6zi
nbvHKa5RELG3FTrObU3Rz6NOyAGQ94wfLhIdFVZcroxsXJAzqTod6siI8rpUplqulxl+XgHzv3Dn
p3mQkyqBgq7228QuZDSCoTTmSdTPH1+dLZdkNEOMXT9RBE81JBN0FiHRNICesO+simQ47SuSQu04
6hL/kNlS5U0lndyjDzLXOV2CFmCBNK38H3l+49LEwk0l01wJ0nHT4IEO3fSM9e1QfF0TlrS+ijyO
bfy4dOU66Tp0HypOavEDTacPXrCbcVcBrwqxtIweisN4q/PB68ko5XyCaXyXlCslz1qt72yxgnQu
juhpzl1WTBgG9joIFJ2mo0SsqmRgOlBgi312SlGmlPxfNgTBoX8CG1Rhk2Ig7CsJO+SrNzKL6NtD
9qDm95JZmBvOfJtJaO54V7lCRtvgYTbAqPaDslpEE03bYXoDdZWwTifpeZrqm0yQIjbHnmmIkfq3
EnVpB+nhZ1bSbUSGc00I65s9g/sb2qcfVa3XSVzz/CRvBhfAL68zEdoR6OV0pS0vs5In9ZyI1CuW
Svv/90QVUTieVmk8mS6biDUGwYQD5mwO/DLFLB5IdcRpYgDmzDA/GMt41h932wqvSDqXuCG6BGJ/
/DC+I6O0oN1LLpXfjzBsuP9TjfD0pO6aHrczCL5wFtUZUcSSZJxZbR0Q+srd/h22eRWGJikM7SlF
HSjHv68UN4+czVqueIF3zpK9lBokfH22cUroo4PfWL21kLjkzZZHgnDrRLkAfIjDhQZAOnc0s6If
AM16wfDWuwNgfUmLhkbCSarvSsoDwPa+yCb0QSjNVP99fHqkSVbHuO8VUnFj5/6cg/6XLMJX9r7z
BlT0ls72FAzngWcDSpvThkN71ulA0CvPFhDz7F+XR/KCkJn0HCqrSIcxWJV5xiY29VimfQvQT5iz
thrAKx+gJXYVtXLV1CfvkchW9fuwC0L4vv2ABnoNw4/5jRae/1WyJC9938BLyfZWwOpt7ltCQWiV
1kDNpycEEl6OBF1gktdKA1U3Yn2F09mnYlbMqR80WVkXQ64saeob6MuYxN1tVDHmUEnIwsK5JTZf
IIbyj9doIKgy9zCLANEyEcj8uq5S7x+tQ7CEdhk1tZi7icPb+bQw6Uc3ZY16hMe0xoWUV+BfYeoZ
/OTLRNlrxR4qIlt7zzB2T8NFC62YJdyfoCoyD/eSZ7l7wc1WVqLWeBdcEGKtQjLyjMzOljKqUdoQ
SgDWrBLFm/VfiNDH3wrFUdO7gcikXNf85oKosJ22iwU0bfOClH96X7SrcevybnzgXM0+IYp9v/wM
uMbXPGl4ULw/o/l/aDm7oMh7wfRnW4RE7PITSdcGBgW5/PZG83E28uvnTMwFk62XXhp9Z6IapvvL
o5c6Jp42BRKkJ5ZihXnhy/m2zEV11hdgD2wkRfJxTVl6z65o2/jA2n0nHZDL9Mm00+q0zqvtUlqy
sfCaLdMOfr4aw1v/OE06KWpw9T/vmRpxVx6MHN8TJo9I42UB++I/106R+GhNP3Z2p07408RShugg
7hqxO4/coMDQkBim7DzGnZMhwnpk6rps3EM+ZwW5QVFzg352kw32JYGrGjCTPkXo6VEUc8UUrAy8
jz8/jvfu6LUUKP6k+IUfNP00o/W8EJGVQ4gDThqn2Gc7v699pk7ZfFYeBOioomsneZqY3N7l7lMM
B4d7aQQyYjXRLlcZ6z9Ev/brqen9NU96O+OL42j2JiaW0BOjiSRqLKcJ4h59BHGJ0Vp0w6hZH1PV
JlHRxlCERPi5wH6xm1V2yraWB9Z3VtgL2c5SZzszs4zL+4BmNNsF4A6hOxiF5RGyaco53k/Q8eJT
FxcA+Ad7mvlc6jegXd1gtkAGQydv/ckpTgLUmzmfdDJtQ6g5w/2KU9zOyKpz/Q9Xi+5vVoFjY3Qj
KJQ/hPpVKQbTEkn/r/igUxlvXCWgYJxeig4tsGYqpRU/RnaH9Hb2j8f0JqsHWd1sywPK5sZCUZP8
EbMb3ErGCEUJq1OS2Xo3LOFBvRunkAej7S/cLay773Z+A2YQu83sxBBarp0cjQBBQv8QfTHQCIra
duzjQgPB+86T0m98p0Or+G2ps1NG/fHhFV73ZzRhvrFXLZYM65yV71tKw1km1YVS/N5WF6Le3BZe
MRpWdPjkpvkFhiMu26bUsArn3plOrYlqQlER3jLCYC13FFhxRnGEVeP6u466k4BbE3GKhXCDm4aE
6dp0A9fQ37t2B4G26MYx2/L2gO7Tq6h59h5aWM59ddAT9QSLx8r08qTYGYEbrB0uhaTcQFvAqQfR
yXrmfQJfBVdzK3sDUL3fBFmk2wm/4zCYpn3fjg6V7uJH++iIBP6ZbOo6ialtkajqpWGyfhFtEyy1
/nZhxBcEwQJVsTGJWfSryxq8WhyYy3MbH2usR8zORehr8n2AdWqJgDl+9DIgnj5EehpLfDqtD4Tt
N25aU6kbL13k4jJTJZDMBL+vDwo2rBHGiGcpP9qDdZBCDPg0NCHoNZYM1dJSHv9G1Gldsp5yfrnO
t8PW5NReJC13vAQGTFnMshhYgLTJNarNdoEfQnWzcV5BstHQ+N5gmHfIYpkIbWG8yHS6dkWaoRwJ
TmKiXQFSJApAoXiJ+waauYOKbqXoOdjBb1AkEvBJXJoDvFnSapYG4Giji0pgmQ8+4z+F+CWwHsI8
l6oOpA8+e+jNN+9pnL3dkt+fQD3o3q2a4cA2673hrRUEPMGV4homjdlRmaOmMjAuJIttUnZ7ATd7
OdGjCjqSkGMAxtl8KoSXBHPl/Ch4h66WKrd5O8KRxMf+M51QUORkyvAvyk6KpE7fCPYRVscnFC8b
w6jFJwCpGwnANa9SMa87yKTfr3AusvVFixbGjhA669ElAYZV9T4cCNdZpR2W4SYEKXrjxlHMblKy
Bgg9NIVCIM/FpsDDnAFdXYlhn9bmMKIar++hDwMKZeuxQhBsDivCDKCDRMoEPRLXQhA3MwzsWIQP
Zqa0drELWtn5GOtBc+yrVOptDCA09Bu4e50oDNjLAimbg7L8h5RuFes/e1gaE8cEC2gCIuogbC+v
PBX9y24j+9mQQkC6H1lhCayCJTb53CQ0wGvY9767wF7megpLZIXUqvfNoNzt4Fx4C9ce7xXNOsvD
1h/+sI+bxbL6NfA0zV4z6Sfv9YplQtCW4m4ScOHkex1eoJf+z9Mkp1QMPZU2pD83O7hvcjHWZlL0
TKs7m94TuUyLR7wbow73GzkRZlneRq1qZgKb3layQhHs+mpaVDGt0o1p7s++E7TVQ1oYU0dBWr3a
71VQUIVApDksxywkAYKsxuuGjijrzzmy724N2q3rBc8+AjIZW/naZM+VyNRjXYo4Y0grY8KIlr+n
0wd9BTNpmaKAJtVfmezsVuNQtRRcAbb4rwTzEuAOl/rMnYIRAzfXOwnuLTMH3rYw4qvsN3r7dPH4
8CdiBiuHp9xsHXXk11cli3D2QmpB+1AakYVHnPzWX7FPmyHWFOX7gHJ8i+kqyNjbj9ACrZWkH/E9
DOxmBKlOqDLlr2AYv37boZFzdyvHEU4hyrs89S1TgCm8z+WUDYBKLxPrbGY0FeaoRrccDWe0HX3U
Yl65uVBeB0sLbrriiieqJCDuK9k94pZ+oxtBBBU7iIxASN82Gyjhkso4yEiQBwH7Y/DV5vPNVO5R
JTmy9CqkIFFUib9nNkV02DyVd0C2PK56OM0zDZo+YkQRF+VPfLrUrQbAIi9JH9JRcvNrbSTR6yCl
6+hdoY8Q5glkX/LuwDDx/VgN855pIc7JX7zCH5wcPTdUayMVa6BAg4pBgJMxTdtAh6L1Z0gIFav7
KiYkYb04SrVeKhC/t1HDS98MsmXd7z/NZI05Jd5myyeUt4Cwl3CA4yVVa4Lt6NycKZdIPmzw4CvE
qq5xdc4WBMbjbSrzYZK2JjnTvuLt58VLsv5XK3jFFGXEiHRqQSu6G+Y84zEqxjqyb8Pc4eHNp01V
2aSXlmENbzm4h9NxC9F2IJCJyIA6g/GOUTUSH4PY8DewLZ5C4U7zf/lD5tfsHMuAIIjyC1XPkXDI
ycFPX531WKp6EvdLsX3p2PbP1GkzUoUKI4obtMuMuygMsDwVip/w3/N87EoUi9N7i42OQhcvzFHv
OGX9f8BOtf8aIYHwiztdu9oKPV+V0rkLBue0QhgMb4mZHsT/jrMUxKqOBsDh9hXHGGFto9zIycSs
ECSFMvz40sqgb42DNHJ9CKZiyW8m6bbq40QpmMpvi8/R9ED2oNxGmVUjmQxqpGPQkBJh6of7SBak
fd5ug5ufX9O9qCflCYfj0I9i3GkCF+iQvujAMjjDBi6SfcWKdt6Y4iytRpC+i+PtuOqOpg/kU0V1
laulb95jDVjrBdAAs4UCRVGMSEAbMZdMDPPUyzTELhEom3mQtLIwhhnjC+pRnXxTR+gYWCDA77NM
5EGEN9/xzV9YBoOLI00d0SfwK0e9TkVQ22xiQRYGXr0ILxZHGQ6k12zhzcJfgGoaj9kuInbrzjrM
iSSZl0vx/LCIXvUXFJs5gykU09/Cln5RA19CAXDkg6Ldnh4ss5J/4fLhMACtSTtafZga5urYe6mp
s0cxTZWeqHP61Kq52Y/4Y1nrzlcAkojeJQ+41VYBLdw5DxFdyYY1Z+6PzCJjrwqAlFNvMfGJ7+dq
XEWab609k/pwbaMetZTEAVss+GGP1RPacvC9r1b2WRtWi2wRflTvPOwlUnFjb3paH66Tzkciq4AD
/j80BKXEgvB7/L2bC2Ptyp/gvoKmbrN2b0r0ePgDU4Kp4QX1RRmw4UWAwYbJCjnEgyde3KzwEMNi
meMK/mU+mjdfWsGTPIpBY7IrrJWVvmhQw09a4BqmEpTvL1JrKq6Lr0YIXdOkWu6vw4cREtjZs24i
4HiLgWlH9dPJJsAW2sqjBOv/JT4kqr8fDEn+PNEh6f+/H699Rcym1HxuSu6LfzS9zHVDiR2wgyb2
MVKX6uXXFyAkLpgpWxogGqEV17h/cycq8XHp5IOWD/7ySclBj5IJM0LQrCU+9LhA5oGKHaAWqTZA
Gpr6S9pCl+K9AyT4HqFdUpmmz7fs1p6it7FHcFySdohcgVDaSPc/sPpVe+FnsxvopaHKIo5pXWQu
6FyebVHG/KA9sobAG1ag4yYCHUEAYavIh1+Ojsbz/nVUBLayo9ijJL1jlwoXBc8b48yH5dELT/uk
a/5fVv2F01zTx7B7L957Qp+gl6oH6R1K7OlgLWlKZUNsdn5G6BZURLoKHXqoeVBC623B4KDTIbm7
Z7f295/3BcDXd/Ge05Wu8kdqsuvZLQTrvNKO0MNqVAF4ds6L6KWFvcp2jRDcd20K0+disMG2HYaZ
1AFVljfzHmqVtx81VE5KoaxmV+o45Irq1jip+2aHOACuf6dBQRcBz4+lQQiUG48MgyMm0gyb90f+
mhWdZijx+hOFSZggNxSiYsNDi/Yih5YMOjDkNRLdfyvSpnnqyI8oUvdoT+MwSwE1XyWgJQVmHnXw
yEEAnwAs2CimRDCpdoPq0vZH8XB/hcuFHnLWcKbvwJSOBZEyUxORfT4vcF6gTuqcBugf6k9skpE0
pDQHQ5GTWVfQOaqnj8OofsCvVMOd9/1Ij9h5vG/R8yeBVfp+6uzsHV2zFmABdFnCpn/czKTIgXZF
9JdHV1qKAu0ZaQzMJB4dYsyqvKb/PjZmynizr44dDvGDdP7PaSThNjOBPu/h1/86uFgMlCvazLnM
mnBClyuVFM3JLcfvUWMdaj/PQ5mwMkNaVPfAZCE3V0KEUwrNgZm0oiL0kA42drfqDAdGLJVvSuZ7
s24dgG6FYFjONVU66N/f5PDLG6qbdaD5pRTHtsYPsilgaUwFvQfGJ/XzHmhQ33OlF+vbGct+CpqC
cTsUj1jknQEkxeRq7BD0avwTveoewPMqEUNRGK/ke7wn0ucJ9FWS+vdWXaVaMfHCf66FMGr0rxyU
enTHzKmnlOleJskVyaHzCaPtaFAsFSyKsf8CokdR0j9q8TwoWMTAoc1oV293y3NwsCUIKL/Ivt5r
YAXmhD+uEI6BxpJMZsQwtPZiPIOCoixGsNE0C/43+R1R1IkSznbjuFo+ki6AEFwwUHfbiSrmhoq4
ZO50eWBrn80fbblkc92Gx67OgX7SrfnBUtgMyYgpWocdEE3S6LgjoLeWalflG5n51bC6qDeTWbkj
YVeaLvtPAzqCqXT1VTxYUo9a91aZHbYQsBQBW6/d20hGXfVP8e9HoP4jkR8htdqlWW94Fw8Hc8H+
6TqH/4jYS7n2WKREpiyqej/V1cl62RUUoEqPrvLUwow19wVHkPoM/pHfVm+3Q6sRxCuZyVmKtTDe
baH5daRCQ6wodShpoxVwJKdS6zGIlt0/3lx/6fEbJ07x990giKW7Zvtb0r5RZ2v+axxT4YgpBbYN
adNvVqXyZUx4v0EI5NzcOtamdz+yAdMyGj8LNIuXnkNAJRHyxUovbFiLYUghIZIyawdzkuFRoJLr
sMyM0SirbpcHV7P0ItJ0IxW9TLkgANn1yA8GEtvXkqEOdKciuSVBxaBE31k/h65abby0UF69xMiD
SxCZ/8hmC74dDucMVng+Or4HtSSgLu0+LlYZlMD5g8uuEhuACNNmdF8aRhmonVDNd7pTDtZ+x6E2
kPi2x2lPLG+lmoBt5TUkQJX0MEwIhF2M0VPb3pBJdWFs7UFebG/03orejpGA9/AA4ojYYu+AmTnq
iviIO1kH0dyl0s0KOQtfjJIskX9tJa9PoOqFIK5YnIKBXU34VFGvliO1si4qIlsMqZeZcDqT5GwH
aTYd3T1KuBG1C1kuKCh4pTMlwzkGR2nKKcGvDZhFmvc8OAfZir7wT6ALp/Nn3Elgn+JeWxPI4Bhg
gITa0q93baNinQ5OvNWOPOB4K5o+As1MtDa/qSBJhcL2qv1hfw98ilFhKHuyWc1usXEwqCyBjrSH
Eg4p7pE254JKhSSKcuVABydB1aXWLJY/0Rt0BhAWN1jA+ZobDMcMPtR5ja8H8AHOAIZ7xADus1UG
6aSYAA+7Ur4mKIvH/RwMTDP4w0FOIE9XNo7mLlZWrIZQms3WdiMq3J9gfL6rIM0u9xA3UioV6OCw
b24rjm6XHlZ6VpdwE6Wnwv2YQfO2trwwBWFOFnog3IiUkM+y8LBALBNBVg0UJnhET8dJwmTCP3Bk
xaPMUIRcUdd5MkZgHK/rb0W8oOPzzeJo5abQfJTmvxw2crhz6nnEL10DpWIK0qaZS9WTrbXv/Iil
WAFbtQyBN6uq7itr4gjQ/L9lCZxP1BfbYidm/bRjIovJP0qDSqG9LypqfuwWoe5LC4J53DeSpYgc
1X+bCpd3xWK1blRoYLFNgzL/FGFImnEiskH41WLifaRkSbI2iJtKfy5fTF5D8OZpIjkwZvN/e3TT
e+RaQRuREIKokd9Nar4Ap1eFE0gR7hTnT9F+Um9Utu9xlryXcdfWOy2z1epYhayKz53gwLYRa3pp
VMaVhhMnz+9BREtQHpHwD/VgV1xbxA2b6ukjz6ZOu0K8OYjwkQL00YwsO0vBjKeDvfLPSXo8YIW3
2BeZ1Yv+bYV9d9BZ/s10+8wtQb+bBez6X7INPlc6aLXxMoFY1YG9S8NTK6Ey0c09Oue6S50GtrzR
QEv9EixjuVy8sL4OvtiNHh35zHUbsui7eaaFKmJbxiYuxkV6idz1K5iRSj9kZCyTvBC98DediufV
nzqfM2QULn9klf9JSSzomJbIV645a5//0pfZTjcBv5Y2Ysov8E6xFHe/YsGs6yf1JhwU9BXwtvkH
+gOyD6RY/o0cvL6iYuetpAPagn++GlZu1YSHCAlUXStrpv2mZeLillnyluJCl48VXXsHQYexkscG
CIXin/+kSEse9e1ygzoCEON4N/nUMUILgq8pOpEyuaN3hk2Y1+XfGm8TuREWc8Dixtye+24q4AZA
eNBkqpXKhaJmzdvLHjz9tHNroTXfgS/U963Mj9rJ/OxC6a/xCu+/GeiSf7AojafzZqVCot5C6e7s
CzWVo3w1fBZ4EJGLHA+Epv/y+pvg2v+owwkhDy3O8EG0iExckCxnsTImTrCsSUK/9cwtv8HFv4yE
Yzb6ggUhrzXja39bulaWi7/xb0XOqfuqCYo/uPPgnegHczbZZ+PxPvf99TIb0f7VnKdmE7YcyxRB
R0IhCfOriT7pYjcS1KFmlGss9LUj63CXXAKz9qNgFgvXmw1fHl4nPla0aCQts2P6joPS5cBfziAV
fYP64u3R3gN2JQh2vk9Qbs4HaWFlqlSriABJJhLebsa0eabKnBKakcESvr2nV3P4p/nLHESkgieg
zFJfiaka1pvXtbvOV+mGo5Ittr6/YD8l0TufmE0CQGZGGWY1CHXAejpQKsebpbQVEL69CJTNgTk8
IGFI7vLOm1oI2+iprGK9kakTdVPLdBgwYPTMrnvZjbssHJtU2IQKSKk+qz/Qamkw5TwN5bE93Hq2
/pEg3gx1EgHYK7f6TwnIWeSa0csdyUmxxQSXMAE1XYeSOTleN0Z9pskeYy9KBDpr84XHU/OUHhka
hnGWUXjmcKO9CJAq3xURxoOJgsmbObhEl2fkSjduYTfx0UeHZVSgRgYCAViEUtp3pgyPRRRL4t+f
k/ZdHA+RUOKz21z+6FOy1y+hW1gq4hW6OVdPGMf8UHwrfdGM05V5GcF3pIKCnYtPQ67LfgMCYHbG
OXhg3/7EwrLukbV5hcqOmfJxYBgRmlYzRU+4t7xOlx4UxmLpSr5srbTvt6sObA97lFcoCWr7XARM
ia+mwmMQiqvCqBFOy0FdlzrMVnsPe/YIpJ4G3G8o5hMAt1bjnuYktQYb6gjzWjp+PJDxe6JRHPRB
rD+y6ZMJQxs/cfMmm+POMsKmLEp9z3VbjG7B6picJmFAMx8nWejKA09lR4UhYKYpkTD+zF3PHpIk
FwhW8Cq3CqRzFQOhZhG3WTC0OEMgulXVyOyPXnQMQINt2aLqb7byeoOsUgbHO7HjE9b26TV6qQ81
aEarQKjI4atW8XnC0dL0H/7dbdHoPDXLgzx0zc583umiuyACjXQgxJlVVWd8NnQeSuE9DhIaWYPw
VH68NtJ3MtDXx5kQjvUZ1tFXtsVsftG3vDRgi4m8qozyHKRa1aaDb04TfGMhJMO4rU3Egv79QB3e
PITMOvLFjOM5ceaAJTdZEOXbrYbDagTdZecamFYlFocBzuUn0ZWMzCzCePukKj8WQRoB9/R5eZru
w2sYK5Ou/TXsWMClYOad50C02gVXyEv9JN8BJgZCLMEHVlV33nXAegnQnP2S+R8I83CW1V8PTi/1
S2PNgAYp5nmF4QI51Cs9VOdoIEuW63IBHPDznpoxKAwqeVpM5FtY7u7pGDlmJQLibwz0py+aGF5j
BfTd7TBoRfo9ZKyTXKWNN9MdEKIxun5OjPhI1EIscpXRFASgz17URfzEkgO+pUmq9LB7zqBoHhkE
gQhQZlpQ1XV9F1qoL7PTSNkYZOUXrVLGM06SRZjRG4X8GzsEJErvsniWWI6AsjSrwO+wimvyr0Hg
5YIciYS3X9klnjOTFYqI1KCPURQVugYoU8hByYWK+v3mWXWef4LZCpNNZ1ip/TaqbG5AADXIgXzd
0tJwEiYZg3C+Y2wemnxoge98sL0kYoIIFteHt7Lh5gUfe3Tfc0wJfLnh62riiqnvTpSRj/a2D+Fd
Z6h2XQdYE49lXOphxzoeG78TIqqsSQvUY35g5f5A8FfJaiXlJS2DnmrPMHeENDEviKKKjPuTl6CO
Gg9arydLJtN4DiG9yBtcUu6mAnmB01cVTM7w8w49VPGJI3TZXKorm4OE3mkYshZ+PADqT6NLVD2X
1P2Bw+G7SRajE99LVnhoLqEmSen19hNnl6RsyhviLqh95acINQsvzqt5SdbJu+U2+4vOZUVm6MRz
tzimhSLLl5ryTsacCliZeuLxIerSK2WN5iQv1n/rAk2TjfbMHMo7G/gl4zWFTfMCcjhrMeZtWTVu
1EZeO+wJpWmGlgwR/mlHP5ohAWZB0S83RWFnw6i2yPCZOXj+UxfaDfqP+NC1Q9jk+i6L9D6yJQvC
JExK/wodhOKcQt6o4qXFKbRt0iJTnPa0dtvNuuKuazyqupA/U3tLW5zULsOajT/kU1/5VcLOAZwt
MmpXa0NoMJ5+ysoFtbkHrIr+0+N046hXyV3DjxALNJUUKpCAMn4R+veZt3yX9NJsAXt1DdZshfey
HSpYDo5EVjcnJ1GbDFXVoxWb+VFwtiCDqWTwVtiNzJVWQ9sxHDKnYKwuCE0bdZzLYB+hOET4jrTr
dOqyCCQfZEkJB71RZAzmf22SGt9fBm1W29w4nf6FsCTR+7qOGMwxCNun6ivQZ5jqbfZinPD6bwTq
DhTwzIsJC6lFO/fwkA+cV5cjOvJYT4HeQ+aP7Z2OBPCgHHO/3fc7QbK0ZxVPM3ZhdwQvu+LSA85W
m6p2CH5WGYAVZMmLQZAfyua0xK3mgDvBw9+4UWKG6YnQRDpILmhD9mYC04y6Jwh2dmzwELWcZmmw
UU49otwtly3vTOU1btLPeKMv3Lnx/KDyt0l7+Q05D9QdaiWdFoos+DK2IRJ02O6lEKW1VOTIuIWI
IILVnAj67A1u6nc6jyCSmm3J6uM49Dqg5qjEhRr92ebRM4YIczvHwcQh4jjMydnZ9yYKD2KmTRGl
V7ItLaZhgmumI5AvwcXYQtldW661lE5sFeUoMyPgpCFqsi3niqAdu0tsYsBJHrHplV0oPKnAcm13
K0bhzrAHpu90AzrvMuG7eLHzBJG02oYmtmRAL3PkP0x3l0XgmHn2PmxdosaU2nlDz7dUKxsKrywo
7918PAttJH4GsZxy8xNjtjybVWYJSK6dChiBAtSQ0t6i/AIsngn21K7oiz6O2iW9J2ZiIfpyq7ZO
TuNWTSDzD82ul9AhIPOOBWNaV1m3/WTMebjEYmd8rpI2Y2LNVKYrLDo6h1WgCLu5VGkFiCeNSuFs
wEfmTBH3sOJke752xYnemzhZXgeKy7oaxqg3x6f6eCYx9m8NwIBOHXY4XeC8AP+taqB08rC82rbJ
pbaLdYWzMY1l4I1xuoszuxA+q7r3bJMKCUiAYwzzABFqsdC3GuvVPCK7CcneQiNq6mRQ6GWaej65
5DYEMyVht88sa/eaRiEC1D+pnWwyUQx3mzk2qqfV2iRoKqI/mHGB0N0iQjAG2kU25+9gX9AZwD7P
vd/eVGJImxxBRjsV/6G/vYAnKgbxPIIouWDOAioFi2W8inmoJHFdRUKye7wz7AOTcs6CoPCsPXls
H42dM68Us7V2KvDJ5B3kO1E1a2s84XN61qsLmUp22EIHHz+RZln8yJ5q9AgdihSKh4YZKMUPttS4
QmylhgU3JGeRb+9fqB6YDV92aEEi7yrP+yZptBIwx513vljEdCLVqhIkRcVh6Fyn685YL0C2GLrP
tpTyT51ZQEfmSEp0wOPcius1de4HagU13BC6UryQr4c3pfPbXxQGlmR1vfAn4dY1H951ZVSkwY7z
JvrsppbGlCFSMi7TvOa5f6P0pR8Mnj86Emno2et+TAFZ6lBmqAUFeOsK8uuXX+FDvh4bE+kvKQW4
s3ULSr7Xo57H3YwOZPWPuER2wcPyfxB79wa6Ms9jQlK9Og+84e/RkipPCx9CaP9/CZI18mm2LqOa
e8xN0/7+NNOIOsz3KRdXT9RAMnTEc4uoSCfssbVJusFh3813zCJ0YBK5G7jgtmd0FcLlGeVxa/8i
Zw+ewbpHBVYqtKAYrue4PeluqoYAHr/paUDFS2AtC6egeFjoKLbz9Xz9ch/Ss5f/ZlrTkPzYU9zZ
VolhhXPaf6T2xa5nMfYLCSut52Sw/MMBSqetth+p42FKyCaDhb5SlAj4iFN6h3EIK7lzWn+jxzX2
cMMF8hWyfjfPhtaPHAWdcH0aQWYCAHenkye5ep7XuiayOmIqXJyOosL8PhVP62fFbFXQvPS6zBKY
d1zdIynojUYCrlcP2vU7dpBQ+VovhO9Vnf/nTL1M5O8X4A6NMS6zYHDLGRPAEZHutVLxeKJQs66i
7ZSUIoYuBPiSnGWSHM7k8SoV2tYaKIF6JYXRobyQqHJoah1LuJSc8TzM8UbhQMTbquIfMlMJXrtf
us27rdppTmEAQR+WwMpOTxPCSAF4b4KFcxs3DXcNjPK9m2Dx4MdzdpreCu+DyaVsmYD6IbSPsGHH
ycB5b/9yvBZigzTWWG5F6Le1+TtDluOkXwTO47jQdBspkxj0U/WzhCRHZteiTLCvsUTG6hMPyRVi
5Vs7z0ofUPZM/MUA7AgRJsEGbbWhEbAn4LLkU/TOXsVJbKrQx3LBHP+is+o3sIjPbbJmt1NiLLXY
4jr/6uH6+lKyTnOhSlgtRMiok6wRI+E1t5iaiPPCzie2eXItQ1Wu1ohAzh0t4cftUs8+2VUmSCbt
7FDVbbZB+tpnWgbQNDh8NWGodFNT9fIoneN7c0H2a+pjT+jPoyYo6LxOnP7Wc/Pib5ZHA7Lr6W6V
PzCKb2I40DFU0KQoTsNvf8+V/ngtyPFSW1KAo9vZJeUVpmR3l5V69DdImF1GtEZeIUX1FGQbLOjJ
6eTbvPXIE6woynzehuq/jsEFhfVkc5neQL3QEtfhajZS0MJQSiwlxtllLteyvA18bV+osfFOn/QH
TiSiJlUm70fUjiwrPnWUQIW27oPXyBK6YmbhAMBafU4MqqU9rACUk3MWe4mPDOdjhlH7r0QyMo/t
csDy/mLQ8LXqHFtFkeOS9aoo5WifR4yuZys7hkMDIn3Y0ZnOg40GWkCWgQkxsRum9oL1gwRypDH7
zJHnYrAjNxYxtRpIFU09hcTBTCO1wj0grt17cOw/ismOwW4WPMULoFYiZrRugzIoBum7a/utQhXH
/f6DOPdWxQ942V4g6Db2liyi6QI7ZkN9A2OKG9FR91S6xN98DzOfVUSf8E2zhCo9258ofLu4eA/j
O979As+07KZC2D8uh4LF2AnRDPEwyrPJsfZcwMKtGGMtD4mEBDrL8iPEln98wzcjPtpMLDiZug1Y
kGYUTBkLMvilGbCT1rIzkedZoTQrbPbpzhln/Kxh8qaBln4YMlO/mrH7OdxQkbk/l4JCinKAEyqY
vS34V8ZEwepZcCgpARbvmvg4QR0HJ5L73jx3w88QvcP1AtV1Jo6O654oaVEhTUrRPmW1GgXRXqaP
g5hVerSFXi+ZVXmetFGnHUFjjNSe/xcOQho+IboY+FBxg4zFySh0Z/Za6xZDcyp88h4Cz5gBgGD0
gvpKvEoXeBAllc673aAHoBg3G4mNYo0fUMVIAUguF0ja9yEwJJRVUgtw+teN3Win2q5w73xqi4Ez
7BlPcUw2VqItoE489/ucvj/PmPq78XvjEFiQRPau+2HA5kFhh5aDkALFl96pwMFmA0DnBQkJbwLW
ljMwkyFTXOnFl5woxo81buA4smBhfaLLnEJQO/L0toHH4D5bRoXoHFjoGtJh3Lbn7f/zbSXIxnfG
/Dg0eeAjbpDW9bgMyE6pNk2YH1d2YI6/cty2m8+2M3V/x1Jqj04gdf6ubMIKpOlmzULdVH6gn5Qq
VQ6aoXeyWA+FrFvn9rpDjasapM2310O+gp+7k51Qv6B2hMVWJoh5BHhWwMue4GKoZ+Z6gD/257lP
JfMPTh8IprXvDjSdftHFw0WNZkEj2q8a6m8H2fYehy/w2kZTm6X3sFyECpz+ku+MtfPOMtPviw2H
52ztzcOXMCtty/pYWjzlwcGsn6JhCo+HtdcuGYLHizseH8I4JQE3aPZIAtJUfbzL712nxQOpGqdw
Lpr1mEOZ4yJdclHdOYcoel/oX1uh7EX+gqgPpjHwEF1TiUlV47M4jH8Gp6XHFviNGCS5dfbWMo7Y
VlDmOSq4NudhdbZkzN0D21p9jnp/tbBs4tXzijR3MrnasUcjRJpjpUSL5IO5PdRJwIimER0wlrND
n1uX8ZZH6eeQeV1onmCZQNpleNfbKQ6do2zb8TlhiAcc0iOCPm/3AJS4UYV1ctA6qOfsjn/AZxLj
wlXhtfKBhU5uQULxGE2mGe7VUqYmknNWNfgEXOcIil/hyKmxDA6g0wbovRJvwEqa02R9WFd1lfxb
0lUg5X+YrHFTEYgTOD08Jd+XUPKyBwiPRgu82+g/woqUm4aeqxCIt8BWQ20Y8vh+9N5rbV0wT+4N
IPkx3daVnaiN8eP2KZwZGTTqjvaYJe2cYT/O33FH/X0tYOSF7S6Zo7xBaqWXxJb3rF4pY/zaq/N4
N/1XIMYD8vPvw0sP06Hoog2hZuCQHnJxv2ifP3MaWXARv4L+gSm9g+ZCSKK0AkRHy/8M4FGmlEPB
Tdu9Mwwfrr6DcW8NS2dahSQiGdSjROuXbSzLhgl/07P/Pr7iGtPQhtVgW9+4M+LB2BmfnsblOo4y
GHSsPlY+sF3e4D3NYoHWHIkd6k/Jyx76VbgG3ZnHyFk6lWlCpL5+78vJnCZ5Eu0iuzRuasgWoe8C
YqLZjKetI2PPkKjSc1kMGo3JzFuZI9SmHb+hIm5mZSnCdHgm5NQn5Y78f4gSSusEIbo3jg0JbyCB
a/uge6dSPuht+fRGWS2RYldithdfaLRw1A36WoLqKncliFh5p5zjN6wd1qvtroDYhiHN7lbagpoj
Quh0sXL3Bv4hPLV0S0nIxzOQtBmVrhuSHfc9Igr5qqXZtRJKONeeb0JQ07B8fEIuDM/4CS/6QP6t
dk2BN/Rw5HOcdEghWInZa6myMaW0G/JMjiOtaIAvoQv37wRAq/JUWBAH1Iy2YPV20YaxptpUZ/Y4
5/kWAt5uFvb88LfjlJt7lZW2XOoMt4/q8A7bYoFd1gtcIb5YnHrXh9jYd/m6G5GMjajvlGyo8nHI
V/z8Maworg1Gle+woLMmpGgBD0Q5hS9KPnkbzkl4mq+Oy1PEG7FiXmK/OJk+lRwVPa9eIv3NlYeQ
DbR8kAGxMmQst/csmAainLLPcbQ0+cKj/AcrAwvfTQQcr8sFPGHe6ynoREwrf0mAOi+Qqj7OnNXl
DAUmZPSt3HxDHFHcAIjskkUejNLTuouXckTgzhD1TFQPvNrfgy6QqQyuZWGDrQhOrj2/PERs83hE
LNIFqEtovNx/yB2Ggv12lTtXYeKn6PjiRQ/4xVh8e1YM2IELj8wCK2B3bXa4GSlQAiXP+iBFNP/j
tzuO8xuUrJFNgl3A10Lxrqehq/JkYy9H5xCIKABl3SopVel//pEzkYVvfU2/Un2YL+ezsgMAy1kj
BT8RW7RjU4ej+Pk/twYeHw/rEkCtk1qHQTE8eALH2EiNRzNUlapm5WtBW1r/99GhShai3HhwnWTB
N1zSn1NcmE80a2rQ7DfXKy/DnuGc8WAxldMAIba5RZ0VzzyMKp984a2a328mE1JQXgy57nEQvK9V
yHQm900RyOD/1Q8fe/6RN3OeIb0zA/Nckd1mRFzyRC1bTDg8Kt+CpaDzsLGCfhFYfhehKkg4gIVf
YkwWwpvodO88Mk2GRofTk+J2JG12QBv3rxXXhDAN8sOD7/sUHLxMALc2p4ttpIbnSb+bjf8un/ZP
ri5WVGdKqlAyKgTiLXarD587IYZF6I+sblqlYvCV3NgPCEl1Rm8urtEV9UFREuSyla94GRPKzheN
2j7ah2QAI9MVVKmPoxayFYCJm8fgPfCMAgtZddWUmDtpUX7JNgdhz958MysObJexOKQfRAFbT3gD
mKOZoPIYpHSlJ5L+uQJuU1UFaDq6YYsJ8qWNXJKAds1Y52wBoVLws2y03YM8/cm4gwvAUg1m3pxu
82CQsry511A/rbpouFX6gZbORKBT+mkK5UHLu9NbsACYXtI2eAS1BxuBFagLYTD79mjZMWFw8cGs
CTTwWHywwAOctKDT1VYITU6c24mOO5nV4agj1e4QrRnjsurEqTVm7RTNtcyTfJtLoy5jnUo+e6vM
OGOoHXL6vFoKaAEC8AieH+PBkxEPRUf7cwBtjgMrfw/c7m/NSL1hN2fixPA8Z1opShRDEt+vAAAp
Kn2GmfMITZzYAYJHFo1Yv2xnlB2MgJrU9ixfkt5RXPnpMFYYouMKX1iRMbttz2HIYMwu3vC9GRNZ
rrRZcATVgTOJ1nB2GAgh2rZEi84qTOkkXhTezeT3C7lgf3TV3yMDFgjlFbRJRWJpHzPD5JQj7vzh
q7nrTHIrZZBOMYCzRNCrsbCRg6F0JTJZr+RPYRdkcGl5gi9NzOxJaVAF0Lk2m0nqMx1mr+RY3gXJ
/84HvazUYDJ906yf+9rDPO808/NrQt1vRg8VTSfwm+w3/DizI0oen3X5VmXTMsRJ6ULdSim116Kf
PUabMRGoUj2Q40T0LGIYGiUHcCDIgdkmPlGqFqjs6VX84GPGmlthl7Srjc194yXejPi6gRMtf6QY
hrqF2WEPfgvZXm3Cwl1yOGh+I1oxKxpj8aTq1wTuoW8bnJWCjGww/01b7aUkuW97nyT0xW+W3EKl
N9X9HIoGg0Phbz1GcL7O51tPWGLQZEEQX1TZmRuinUlSK1bhZFCkYOi/cWUXrOkOl0jgbLY79YR1
5wXC8FQF8dkyGDX0DZhfEn7LrlQ8ZMOEKrQzxStJdmgLXzIVD4LIRwYW48bxIyyw2o43J/CRbov4
m5ryP5IdG1ls2ofKBiZ4KvBC/1MrCJtxcQX8srW/LJgT5LXCGwk+V1CbpmBOMJd8pVpGI/N+2K3V
ly8l8dN1y/ADvYa6ZIRk9zPNvVCWhkh360BEtmbSbIl+N2Y+3lFFmO+Vlzo4EHuDfARmHKT7Zu6L
jytto5CfWcH3OeoPoYaK5HGyVi5+5Ta+y5T8ITg6rgMv3R3ZR1TytAdS1abif/TQm+IRRerIRPuZ
MADfOQVG9JD4oPo52w0LMDk1BveuHDTkQr5eV4WEMwJREcbwhUa3B68fgIdvLtn1hMYks5v1/R0U
6LUwtcUV48ozVDKi/IfH6472O6Scxhd5Od0XDAgZc0bD1hxIVNqGIXsufNlZX3a/udfADgAPNSdt
FTpJNQ9ZwtbYffERlzWsYe9F+SSYPLNzWh/mjOWvMq0jCLQkeGVJEAARWr0sk6vvxUbJXCKlkjei
+j82UTmrRT7Q9ku9ujSO7nZxSOynRpaqwIT+SfEkrs7Ckrbz+ETDmom1+P2b6MTeEyexumWnML13
zYvIou5R0aDjzfCzagjZfnxAFo6WhPIrAPlC+lNviEkUM6MJlWPd8mWiudENvXppGF5bOUGV4zrf
3AWHDG/qWcMvcEfpJ8aejQUlTniQ6lNaGbBr6c1sVxEISSXGjj7iXbX7C2xRSaG7NaH//gVYEMZ5
tX4PiL9UgGy55S6XO8PDP2c1DH0qSwgsfnIG3I+eqti4RL3nCUjsCn+3KrF5g6sunEdMQ51B0DOu
eOHWtPu1S5exc0P/UMh7iZtC1MSDWkaLucGN0XvdY1Wg4WFBthkpq6UA2obVWTx4XxUeqE6e0AXF
zX+JWMmhnU4oH7IDjmV/7dYeTZpA06eNS7qRv3/TdMIezdBovKurgqrYjcKO4QL42pDBXT5WiOFq
4vHg5Jn61gFrBk5IDDPORRdyxNvZsblphZBoWxowr7ipzcg+KoA4OYnuDE1JFuawKSViRTvv1Ruh
NHceO1RI7tsH62M2iRfRwExpgsJFuVi8npC0lAXMkYviRA783lT/yI6VDBOfrbOUbeLtAGuiOBVo
65y9bZp3V/MBpwZY4SkusyraNhdYi2Uc2Wi3vIwFGTdmEoH5OHw2NGG5KWJESjCQ/cHTySmfmNE6
Nbx+ZIKnI11F78GGF38knWkqv0bK9eF9HMZk2WtKdne6LToJYdm60JSq7uadxi20eA+jWEtTWwNn
lUAbbrl2EG/FsfpW2efKaWT4L1xRDSxDGXUuC7i6RU6JMMF4raSTW6+P620fOC5pUj/562iJAki0
UX/zek5+U9lI6v23yKcwE5pXOpO2DGeccXifHq3j1mYOJVp7xvdajfnuuQY6XIxSlQ32ZRca3At3
rKMYnCYVGFIvpTgEIhmDsvI9Y3J8bOpQvBfGbUROiVYZjegqSKb5rN5Ix3XIe2KRePGdFd7f3vuG
4uCHne7eGjTS8Pkl28UKVJTBBJ80xfqqnLL+NTu2TFZn2Mpb8lVn9S8ve2peX6WFVxG5Bp2LcDsK
7FVl1Pub/IniQ/GQf96OYV54KCrs0hOiTTH+9/MeMgVCIwv6CdW7ZNYQ2coEyOQvdUUivnauvR0L
uPn6wYbcMrabrhtT/ofEqr0f4UiVhMmdXfT0exRzI5YJjHjgzChkxEcXRWk3ns2vEWUZB8esObc6
b5qlJ6wh2v3+A/IO/+9qwuheToOg8NGqw0Jg9OKIWFJHC6MUMGlrFsr+lke/pwuRFY7xBXWmg+91
rYzumFqK6uFRwRdGoxB1hE2LLjdgFItX8nfSRKNjHkV9gFvwEAp1lda7aPXaovpJplRLumpE5HPZ
HgbW8LCrdNfzg5AO1OxCiAFX4hle1PPpEw7OYt2ncRKs7nDjP0+wop2FPNJqojYhTmYQCteY+xIQ
t839Ks/b7YyTXXzRxoerbUgVo23A3JlBZMZ4tu/jjTaV/uc29ZxaijDsw655aEpvuJDgTusBG+gS
VxQSQgPM+pmGRhTH9tf41MLazhTKXpCRyzHZTIibByRxfTXFdfGpNOGLaZkRkM+dotrwpUBu2ov+
zoCnDSfEk1pX76VziqcytN41m7biFvPgf8HBSdfEaWGD+FeRq545eKW+6KHYlfUf3TEbm8mCFNOe
9G2qQsVci/zfJ37y3dbo842QNmYD6miHoJhG+xMcSv0Q4gSzCofDepf2T7jTqIIc0/TvN1cT4ct5
PJo0Df+udlfTo4VATRB/8M5T3vE/uXaWnJ2gHco3biwzIswp+XR6AZpZuIw7z7SOPBPJV3Hr65Tl
UgcOJ+7z3Cpglq3RIl34qi+bsHvG8AywxA4IAqd7Yo9QM6quBpGDBT/bKLwnJu+d679A7LbR4fNq
t4XKJhWfhbGyxXRzOWf6OObz6FRDTYZE9x4hOMwpOCOcP5mB9NaWDP6seG89sMMDVApkWwWKpCXr
NpdrfCSnupjv9XhB0UC8MN43x+NaVDGS0zldjhRjlBGMjCZWb0u5lZuyPBAgcLoa0Tj/nBJE0IHF
bxto4IPwEiGLXvLxKyJdYnytNdnp3Qi4QcJCoscYechBm+wNCiAGMrenq2tk0Ocsc0HfoBXse9KT
L9FLlYa2mWxhx+/GuszvXd/yN3e9PMDZ69eXybWL+hvecQepq4TfuAP7i0DqOKqYy+1WmtljQMLR
WE+Ys/DkyUXAG1zGg9kxvcEoeu4hvsPON6sLxf6Cw/BDmLLQegPlHKQXhLIVDVNWJwXJWy4O7IAI
cE7TrMYZ1ty/PNRzSeTbuhorX86havS2HiYulf0IjrBTG+d+MuDadk4tp1v/qEC8DRqfpEdbwQfa
1AwvBt8t5CtCoCd4SGDapO/EwnWahDkIsgUKsbcjz3ivAOTMmtkmK7E+kEOlXOhFayowl1pYjtfp
4AOGzy7Ola87Coj1yejTxYap/07wTchwusICUb9P4VB+SdcbmDj3od5dktuff3+J4ILIDngRcJVV
/OZR9AjaQPwSOIxARqqfxDzN1StvtKOVQRLhPTWcEjvJmTWctjbCHSE05/r4RNgBnTc2dWme6VKW
7j5zyh7TIR/tG3HGCc+taNzXX3IKrazzMvPFJRUSXsv2VaRr6Am8la1Y0JeHGvpPs6VCDi3jgXwB
dBENqskUU12hrakkNYhvwFbjYFA6JxsbRTtVQNzZ2StbsyYU5bzJcN1V8FGjNduGhUWnnNQUBA4p
HVKuV772nV0Ktl8GW8B5ubTGaL3VIdj4L5j3rn54MTDTrn/0dbJRjA2V87VDV85GIa/YWhir4rdA
a1LWUaHLLduHC9Z5dE0eElIp8DrJQ6J9pFFtOPp4sEaV01CBUPmGcouKWeGfF1kONtJ+vKZqz2J6
/3bjXfRRxBi/WjWPFbtGi6/Bpkr0DyIjWLcuQTpUimo8EfZkxDICQVGMJcDuE6O7Eaj8O75oxlMC
un3w7wYUCFP2TdAD2Av7oOpyDsGyvCYexnJaPj5m89l6DBUn6mK3t6jxHEOl1a5x9EyT5Y3m5MpC
/GVguQasoSXNCpPkE0MoGwIkHTeFda5rfcLBLORun6n12fNMGoYtFru36I5tDK2+kNrrem48ZqQh
NEZxdzxwHP7K5ZoGjO2a5UJFGo7yuPtrPYiS75X5tsIonNO0+e3QEhK8AUP7iwE5OmujdnnPvuCZ
qyRjjzZYP+z4vTJzVVJQMEJ7b6pp3h/GjpL45L9PmmACXbEgo9uD+bUG4V6RQxpxmLSZudNUsWMv
azBsHGmy3krukm0z7rijSSBDpTeseHzeI4kKPH/zqehywNlx3tuvUbpGRkPEF6OAKzg0RgXjpExm
MJKRGGNARstbUZ6wXU2vAOHiv2MIiS6V8EUhcGAZ92B9ft81OM0fn9O7Il1Y8Xr+cJve1xjs2FM4
KpQNO2f1G2TNVqexYWo3rxPQosUyiceP3tYR3JRl3iAoYuMJnZ27tUQXtBumI4cObxoExjs+vGv/
fDgoN8G8AyF3c8x+0wi3vBWvD7UrND8y1yyFKHSkX+2xiPhboaKsMpeO3whU5xSknQokpUq7Uoeq
vlXgUk83bsGoq3uMoGIg1c8CGLrOcnfdA7HpnIUvNWYcvjz/qJyTrxAeo3HXwdQ+x9qXiCMSz/5/
P9FZvfNzadaw2L6qNi48Kb/TbEUUFbQOijwqb1MIphg/eOyAPwwPbowSLZaVCsAVvRAcusXK/ypQ
UF1bCF6BG387o5vssprt4uHrKP5JFVdhZ5aoHYyDJGQXVvZPiCh4hJgHQSHHi8Nd79dS40uJuWOZ
L/wcwC6sXe8qG1eni5ZkcatLuArTo1ZgzRS9kcAEecHuXSJ933fqZF/i9a3SiBPwsr9UB76D24yp
yV6sHrMvEtpmjlMD9XOaDPtBdC+wtyPg/ax7/7aRpGIvdM1DD1Kyq0MSRyjMzmmRBXFzEeT6ZycV
D/TiARfd8ZDFfmCt271txvBVDirJalU8Ocnq9Jtsz8r+uQ6myt5Czu/h/jkPLUah5L7wdsqnugTN
2LtutA9nChCmGLiRdnUwR6lKG0tsvIoNsHFaBox24Oh5eVr1YpU6lfhmZFNmo+WTmPRaAXEvG7ZN
FAAwoucvR3g4oXvpWPeGvdClEUXizZs6EY3CAvKiVKtWEoR/OO3ATjxM/gMusg+grjkyv8OVk7mz
dyh3rAYOKEw5WIAcUkqePfHTKQx9hg6HA0d2G5Eoc0vkafhvm6yCAgBQfk4rDZ1AepnlSl8x0dkt
JRHFjpHZcZ0WWll2vXnGtbBpya+6tpHP8dIW6evOfCGDLo1sWry/bEzGlhXLU/lfZHZfEXtsPjbZ
8m6G9gH0tLdAZUQjxMq0kMZx39bK+51MYfWePmNKMqqMAtL/US3n7OOL2TqrMI9Bi3ZBfnjmzCQW
jhES0/7mnQAvVgMk5PgV/OsAZUKIdj2qvcH52sXG83twim1smMOziVeZKJmU57WkG4V8f+NOw9HP
xYVnoQJS9iMp5rBult55Ws3wvuVWL5ADCG4R8xb5ZiCr0cN4QNv6TRLsVNqoZN7UJERVVwhXygpJ
rFMveD9+zUof98dnkBB5JH2Sibh0UdFbSGWy2RR9LHAYUOPiU3pX83DtN+6OAqCf1bRDii30A2qR
Hc0FlaATLZ7f40P8rJ8lzSrl3ywLz92IgQxeCIbf5YRvAeNtHnMDCwETxWHzjiJ2MidzU4paqGyq
4LRjWKYutqxYEVJgL6ezwAIncUzKtxnXYxmNnN0U7OxLxxyQD8FHAzj5PSo2vxD2zkr63a/4fRUl
uGvkamv+S8udwFxNLv+8KTWTB6a/rRdE39xngg1YPLLtRal3vXLEER36iFZmQcv0dsXUQm4+vHN6
SiYq9Y/UWBeKbge+CAq7uOTy0RCqr9eTpnustdiRF1qbPzEg/5sHmDrQe9wB+1aRJBc8Oe/mv2vL
mVqk9vPMpz3Qm+S8DxHpcCQQyCV8A/JTcMfNNwFfhv02E/1BFC54+sRt2dICaMszDiRq4SaJYeB8
E9JS2MKa/04+thrRmvQPith30dBnuPo53ezqco1RM7cRR5UKf8LusTJdcThMQVd2vQ6GG579ri0Z
tc/SJsdwcrtgB/xLHDlgw8mcQFXGtVLCGQ2AhD92wvzoRvvheQQ8hWWauyPCmYyZk59TJ8aS/nz1
fTk06ul7j4RV94FLxT0hluMIXNQE8fGu+zcHzA1uZe4W0cy6RXqk80eYOB45GdKmOSR4h3EcqH1i
l8EVrYZdBmNHg9zqMZlrkMs59tngnS0IEVD5842pPsiVicaiyjAzwCytDxDgtKBuLm3bmxEgqUJk
xjE7p6un62SnZvmohAjyOdl4f5hniCf/aS4xoVqIzeeaIB7gW8SAb4FJazWOiXiG9aMgdlYO2ECr
1olf626zYYFdaUqS8XzpaEUrtazIKg+r2Xiw2NGykVSyL2PoaXzGMyyI4kq+E/Hc8as5XM/jeZwb
rKhmfge+qacxhZTJoLE1FpYjJKJ4PwaiRjCQVKq9WPfQm3V7z+1XeTd7O4meXwURK4c7yj9xO9L6
LBsa/DmeOsdUzjNOHR1TBMI9KOUX3UlW2FQ683vcy+glXWWTNBxaqVCW7zqrJlxqSKj+aM3yZ2wF
SoOM1+EqDuJKCBbvDrqm2kllGAOAWUBfofVsL89eiNTZIzHcEIGRUTMQ65uwr7HvPb6ibrgK6t/o
2l8hu+Li+3CUD99gGYt+ru0CZZltw46/VLQrHuCEcKtyKdA/hubQBQyLR4smzcVJLWPVeyhsR126
tEIcriRBDl9K4hvpaTWHvkwCK397QQCUHDQVEKXvsLJ3s63n/3/myXvGZfAS/kklxqUipKbPmZNn
2b3NwhMi1Ev8RZ3nidCFnL9FyOuNoC+7yGrHTz5mtSdPmj9ZRGmBZ31/MGE/qQkM08jTvfb1YNgv
PtnVSq7qJWcxaDesmq96e74KYQ0lMlEhYcCkoi+p8GDjOj9G/K9GVBh70IHKLXofr1zNr8KHec+g
zuA6ws/IXy2G8zFt2DKa2PMYQu3y6lASZEswBPycR2k7ftHbzkpdZ0n2oTBKB9dWSZKrO/Wi3O0Q
tK6oOznJ70KyNvVWRgfXCHziG6y6TFEmBrp2Iv9vhCO+0FaIn9SGJDUhrP2+NRvcbYOXa9BWLSqA
+qSmbHYtDYDoRgvKcjYfM6Cm+KHqRts4V2xsRwQHZ3jw2XEq/QYmmRPxFYFizGQOD3cyOGt7N9ee
qx0T/W4GSXu5CcV7sPdRq2KNUAuuuj0ubVkrLBghs1rxLuO8zFo42kuBGY92Njrhm+j7hnHL+B/W
st+eVosNpQWiiJY0wkEur0PUhXmGCYUe1o9Fzs7+4ckm4By+mAUUGzw1T6ukZDKIJp5ldjGck04Q
UZTQ5++X8pAlZkXavR2d41VGB+FuU7oTiH/ra/uhkaNkqeM8yM46cZd2lBzIo+pkfzXExh9aKlu8
8yJTGOg2oe1x/0Gr75zvTZ0F02EOKWXUtD6WSCMYaD/NXUfHRk/VzhBvlBdpmkY8Fqvn5pkqQVdx
S96ojSfZx3fnv7gQqRbaROdhIZ+V+rVXvi76Gr8IMwyLTvlPdxVu6IuzP6rKnAybdvrXFDZmiig6
SUE5c3gOwPPMpemFB0rDvep5PIiu01ZnUXYyyfASSizcaGnd6o4kiLaBKNE05Gfae5jLRVf381jV
QHU4+pkrwvODM8WcS26O46roATSUd1U5KmoXRoOMCtsVGVAP6sXUP795174ZlsTvAWfwIjDfJssv
WPLfUPwQoD3ipIbbO2ED1VBOQJoQKNTrYG4bTZseyq9cWvzeM2wlcIALvRVpujqC5liY9zaSm8CG
JE8Cm4PY8FVd3MIpeaVndxTbKZMachUArZsxKLDgvZmNXhRANPKic3E4IrIwhbkZaGWlTkHMDBij
UHD+1cqGYoU27cvnYsDqRLcxbkuSlVXe6jY6jpoJsm8xDh4FYfCjjKdZTDfNYkF4WGphNEbtO5p8
HXBPm6eioFQBEK95dgkwG8Rr52AIOJcKGgSIaS1eeOB8rxzk0xUT/NibhOPysGJa1PTTZ91/Hhih
8MbU7/OkOEWkWBtd6vpQHhItPnYjKQ/5yY5vMJqP5/Gl/srHyOzhwpXAEGb4bpfGXcofyZmZOqZF
/89dy68tw7hAAb9DL9oihmAzCFZRAHTeLIRleh5JF5LCE3fAHrrbqEgGVP/bN5TXSXCDwRli5X5f
4rsP71nYWlviMbWf3XKKgHYsI3u0HlFXc2U9ktVm2bOK36uGraVRhDlJYZtCchd5/bi8gWnQwPUK
XLiP5ZgW2JsLrVZbcOER0FyjGpean0ZfSNVfa0Bu8azIgL6hbdDC+7otJYqi2uL15zho1mu0vf4n
SZ/RX+GoUxfVtaWGy7ccKHvu4HcY6kIg8mqZCT2FXfVydtZvs8iOkPjcGEAkyokPFI7IzX4tRot4
kL+FtSsCy0D6q3Sz3LbmUlAO5YrTyXLfPI589d9whYu+isVQq31aFaUuL1YeUJ9MQM+6gMovkiIM
Sf/KEhq8VfiqBeoaeCB8yRSJHRDtdbI98NcKvOql1Bulue2liG4Uhk3a6h51uuWKTkzTBRVGB1HM
yQLHHCb5Zmj0fenIz3N9rAKtCakbYNU1TyCGRDhAQl9rTSqowQ8TQTWBHrm9QQWWzqtrSVDCoh7G
HX9Bcd9SgX9APtrD8nX2fDiJd0ONiD8khUeUFifwRDGJ2jfNB2SQiiUsdQfq+R6RE5cbIMPyU1qK
HcCWLyFM+JIBaYk1BsmbOFE66J+gK/tW3epjsAQzb2Dzozx3vVN48LN0z0fbDbCI6B5HrF/BneSN
s2itULO4HV8u+rE5kDjT+bGcvvWgCR8rEbZW1XJdJsL9IfY97vLdKZXSnQlyFutiU0bBB78eJe9L
QTp93X7nUPOulGKXBWZqxq+27DCj3cPt2Nui1sSZAT3Orsno+fZBqtSlGg+I/SScUST9rXC8DPTo
27uEX30TiAmPrLrsV+v6gQqYduaRzrVwP0GFLVTATvQw//B5SCD6EEMmgB74czMwICRVkwFnhSD8
lSD/2vh6DTHRqiLDyO/1xQZ68dvpneULhs9DRdpmKFp1s3QIycR+tvgBgG3w4doPepYF9iSzkT/7
NivEyfsg6RMnRLtHfEzTKDQFY7kohdkEYKd6at8iLxTtR0Ob1TqE+yMFXuWWMtL1qBQ5Dj7BT6BA
2gjaO5XERtotswIi11kD2ORhNNGDGa6MJ6aFKtsozivcZtPG/W0ZesdYur9bwOulkv7M5tg2YS3p
VJE7ujO3k/CdY1eRtI0iFEcR5cR7MsVuQ+Z3yWN3kmAjfMLjQE+lmDYApE7EziVasRt4bBUZSJts
7WXFL6AQ3Ejw/a+IpnsGQy5IXkGb0z1qyUjKNWJjp4M17c/o2w7ikoOJ2HqLVx94iRp52jz29Ic9
jEtkxMHIXIs9e+aUcqjgCNjEOHPfpnfuaRFr1rggTihL5v7CeHNo9PWGpidKTdqEnJOjiJfv/Wcs
8ejkX0kDFDBh3Nxq8fWV6uOdMcovm/vOVGv4FbjjjfcTDu9VhNEiXJWz/Gy2SQOu5m1ycy0Th+gx
uFcaQ04dH1ufu+q4iF+79Of7qkd7kl0YBJJ9eiddJnPsyjQaOivvb19LdXRvmJ59zTGIdRvD0pZs
XOYp00qWxEK04hzkbOeHZaECwdgebGRyF3Lm6iSoC2ZTiurOXNKOaqfR1ssqyB390ciaGqjcthJg
1fGljKSudjDTf3pgBu5XQsjIXl+OdpexLXAyCBfkbIpvzzDyipm3/rW8phOxAuc0niSdQa8/VPR6
dhdZ1gmEZmTrdc16z2mU3dEGT7MelhKnF6fGb0z6TqPNaAEtKwLU/EyjoHIEkxu+0Rw/H1B+hBkh
K95ea22lkuGX2FBdWQV7Fu2wnIWlMhLUI4phvSLgKUqvmR7Ls/hfTawlcnZDarKZcYtiAKVUqLc6
EuCeUScD+LAItFQ+zmTk5fk4Ij8ItwCLsUVboZ4S6n1QH5bo+Ls43rrwmBqK4mHUjtSF5Rvp/pkB
l1wzufnQVlRcPmX70wBp4sF5azMJXi7TraWfNbuIFSblCDTuYsjLZGYqDK5rZIuNTIi7c1LIRUvV
2NA5y7ImUYIDIytMFUXlTgZ9X0ot72AGwnKd37utY60+k8lUC+iDJ6VNWPvLMmChMzOm81kYR9QL
PikDbu9xKlq4qANWI4vMExVnCjdM4A3jcr04UwkVwNBn6Z3rErB1KtFw+sB/UUoaK5BqOAnX+mg4
rQHcg9Jn5UsSmS5nq2qLFlDtg1NORfdN8LwHvHL6YhjFQ84H/AuoWPVZu4fmiHKJr9h3FlPm2Uya
W4s55sF6SBzJoQpKfuEywC09NT/jAULlrWTr7Z+B4BL9k3xP0edPnMovpveDl4BiALri+uWnPz99
YWoJCUuslbbMYlf+v5lZxfZdNw10VtfSNxD452pB0ngGkldq7c6FbbY9MyElmbYryFIuS9zVnoR8
cliPnjvhHkYKKwfqfxWIEpZmbuJSnMkVoCrFuytGIAoV3GrnUCTlJHA4cVarTaccXIfu5TXIVDwM
Vpg1VlbykwmLegVJ+TNFegijibDyeQSFz0HwY16J6+JhkZpzMK0ElVzWQGl2zzidyLAGWen/UBfV
2i/7QvX8i63MzznTtf6TGv/GSy65DBvb+Zf/XvuX/v8wlGgkbGXVwHMAawyauIpkIu/+4wYKwS/R
uaV+2TH1MmWedxxIpoV+VHgzgFKPAwMpsWIegpkCk8QZHVrhW2L7bDJeC7DFJfQLg0qQBs9Csuxs
34Bb/yoWW22LbxVoTC4iIvOsoRlHtS6+jAk4W4aUYKaCt3zR/vRhTKy8QKrRs0q2WM+20j956n2+
72uHeBAIiwPtVbKQZMhKQDBbp4Bo0ZVmlcsaQjsBiMV41YsMMwT2+NimSsFHDpl/zm8SUm+VUnB7
ZrQlG6HgnLKF7m5be+RfNWFQjNsuWBoI9DuMl6GLNz4ZOAIkyWWVUkWqgR0lZk4ZRbY8Re9XL38e
qeSJdRmjcXnYq8aHYc3kFLZpwmcugTMLyAV1USj0K935eL/z8hFRB1Kfwe0Bhlu6azRTf4mhj5kx
IcIf6kXgn33W628+afXK285sVp080A8H8E0wnuaP5WB1uMtiH9Uaxy6HmPqZ6aJ6eeOOc00bE2Sa
tm9GgD+OnETdxE2ji0TJFpugI0mX4N92LQEZB5Y/YEShgqOqIMfkZYBHJN8YF113a1jH+rUEBl6P
GeDWdo/8IIJDjCRN/DtAhRXixQuQ+NSw816cBEF0EoOa15MC+SkkIfRLTWWqLeEbUWq3Gz4kgPGc
VUb34xlUhGTqp6vqNL6eGQOAVfwQ9QR895cmsgQ9SAAlfBaQapZqA3d1Qc3cWbA9ySec4CRIHTjR
M7AYZ+zXHlP9jowMGhBE+qZjoxavxNaNJMwWPGeqgRD8IvQgO75VMykhy3x4zgSG5NOdV2vWd2Fj
BbEQMGbKWaXWrMQZ2BCl5GdPbLolV7X9EK7rpoe72GJIVHwL4ToBIglTBCcnBs1LOYNqAEXCl0e1
30vLQBWtoGKfEQAirKHR5erKhnP6+v1r/XzmE8PnNsTTTb9ncmgJS6fQ3zRb6yu+z2jM66091mXM
+wUU5QyhTdYMSS1GQCIekTcV8vDHfmrIS5wWRgbH49FOY+mAEB2jUkXsXc+VPtHjRykuxnWQO78l
ocn9EscXTlIj+p353kehyDxe6iUVCjaujFSprvoEWbNDluEB+QO1MmSvy1ILZ90xhRVEebwb9QmC
objrHDIK7GEsr/RJhh5AZ+oEMMTyJTnZ9qec4aNRDcuyj/vlfkBx0xFm6tkrufww+O+YN47j2fAj
Ki77JYkmJBz7ECihrMkQqQ+sADpUFo4LJh8Z3bKqI7ysq99fM6AZcQOMMVp9SnPh4onxptWyGy6V
kcBsJXoBmGL19T3HSVCkuvxnSUsu8omu5KyOMSbGuoOKx3G6mhQ6QKZO7kESyFMhQ1wPSLyM0Qhm
vOk388sujNx77AV00F5T1YuhRBi5Q+84PHus02TDEPihx5qSYS2F/9eH+82iFBgojm9SeRoa5041
oHP4msiFQfpZqVc6S8uALN45AO+OquokYBAZwIrARf0753ITjGJufwZEryaoRry3v0jofdHnjOpw
pLQr3vQGvInONIjPJwFzKSdLKDqJxKv8ZNuNtR/I5Xttgjl7sJDD+Ob1g1J2zRTysEYQhSjGojxq
I6gQ+t5N45l9Ss3QnjXLbZmlOe0Hs+YjS4tpdjrHa7lL95TxaPSE6cwZ/zR47EYiLRiMxxdBfoRn
bQ97h6YPEqB6ljGzEswtqCv0jLoX6T8bSQtIghkJoMoS24w+fWfTMndayik+H/6meH+rowlYbS92
Dl3At8PI0XdT7HGeSrrsHLXOeuhsTnPlijGJv71uPtb3ZBZQ46N+l5HevaBdmjQPBQngvmFr0pKi
lXlovdcuvcGSNlqx2jJBpscF113Jr1edoOJ0ie1b2NSVjiGS/Xcym7N0ea0rpKgFgvOQGySBjnjv
WkLRyoZzY1rc4psHi4jblpfvMuMzAj9KOi5+PJ7sMWy6GRtAx69zkClj9Ars9T2zYMscRdimf3qq
4Bj+Zr1pDHdIRh+8bwwZn1fbNe+w+xPfHXT+tdBhICRF5mE/XL3zZLTRsUrFCq70JQEsfy5PdAbv
ifEdJPEDB7Jdg+0Gznbij5GeSeMLY47vn7cU8qMqif1oNeSUK27L3U4v/9eBizOM2TiloDDI5JPC
FznL03aQOPo1QZ1WLOs0PJTeiTSPzjSQYcSN8BstM8bX/mwgPCtVIsVSvMg1d0AnvB81uYxpK/X0
zda3dvsMNyfRkGMwImaOJ/NK3MsjT1loXH2VGxkrbe5kaKLPtHJmyFXOfqL4ItLw6+B4BtiyCJhk
MCtn8Tcjmn57bv/VZjW6nZHEwIT42lIrft/5r1hcUNLFMy9kC/xwAqQpjKzVw7atJzc4fmcuQ3sl
Epx0ce7WLX8zuvOp81luB3tKvQ3XMOeOrETiYu1Mx3NfWcVes7a8I8ltPDglavxxyfNaUHuqUKpa
xo0dhDOfzdQR1XS9eGFP8zrhbF2cqVAhnjJT3vLjS137bvkBzCSxtNm27pukjlI/BH1A1+AzkfRG
zrLVw91dkgaMJs0bcLzpyUZpNphROICG1rVGsUbVcAeiO3x1mtX7Ake+0suw2twkXEv+DNK5gY1m
aZuxV7Sx237uwCXAFgGgnpQ5ZOKynBHVay8VKwqFY4jecEHZvMILCWGoLPmCQ/LCPSb4PmSGGGWo
26kyI8fe6Vk73WPKKn9uLWhHO0Vjad4V/u8caqXg0KzCPPe1qA72dyB5XNlhWHTc1kijdeXWFt80
qyHxC4aYouyN0bTwF9c7J06qKyfXMizJYmNetDx1HBq1yma956TNlD8kvMQfvygHD7tlV1xGNVCM
uz6WuR398bpv3MdjYxdXVHvksyF6ztxTlnRWBnU/7o4ejwcLEjdaCoHghjKu06a2Oked44IWw9rr
LXHc/u7xnNOovwgVUEhaqWldHkwTiBVIyn1s5oPhtoOyQ4xkt1LD+C89j7tp+QferBFwhjDfPuGO
/fSW0aimh0cg+4emUkV1naJdfBfXv0iov/fU6ARBqSwTHTOk2pXKPOk8JY4tFtZmFCAYpqkeguRQ
iJTh00Ra4qQyknXqlF/XngSWHjCo+wRK3B5D91QxDvac1vo1RdrraQuIvTnNVMWkqeobymINTO+n
xTkNPT+SsgMuuCBNMu+wCI0vF12Qk0ke1vcDeszZUobO7BdQ5S+/jmS/qeWaqP7wgIdgbFkgmE7j
c0xbPFzk/7WT9Tw33RCm/oPKVfNX68/Dv/TTtyIr71hJ0NqqBFzmrBtkLrL0JM6dFrzzcyz1PZFo
YOhWjEGDPluZzLXa/SQ7tsteF0/D2LLNeHh3KLPju2Z/ZoLADB8OKsJ0jCsnQmC1Lri2+qf84Edx
fzed+lkxhiGfQX2jSbr/a/l7VsGHRzuTIQYANWQoCLRRaeDhHZpSTIerWoCcu6Itkob4hcYJybjx
zKFyapqPZf6PwBHeH8KF+4JMs8SWWSP8COJG2gvMphAiZ7HdS6Z5sqs8x29IuaHMoc1jOQaleaya
aX9/31s94qbN1K1ABlmBzkWoLfexrTYC3Hqk8pIdTeAo+moIkB0mQk4ovoMsLXcSxEMtwFELeOad
fT4RxLfTWBINYr3U/qTcWeQsjGtc8VDTZc94734Km6iFwZ8ImYdGBbd0PsbU/x1rmFljvBOlKqnf
HlBZ+nfVISeUGyGPKQAJJy5aHPEWjp5UOpWwiIRjefxXG7kdQMS5oNYbjauVX5lTQQo3mAEf3ODg
kt1rgqipRedbj+sZQM7ahEDZU5Fl/HpTSZugi0USlJz+XjnvLrOoZOZAMBD69nKSsd9eNddGAH8R
DJZzQcp/dOs68ArgqH82loKX+YerHKD9a+9K1MvhzxQh+PhstdDRxjkuRxxKFrw+e+Cb6dZ+iwLk
RnlKpb5YNGMQAVgPxGizqjsvN+OOaM/EzVPlPn/pt03OpNzxh312FoObcElRXRYYN9f1CwIOOArz
/uFxPRcDz2DgJeJ090ZFsXRbr/zX9JhaPAeFMVXSj37x51Eaidit+nk+nmhsFNY+ZCkqBFKjQkkX
27ox0i6xy1KIoBl+HdXTWa3WvomiXOtfgnq5V794ChCGrsorbeJxcKoCoTv1mKZnaiPbVly6bGHw
Z/1ckJVvQ35bFBAIdgK3a90zfiT8BqSQZKyR3wBksMaL8J+hsbk7uWuZexiLzJBu7DULElIxI1kn
1PuYLLVXHeHa+RTC9Bs7QrSHXSf9HPpFmLRwzkshqCDvc3X0hqBMr1u7Fmu3Uk2Rivu2hqSvvJcb
QirtQe2C+vB92Aba0ediKPNUwYOgFVNiS5UssNSme5FXvqXl0kWIpetRTuxFeDHtoa6u5E3CTTbF
RPwEr4B7rHawb5dKYykktP56jZFFUYmsqK/5Ba8onk1O9cpP0cGpjzQjCyczcTqOVmAHaHoTxAbU
5P1NiJ8sI2DoS4ALuSwawLDcxrakjNt8OA13OVEl0naRF6ZcyQvp/IodE4WhWkzCii/fkOoJR5mp
UhPoZclu8PkJ2fWj+SX2h6IDBmRAPH3YTsVpbwcV4Axma2QExPbwkzzITMTzyZXAF9/TAgfo/rqv
ag/VWid3yIQ8fpebHoRc5JqKNdb085GW4Xn3h3pVaQL/ZYlMmqgxTB35xj0BGurmTU/vjoSgRS2G
jhZfDKmbBKzydb09XiJHRzLdU6rW6gvAooM8+jOwz9cgHTa2FVLfEnJqMNtujiTi7zLv0q3cvjcx
hlZVEASgjZSC07ORpvmQqkueGp6fxsjQe4zrzBxDLFfuaXoLZvOU+hgvTqufAOtA1j0LTHP1zZSP
LPPnLmO17leNGx9X8NaVSIa1VWEMvW4EjtSipCuPctNirVr/y1Fzi/la3FiKT2CzdqrmlXG8+T32
+j9IVQGPCebAUP1z+E4EYFjXRuaE8wbGEkR67Wwexd1rgW9mv2cPzpcTGkhtYeQ4UquzDoFpD6CH
/T8c4bYY5rB2WwEvS9UIdDLZaGa3pftzNk59q/DNZo1yylWXrH9AMCp/UU17U5qcBXLixDfjBK9y
NUNMIX23rBt808y9vfu80LHfin1CbYC1e43ZzSVLYcyzFcp/9FAnqqJxp0cJsslemdbQqLM2Zv6f
AaXgbvUhg93onJua7LVTbJR02Y7JNVA5zRRMUDZymvN/6LdEBDnKcVeu4yYR6Z55jZqvTIW3VO9T
ZpkSEnKfFsuoddTqtR+i473i6tgymAwRF2QvLC1/e0Y328v1l3eC8SYJU5wGDZ0q4fS178auP/M6
m41am8p0ku6TBYYMH5vewUZK0dni/27F8vMEHVreD2ZW40NCdSEFTwe9Y8Nz/DRM/5/ViG2SObFK
15wnxA5SKLX4dNaFtjwkd7tNgd6zKRsnXLbexy820RSEJJEZcPoicN3Rhh/c2oJJ0F7uIOe7IDi/
9VU7gWnx1vDB5JGJQXcUyYXGWhh+wG5qekZypDedhthzebPyiRlQVi10XdO4xRBruLjaFl+K7FJq
8x+bTX5Gx+q45FXtYjL8LfZ1eZiUCGddVehwp6phQBtVUjN3gJxXFNqPYtQ050FHReloW9yhilP+
XAcaeI13HZ9Vx7lXiuUb0iZIkyR8H84WygDrqGIM2RzyrFj2/edYoDN6kJ8jp68kXcTh2bQMaEMO
37qt6xxNP4ME6Q4x98MnVVsX5fw+XTqDnvt7JvXTrzZlnkl53df+VFw6x5iveVcak5Bh/G0sh0V9
PGchY9/MB8JNMjBGppdqbKGNceedg9hpp1jAD3LJQvglDUkkbDuYWZc4Ufykybzm1Y9D7BLIxwBW
m5dWcYdf7iJpA4zqsiIrRfjkxYAP2ZtGqpPcx5gEOt2AGsUwkjESL0TfMxKgmJjl4poGCQRbGxrD
poc78Jxyorl/mXZPo1/sDCm3+erucxjyaJk8MnD6azMHDuUxcXYEPpX7f7/PIpIzlseuFa/NEikz
VW4B1BgBY+dLWMJF4Kpx6t+nZ4cgxWjHCc4n0ZY1wfQ0It0dMeQLYbjI5aY2dliCgHNu9plvaGjA
u1j/WFoTenO9Xcvw2AnSN+p7kmVYRGk9aFULUH7hy8VP24glxC8TQ2XDHQ3O47/QML/tnwjsxEHb
8CK0t4TPUQq7pvaUXpFAo2n98i22Rr6BuXrmydGYnK2kmcdshsVV4hUUrkIc3Ylgp6OarxA0oSox
0GI3BFHfWtLkJS2ybwzLLyAgXTX9DmGUbWQumieqn3E8qfnDDIiQTqTGbZJfaoG9GwU2yU6Ao2Jw
8BzfMG9+iGA70FcMWmqsHlIFFpURMHn4j38ltKT9NWi9SShj6P18axUEeVf6MjN3VnCxCBdvhVwE
WYl4rvV4n809Se1hzVoHfpP650ZCDioYY6SH6MzgObitIpshA8oNFOHEmaRLRFjjGJ8fy5TIHGsP
aFe8viGRcyWhxehhDHoAv9koXPMdARvxCePLxmL5yu0MYgsav+Gtcr9C5mKJMB86AUZJNZ/FiYD8
jcLbEAkR62qN+qTSjv314P1z0qFYtuinmKps61OlPS3lTp14uGis6gxkvmZfHPH/lMJW/ZA1Ej5K
sPsTVOe7pcdTsr0OaLjjjPnTinjNS/CoGqo5SO1bY8GhkGPZ+iPO2wR2nVIL0C1XohrcXtdfSiAW
iIbDeg8GiXVm60HWLBcIoOTkk/+hwQaFHT0wrRU1uucBWApRsD/AnDg1Gb8PfsgfWLpiQkfRjWsY
gAnScOa/hCYi+OnSkJgt0MZAGwxiqQJ0V7CtR862z+QkcPGFXvtJzPmcZbftfT0sp/G9oXeUXLTC
Blm5CzwUyQo9LIV8urfDbPvIGxoIk3MWU7TRnxSyBo0YXvRrZ5z246M0HSHlNYPl7RyxM/jmJpDN
CFLdM5r4b7iN6LTjlMy31VrNa1miBSNkiG/LCt7axbq6WBRpFizVyIgUbhIHBwpRR93gSH9LXdWD
r6+dWM7eheU4zFvURqmdfmYdWMKjXljaLSL3vMzRDMyLziysctRoex5bVRTQIEmIxOKEqqAM4bu/
OEGLXaDn8pq+hfJClw6SrWfVlA9llo0aMZZEq87c9lyl+7kSN2ldPs5Jviur3fIlGQmF5mCTXerm
DOhqsa9wGZeL7A0gV6S2tlUU2wRa7LS/Bn9LCnw2K3zqocxLKxxhn5hfCBusfnFFmyOyBbvpDZ7w
yvrvJEJHpdHZUrRWV6TGMpMeiU6MuTpyiKi4mS4i1VCqWxTpJirXrXXE06GlSv8gyjdVxrFzau4I
y5FyJ5Y6AyImiKVgi/I5HOVuYFPQxzHh+zPDw1TyiEAM8cWuQNp0YU4NFwF9qP6CJoYqGz1YTnLO
DPWPrJcmpIfcJJHY2VdUslsTQ1qY8uaTr2iN5AldF07hlWmRg25jj5wn5GcHbU7IO0yLIQZzym7c
TUSsrFF9pQgWjrpIb+y894PETV7Qx2rKfBemCWIbDDqfw63DJOCYKoNbRHmi66khUxdg2b4jJ+Vc
ZohY+WXg0t3V/9TCrnBfukX88UWefISpuv+8rw/eTbQHJA18cy07d8/cUpDLMnTXB9HHRYAH0hq3
znjxIZn/EVjVvi1uLjsH/kvKOWl2gg0FY05j7B7waFqNKq4TdXFKdSiU+O3KNJZ/2maZZy3pBJ1b
MscVotQ5Z63XVXzaHj4QsZ/YXwWapT1OgRvwAyWns6GLHBuZSUnEmib6kHwlMt5D8l8hfRfh1ErM
ciMuIvSenqOirrsHDzQkrULYPs50fjDQodpZQoecivvgMa9iuScCiWSjiOJKhwHFq4cx5yHmlIK8
nVMYgy5DVqNArMHr2mLcqk3pznHKIusumteDmF8o747Q0zOz6FXKDqySGcFnc65f7tr38gbzdnjK
+ROX0kxy9RQlKOR3qSrvXPQN1pdL6dpIp/AMDtv6c9RE4XdEGid5Xvwk4O0a57mq3IF7DqKScR+4
fifCv26+dPeMW4QCH6RmY48nJQtJ9NAULY/V1GmtoMYPwbJE6FESJjfTjJMiEKv3S8sDAdSHV6in
I22ABkqnXM+YkTqS1UFlT3V0nCuuel2ZBMSHaQu6VZqiKil0LI27cbPj8NRmuF9sVPUWnoPFGA/F
OJvuPra7BNT7ml5Oi8nUFOOVRtCDcDjNCwrSWkrsgiwlD6Oj323IAAsqacLMLKaONV3MUTzi/Jpi
MimObGKr7fz8bmDeyrJrWao/nlvgdA/8VAx9e0F7+r+4apZLJXOXV0d7mLAfjXJ/ZabV3LCmVuzA
Iga45CpQlh9nZLAQlhHBbaXseDd57B/ZrENZ2Eq3mwcP+8JoWROpFKmp3P5hr6yvvkYPaW2Mw1Oh
bwQ1fLUgRvkjtyMZrgHDHxyGO9aB+RBZpC8MnfAtQwlFZY3mpq2854nb8kuqCCu6r2uhbXhAnMlp
UPqfDEq1eVV3kWf0N4I1+H/Xw/6vMSfI93GeFFXwj0NCujpXrznQsbB7UUujBJbtmVsweLX6dC/W
qKDSa7Wih2M+VLc0dg8P8nRa6VgoIdbJny6bhzLQ+B94vn8t/l9dFoYeJiJ1Nk1e1Du5MKRxwNRn
+VDXiaMT42msQVO0yOJzVQjWIaXWteMhyAIAw5bjYUNQVJAGiKSJaBF4HAS6HFBc9EBU6+KSXDAj
O4UI+IhzGsFIriywsHQhNyxOwPMSfbM/R3/FeUodSsnvi4Xd5io11BtP4zcUUzGdj00ic8NXTJ6B
pxsoAXUXqndH1g+GBxAS05xO8brlqIS03Y1R6IQ/KoY1IIuFjsoouW6nrGn8SUEmu2GrflKUvYrJ
Zd0yS22UanZmWCzA70UIT+z62wDHHMUsA+elSo7BrNl2jC/HRIbN1OrXa7yWcuy5XhgzrbXGVXJN
TJ3bZoabFh+tI70fhdnjyFJWskKKSXHTYmIpcRK+t+p0o/cIFkSggNxhtytZ4lRVCmp0IUsR/FKM
n7JoySIgtVI5g+K6CoVtDzBnpcPx3LDIUv0Oqa7npgCDo2viEXe8y4B/v0DHJ69Ie/3Yeo/aar4P
50G/QdV+hdCcGtbAJCn3yFNh0Q4qmg1sUCa4XuXP1WPRuCMTGmUbvHUXEWHs7vC9PPB/xr/QHRSb
hVyiPf4svm+eNLuXX4eVAjwJeu8aVch5BoVXqb77AKg3hebCBY1rom9dWt/Q3eWXeiGKzCNmXjf4
TIVvAH0Fxjhm/MmwnLtJ0WcVaVc31bT5ikSxufYeAwQd3H2/0sJZ7ewc63fxRugyH0w8b8I+0Iap
MMXwMeh7haFDMPPkT8HA9YjX4QLSza1vleA5B0FRxVySAGrGITy8GudQOAGCdhMzMy4+Sa8z+5kJ
MmJNTUsuxAe8x46Z6MFCpTwQYPjFadDOWwpW1lZxZtPVLI88M6kdSyX71ika9AGAeiuT1er5Af1D
WhmlVY0SB7+EWENcmu+vkUVkvtL1fm462o1knZehWo/n6v7R9xBGb4i4DW4KgM6HvQmcl7Rlki+J
eFc+xmNUhwWuakbr67ZMrNxVzqVMIeveGq0nQMQkmaqijFTc6kdGVyyucmNWTSUHRa3BCfAQuVCZ
fJx4saZ+Of2g6p+s3jiBW5fYPa9tnguidk6CuiLis3IuSifkOiIYKeUzw2f+w0bJ7YW7xDvotwVg
Je2A5O+isNXZIwnkZp+HQAbHjZrLExZCgC74xP+aAy2+pg9ZAe5aZLUnH3khJJnLpk3IMtiYF77M
JGpUeixem1iVllM7YzUfc747rueoZtcwq5FtZUP6j3W7Vja9RWi8EypBhHZBhxmd1VTrk2EE1NIY
gJB1fBPFV7IT2MDc2MijyxOzUGfps9tAC7rFQ68eS8IPdkGNbTl8CSSeTxpzDe+RkkX9gDuxbVVf
6eM0XC2UnBal2ZvidbvOKl+zpah0xodBcXWdE2448u8rYCjyKIzvRY6yTGgfGFISZzyvCcw8Kkt1
JqNn6eorudmmZgx4ajEgwNlSoqKRaihD0DEVnsGcAteG20vTZ6oX7uV+sNgOJWJOOj15X9s9rLJp
HcgLyx/uodzGhlTs01IMgNEvy1xFWFzCNsn4t7Z+XhJKUcEf9IT6Mbao7aLk8SBq7bcq3isuG5pg
6ApxrEpByU6vETNHZCdI23DByCfYy8tyxz/TIzrO45YYyoJKjialmlDj39B1nrz7iWOe2wbgiDq0
CEvPV/HQW4hGYPfioX5rGnxPhZXc+kwimMAiLwJy1TPvBasq9BXlgIxFkYdPYvXRqhu3QfRtEKhw
UfpYjIM5ZT6LEkQHuUy5x6OVilCtSyAQgTjsE6T9oLxQQlZSnX3Taxd1ocy59LaEGuDTpRJSO4Ht
Cq3YXRGHcVW6+dmONcdcIxEoL+TMZikWHznlOIFd3sRmCVuVP1xQqNAO91DbeOpoaB76PunB5/7n
yanUVrqi0Ux42aaOlqPg9eOdtDk6nn9LMjLAC84//zw0xE7458VuixdXdfPp6Xq6ifsKg8N71eTU
n+BE6RilMhBu7z7kHa5u1W9ngs+H4ny1lAiWMV95xdI1SE+9SVy9f6xyV41E2+nCFBe2r9CGTaMU
z19htCDThk7rMDuL23DmWVPV9buSRVU9FbzpJg3ijZhIA9sUDYYJcvO3+euDYPmGu25yyNlbiFVj
RMQ1Vdfnfrw4P8AEShNFvHo6LF60E5+6jwGAgqeMx0Gf+po71oR+aWFTAasih1S6mqF5Pjtu2e1M
QJFMEaGLKN34TxZpPHCgA/0VEAMiCQ56cHtl9BAz0qDWIWyoxDK9/eNK8aO3lkLKaCKq78HDAgjE
9x8r7kIeflCWRQBgE+86MD0rDIaHF5omLmX3ICegw7C7/XEJt3TgJ/LDiZ+noEhUD300ouekWSvq
RzZeIysfT4u04pn6FhvnmPTFz1ZhN+VL8ppR0sjfoNyhvXOKYYVjqt0JBmh07LRvxPUz+uyxeTlj
81myFlxqaB9uNIpIGbMHZn3+gnYyFQx3IKCBDDrDfaT+JwL12rzjm9x4UFf/Pq/FXJyo0skve/ep
4NCiASPLzMpXeWOCLP1w2fF9vxgL/1zOKpst7BDm3jSEiMRF1Aq0gX+ayqsiNrPp+eziQMZrvE6B
C/be9YljZPoQVS3oe3o/2yYYJp53eXCdD1f11wTcebG8uKixGMLfECkDQbKKI8juNedRLddVr0IE
2WK2MiwBgz4FGvHaHzmOdSzerWtMN1D391P/3L3OUMS/7MKQVmX9N9/Dwe4Sz2yXgyed7D3/G2oc
JSrr3V5Lr0qJVWveS7Rg6zNhcPifIQlDuyUdAkFung6Z9mWhLbMO1p9WqiIisvg7Imw7266SdivA
pxO1syHt2bG1dyWhgA/fDcRzZRLgSsgH56+o2kt8qEU403Z0yP9QEIojD9MikSrIeLbSU0ndN5mQ
d2VOg/fHV4cpZQfayRNHd7yqVm52cejBmehmW2yYSpgNZULqWC4AvTc8Hb45/UVhmcvmosnMnSLe
OyUgse/QjIHzKzAlygWO5O79zn9HE/1ZruvlGA5pVWmCif+d3gxcs52HbGN8VC3+g03Tk+ufmbrc
jcepfJoFSmvgcer3T00rzlt4YWSIlXPSqX4134pZTXwzqCxGnbseqaVnRndfBt5+cNd4cxVf1Leg
uHAwbPqzPsCQs2lr7EjZ/BlKJ1JBwJhgxfQc8pkSdfm2pXffRNReDwEG+GzekdacDzrO2moMSQsE
HWox7N80K6ZHfMzor90hULDnVRo/8RGHViBaEUPXZm4XktwBB86TyfKD6M5/aiSpTKf6PZjyRmvM
5sr3qoncVxA1AoqD+qbtJIicz5Us5OBpHdFMIRPSRwWezhzAH+W2aqKb1UTbVMzD7PIipFEAkZbq
lewSWtrxDmvZOQC4GhEhY03H24PkvsceHZsYKTLGNDTS8KxWmC8lmQu1pdHzfozbqiGnleUKWotu
HeZLqVp/DblPFvbue+fv45xYQJ1VDVrXGbZY1z8XpFDUFvRBPNb6k9XNeEQs7acNPXlkAWxBGisZ
5LSnkGKrUDDc0+ZNNAr56f4EeCQI3y0VOGAX6yG1yA0kaNWayaQg8pY6Yr3aBU8ijFIIMFLZSNqn
Dx8gITtLqgIaEf7McKvznJZn2sAa4uyU2Ubwo1vYmOygH5LgsrZaI+ljpyS30kJANzbWUFcdXJ8h
jL//xQpoQmhw6XCkhcITLcOfEySgy3QBDtH5PA/mGtk+x2e7gVWlfc6M9gumuue4WMHB+5vAXqgO
waao2UINAgVR2tJpt5bpDRGR8ysg8Sr3dgrJbG9J/2qFfryQhpZjJLPFXGW6V639JXiOPqPTb+Is
ecuEGkyDH0aAxZM2PsR9C55c6jJXms1loFQBFxrQllV01/BP9Ff4BxCeUDyL3Ff0F/u0Oi/frIN+
JeXZtn5g0eL/n1Q9lMKk+RvogHKH0I2lU7PHrXeioPZmwEFm3/1mRVWS9+NWPEPnl6IWB1SYyJ4C
A4G4TcWeH+PkGrJoRSeuEJfgKTJwDPdIdPD47+P+zRV8RLGK1eZX7cbNd2ULUL9QJpZl9OWy0VEU
LkGYYmIz1yYXsQsyWS6MWDPfBXDNwTfPpTfJGx3vE/1C+TiJdJjls9jpSz3kwflg8e3NqMfXwSvc
wCUoauT3fFBePzIyNpzT5OuNmdYuKcB5WnR6HgKaRA1JXRj5+0cD2HOyh67rVKAEbq+1efFpFOxe
ctEG89ED3+nb8U3nkH18Szb5AFg+r7gtYf4SiicRbiy1gITy/vMHZ5I/6ov0Qistqp0wBpi59njZ
lKRYmS4FmQszNY0lRCw7FpjFIEF3pti808piwAli9U2NiPaEh5x4nLRS+FP4mrWHAUkzvAbkTUOG
nrBYz9KshZhk6qRQ/dAt6WihmwILwVVIkK4U9ioEZgaZJHo3sAY8ahlo8ONwTmyFgBRHB0yHpwXY
DKmZg1F+dSowFc4cVXOrnvnAGEUh0HaCzEHCEdPdNhA4K4CYxiA53e47cHsccwtt229ln0z1Assb
KgyYQ05CgfIDOHTnYwdaXKobiahp/pugJ48tYidsly5CqvTytM4lX1IR6SHuIgwWaKAv/JF8PPTA
QZoFph0a4ZIuYj0ayMR7IcsrUoPl5pLSGXqlTF1Z57EqOgJsDzgEAWcpylHsFJ/QEgpAP5DMsV/w
aYD4l3EMZx7wZBNDE7ZdcPk7+VGnL7pT+CSjcchTRtuO1krnUD7iaaRddC2uHu7TyFS8oRJoNAYf
9M+3ByS0l+W7L5yLDgjjb9yGD5Lq4dfjojhOseRL9eKn6zasw379AraDeGqqwrIUtcPRzQ5Nd0AU
m+ktyBnxqGCb92S1W/zYOdNDxPJz4z8AVfNHpGciKpCmLg34PkJeg/wOsqP1uFgkg1JGxw0AebGU
TzcRh3xyx7jn0ikIuTAFmNOYLTlnB6cqwUmiBcRPX0YA4azA2FEkSmNjFjpqcHbf6hSxcTtOPOc7
7XdBOp0hXwX25VfR91uA52xUE5ZFS5TuUz0KtKYSoqMqSmCJvwMy//gcEGmSP03P/l7uMS3WPkgN
FkJo22Pc+al4dvCckS7kN0fGu1QJnqtgu7LaBFceiAOPmMAV/1IIC9X6eGtu+KHsvgVe1hmRl2rY
LjMAPpDmDSkeGJxH+ORArnxqqOVnhCg34UIud3CUCwy4i3Y4dRheu7XN2Vhg2WSugHUZySRzf/Kf
IE/MTONqMbFEB/7sL54mx0Wxm2RjvNFpCxXxlHMPYPU9REcLIjlzI3pBMyIt+EWIXjy8zXB3H25L
/HOGntvuiyzTcW0Bsiqxd8vdJhxlHQrrOVcGDMxMkCwSbvjs7oc7qbFMCPHlpAxjqFu/eG3supVL
F/ld62voL/2WVrPN3bCXANHQr0MWhxCxdVuegmRqYFzkqZ09N52GODAPKnpSBjbXCYXx6Mi9V1eQ
VU07ZRnZJBJ1rcDAoWOoh93zjlWXWeQ77jTjoozeRqGmiDkiKw1dhGm+xtgpJ1AfsQJd0lTP//38
5xmnzKjxze0hnO8wHYjGhyIxhnob+lSAXuxS9zD9MgHjXuzuXdSqRvsL2OAmGcumXxRy8GemDP1K
HGIkiPDDKGV1LiFr4Q6QZmCFMLMeuXGcE4VdGWC8Bg5H7yavYLNgWY4kOnWZLfQ40h2dYTFEcwvr
asnk4qq3mQdPq6B2lkUel2omnQmdXsQ5aXui+9WBAiyP0kuIkwNrcLv883CZyoKFZwLYLnGgFio5
DZMT92+jRl6yumcEKXhT36IdzOL9Z+ErzUVd2k2/rqwWOgofNE3e0n0Kh6iB88NAKs3qj6VXJi1V
nbqYye+Zs549XogJJscFsZwDwINxS11zNc+nSc3rL2gsNVciOgs7b8iBltrngfJAk2HKqUc5uoxC
XhmCtXzRFb2902EPv1/s8WhEvUc+oMvMfX5XvcsT4PDl6eoffL7HVK+iAzRC0sq9YyQK+cAreHy+
GCa0twa1AX5uClY0pbC8y+o5zvCGs6wt0zYRg8SWM6+wJIsFoiHdxXCrl8Nl5d/XDcZaW0q/thtJ
KpiwB38TVVtYqSewfeKfKRuX6VjTsFzffSJGw16CnAhZYJUdCeHR1lTTPj2cJ2Hj7f6n6Oz19aGd
LfAqw6Ut/vs1v0DEMcl1MxXu86sy7WILDLAZtC4N7uuxUB8+nrrNbAJ4xk4l3SZzlkrcIY4gmJaG
EvmPFyQ4SuwJRxZukuMoj4vUCTsehf1Al8g9ePszO8s2O3w1LI8ygW4LS5EloG4mNQAtmTAE/2Yd
S6QTfeahMe9+jMALIY/qlp6KGfh63xlnytC0eHwNovzvKppJaMhzWyrporrbsbg2OISHMA2Nez8E
559fQrEZpaQGMluWUH+F9TlAyFENBsJ8c2gVLRrhKHzp2xyf+1ifGVxcnrdCCjma/ioFh7QZ7C4c
/VGX6NGLU4BG74EVgQSGYoUPyUYTyJwftR/4KqJchF7yyb14hoStSXfkTut7C4ERqZd6Dg1ludFe
Xj9bXsd1/hll3O0olN1MGOtdP2f8G+Y/ZtKzJvSTYKBo/myyOE9/3oawY9KLWBZIsJkVvxZLHw6+
8PjC582felFKEGdMwHWd0/csyxJsNKnS6yOj0C06q3LEQ9h1I6MbGSDWiwLS8UlBXkcGdETgE1FK
qNhS7OweUSFyGA6VGxO/0QPrsUaMXj7vS0gpC/fWKQJ0Gi5SmrZuKQcanCSEUWIEaL9WSUu0S82s
xl/1JY+auAaQfx0xg3wPIsip+4H6GXjm+fBlGWPqPOFxwb3lp5uHruEjDggdrFJmnXNZS4CT2s1c
arwRZKEJixBp0yiqsRFvp5xyftJ3BHRtbVt6+k2tzsSagYUitauMhjWYNWODgwBn3g9YCrRROFu9
WbtpX5IaJhlFKyuGqu2+PxNbaxJgg1PlHwLcrIFdVssr6UV3YESj4nOUdhjpJ3RH+f7vichrlAyA
vsvpOXdB/CXyrMHjLM8UH4WReLt/LU/htLNE4xcmleDVwFpif2oLkY1iuRQsHMjXVxrSUG0lyTns
prfypfDmHox7F9KgpC8CQ7sZu8uc/R43VDMmnGBqpsbYzQJaUv7C8aGDH3C7fs7TKfAjgkGkpNhb
OqBQRmm5AkBHmpoKTIXS2gJU7+XUp/zH4Sx4IwB3/BRa0FBcNS91BxpVXmkbPHwvfatBd7SHh1Ya
FUQ7cd6qd1ouFyTJw9SqUqtpw/COKn95UeRMvLToqLWjgcq81XtdHbMP+LWZkyGfpUF+feG9xDRO
jX3YjizMflqFIQQYqeWPwl54w25eXFeehJGUk3LKZs5d9pWBM28xiAU00RBIQNrSjKeid2yxNyD5
hklJVK+sNHbqWLLNbjjIkKQlqln2kvuxP9HCh/1W6gJgkQsCB0pgDlKjFVVgElAkoBkplvTDKv7N
Vuo/XehfcqNeUNr5K+xFlZHsDsYON4wrXPMEz+AGY6C+pnt5UKh6gdIaOAmxHmV0Th14/Smwtzzz
WJe3NFgtpXqYEYD2E6kwDF+/IncbHJ3E0tpXuDSipMJNC7nXpya3YpOyjIgRPlJGf5q2NGYXalCE
2fi3nltbyNSKTZAvl7j0oixeaKsUAEGTIqvkydQe5agF+em1GT3VClDh0tEwLT9EyKpQgSxoVUOd
d0x7kMXqqWDIcuNZHDQdHhO97ZWKPoYHFzZeXD0oMTR1QG/dzME0Ipz3fYJ0lJDgcJcwbmyDcFQg
QMo0bg1YiGXYNjmQRZ019/uVRHht/HjSrDwGWoE9IZL3Zf1wm1nszo6dJV/iFjxNZNKPTwyT2MHl
edtEw596ExqDyMzz+wnLo9hw8z8shz6LBzFgdMvrDQNXuKJDN2qOMHBn8LnTrQRNArjFtIe/Wtts
+Lc+YvygGU0IaUoxGq2tlCymARq1/ILnF28J9t+ktHMU40wdNRqxeZuvwAcQrCpURaLWCklikbom
Bdhj185Kd353weDQU/DGR8CciXbozvOiuN2V6HehN8pIttI6ouckCWOQ7gZ3lQpDam1BS5diOq2P
nfbpWoQk3KUJZn8VlcWzDQq/sJmgxRwA8V9/fkwjfFWh7LGDGrJikB9yIQl3tVDXDKgU7fVUqLNp
aDd7JoLrZKvrAF0YAsZs1jT3OV9XP+gpcmPs1a8khvcZDFDNIhjvbYpFAZ4ZzOlu3ffY9dAzZBDA
2YA/N0VGAZUWnLFIXQb4Vx4kUU+2GGc44TUrBZybxJtHuYhl9dD0tmrz2czm3DpMHWgjkc/PYDFG
5mqT3xaHNrSgIIBb7Z0Z54+BvgEXDWIJ6J6Crs4WD1vZG/bE+1fS3yLbZGGIatjOo0sv4FTjLVf+
STgjoYUiqTCYOFmT3dU4e8UDJ6hNSphsXXAgYjj1afINjwAtaQPV5VfJ8sjrO/iIrMsbvqKFI5mU
1ISGnL8key3zmzExX3h9mnBut+JxHAnn3v2pPVJu7YlRNsIbxnRIjC/PywgcUe70XpD/fBarjNjo
tixMFK4d+TjQQLo957LNCzT9s0Ib/Ew+wQW4j5tGbthR3ycHPvtAbxeJyvmBtl9ooRG+kCKTaIAM
JLpLs8iVZmh04+/OV4DAMv5xFL1unlt3nFlnypmsSvNHJmNPschx9pKjtI6c+vTMGH4nc1ZBJKNH
MZomO54hRFBNPQRYE+WlZxGYS/bxDD7qoI/9vrb/8mw1nYB5Dkqw3xznZUWqKBN1LQuxuWaOL2cQ
KLksUelj0BnUK0TLZTwhqVRWJ1lr8pDJ/XB0g+9c2pcipkgi+OH8UwOOAG5sLPRD/SrtdYYhiIA5
e3EWGzR/UOUKD13GDYZHRqif39r0IUjyib1GZ7lA7O29RyBOVm8qljsX3EOJyFiWUvMhhzUygQ8U
HAwanem5/liZlLTwbnWjx9u/umBJoqd9JKt0CJXpSBDQwiCaGPITowBpEuCkvzQ1BQlcKbphDpp0
H0S1Jgj/ScJa8im9RCUVB6lqoFvFgL8bfMiWS3mEdEqrDWUYZKfU+gyOa8jXwRtKq37jxeDnTOXW
c1bPdCwDeHG26/r4TMDudaRsyxTwb18EhCsWm3ETRg0vw2O876ImgJSxtAlt/do8bslGZJ7XFMO6
LAhDQeSYsixqS2Dn4FO9PnegpH04wVNMBPd+/vGcOdivJRQbaSLrU/JhA7mDtXDjrorAxSuYPaER
0HajH2F9oEeAdLDNJIEcXzZ7YxB1lpg/MggsO2MhReWwzgaQpeNK43pYnpvRS0gDWERZ/ptRiOIu
qYf0eYlvUGT83h5+rBqfhkXwusXSLv+uMtvqiRe2NIho9gv4s1rHYYxU70TTzDlnFogMeKvtoNCZ
z2x1SaN08a3wja7tNQAOpE0fO3CVoa8O6uYasxZyjVQFPqA1b9ZjKU8BkUtTjgFLAC/DA5E2hLL+
wr86ZvhuxcPRvPR5g+HMZ+GPsRan24qDRhqNTIR2YN8Y/sLh7icxTOHxkcDNB0HtnKJrUf5hxrdA
ThoqSPSiqw8eTBGp40BmoNO5JGnAOr5y7H4mnx8WrjKJnmbEQwBBYPHI6AFJtcTb1Ok1jAObHwUD
sbeXbA4XgT1eWdjOUzaVEJ5LF8+1PwFl7F1cMbCPZX+TSHsmwd4g3UZKWTO7Ou3bXqIOY4AwqLI8
dAMQ1jZNhtguhQiuswor5G0UesvUCpAAIUDXdMu/4WhPMgJQW3aS9xh65fkmJC5heRqA1bwVJ3QK
8XZKiO6HuOZUHPXtg12fXVarfJ5VMlKT6BJznawmZkDr5tXWMAbTQ0ULDQIbRtPkOyusDYghJrJh
+H/tBw2MAP0KOPrxwRntYLaWNVljjBlC7DQrmQoxDU7oP5y8JSZ2wy8+5PY4MGz5ramCtcEsJG7+
wcQeGFJxNXcUdj1nHdCeIipQyFTzQVfJOipGVMi21Xyj3FPhEh4GULAUZLvSeBxo/cU/hXkW4m9M
3y3YrCLGe7vPXWghu3AE1mC1y/NWPvMYDFu/TQvqjlQWxAYzdyCAs1PYkT+dsJku5Ti5PRHumAzq
Bru67bJRS4CfGFgHLZh1Ojv17FnRRrb7SkusQjLnEobMMPiVj/fP4Gw1hlR32jT5S/uzxtTVll+4
zk2VTlpHUymuJUvv7T1//kawswjZJ4ORcRrycu1SCflnSabCnGh65qT2NbOXaua/I9b8Swapsvox
1G13m79cKbIX7w759+8sypfWzFo555hvZdEw7tfgTSfGTuKV3FkQwHYXE34VhmOT3pxWAQbfr2d4
8a6Yu3qBnPsrk1HWM5NU/8s7+QKgw8oUHIe8smEITGhyqK4sfmksMjT6rJ4IqtSjnnKGr3t5mpEg
+J8N8XOcbiRf+Tzxi1SBHQLJXHZG6SkarAyxTqtDykHi46SI8x0rHQQwG173aYPbo+0bHhFbZbAU
Qj57jVRdHjT+NGCjVsP+0thLx03LJ3FfcdUCuYud+qsM5MViKs/Q7AXGsvPeUqfHaGnvA8m/2nNo
DmJ1mCLL/SRnvycElyzP725jgpAMiI7iRm1JCJXRiOxSwqBqAJ/WncckguaP8NQDSyWCRqHNNboO
VBdRRg7kq3OGTWWA4upzGYfQYIJCUx6HhV0DTnVtqtHDQkTdOHPiqK10+FoFc81v91xg4PQdFCMJ
LbXorFQVJD1ooNTS+d/DDvGMDmOIWXvA3TtYsKB9fpVwx/hPZi6rOl/V9GfcGH7FlJsXYUV82m87
qMHwpcbFaJDxbadNgZwu7Uq+HYxGq84R8XEVZC3Pu3aymxE1RS5Vdz2nwadxoEKhY4vINXEUD1xd
upMEH7Oe3ZW3+AHrwRr09IdfJP5RZQwK+kqz9jNZ5wm8OehUmyFtl6eFeLkjfuvADNTnN0Spy96J
E1+Fa2b5wtS6L+MXXc/m4nsgCN/2u9Rbm+xzpx5mcXAF8IRqp1R3dtE5Sb6HXNpeZSMyWklAPpra
LCv/PXUskH5lXgPgzfvd8xOLj8w/yIhwJG9UOaJ83F+/At9bRAy/edeCAyyu9u/zvuIqMp/1cYt5
8eWBcmwcjo6S6cKZypg890dDAUF63l+1WNoLD9wRyacsU63dUn8EGHY+VzxjQC3eQx5HaUBH5B15
XyR0oFCHwHG42iYSZ1t67JgeTR1IuXBIXK8TZGDApzLmd4N01XX7ZY/gXtv4g0+QpyL5vtPfo/Ni
lqI3elDcdSCu3Zf5vIUNFb7DcxAaKMshlpK8zMzo9Yc2zf0DaC9XGfRv6aSzqc3JSeFpV0mg3hgn
lG+2p+XooVzpVG7GjJlV1uTMvzfpPSCEfCV6WLMIGJ9coNBO/Jm20e4S5mvbuf7rW7sQA9m5e8Nf
+7b5KAC+Vgtmb4JBeiaBciNwI4aDn+jKztITl7x5j4VOaPglsmmEFdRWcIS1iBmtzruuOtT+kJs8
5kLdENxqxdRqQxVsR5uwBKFDwIX3CGzG9V+pYyg2/ferLqa6PNN8dAGYCciE+6lTLWI0y9Lglx0E
PicVf727QRIKATw2voEX74Nb+bjSenSedP2PVf/K2ROzb4QPND4oZL0aBdRnRNp0rZgbunZj7KHH
w4SqyjUx8uXOSgEeuxmvftoWQF7OP1o9i82x2k9xwp+QoCWs76s3QCQFb6K3GtOudu9aXei1Ijf7
Y3TB2sa7OmoGSLTUa7Z3UDB73PFXm0PpB/X3pvxbT4XF+ptGdeQWE4JgCJ39ewESoDo9ShoGwKIH
sRh9WfiqOR4yekw9knZmdqz5Hk+MabgYgkrwwl5nFwS0Gj0s1hGKH/kJWtUvn42fHbmQ1Pd4NfS8
FDpWy4l5mzKkF/i5MfTeZB0x7A7HfQLHR6XzN/3ORemU76n4VRU3wh+VOZUFH93b9b/gORrXlq3B
x/M0XYFJ+Y+QDft+XSOwYT2+iFPGNkAzXwPHFWeE+JN2/G1OTa0mbSbscyChd3W0pnpbsL/661mT
mRd6RfdlDkjbEBVOpoyuAmLE5AdNipqn6309LLlY4/tRSDnOWDNaXnXDKzpFlz52XGu3SyL1gyq/
zji0ASoAjSFiq30Sl8bFX7xx3rGYRt54RDje3Cn0X9aRkham39GTkrK4eEeN9NID/NJ8rUR5KknS
DU2+/2d7T3Cg/uPWZayFbUdvaxiaYn0/OeFYVkAy27dg8ZinUqiVzQyz0TswzsYYKsHimkd4/55u
67rGVzXXhzIaSUZ+/HKLZ9n9Bhyxk+a2Lj1Gmmi2FrWE32kNvkiWwKL/lfPFfdPe2FpMrcXCutBo
kRRXOEypVjkMER45mU7H3veuhDDNl23ayhC/FBp/5b7XyCzDWq2wR85KK61HWrL+bEtxBLU8Q7kA
AW2e5y0sJp++nDOCBLzQtaOSfIX+YVgNqlr4DNABzvz/I2ebNIQereX8laEZYkm5ySXr34eKCjqJ
IG6TUkWXYbbc3TcYWSxSs87TyeMB+lLoLmZHEVk8uJ74rWheY0Tzd5i3l1YO1n9xpQueKNte9hED
W1hDlEefW3pAziEe92yVPM4No61/DZ6GgnNGnFOIsaClpg7pARxfZ95TitozYcGJ7UflNSnDLPou
ycmZL9RVW0gIB00T8d69m/Qrf/arnZZskTyCuLKZtTo19QJ2w+dFgiBEm5zBaewpRW07hoga2X2s
iGjivn5YfHvPlYNLi0CK3jzYTbboVR3j0hubx+Y0zw7qCBbdIVUSJE557DKUEc5yfmnCvpOXm2j/
uprvrxppp6cFIKt1Sl3PMLXjuYQQbNwUP5ayDB9/D927Y6ETPnKH2oo35m7qlWhJN3b7jVMA/5n8
QQHnzKK6xMVb3VU3pbsvCYy9O2knGsKz0zWK+CnfkHQtGc7LkcdQG33C8bIChbVl26qXEHNGBZuS
FwTv5+oHYPm1YGHUiUydwWEasucp3pqmMcw7rM2Y2JH8hyAwqB2/4ArkvrCWQzo9AcJ+yiSxcTxW
N9r6Iyy7yh6j009ZWWPhvWtNjv+1p24HKu6MZtiFvShULKheXwJ8EX8RBsj89Lc1F7ZoDDZH1gsR
f6qqwgHBVdm+yZufKghsu9rCL5jekbyVHIzejStXcm87wbhf7mUBVdFIN3lxO2+sZy5I8Fx/Ww2o
wShnC6Bjn4kRWzW5m9ixX4igXszYSIOyPcPNaciq2Bw0VAAQxlgWuhYrJd0PwguzL2ZcEiEbUEUl
cCRfB5Kgohj0gHQeT3lXTkiAFQmT1jaqvdiN6LKz9GbXtHpZaNydwcCmfYWw9oFyoUr6dQG1gbU1
1K+3CQcGh1axoPCUwFoGE4uzkk8PBsW6TuPlbacddZi14zS6/wVgjB7OjYAjHiQapQJwVyaTh2mp
WzrGEOLksG5vrfEVSmG5uyZLvl+EvFlyc6m7kpTNDEoqvjl9VClPR2YHGeEp9VaXEalfghIHvHAM
qzIfC+1R6dvtMIWlOh+DD9sQbuII+AXmzHtV2zqTmbbf4t2nIcR3ZCrPArrpE9XteP7KuF5UTWRS
zwOxhL0HIKoNMukmSz5SjswmCl4Zu2R7N15rGM1ZIG4Dq1y2iMU5aNtxvEUL+PG1XmUvzj/864e9
Nq7Y8OGiUDGo2DZUtSQvV7Xi2/2h6IqedoBMvU307FX+6g5ovj9964q1847WBieVkIuwphzscHPa
1JqWlTR6qqqj25akhk6ardgROYGOwP3OWfG018d8jWASISfHDvQQPMJ6fAAtDAGyHIHKr3QHwSS/
skyWcNyGECkq5pu3Puu7+TpFUBIP9mG2aVRmLlbdznwgEVVqmKy+/z9SeFCaCacgp6+Yf0KfpSSQ
lrKFakuuZEiSfFMxOo9gJww1qnpjD+YxMlCtiLcQYTyOd2SRDdXHiabg3pzm81lNi4M1h9eIedKO
QuYQLX5vWtZ3nOV0sV5U1niIz++bUa64vzP7Q8phsTWv5H690XVu3WSwrT0BehDF2GhhnPdbCXMz
2kqe9B9QVYdHShwiyhH/Hxciqu/wOw+oZJmwsAUb0VeerV6YmKl/LrMy8TWd3R8CpC/vWtSupb24
ELv2BaP8qFbf9n54tMpmqalIPzxq6wHeEgDjluvXKeEm8q8zUakQqzOPyFFZzEdJ6gF4pnsRKv2c
oYwq5tI3zdnyX4JbL6D8xOZ73R0pfP/0Jfa7V7HOmv+EFOZp/080C53BhUlOWGVYCtoUvGuMpq2j
FZ158lL+kkKKV1xVTlqIaPTaf+TWpQUGViR/itcA+LF3PN4jqN9Wm/Uco+D5qkAQYlDi88A1xzlJ
rKX62fQJgboXx2CnHqS+hj9ZbcGMcoEkRJYgz/VqTzvClgzEP3Oq+3hviRb6rUkQiYAkKOxjAuEt
1B0zdRwTC3tAdUrIxH0h5Bxc+XbUAwPKECuftef9EdBXFO9ft3v8YzzrOhmu7CfZcfUMgDxSXJN1
ePCX3jk7Q+r3PGCK+Z1IY7M4T7F1KYBsgnfa6K+YUjXGt/qOcQeskLbk5QCr7+yWtQsRCKPl19O8
DWm2sJpT975hxrTnY4e3AXmLP7l6S4PNE0BRXWYWfGqPaCE68UefVoP2U5vXJCY7vhnZJ4iZ4DMg
oMU60iFhS/73TzRo+Vw0QkYJSg1wGZQD6kLlE+WzW2RI4HBz3Qb4yjIE9waAhIwlvnJU2JFOmZ0q
Lec5OfAeBhrYezGkK0QfrKYSXY+3V+5BfLZypO0y9WOTkJQKc13fyQzjcBZSdbgKVzuYkuebPKmi
TOLj8qdNAmzU+OlZ9EJ0nRlWFLdIi2upJdjVrIV+WKxAZ+YBXev/iS3ZHNiNu8yGOAUHs5XQVcPX
6AqQf7B6cQ1qCMPN5MYa2SrERD2uaTbab9mQd7WwgL7H472qkK0w47k7pb3AIbCZrwIetsr6j4AH
d21tTSW5iEjFHVszGxmRW3lJ3W1ABWVhzCrcFcUeXGZUad3MmLomWZvDwUD5kL8Xa2TQp4kVEVlv
FzQvyvIJUJiFGC4eVxheU9biOrdFD7UhrsZRdPx89ZBFvWX/zDcbVvLR7JMepiolCBEPg0BMdcuC
KjrO+yDHQ5DwuKdDW81J+XQPyhN1zXdbTYliABP9EXhZpbBE3O/oEaYudSq1k7Azmec9BPFf0ggW
N/9BPmKwGfKxkSBhQDWP2yFOkkBPrvcWWBkyyT0i5VTbN9W+xqPOfwko5wVsDKcscwCaXzhxi11K
m5pbjkmNyR8MLBrlZiNOpDINk5sR4S75OjTtDyghcc1K0Iq4tOqhyTjg8rnemOyN+BUZwiqjJOm4
6o4wTmHdgK89fi3DsKDM2l4nJooXWDeYIGdUEaNLJSQ+q/tuIh1EhfhiXARMXzVXj7v4HNrBSDbj
2OFDlrsfumpFLXOcIMxWrvYUwtQqxIafTVAqQKW5VCtqdKbW8KmGWjnLyZkifJaqAmiCP+CfuEMz
O0FDooQDlMXyHvxHDLZjMtIcPNucLvuMsdQEAQSDJOBtSuKbaxcFnH2XI6zQihh8Ksyr5l9trDm4
5lysC7WZYPr76llrqpudwUOOXTM4+rWsSKIhVFs3J/31Tt1eznCv7lLgpApTF9mWqt1c59fzO2P0
KOEG249lMllcHyCS34fQTlBEXdBBFvmLQqZTlf+EBJw3C7Jg/AWpT+xdA03x3dxUxrfHnZi7ykLR
H3eSmW7rnh4KQyYAgUztSbd6fPUak0ToQeys7SxGR1ZnejBDjy4aanysocR9+nA9QDDhVfVWBsFp
VCpGc/9WC3HpGIQoG19RVxD/aLj8d7ezcL9mHk0eROg04frLwHRPPG0io4aRstCcWIHMpnH2/gPK
F5zaeWf8WnF0SftnR6HlTlGz5zXRWfia+2NrUFyR6ZuVwwz8GV3n1w/3GYCyWjWi5Nc3RiFGIXtJ
7Ulzta/t85yvdwRcFuFWYd68Zu/vr3eVaE1VfSLM7Ul8eEZmhXfXcMd4Tt1TAvDKS6/pzIO/yzSS
ZZ6VDnsWovtIhXrKfjhpV/zJ7JQu76sLggsoW9mCvPzmNOrbYELR0medcqHA/Hnm7LofcpbY2xhr
xT7K+oBzPRZrcYlNu3QGBGtWtDnMg31kqPuvAi2LlSYlm+U+oEkAcpggC7z+vTVlqVxQ5rpz5/sa
lmoZ9Cffr5RVFdL5RMLhgscB92Df7LtdQDtigOjuU8Af1tVUnY7dYc4d6TRxsrAmWWXuf0Jwz88r
Z+fj0Tt0s/ky6/e1LgWk9yJ6ChemUdgbGqNRPkxmDIDZR/crQNaoUydqCa6/uoUMYJpLiHJ/vv2w
EmplH7YKGmb9teZUfVOnPVN1Ud6rVtci5s63uCYnz7RNZAXNVkuH58f2V6XNGjKha2PBEsOUJccR
dqNuE+hquNHVo4wnSfaZZugR/PMTyeT/VmdbsIbP2mhYdePgceM/vWQQ/TfT/zXCUp77pQCN37jH
ceAWvRrhPnemMybskopa9rKntl2m+kgKghoh1fLW8MHr/JFytHjQLFhK/ENjfaPQbPFvStIOquok
iRkFXz9AJzfQRavZwyJCv4jk9y/lz8PwP1wXHXQqUlGUTe36MAsvlp0xRJFDFTqTy2lKvS/6JiGl
vWQw0Chsf4EDa9zlP2HkxDp+OfGPHxim5hnDnzQNS0jbuljEmOUDeJoSOYs6iNVxFngA4Ll1et9v
Yl4V5Klq4WFY7KydO7YhMIIAwUqyacUJaGhjzcxE8U3yFC6wHARo1+XulCi2ubrRcYFSNA9xVfEj
6N1mcEdSVZy7RQTqSsYSvHqbzncAW+HCn1QGnYsrmNAlF48U7yOVKW1mlJbSVfQ7VOmfwZQA+Xw0
JEg3kMQUbK05M0oZwytkfgceCDAB0dpPvCAIWN55/Q9A4HNJ5rd0VIh9tcFbziAP0Cr24hfpOrFb
wpKdmR+k0esiu7sJwEHGNvbtgECSwyMfdHJhQ9T658acA4WyJrDeRbXcAgwc34xImTDmlP/IIy9V
O6VADfgFHAUNPiUgdSqViQGLiH+DJjlKlAkeP9+IZcGyWKbTp5Ctek5a80fuzAtrOMW9p5jK8/uI
GM5CB87TFp4jCuACQGL/86rK/bbRI5vVoOxvrQNwdGv3MKrgdwkhSDQ74pyj8dnPFeFb8BPR4e4v
VuvdmE1uT0MEWKk5sCH8M/yqflF2WlkDSfR2eOqwkYl1iaKTkmAv+ZglS6Aiio7SmthK6oUdg6OP
r/Gh5WwWxPLlA/FUkyd5YXRFkY6X/yQmvdbT5/k5wO4qjyVzN3s/QCBmgXSWzTAxiTdGh0LetjOK
TThdF1vfovmQzOMlk4zUouO6YUAMBKC7GSPibqoDL83bzKbwACTiYMu12WE+zB7augFXrru391o5
OaCTP/swK1ZT/Mjcc5FfnkT/UyAXk+j3SR6l5qJeorVF65dboL79tzXrsljVeklSvk2TAywq5GS8
RlnHksmN0MvFr+26z3/x2kcnC3LFyE817qMo9YBiZ3k9Q3rp6TFOWU/SOkBk0Gi61/I+AudlPfei
npGnPXIQUViR0cvrnw3Y9RfVxS6R9sP8QBjmZIC+YJH21xoPTPerBNqfx7SW0ej5/IN7b1GIAmz+
EjZLW94b7jA1bd4UN0YycjBzrQsjZE/i3We1AHgyx5bDGmALZvHQR3scAJ7ZYJpm9+KJjGMM5upD
Mom98CaEla+cxntFu4vLK22LbHLrjxcqAyAzLAL3Lz2E/xRarKBbpH9w6Y135DWm71ql2ke+CFwd
0DmoiBVz1i3Jq8e50xIps+trWy4D+7RfEEXJJ9ZSnV0lysnG4ukVXhVI4P9pdMBveGZBRGlpO3Cw
ajaG3XzxcT4nKvO6BAkrDHf9Te6p85tk55Sl6cgutok2v9iMdyeJ+dTX3nk9tueahrzbtR5q+NyX
Zx2ZWYgRWH6/AxJlxtYbVZPYxiR5rSqsR2Lz9BdTMpgi3WiaJ2JeMhZPWIHSpIJxggwQ33+G8hw7
lp2ESX144qPqmSlwoaMyWbQ6B7Q15g/iS3axPXEJdaM5u0U0yCCgQZod2S7a2OVWFD+2Fhr+HJIG
VIa+oTcx5QA7E48A5eEF9WojwrD3sQiyM77NAirPV6MJCT4Hn6yAVug/hPMV3aNg31mX9VybVDvw
ODbmK4VwlnEdY820dz+In1YyQq+AAm+uCdRh/trRC7/y9Q+oJ3bQ8vRS2RUFXiElxxpFCFCN74ZG
meiwUZdxtfwcUjuzA9oxIMcozWFCh6I70GgC5HVkesQSeRPu2waqI9cAiKdL3zpits6am9NVhaNu
QVRiUPid/vE2p85d8vJ8X7uWG05X0FQb6f7YeYOjiIQCnZKD22j8+EFqzBNFCzC7Hyckw1StrJxc
EFRTYAwFhhDIS/rrrNOwsv5QCmJSDuNpF6df+urvoemgn7Ot4eHx4q0lief7OIoBts6gzhq5BpSV
Yny08QdLMTg/i47SsdKJE7H8eeiM6kxOAGFBWcrMsPlGKn2dDdx2A9DMiPYIPmX3fXSqZXdFxdxc
TG6+UquJqatiXK3s9tTW9P3XOcIjDT2ON0hLOGkO7Q1oIzsAM5mEAYkIDUQ2WfgveaVm+3XT8WfK
34upsZnWoHM7Wf/XPjAaRFvLsk/4OJhQh6yMy9Tvxw/NeUkdhUszshBbCs2vD1CEmH73MJrTBQ0d
ReOuw4NYHeogTvWvSjgesHxnI7WGHYECMx7H+HJ955PS6l/sycKtjOXqh6gPhIE/KmpuVUMyODWv
6B/pbodsJlkvog8LpuwjwA9Sj4xjDRZkQMlCJqkMU55GWn9mcXyKeAEwzao1K+7AUT0jZnRh6WbF
dIvKZWxqo4MRKlNJsDEUlHAH/HMT9nM4Rv+e2WOK4AARbxt2sRpRi2h57rICf/0ykBrjEEhHwQFP
/jA+5io6LDQVSd9V8Ocn+oD3ZzI9ek4dAa/dQNZPBeQJxM7OQfL0cZsW9ie4ol0G1KijnD7DjMtK
yOx+PSgjHbu4mIxnroIkt47am3UVpPH6oPOx1ZM3G1UQMvkQs+rJqLfNryjWIJnk7AdV3B+/YoQG
29wJov/mXsnvM0zu4ts+SvXca6nkTNkIC88R+TMMeAeWi3VokS2/Mmm2yoEbNUYrpWZLfn70HArQ
JmG5XKF3kIynX2007HB8OmSFthIDJ8wDHqvbdZVamKvopKibBVUGM+XV8qN74UXJd3ceDGQNSFqD
t3uhkC0lEV/L8uS2DwXrOBDD2BHu/VY5avblq5eXyjRBwERsv9n6H7MUl7gLdj0JUDuH3CqTixxp
zihJ67/fX15/LGv+JduNIk1DRs4OO93NQIuGENs1qt0+BO6mzFlJrtNeBw4Maeickfjd0Nhwm8Ne
yELMTkifSOhauLDRYytIYcwozT9h9EeVy3pp1YkDDhJxBIIZtXg9nR36OfeRT2EDu+aIkvXBUvSP
Wiqno5xl0chYBu3BEc4mmBf16PHDmvSOGK/275S1fa/zy9Y0qWDzoAp9/BJ4CSkRgzicVo0LQQOB
s+ZN0uo7GdhkDuHJro36EBI+BWIWV5patuK+9YPokrQkaBaZXMwdc4cwM6gFnp4V8Z0kgxuiu6ji
8rqGXcaRVr2nN9J1NOsUJqdT3hvjtKqByA/Axs6/QfNe6a2KCvul0gfUZTRDKISFv2xV5tKWgKjd
RlzhX2jUWPc3AVd4VjBdxfSgR1q50yd4JuQOr9YQnk1HnBWuRRmNk7tVWGA/zV1Q4L9tM82HQmMo
HeJM4EBjQuA9NNlVcUlTOoZKYBE8RzNzH4QLBHnD/3cvX9T4lwnuh8IEPVcVLr0OHFtgstfcbdTr
v7vXmUKga3tsGlfeiBrWNgKj+NCWDo73qH/hxl//6keHM3i9jcU4xuawUliijaO39BrL63n4NCOh
fS4U7LqxaD5HclB4oEGw+4VvxIHEUDq8iXpT0ThZXL5n4LjjnhoCFf8RnAg6BCL4ju2g6mSWoivM
8RBg1uOnm0BvA9duVp0Yy3ZGZ3DYjpIDcIyVdv17dSPFyy0ZEQbtvcjNNrycRdw7C/uIOXedRF06
+i7Vtu5qJBA8Ypn9DzhySYv+aNbzzkSgjDndekcM+vMbCRJ+QUlxuwbfvi7sYLW2yq0e9YcB0BiN
PE0VPQvY/Yz9JEIVGBKI+eY9MDzN9jFfM0P0Olq0tb8l84E+MsbRPLNjZ/KCKyv9e60tWGESEFNy
DHKYQ2kdz6J2MENfbxlD9VA+UsXVe5f0ebCe6V785kCVeE4LjkO3jzLLHK2AeFsZYvWW+ehs6bej
YP8kXmdo3EB60kV3cK4NY+jiHQ8SGEWk6nu0g9yW+ry4T4sqokoN79ESPm09mrh/AJhzErkObUoP
wiHxRfR1oZdRyxehuHqAAZJeZBrqXdSGIFXpXop/eBocUBZgxPXoL7sH45yLYGZuxwGGrWf8R5gP
U/9p9cb+xsgzBpSK3bv0ygr1a71GBJxNpyTa9NuGJD3lwB3ObxV3eXg/dIPuLSXxDgyLjT+8DfgW
Rt9ahsVS3/GLgnmowjMMyS9EUnoh4M59P+umZduWpvBRCaC2FA7Y2W1uE9bqW8gCurtYZ0TlxzEe
aHD0EumIN9k7gsDu3AQ+dq5l015dpe9e9L2yr18UoRP71XNf7oP4Pzg6uLcXj+IX95SoEa1zODQ0
vXdkubpir5wtnMSFjL5km/VYXYadspxyyISP0G71JXW8zYiV5y4qLbLk5BV6HxDYb9zCskJLIUyk
+LiZ7pidTzrrHPFS3GaMT0yGRa9PrjjfDTAMDW/gy/DaDDCb+MR8xKK6cAWTR+zxmoP6fRzo7LAX
0VhsZxeIfMEN5r4/AxsBYdJHorPcmES0jDAUEtwVOw3+bczjelmQUdlUQ1Em64uB7wyWSuVGWvnl
YLFKj+vIYMk/h6b2qw97QdlANv8Eu9vYZbUScftUgZtj3fpojd4JLbYorxcNYP6AhBNNraQgcbDL
3Cczpx+n84oXYvCaazYGn5Mglv1FpmQ+AnDutRAd6HEOSonti49zNT9VcHzKfG3eCANCSos58tYR
5sRBoytEBOcsfAzE4ToDVLnvrhS6k3OSzgQnWeEK/IFfMmBP3gTy8D1QUBfWpm/lHOJVW8JltNce
KBC0FIncBbNynsICKg5Ht8bztMfqLfSbb1B5PRAF5/Q0jt18VlobhRBA3WgCem9v9al4lpfTKVIK
eghifuaEtHv5R1CsyH1wOZ3GFwf7TH7V/IUuLPQb6e6Y20ZdfcaFQo08ZpIx0BK+YEY17xnGsQXw
Fy2zrT8ZWf+rYB0rWJAAsFxBGnfSwguWh1q7xQw+oxtJEUdRDYe4ZVbKjTX82tJJ/WkPKzmDtfxi
ZpQfSJYJ+TzZPx7WJVOQEb40SJ0xsYfv12l8wEsiCZ6am2gloSuWqmHiMZbaUpy2S3BiOY1G6/E6
tLTVzW7fFYQ79jwzVksE9Q5P/apaihdHo4SL/+Sj1wfm3P8uroDn5WpvW6x5yEKZ/TsNsJD6VKEq
x/o1tpAXba8RVnAfZ+GZGxKQemMHrmQtTdG86RCmIL0UYPzYb0aB4iMPPUj/ooIz0kLct660aJLE
/3lksbya4fMmuu7ENC3Y+b5kISOnutxc5gabWHyaiaON7xULzreHLqF8T63KjB/5hewJqTI8WcJ6
awlB4YhlCDGK9rjZm6QrqWH2g8RJ/zo8GTWMvF3qsx0zzWJID9ySVl9Ye7Tv3GhMJ4e6cKt5ojM1
jfATGB89KD4v/XiTxOpKiIYMnIOe1V/TznPDQ4zp5fi7h7GrS8kG2Ewws5EM+VCYxYdAFsw1/sQu
vnUASnpUML/j9Uis7BG3nfirqLJKShrLp+cedDujXFvdTk50Q/IlO1D0O/CFXojh5a7dGSCDialK
4B/K9M6Q7eZzSisVdUQZ4m9Rzngn1J7M0fPqYmBT6H11MFGQbVd6FNkrcNN+XVNrkla7Xsmh7rfa
G4I+bGrpjwi+x5T3ijmXAOUpHAXgy9lErDDNusmeHQvyiQgkBmREq1QmpdDKxvVgFdK0xIR23HZF
b51aDEzSWoy+8+addrWSrEKIS3KZVodEFRezWjaQanQf7WxHF90vzWgaNF23MHAFOYXhzvBLn8nN
NU28mJBEGzc4iuqK6HLYLmFTWAe5XfH1smMba5eFLTMH/OwJRzntaEj6fGfkFTtNLKJ9kw7mnjNL
9rn7kFYGOkQ3lS6+sm2gBqKkNAM4KsngG9nAtuRUI0a4EVIVETynZ10PxnhdBlx2MZrFve9CRE/w
v3ZAUY6c97Disyle83gWadssU8z27Uiwb+V1LRMqVR3tEq3FqtT5JleeOKTuwwCQ1cfkX0bRbEGB
kaNuriN++W+W/8rWfWwme7sPgP93JTPY4zzteTslCChq3YJnVhzWE5DjJDmz5tIuYIqIo/iQu5PN
KkPv1oU0PKHAYMnm7yoFNE+i1MSz9e292Gq5kMjOQ796R3R/l8QqNjAi3bo72z+wBLP5s1/5uSTl
X7xOZ8s0+OKTSeiGZOXKmqWUWPGhXGMr4D884EeE+9rFxg/c/GKfNdFEel814rATkbFQgjYVQgoO
iCsMzOyySun2q5Vwe63YKEpGyNkCzTQh1mQnGU6Glg1DuaTRB9tfAI0QG+wX/J0w3n3AOse0ck1I
P8YngYQFPpQsyHjfpE7IvVISI3SCjfXxN+69yKWvnZ5Q1VPa2FpG5StFqtYzoAIhm4zla9XM3E/D
RzCW5tbNnxE8OconEU0+sv5sX3uGyrZsjOiR2fKoGxeyOUUFZHjPhQUh22w0Gp8NfVYpNMMIzRRY
vQSav2lhJU/uk0kpzzos1s0uYRWe/VR3R2IeIxTXvDQtw99mPoNZGNntnSbGDOxWTfivnH6vvqPZ
DrKB0o0mE46wkNmizdX6K9v0mD66sZl2aQribS1N/eIcFxixDJE1PfqG6FK9cwsz6YgYd3OPZlcW
pmHqyWgHGbVdIASpxJVOtI5fS6m4RqfGpLsyHtwamXpfIXSEKQ1YekEqult9RypxqfWbhRUhDdIy
sv/NIue0WBPoh3gd2WXutkc04nPYTeXIJZASmZ6bOTb+z/rxb48LVzzf4BBx81Xj+59x0WzfT5ik
rAMbYO0wjVP2W1s5KEGL6TfAc4tRalIaBHh8u9YaFMjn4THRUjzjIvk3ZkDhpcIfIq+uDJgfI5q3
B3kAyM0Ym+1q72iFH5Z62IE/K9EBReqgQ4FXTziqqtLjFrIkIYK+Ov8yBUYNVM3oLLeTPElNiRPF
LsGNb2pYHQCjgnQnKmhaRzi0LzvMMMVKPyUhARxgQRJnr6T3UPKetdxMPQQoTenfyZC4s69ubw0E
GAiK8KG1owhpQDtpwGZwhGg5MijfzZLuKAZDKaAPYiHyucn/oW7coi2LP7go0BpU2969teumzMsu
xyfliolp5FA95y9shYHOalOYallBC2A82vuOfSS5x5FGND8JhX5ZRBq4zhsSo4Ob0mGUr3lYixCJ
Wm0sgnANDwWvR0E9RcB344XaN5AGp4lJMcj+HsgxHRTOHZF1Q5MW2RybFKTy1XrmCKJl5JwBmpZq
1C+OwIu9dABYMnv9BfAvAwrxHEvIIAlkLG5ZRW0D4vYMBqQtTFHr/saWZ37C8Uvl1EJ6q5ymNoeh
7oJN2/QGz2JMhR2/PluW09xU/rKAZMRkBHWNU5WpGTgPdhU5NguOahWXLy4QkNZqZVhleOO//Y+k
jlkcnfuK4qLbzeTJtyjEXUg0omiyKtUKg9qTxtDXoRzjaMiaSkvS0jFBwmdalhpA/0W0oXF4z0C3
p0LGkCLsG28FHxMkOGOuPGl0w3/4qOdqJxHqVNcQmvkxthskOCU6X6JEl40AmNiuPxqsAjRblu4P
NKD5lXyatf63h7aOqX8wrexqxaBHpEKOHq0wMxwWq8KaOV2dDP7uJ3r5lAzpRjkGESDAX+Fd74oe
SeIcAwjayJ0oBsZnYeqygflS3jnt+wLFKVWa55bHqx0XiCmo9xNJeDG0FKkdfZEwUof8IgFeSHFs
nBj6kg5mOs/GaiOmqnKzjH3t3dVTSR3PYJLXMVZmdo1taSgbZ3XRnv2VUfZpifCzA0ZkYCKps5hl
GW0Zl3TksKPO0Ci9PcknNV/oR9hxuO55V3zjqDCFKI8O/kzNZZO2E4iZqXCzhltAOJKS01cd8aGA
vVC33dgeiI900Goxx8mD9GDkTvyhG0iiA5SaR+9Ow0Znd6JmJQBPNTHpFLoegGID2PAN5eMj8b49
ZVuhLw5SjE8C/1s7eDR8HodC4+4t55ivPL8qpzsZEJYGFaV4lRuRnVdoqk8w+5d8o3aZR/1Q/+G9
fs4a27sIdeLSVuundAzTQmPz+F3WVyyJCaCvRIvomib1P+ME2hHpqnAVvG1mLcLqvmQKQ/9jEdHy
aMCPSJz90/+0sQiNEDaX+2fyeYAC0BxWeEF5la6ZY/X90nMDA3F8SFBK2B71zKQZRgbiJIgf/4r1
keXdIQ9Nfnd6R33TPYiHPwZ+8A2H84WwXzhfeQ6cU61hzoL42yBECAYnUhCxeE4fPz4/9kL9KYR7
HXNVNSLwRUM3NVYxFuaC1jQ/FCxf6enmhzka+/T98XMkxk8rBMk5y4CEoWl1RKbCFSjN5520TxtP
BG99y/v7hhhJ/LHjRse4K5+HsKjxoToIdE1zm6RlURtjckDQjUwcABHMg3wdJId8u9bUu0lj2han
GUUwO1BWUu/Ss1TE7qy+bPg5d1DfCYD8MCyqAgTR0MHWL6npS1jXrlKeJTyHzl0CIUopFr0UARln
B39AGbxLZOCAOoQgCvOEt+v9R72IqIO+a+R8B/RGHHiHmlcT5Eg49uGIZDjEhUPmt0Bf0+LaSlNk
IxeCUvIsCDY/7GXo4EO8TPfTU/ETJv1vDxrkTOMNB8RJAThelBV0ohTH6QqpFMaxSg2qr1tSfi+5
YukDlTcumF9ARwUht2ZSm4mZvTzhUf552A+6WEZtHwsl5TBwgGgPpN0NL9DZugdEqO/mdWFe7zV0
QEs6yIiRng6KspKTUaI6IUvdx6VfLuLwIhfsvZaXeZLI8cVWHv8cSrrOBTHk/2hwXQIW3vWsV3jZ
kPVW5e+bVOi74u/nPNzSIgcIqVGLzkzk6xk/wSDxV3k8L5uVWUxbUiOko+LckAP7Pfa6nEq6gU/T
0cekzKJz2spJmB2/6A6lwItU5QXdbIMdMRrPyvem5H1O7PThIvl3+tBsX1kamwFSO+hwrfVaV0yS
19cPgle2P3VIbWbowYDZCZEpDs9wQ377u13rwgmDQpuPR7o5jBPjvUikHwF1IN0njocJ8fTXv1zn
lYWtvHwvXNGarxh17E20s46zohBAkuzEELPu+uv4rlF2HFSwuuRjmqdgaKNmc5iLGwEZQU91RZO8
w0B8r1lLnQSbJxQRdivhUJWjuKbrVZ+v+OGhbU2IM6MxDmpa1twQHfkebh/5cVMJfk0H/C8atQCG
lgTMRGMwQ3k0oe66ja9JqzOjom6P+xWScAeDVQJZT5xEao2gYFQV9WNBpglHwPQ3+2v3oDZeo3Sb
ttDHZIFNO2XaNLwSIWiiAZ/8PrUYPaqZcvJ27y9X4LACAV1aFoI37p01cP4BShmdvURbrtTLJSZv
OqensEvs1wOHPlwS0sLxlAXNS9PBo+W3/N/EIwF91SW5YQzg+K2aywWK/sgmSBOYt5Vhlg+BIC2y
fT8bkZL8/s7daIJtxagOfoHl7K7e7puU6QZKCPrMU87JBxEoYWWj8Jgci5BR8OKifEhnQNw6NVWY
J37lvtp9LawGWx+kDD9RRHJUz50zrQ7a7HQJOz9Z9BU27JX/QqYNiH0TnoV0Nka2KVhyWG2ODqa/
Da8hLCRyMebL+qaln9+l5eWdFo1TdzX4djayLKNn7xQRcsp9iMO7A4zwx8k7aZ6qpFEtTB3YVn+P
8a3VS41EHynhXCqR+6f1hRFBRkUx7jHi+dqHgvHPHMGde4FgWPQyjZvZErToXjgaK5HATpgfciT7
QGCvEjtH3dWr0AXM01aLcNFWDaZfwQNA6seleUc/FkCZN5eM87dCbS7UFBM8SqA7gUGQatvT5NyV
f1FEVD56ao7u3p7Jw+sfm5KBsKeXGku6N4V1TUCutoVaqVcuyVaRTz+nK5gwuAcsi4lh+N2Mw6jh
P2pikpxSjzdAv2qF2mQY4gfiiSjwT9CVS/6vcmJb5zNGV0cfmuReAI+XWHuOI8BycWKd2fa9Vd+f
2bo8zad7w5aMv1lZH2m9lREeu51JbksaV+Mw0yMzrDF5mNIJRqhZUMxr9U5gm8ABqSfqcOeAlelW
p+k8UpWBd/dWd2lcbFjUHmGcvbrnc9SE+oxTAbLQdso6fVUZvcO9Ux8sL4BdR0vkVCWQXpDQXB91
vAdSvxZBQX0z5cJ2a3IbjU3k7crVtDCgwGqYJIVwEJLsauPK7Ii4fOVlZ1OOFizWi6Ub9ifmQLAT
vBnhWebVNm91cOj4lvcUxxm1KhfQhAP/wJ/mDti8Z/UNQkbTIemlSEOcpyo+kEHjNWHKHv/txN8u
uGg81cPH9TPgAxVGYQoTM2bazKB7/IoCPgQH/4S2rsBM/WGp3Tc+mfW8LcACQMUJlsfBYZBJM+Ea
QwYqmk1cdo0qucxmvXzR8VDRUVz8q7O3V5fYidD5r1jyibVKeiTjhCN3XyMsR6+6JHpyc4EfEZQt
iLo1npl8dP2Htz/XuGy3ojSDGcxRuwjv68Z+//7kyuPo8rQMIKvvaKACKJ1NuccJFOPWkPDoRTK1
nP2Q1HBfaNFsIUQzuMZB9i1z3TlL6iH9jpfTkXB2FIvD5eIWRbjjn0I53oLz6Op3kwSu/6LwFGMc
w5tlmROaEAt2btx/IHEZXQ9UzaL31ETvgX5quwBQZoC/u+EOzqBPj0TV42noOvpI84uQu4eobSgY
JDuN/XOtCvxzTP6NSd0lvq5LmTEIBykvQlRbP3XMq4I6+hdejb9Xyrg5SvijtpxihPsE8qe5Aa5w
+47jcyOdU7mwpq7WBnBvZ6p1NvJpbhaHJHD2i22UWHb665MvCsnxvhuUUVV61BMng3ogyz92+taY
1hB+Sw+/V1/bd8jHaGr7CeZEjt0i+H9+qPLywEDlDPFKvNa74cr+KPMaRv5EMONjwm+2T48/9ldy
bSQN7fg1TIX2Viv3fYnWHPVk0sF4f74rmfSHHUCvkwBEIb8smcdMZKDt2nHEkfq51F+ADU6LoI25
7cYbuOgkr7cDTfc8lD9TZAeZQGhetBUn6FjFO1qw47nva0qI2G53Q3vJxjLMqPB0XKNrqKo7YLYf
ddetLim2QQeiiYP/Bxh7h44poOK6Ld+nlVzzFGrM9+4rAKszoFs/AyNuS9WihC2uGGwY4BHZY00w
RW+CqrsM/fvdgy4VSYJpGVCGIBh2sAYpe3Jt7hC6UodONbcf75pQ0/f2zUiRTBKNLapej/gk4qXL
M39E0zwHWCVRLverqFCPNko7pHgivNVmVtmGSRxbYWgExWMlueXKaJcDhF8zVrBk6sle/e6BNxt3
LKjmgEpns46C9chcdY6EwQsx3wpfHfm0wqYT5ra9DSehoxujSCuQXXXSDEJxgdsfk8d2kfOpFER/
Mwu4WSSQlKU8xHGxj3MIz2CXP5Koq4hO9zZR2gHjqMSWjlAmW5WsztickzjtzURNEl7hN49MBm08
Jwhg8NBW1dLThXLaSQNurxsAQIA6ke2L4zjJmm+O6FLHGGENQmJdY2rG/Ne/ah6C7yc2NcgxWk8K
1HZrHh4mP/0sler7OmSOPTXBOncC1KL9dgWK6RYn0aqWtvPCwIAWIMnl9VM0dkExT3MLdDgBCqhU
ln11lhjSFgT+fOF7KRZI7A5ql95wb7x2Q5UhZVtQz0VvVeOvYAXn0lGHweQAoZgQe6xeaZVKW3Fk
vYmzsvjxOB+UT8LSRcClOEGPwrV92zu51V65UjhRuDbYFmlxWluldjY8KDYh5uSff6JIY1sDZUP3
xcr4YAOlnbRxZxFtmit+7iPelvPYLfthX/dgsE1GLVmL0iPVRR3UkliZJMo0pWBwYpc2JwDSHNXZ
+nioaDX3FKDid3yImXK6EXhGdH5irlCPLh8hZC8Zd5DnVQuN8Og9UqB4mZIkfkW2VqpML26yPEUt
eHzaxnwIvoHtEwYOonkg0P5y5gCE9kFwfo61fx2dNNO3TLEUvXLLeXG83pyvZd4I7BeP6BJQ56vR
oezr+A9le7AWCYoR9xzzWg4vErR0a9a84jUKQwPsGCx0kBF12QHeMrFMgbpyWk8XA5ajU2o3BBct
P5ntAb7ZH8FgKqITvSJr4MyaJVgSh1QoPqY4IA+VhGxz4JheAFuotxHp9vK2rYcuInK48z9P/emv
ZbYw1OYImM/uIM/BQ0lQazkEBTxV80rY+0TG0U4fH1vMkaUHZ9Ywro69jCLbg39GxCni1UOAjZpJ
DgQrGPwJqfPX4BrV1V62z6SS9ILN0WXv3Mf9+vgcYBcSfRUAlQUpOZHKUK+7O5ulFJCF22UQuxdG
w0BikEvMKkWJq5VtrsRMkvJWoS10wwJrhZBc5mZGTcVnaUyne6PNQ0goxlh3s8WN2Kd7r1f8vKgV
BePLi3ZWQTawdWRoJhBr+PzBiAnt+nAWjcNXUc7eDtttB/QyeYXxE8n2pUt69mi3YDsCj6BWNMZz
faV3kC8DEBYbTC8V2VDy38EqzDcDBK438YbaH9NwfTweV4JgKhwo9dZFUGvHwO+lIrvrSxLKN2Is
l/2mf+RmgiviZIc2rFcsp4dCkS+hv7StblykrSGdT630VrDbIm8PZmqG/c6TeD4X283hT+au5mPW
iKJv/YgqMT+qBX+F5Tlt5ilJRlaNP2Dnvbp6orAn9nh/SMWb+ZrYmI1I+v5/kBLXDjkHXwbqFPW9
EBW0uEI8qi4EEFW7c/IM6lwOV+Ayq2A7AmRqXFjI/ku0LUod+ZiF1cO2MFtiOAZwPzqobvype7eP
/7qw9R8wQZ4WjZcfC4M19MWsNVyT7oCbOdXWXPMiTE99oJEnItPNyXmguJBFp0uNqy4ar41lGJ+l
Pyz5/0Wheh/taVyqmg0QtkjHhZ+ong1uaKizrwuMGruBCbcABP2IX6s19+ED8Cs6mnMu4g1sPNly
Iqp0MSILMc8otF6C7+qV9BhnQV6UczmikBUxng+22fTxCq0W3zKVT2tDXoXUKZWFDVIxeRcLGo/a
LlKMynWvYYoM8nRxoE4u17XC/gs9ONYrnrIx/tJhziVqg7eBWgApZ0NchPDP/dZ223FpD0gB1JrB
+8cV00VScq1y3+NEnANOjsRPwi/3h+q9r/5MUfZ7OpCFYWkk3BtGNhnyUglI3k2jtE0GpIYxOlm0
E5TVn+DPPnTHaedXvhalzvcb/4SmWbqrCwIh/GCq4++0dI5STqJrNESOonaUpK1ZRlMKEJjFrHrX
smUM6yJFodXJf7oFIpuvqt7Hy/IA+Ok6LrJhcS77HPPqw27L6iovY99wrySvEOifnXB8b+j/z7/7
umQZKuRHb+RzTLjqAizqzPgSXmOSGujPsB+ZVw633ZLFlUC9i+dPxNzrsnhSPsaKxgkYrerj+BE/
bgt3u7CD5D+7LEsAAk5/lHUteTVCtrGQ4cibhr7S5z0Q1vv6ySXMmzyPZjyGwsY3zFw2oasNFABI
xxTkjCe2v3ta/FJA4vUxZw0+6lRuiYXeKQ8JYZwCPL/TzQg4FWXnu64Q8Fy/6CwoDwzgeepWCO8b
NWwur/276lolVf+ty1p/Cj9xbHtR3SU9bMfP1AwFWnmPiBSaNzq7PooPw10A13L9a8OXTJidYTeB
r7kJQFp1WwGzYjuw3NwXy1Ccy40hLgk6co+6IkBJ+/Z28F66Aq4QgMzjOb49fkzE5O7AwVRaEXe9
Z5QmVGdZy6N7pEdf4b0dEEGwggxACqoZZJeJ9Pe+isuyoR5Ec5ChmjyZwpOqBVYzfiE0+MVUrPvK
3P0yQOxCehcjLSXD9yeI9ljCU1lHJiw2Uzbyz0l5IdM4iEFt2hdVEhiBwOwAgW73K/Iri2cTUn9X
JwISE6i88jW6QggMccyx4SdAOimNFaEQcJ8rYVzbaUlXcTVfI9DFWnuzeDfiD0oKdI3/EKJpMyb9
KNNJakXhLHiJ8CKV3F26jjmZ8PIhqJ0eDlIkOKPcWFhz2ESchvupysXyO0hLSTT2AtRQ5otFyEuM
ikAEz+igxqDy5zQhuuPNBHbdTpnq/bqm7Bm9YNUPhYF2G4D8Yhft8SssvlhaiLG4qgMOP63iHUip
ywLynhctYOQ4dfScY47LpQsMrhR8LCPQDxTQMITWKa8ybXvcMUwYl5/WZJE3ttlzy1w/B11+xxFx
/rVhXWrlQ7rNuI+BDds78RjgM/B3IScbHVn7zl2Fcm7/K6+Lq/F9G8/xXpV7V9ssjmaL3idqkgg7
5TAml+9v4WjKJnxRJfQ93JHCRwC3iRBwO503wpB8SOlrEdZW+3n19y4JnH5k8XcwmYGIe58oZAOU
tpDT5dJeBO3M07W1xvvKARL+Y+W93lKF16bPQfeY9EBgrvcchCpAmpXtXIy6zFnHh0ybUBlvCRBC
f9CEkueMTAzwnKXrG+HQ2RHMi6guP+mUtR0LaS7dRMz4RJJ3VfWsuTV8gw0MYuzRR2XlLzKycfpU
1o1BslP7gdLHdBflrVftmEwsvXJy1tqmaWW1QPww7smcEmMm+0WasxF+Nxvr6ZR6zQ5rqfps8kB7
w7m8RejFFCzGgwduAPwckZ8RPTaRYI5q/I4WqPKYQd6OqrtDDU6AySEVa4bT+1Q58TzG6LgEfvVX
IxEa1SEoMEuM+o8RLPsi3H+u3X302Jdg4IQEKXongFav22LQ3dE+MHvhdEwKA2TMNjb6Iol9AowL
a1uRJFt+7X7axF2ZTN84rNbwXybpLyxEYtdOCHMw+oVu9YhWDe+3LXZy/YraNuxHHhbH3+imx2zb
HJ3hag/ZKd9tpXSwXLP+z0sNLhKAQK0ooMroSyaRXJ5V1wc30/tKMMX/b5yuPHwd8S9D0DiuED4A
4vdBh2HG6wHyU4EW3Pl/DFXVtGUAhsrd5cd8amFIktzKgENjQANExVUPNnbQhocmHhw+iGHrwoZ9
E2udGW55oRljiBIsNbHG1riZhbEKZ/b9g5Fdz823nd/ro4taizxxrdRS2kmE5mwd4JalTGBHcjZP
hh234I6STr9wJTB7Ie86K9IHr1LoMvgdZgPGHfv+BTao3zY2vdciH9zIxZAvDXfHLw/9y74q3Y2r
bi+wx5hfSKZZccu8zczQt2m+rD3IQqlHTTlLrBKP6Y6hNKbYb7Z/BZ6qP+djN90lQCS82oFZnmeS
u04ETQhtxroXsyt/pxF2gKCVqYj+aqzuZD/x50vXX1EasIcgcBjxZf/S7hORvucCu0g/aTnYHXZo
F9KXGCEqPB+U59PTeZ1sA4foPEtp8WnV14MwrgbrNne/kDLE+Yn6NSf9HVgsuVTIoRQgYQxuVgM4
xS25msBoWp+Z5UXMcysou9lnGEq4U4LuFyw1UMYpRrFVw4ZVeoXTMifuyR3ap9OqF2+x6vNNW/hF
mhXx7PS/U3AWkUoUXiBDgC5rWdC8+drvHEXpmv4C1MX7jTEehr8AvOL9pwl573AUx9uvP62J/2UL
w62tcwo5Tcbv6Tbn8j1QQJWvFuOhIXSCrfW1ArNPo05C+C1w6Kz3drXOvSFnJ+LZXq2h/zQZAwqV
RSaTryP1/jhRARsbLLi7wrfmRMpgPaQzm4q4suDxAyeMtOo2riQRYBnAWduFMQDa/3ZoP2+U7Bp7
0ZIC62pme54RXtwQNfT3Yy0asweZ4kAEWm2vDw8lG/ar/19EvvRp0witJ5U4CMtSXcUYreNz9k6t
srCQA2nlxI3Ufd9/lD1X6DIx/dSieXMd9qsLp5pkbJd9LpMy+EyMlrUxi0Bv7z7HLJJcRy914ALV
Y+ogF+p4GMGvg1aZ2LJjzSt4uVvGX/v08HIl02AcHv2PPHbenjQ7Z6nv3y9weIEgW8UopXwB9Wa4
LKGdi7ddtIOmpH4XkUtEpxW/PY4xmGqDW/KYw3shTVQd2dKmrtFr4L0gZLWtR8LuUZV7SRF097+X
ccCroO4iqT1eGljD2cmWoHLVC4NOmYqNxmlxQHRXdbarct961e+N2Ay/tfgL6j4Ebz5Cgg5r6CQh
3lZlvfZcvotMo9hv4ZHlHTT1tjOaf81OnoJiXvwODLh+eXmNGmAMClvCPjtB4KFwNXIhHI28DWAq
iJq4HthD2VEb6G1uH2k0Sf15hZTahcMQ09nFHUA2khnrijiIiAM5PVGUvX/x/GAa33oJaBt2xQ17
CzRFKUhNZolg1M3zuKFWLJAfVoOFc61NAQsxtvdMxgr4d8zpcq+1zleE7pytPdsUPtHAi9rXxj2Z
j84CPn7UAmi8Z5xxPrpyeKy1E/w+6a3VeSgZkJcxl7VbWdl2s7/O6nzsQ6x2CKpDtc6zsWUTxe3s
Y9Pftx/FvClcqx4x9oofJoR9mFn/8MZDBHloEdC9dI/DI2BCFWrQwkNcEp9LB3bbstSHh9PHAPbg
Ye4hKEnL3U41jKHPnCFHqnDHihZoAX6duPPhvbJQ/pk7RaSoWP4R/I9Op/VyCCu5v2oTFEoMhz7U
svfi/KcEiwOzGHiJpBajDfy5sGWzlcjKsGEHfUVrC9zxxddlMUXw4hrl+0fcxt65AggFz9NdQOI6
nfVzs3dS4754MN+ntP2q+fI8AGJuqBTNXoU094FUC6s8iOYxJ2RwNwwDmLzpnYHqUBhHob8ek4s8
SyxYnLtLayOm4ZZuC+QBBFLLPbgckOmsGkuXr0PPiN0dONANxGfsMniNqGsUXMfKzPEWJrTyyqOK
1H2PhZFx/Ex/iWu0zbmMR0+xMKroi1KhJW5YXumfJh8KnccQk8MIRv7gJBq29wAyRfY2K5nBux3B
0pGpkUF+rDQMuTiQ2Dq78mBTbKDCMEXxIdQPpa6XvDU7Nv5SNovdeuI6rwjlbgtrcujfje+0Klq0
jkeeOKN5WY2W1Xq60JgOayWkqUcNh5uYLyREcMPDZrxjvfUylq1PB6+M8dsxEONxX2+GlpR7mG1J
iy7IjAxk/88Qw2A538tI+7sxZUJbtEhqsp0d1fcBO1sEen/tZPrNuRuX/9hszITQGqIYD+fDalB8
X5zwaVFKRbiZLV3uWHJgMsHctkRul+Y38Bgc2d4r9Y7+5289JLA6tCb7TJl3iqDEWB6uT79eDlL0
G/q90kwxSHweBVxQSSiAJKVcUz+Tz+OpYkDmdxk6/yfDkdWJKb/CmJ6gpuycjQx6vYxys8epIimj
dMG0fAUMHgKuumz0VUsvn5/DxXgGW/jpJxYHWSVOjoDWR/K7UGF9jJiW4R8xfX9bR+RMo62PN1so
+RJKhPY/lq10svOeAn3QMFqnezDjyE9yTqnj+12zz/ufZGp9Qi3UmbhbqTEDsxrmM0Tw1AmS2mdY
8L2zxF5YvxIYReHmcUkr61/4ZAoO2RjyuDRzFU/ORT93p4q5vLp6EoCj5LXTP+07Z8miirEWB7hH
EQ77B8PM9HGy9TD3U6+egodwl535kojDyPJqCBEHExL0szQ71WNn24AnmqCWASS16aVQJHOM8ELk
Y5qUaz67I9UbBLO31V173sF1S1ktIAE6vcJGiAI8T5Xd6ZqA8MougY8KXIKhabP/444WKc52gmDk
cdWZAZspj5TDZAscATJ43u7vyklcCaDeG4gkDbnBHy41cJ5h7U8spFKPTNmVTOZDKeChIsoEPGHi
olF83muDHI1dSFi+yoRftSbd55PA5H/O7E8AFme7hlzJf0xYkzZvi/yj4PSqVg02FaRJ+UA1JtJG
yRaXSoE7mdTekLplhwoGEYwjNGlWgCqvGdQSLquNUZ4AUoft3xzEiV1cjrMyVdZHf0TWFpDes+wV
cdeMOvAeK/gYHVV7jC6BS9vqfhZeUBX3C45smIV/ayyVZi1j9Uu9+zhXOKMZqFda3BmlbCmMDRyC
zyxWwODjUv/BMMPlSkpK/NKKajywMWdokUVa/S+mIftGTsAbmuuMHCdNKiN6ZtHt0ty++dxCXK1p
y98+JctFuNTcP9Z1d53AN9hZ3bbH/VM4ZsmL5NTb+6sVIe7nNOCnHRwaTDwxkdwAnSxTXD/P3K/J
jSpwKGXF8fH96S5fWo8sLYUo9MJJ0vmYQxD+NOgVzD5IgiAI2YihDW9hdHzY8maOMRVNC/DcSw6F
MoOwBDe/IgVM5Dkz6kIJHFcvr6oGB/Mv0IoUlGJ9VWmIvuA6/ywreKTz9jXQNqJLvIq9f8fAUmFw
JNf8OFvasModp/AV0+rFPkEPt4B/fhXiQY+5fuuBsmHP31GcvaY/yvTY6+eF7DlOeYnfpBufbl5z
xD2D/x+3+/zlDnsAupqptOK98DJaSOli4IHkJ7xJT5qBpg4PioK18rhlqIO5Fq9TXawj1XdV6aVy
/sWyxCgGZtbpWdTH58vD8apnN5t0BBl4n6VZuRDsAcTDQtOilfr5N1GpAAxI6BomtfYaDyuf5lwy
ei040BYKt+e4FmOrvftmIxvjY188+Vj7xzRN8gPtzfq/ahOoqJ807I9uZ0JF8MRxtgRq3XVsfTAR
yNlLuSaniRazUaDvq4ku0bjlzdRPtmI4ibjZjgI3n0aC4hQgjv9Wy4nagLQe+Z8krp2f6AIeQX0p
4JLg8vETrIipqqRplh4mHQvYW7fz5VZEBGnmgintvR0EyS3l8vx5MdX1ghEwIrKk6UF5+Th96XTv
YLbEdwm+Y/n3nesOkyAFqgEy7+tW/QZxAvfHoiJpZ9+hY0dLOsGI514TDNHmsDdO17icfiKy6uaP
VWnrfDAEqnNm45Y9yEq/ukIk7yC2wnAwQCQd9jiSOIZyp2CiY5qSJFgNEZ7wrQaJN9XvKZfsi8jN
tM9UKxRBrO/xQIuiuWeQVblVu7EQv1YcB2jAADyzSPPl4ilm+Yc5WP3kLEfGhKxCxWO+8zGD0eif
emutgWg5A9GYOfqCx/QrOZWJdXVS4ICzbK6CKZv64VqGid3vq1HfGU7R8EwCWgb8il1vlBeHpzck
D9OEoFVDqrnAK7D50u1cQbR3Q1DfJ8+0GtRvDVKuhbd15CUXtEnXtVP2skz0aN4WazXqGVXxV9tD
eeRqfx4ij6Eff0oh7usO4JSobdD38bZD5dvtuxe5Vi1UCwLc/Kfmk/U6yHuIl1McCGpiqUlgvvZs
qoSwfXFe3QUrxG76LuTkUzFWwKKqZsYT1MpDg3D7BDydxeJXm1o6Vq+nkfe9MZkkNP+VUJgmOQKA
qvEWQtCewWA7r7vnGdT+Yh3ao210QPcf1iBynm1rBR4JTiKi+IBgNApS4UOPZRhMkGYJaqw7Qohm
5om65vpVlEEGpYiWVtoMNXMSz/bLElIrUYcdOqHfD2AqoQjB4XDoQxR7PhJv3Zeda2m0ZW2g807k
MhuzKcJAzuwcJo7vgABUFgq8NhPRf6CDfIQUnXdB99SR3YIvKpgTHkCsVLK6hRhnxtgynwZqed1d
M/+i7WQJ8qAY8947pAHQwmfJu0mgr3lJt2+0hLKqp1VDIVBciFgwfN1On/bDNw53eqlMHNRSSH98
nG83225/khG1EXcn4cv3OXx4NBWpnlsXhcsjG5gAqNxKC83M0wje8nxFxfDY9IOohJQdOuAiiOL/
TEpiwBgGf0DsjFX4lTVohCt9AAEKvG2RxRlrVWrHRZvWsiffzzJ1B8bC+htoKUl1MIJYuRNv5hTj
iaX7pZDMJRJcKt8AHW31rNgXqDAzlpjX7+1PSnifneZWbfPWm8IEpuXoUSgqRIjQsdR6WGrFuZLW
JyZEFXKzQ1vmZByr90hMQttlbQYC8uUIw3RNlIrDnfhrPetisA+EgwWc3kWdq203h7ZH5ev6xbxC
eNuzfN9WdU+GR/fhR4tipt7zBAyNc4Cnz2s1JOYzD/iXwYMw34PGch/06HTdUchNZKRhe5F3ZQrx
f2gew+TbzjSzU6t7gYwleIHTSRX2lRv7wvKl4hHhx8xzQW+cRMNMAJinzNqJp8nNk31ZwiMPvSzC
2KXecKwataiGL93Etb9X6Y2PxJUNTslcTQcYsi+jJU/FAWam/7cSGTC8c2DKtqdDeypQnvcyVcs+
1CFiLu284nGm+jsZkj7hdP79fbDKP8+crb1FxrVFm+Nf9xkIVckkBkrLs8W70+SjMe1f7j26lPf/
PxvswxrpmFyVjuJRLdIvTriXRV+xdAbYOtVcouaXJz7s803Vus5Qx47nimHWsXu9p1t+P1Afbady
7pfO/GozlYjDHPhpN2pqxNyzRNrqUGSma457CFikS0Ppw/9sB/YVKq1q4mVGH32IHZZ7TfCsenOw
RydKxiGR8rnFsEcxRSrPZU3JWH02FFEGKW8gSzSGfSx64UvDEdbMSKkXz3hm0ANmSTPHyfHd2oGr
6ofdvmLT/hUl7IX+l4sTRo4duKv1Cdenv0WptseYe3qaAUevm4x1nebu6mhaJ4DG3pTKZqbvuOTm
FvahMBVO3M5L+wvfpmz9YuqwqqKOESF7V49Qv1nJ7u7IQKhO4P3Mfi+tOnE3JGnWQexAIXFatyn/
QG/px4ceePCLvAFjZW5qs+o2fK5v54Wncy9gX+0m/hgYErfS15FfQ1jZqgQpPguX9oyBG2o+k5Wx
CNFBGDXW0ZalBEUsljWj41YtIBUNwq6G108q34idD6k2/ErpzCCWogeDlhy48zpG6DGmOLvqSX6g
FQHIki9kCQKB3xVCpVL9WwKMkWA6l7MyqxZMfZM3MuX1k5jm/ULaCtkW/4DkV9HwHu/SoWAmePPc
9HpTTQhD/8v2bE95iGIjzJLzQyeSIjOI8/42GEAVGlVHn7F15IObHW+mBjkckfH/zJ99212fGEku
/CX6DyX3ppZXgAzm5fUSBioJ3WOoDJeO4twEYOnApWe3/WJ6uf4bRLP+pN514N6zNgCKWUwDRW12
zxajAmvBSN8y7/5JIU7CJV69OPgdd6/00aqftcgIEFeATnbraSY4ZBkw6ZT7tq4FdF6mbJsXLvKT
+Drq6+ftdH4xyU+Elr/u0jykCD+mZXJcBXVd9IGC+n7+nlEYyh1RKLoaNIpdO8YU/W0ut9TgbfxB
WGL70jYTKrIjH9bTCRSBs+KROVDUMdVl4gvJ3b3A0leLvGmvWIw3eF4kQs9Qrd5nw1Ep2aeDBmIH
8CkyqFYv0RJ6Y5j7o8NxWj6xN84O0aEUPLrc1wigXGtThOtQuAmd2TMnWWwy8XyX4rG7GbONBAP5
z/xVJlmmLhVnpgHQxI+iIv+p5duc0BO9dOiMXFTKuqNJEI6YMQ6rwhtWjLz0DkyYqq+HdcH/3fLG
JlKIi/uyTxqEJuup5Twg0GjB5ZdqIS7aEAoU2j8coKOPW6AiEK1soDDrXNanCByTXWhtK7hn3amX
UWNqjfUqKpo+C+habPKzfaEYOzrVjH1XjPkPB6xH3go/jCw34bQ96hmwdPrQc52lynFZicThYVJR
GtPS74Y5NzgJIDKdkaro8LlnQntRj/0FCXnprxc2tgSJjs7BrhpSSMgk/2Lq9pb8UoFzj0x0sJD4
4IAa5rAHJ5dHa+Ri+0Nl4Rzt+ZiUs83P+N7sy+eRWdSIT/p8VgjRA5my8ExR8Ta24Z7jP19BjvmE
if4XZYLviqgmVIFNnUsxMZalx3X6SGBRzl2wsdTF9lS5uHpBFtsctLkAMm2rmoWcrkZm/kU5IWnL
xEZjNjjZptZHcOgMJhTOzHdqkFEJM5dW3d6V+hixyP7tQzUbMqtFwZ29+Dmk3dVASnUHIZqUjyT+
edZAPTnTkLO+S8za1K3Of+iNBg4GNeJ2HEoUNqSmR0BWN96Fyd3aM8WgaJ976D/H8oUC+zxuoI0+
kWojvN3w4gU/uJNPepXWrWEtAKHNsO06dnsRxY5QE71JfQrW4YVd8rN1XCnoO9Lo2U9yETMXmvB+
P3t0sg+TUYiY/xDycJOi+pnmcWc906ZhK6/oDFPBPAOX8nP2a7JtXN3B2bL0Qf3ZX1uQX+5EnYya
KqlEg+gmfwZk+S3cGQd9oWCo0xugmAHnKNOgXRgpqhveDAI+GmbfjhKezZXuY6dRfINhMKAtg1a0
TIgKhCReENSO54xPHtdpKMmyaHPoNd5tuE7oouXvr/rvaLXKxtLSJcEl8u5mRra0c0kgW4YKt1Ne
xTY4/eAAkj9XQiVvnp43dwE93YXQFXfOC2J1xepHzoKNtGob7Akuz6tUzm9iRcT/Ntit8T+by7Ur
tKDk4rImfjos/+79CPIqJNAt0mYcxlaW2uN+EhlR6QxXDu7MSw034gzRzmO69uOFRMx9Yz3T7aqJ
N14p2+lozzzGLDXLnW/ajrkiV8Dri7fgW2gQggUCzyPEXSF0YUsL8aMVpus8QUsFs5JE3zV59u87
jNfzZ2ll0Yw9SYGZK0zdlT6kFDf5L4Drx6I2/kdOw5lDU9CLxDJU+V2DlYALJqM4HLPNMg8CMl6C
KZPZOGrqUDwgGNTt3qWUNHg/BwLs2zcvcG/VQIyt8ASpwPY6cQAArktqqz/XPUETpSbdquss/27b
WNCYJQfdcA4YUicUc5jDI/IgWSQqBo50B84PKBPg79TUTZHIzzbzo8sja3tQ2dYRjYzrjbS2d54+
FZ3yzTnVcLoc2TH/YceGy+as+zzGs7ynIxSL2yHdPvjGfJPbjUmSOgBmbJ1UtiIYfUPil/MELFhT
EomaTsjB7QrYXERrMN67pkVhOLLPPTS/nnRTig2de6eh7GMr6qsATZfGvqcwm5NODem5AdjBQbGP
HJ2GHc6zQRACDxzQeOvXELv0z/UzJ+7uotbZESg/X/WEzTTRToY95uywch08qsCgdlcLbfYDATS7
tRaMT5FItsSqdEoUZ4oyeXIy/wE3YM0pvUTFG726AszMawziARI4px2KyNT90l2iIyq8a1Qiq1zD
wZJExEIPjYNrtFoaIPuPrK3fMN0bP370hGwCmLw3h7ptLzdtP/FhGuPDFbk6ElXm8bKJfv0jKZt6
2PjWForshs0hb+3HLekrUgINZz4J8jP/c19HTNB74nMqv1NnAqxpJJmPrOaQCnlqSYCE1mES43AN
HLs/dIKih3a9GtegKHkR+MU/xtejkGEzb1Sep3Tde119awZMuzQCe/KFI4UHdugoqtnT/GjVG5I7
1f7apeJnyzVTi0A9deh+tzpxFSxQbOrXXL3gpihG3TyGf42MwTbz+i/PeHa8RerenABU4yG61qx6
dCvejXA5rbU8jR9q66AiNudZWFJbiqoQ1LMS54dzYvWJPeS/wZhZC9Se06yZW0Ad4y+cfwk6n4TP
0b1wXIwIAbXH6xlxI5KmhVM8Bllu/pmIX9IAAdrCuxwWYNDjT05NshyD6K7r06lXrQbvilA04ZCS
omXc+rjZwOU0eJUHZUSU9QGoZm6DYyw+XPKY+5CP0t6GAM6lPeI78yzNeR3+TCM5GrFTi2aE82ll
emH/gYwOO4qJBbb1N4pQlzrlzxr3rutnQySceSUS8vkwaHRzx4ZoVxNkXH1xMbi4jl9lOx4PFCWt
/wNGj9o1sm6tUw8TLxFgeRaDXOP54FqC2/focCtdSHTCMJEyq/kbA3nD9UWPnZfGY8I95tseaEJE
ulvQXVK2U4e0rAoCsa4BvNPV6h+xmJPh4Xc3zdwmPqcLqwh1KUy8i+5d+MVOH+Mpn1zK9u2zDzs/
osMSZpNXVxqjLdGLwx9/tNnW1TTzM3a5k+cgrPodX0F3TgSZtU1m/xFd/I3BxIYQCN5NF9NfdzCW
3bMqlT32XMO18ttvrWmj4fCYk48jksTAE72KQz7fKBZyNA6HeFJoiTYAmH+zIobAUglqiUavvkel
oeF5DiMQdY37IJWTPgtDe8ig+l0eVh81U186vw8Xi2tiZxtWbHYa8Ouhzt/ZOYcxpEWJfUqjWY1d
Dd0atvwYxKYcgnPBVtCDz/yb46FQyHYmF6XS+rVCiih3UISs4DuR6Dgs84m7VCVy79oncJAA7Pwx
wwEtkrya93H2aFBFNYkRBehcm69fL2+r+mpER7LZhl+rghQ1ZJwl2o5orBo6JfaPk6R9yYuX8IRy
6+vEZA1uH8Lvdbx3WuD88sIdsJn2F6HkkmUg7iQ8KkY18eub4eQYc5YBVzeT9H+S2jtbHWo97KE5
mXoICot/N+j33O9jRVJDAuI9DkN4yipw7pDQ3QfCAoyTDs7yweqUgJSm/gK6mlxWHioxbRC969u2
UlKv3eqaTfMdguyGJgdgBl/hIa/Y1U08y2s2YfaM15I1zj1RrnYDD/YS8Dv5r9MKuTyh9NY9EcvH
4mxn8SjsOAMa9B/5Safw6+IgKuNPFPYu3RS/SmMeBqg4j8fHF9K3gpqmNDBQPpxhoSsDE53S7Q+p
FCp75nFoWZxRhSgrN22CccaFIjX5fnPq6k7sw4P2eSknY3dWowZRqCCcLf9NQ7OYZyHHof8NU8Ff
SAG/8oNhyqpjfqsdRRgEIHOID3uWRinQ1ce14oVohcxrARlaiszIT+O1a2mlsJkK6qp4E+e2mIqI
DsHTngvo9kBDjU8/rVfQxE8mfeZAEMzCAAO8X1dwHKv80En37NTGc2gQz3GrYdRdOZ3n+MO498zb
+juEvPT16inHPEfbMTaBkGsqBFdlj1gssxzmvHKl8a6w2pdkaHkd45mIxXePJcnc90K+n1KtIKDW
tmHXQ3mmo3t7uGo7mR88LwxKIKAJZ1jfly02EaeOaxlyJTLalL9t+ncv4Ct8rhz2oVFZRVPlb9+u
qll7/gBDn8vhTTzB1k9Xf73MjBS3GTRe4hDbiwKQRou8JjvCjWlWHHOs31u7zFwxQnHTTonRUji4
8SemA25Ld6OkpJPfAz7gBLLtRzTxLUQ9uQDLiL7jz5q2lR/vl05t8uKluDAEpqOePBGzUgBbQcg/
lvXD3GKffmm6FLOstOy/4lRTKwJSIghx78c4R1ShHwWqWx/+EtO1+oEJnH9hry0oJ0K+wX1x846m
aUNX158EG6k6KmIu1HqBMRX4J5EnxTn4j5/QY41E2fJhmHR0K3PvkdJGuJVtpC2NuAj+q+/2g7Mc
tKeSnToBo/7UUKWkqF4aF1kZPsvRTVeGFFz3+mX4hKYRY/bjJEvSD9K+vQYQWnfV+PhkZHJL1bmp
cU4YMdzIWjLuFflth9iUE0mnQJQSnRIjLJ3dVJ4/eSsurv3EUpAveShhN+uBs8kcr5ExauOdEOf0
k9OjCY6kBv8/NpYhacAKWAnfpfaM3AhvFbB4bW8fMGfGkKVxur5I4abr8i8YB7k9kJHj3RFAchlF
MRgAxI6AWrGbPIR5gYgupzPn1pT4rvfxGOD25OLlBCwC0DXim/Ugozw9RZWmiAvFqxJO12LDWHCJ
Wg3u5DItXE7VGOrPXjeUjY70NMYuTOftx3uXOMN8I4oThk6F6ezrH9bz8T0zJhyEr1eevYVFsq5S
IbHt+sSbHPYVh3p78+bMy6tgbjNGHj9i0YT5y5xsJPVKrrC6MlN2DNGSu4DC97xMKADp91FS/c1m
Wo1WgVSFSIJ0QXfF7UVQsRinSSVV6SZ0iXR7gW81CcabUCrOuNcgdONW00PxaKrxixs7IeKG7EJF
Z10ifTFF+zP2QtRiKtcgIR5ddQj+ro1iT8fXMGoMQtJoonbTFrFWn59CR/9xJCfCRj5KBd6Z3T1d
GAQGjZcX1W+ZL5gTzSAk341ahbXlzjbOt3rubrQnkO7ZSQOAYeLbeiwLSJjeCPd3LATfCLnt3mhN
fB8Iu2Pn3VAhgFjlwlH2pv/SSGOWXWPD8sjWLRu131kjND9/ucV3L99BoFCwLh7aymbd+koEY99e
VaCDzqMkX+XAory6l0j/eHAR0ZRszeYrjTvLUwyQbiYg6nZjEqWcF8ACYgyOFBWNTTd3s13A/DRU
ERwyyy+Y1vBiyO0JFz2luwoTxMaGSIRbj2z/xqrdstKlfWFRGljT2+hpUzTC9bLxTHJu+z/jz7Cq
HR8cuFfJFaF6sv6QB3wKUlwl90EL6wTgxTSzmxSaHTX2pBbQdqzcgwUP0I4akS+uEOZoNUJhPYB5
OKPiZEwwjoZ+K8AnDsat/XRbBe/597XBMbrmsA6MA3HhT/You5GM9caZ+rIQmHrBk711egnhZKBo
omeBdRCDR3KQzwY10Uqul+yfFpj8RTcNEkA3+pM82rB6F8Dfs4zDN0NQpTNIHCYOjF6Liq2WV/bR
EojN89EGneB9CZISrsfvqoFYZlSyee0huxuWG+Bq5OdsPHIhcKT2CkuFPGfbJHNAda9YJVSyALYP
nao0fCxkArIDaxngP3SaOtL4rdrm5tBaYyO5RjI5Xunld6Fhk8x4g+r04l7MS+8QUfljlc69maLB
bj4Cj1cL4PynfyP0kzGDUXdjhmW8Kmx5JIAS+SWad+kUiQ30GX9AM624lDbpIjfJq7wpWdttoXse
S3lmexRx1N5nm+2cHdJDdGahGB90LFE3HSodEYSFNjUtiS8eYADTeNoRSJ0O87TkTDTN0+5PgYGl
8wxV2/I0CRHgEGNilE3+2dj3QEu+C0a8B2fpp17kVRWci0lreSdAaObCOzn8iMqpzRZSn1UK0NM4
5H55LEqxMDBf0jbVCZfI6892RzaQGodaip6GQilw46avNlHBlo7hbDOVS/ISmGP0M0DjOoX8p9s3
gOpu4kxKapx4RaDZ+WJxPDTHG83ew3yNvsupxWaFUuHp9Y3tuHOf+oRswz6fXAhEXSy/Nu3WbRsH
2jlWoFjMSdjga/fL4ggE4CHz4KYWAz1R55mMI7Dg+VH5CX/phujod2pOOjET6vM7qcwr42Sgum4Q
RKdSQRLogpQT3rQKDSId8LDlkNFLRUerkPVQ1MgvKg+/fRc7+oPhrpsRGlEEFi0hqI4U7Ypv4g43
2a7Kt6snEhea55byiMXrkSVZGmi7JPavYfgMUTWgaHvi5B5mNFe18tKb/JFylTrXP0HC3ROJ3r+7
kNnMuxaMeY0d3NucMBTKp5V5t+MQKE9o448QYdNWZaCqLkjExWdgNUtdtoh/DmCXfRMiy09MXpoJ
kIczg3AsgAADAZ6fvbPAIob3i/jXMcbekCYlhiaKNa2DOjh0sItXHFPnRt9BrqRUWWj0/xUNyIMe
6Ht4GOSo01YPVoaKCrc5MEibID+bXAKCA1VhkK68meKlpZRbEglm3UrRWBqa91E5dCJfh1lnA8U5
Q6NYb7idhmAXb6kJaICm19mncEMasM3GCww5lLd6aWQIvHFr5H5J6HQCY5w+eko+JLzH78Hq9s3B
B3rdIf5QZfa80HBST/Q4f/oQcpzvXhldZyMrdJCxSwUjoFsyb5Ti4NtH2doEcWVZIFUZuzSn/aJ5
VUZK5dCm6jaF/FRKSlS0hR6SjAqRa1fFrRhAW/5cDX4v/kuX4bxKslKXetJvL2XdrSToETzAs0RA
BwIrdmq2qk2jOa32l52EYV//mF0Z+TF+kOE31QT6UQzHpAiYmDERiE96rualQepI0vDts2wUBwAk
aCpLQYs3QpUFuGFrS6REU4yw+2bHLCtBs41k7JMPyGE9oN1e5YAMP0vfkdfL7CojorLoaaA051gB
l4R6mSzEnbO64l0zkn1I5uRyyx6FVgq7HzyCxlwefCYPw7crHpbgaAZAo1HV47Rkh79HlOukuNTn
5b+70MyOU2jv9vrnM//qGSG4xtBgisdJcriXu3k88SOKem5WeStdFJRIDDMflYBJC1yGnItzuTz3
IG9jJmVGEIlGfnYt9rlPIW3hZjr2VCXMOip3KuQq8lcUMfH7kiaxZQp91mwvLiKqLWiyGtwfXRag
+zsvY2Axt+lOSqnad2Y6/Ckvt1zaP3Ik/8C0Cpq40IeVP7idJGEXM1G3Rl0SUBA1bGAndh4zfQNW
0fEXPXCeqxgDNQ7f9wKf+pjvzsSKfvhgCMlO+UEh0OSyxm5j3l1S96cqIM7lQxGe5C2eNVTvKniS
jvOZq0s3rNMv/E1TMdtMIrYTL64wmkH4QdfLXiYV1tGfNjB+GNsbrD5qvsfGV7nJjABW3iwq4FT0
YmsG6tC646qVyitqn5HDPWae7Dg/asqQFTqo0l8U3t4Wy6H/LpGrrLmW4mXm4lrT3Ps/i0XVDtkI
S3fwhRtKc5n11uvAxxb0Xg46+8HlL2P8Ss1U5zb9eB6WMKyl1TrD8P6fZ5pEp2g6UbnJ47ohW7Ak
XicGZRt9sCw9aijC82EWVoCvgEtEkpgVLpq7+TeJvTIs3O3N3GY6EJIoBTUyzLi4t6XxphRGYX45
V0kck7byfIApVRzL+i++Xd0ZM2sKbd4HVKQi/hW/TRIxjfsiFmYqwO4WJCqKS1jXqUVKWb/Jua17
MZVfHpSNI8tZfAu/Ch/oNqdPD6dxQnr+T42dCHoWz5YrTItKJS91I6o8psom3kWtNHI+/y0hX7SK
46R+dkWIcnimVHyaoxcVHf5KtHIz9l2BXIwUvzJnbCiIWe+wPJmfagqKEUfs+sa/sPJr/jT291hr
Frjvi6b/iH6AXECD8fq9a2P8Xq5lg6d89l/aCn5SaV6RKX4gySfvo7M2Ve5VU2VxdDkROwjncg3n
DIVOMJK0LA8ipGqo9bQ39vvQjYFdKzcy5u4PdYehmKxEquAVJP6FPiO0/iwGoE4S0z0b57AFehrZ
gNaw4odzvqhWItueNqWnI/xcuZITV3yeSQ9IU26mlsBkX/hkGzSSqjydiiDe1DJ7uUanqV9BzU6d
m3HU0iS8tQ04vde08PE51LiOWKULKaGk7DZ/R5vS6+Sm6Xrmjc6aZZ02ksC0UDxUji4xjBZEdP8d
zqFwTh1LakcCocYM1FA0TNN7c6LZHR7EOz+0Rm7LwPXcx3jQwyivtAXj/iau+B+vGMhAGYbmPLqb
WC+S5InD7jyYWL9HkDaC7vreLprtaR80Bkw8wo0Y/iZKrlFrXgqhuAdKW/Muc1s2yawvmi8Hq26v
qvRJ0oB71wK/xGTKJYQQvdJekiQak2cwlQk93BOnsXetNuJV5y9fhFPMPNRj2OHOD6ysyK1g57tq
9yvx3azEYsc1PtXDXzAQEJZSFp6LYT2wSWENEPyI/v22lX0G7Jx7BZdbzdfuHSScQryCvQioRaKt
y4Cr+9ODRlG+nWjOAhBBhptJW0rD02XDOnZvKrdiF1lGYH8ArJIYyH3uTeoaL+QcZpBH+5zs2QaH
ZaHWhlLOjLd4bnUXEoPMt7uLabQM3k0+bJrGfpYA7WkH8E9RNYCZAo/EDIgQR1eI8WWbB/KGyeYr
BeBtkVTSEeZGn+aQpWKNT7BMi2uwWEhf/eCrKcMh9LBeWx0w8vRdJTmaegf55cCy6s/cKBEjGG5E
Bf6VCus8EKBLBHL/lEgIi/cnvdo5DGBXoj0nOoi5OzeQX2eakdqsCl4UeqndqrwLo+SL7U2XxP4W
fONEevZ1qxF6GR8MGMCDo1wmK6Nfvzj/pqZMKsaswAxlqb9FHmXDQZYrXaWMeaUd109HQu4cwHSu
mFnsCYNnKkVUn9+0/HcbTySbyvbSepTc/UaRb0HJJ65WnJyKUd1yMLqeVHCT26EkzST2jj/D7vty
UldMMSHa5Jb9ijyVDTFhc3xhDX0wKw3p8Rka48tcSdsGXUc6uOw2DyUq2Yk5y4DyxrkstmoHBQKt
8emrUiaCCLHH+ZOz66cdGfB0dTtO/JBMIvmnxi+TXD8Ekg7qDTEfCPTGrbQRUEs3y41fvqw1oCG2
QQZYTCGKQsIjurBqWMtX7PtIE0/Dn4WBXwR6KP1vVjvfJeStOBiH9Mmlc00vwholXG9r/vsl2P6K
wlGwaauaDPKCs9YH5YZ7Oepx6PGUJ5bQCL8e2AHDW10uyRrxsWh35etOWMvAQ4UnjeTtEs3Mj4HS
d1ORIL9wZdxQS+GnrZtL0bTu5/k8pY1x+1axg+1L75VVrKuBBm3iDCEXjj3k+YGK34OExS+1zcAD
3k0KA+ze8V5CM/ldckBZWaffexFwOBzKwnEARN6FKBQid6hBkal05urXrUqLUzBBAJS3lRxFYY4o
cFaC5oO+Nwcw8prXd5aoyb+p01637yo71eB+zeFxUUKAq4zv8PRjJq2nA9YA2mKuWWa/GrpFuysP
NIC6doBJLS/BuoORme7GDmWRz8oTNGKPiJT/tauRMjgjvZ4dYEhoCJaTCdanJ+ilvUhSLu0rWZST
nNWtL9l++phVcX6VnNJHBVZIzRFhloEugFXAVMU5Uo77TyauCZ+eFJBc1ADSOeIu5TCide/FZIjI
BYVq2v52MVcaLpDWz45oT1gcienugdUMcvD6wrT6TXje65Wflywd2s02bs1hFa2k1BpuxdMe4eHT
Xqi7SHIGnGI7bNBkHp+2PpXrTyg45H/cA+DC7NXszzynCV8XXGCcOqvfmc6DGRd4BRzt6XNjpEq1
Pw6D4GlEybGIAi93ZszeAQBPbzyd+yVASRoEx/fTAV5G4MXq322glJvKDB1n99NvUAsxuHx/KsMg
uA//kwu38mIpdA0oMHLAlHdR52GRSdOlDzxJencPjAn0Tbyrj4rpSm99HOynN5y362XFyjk/GUno
xE9sD933gm2Iswek07E9ZSNJV57mWsQEuJWCiBgD38uppyrivvt5lRhp6QJh0pl7YSK/IECauNtf
WLUZ+e5TZxgT0OfsPaYfQ6WFp+3JQxDp0sArx/kfKJVkt3YR+mqpvRKB1MdWo2NTDIj3MQpi0YCo
cYdTIiZnbr6EM2MfW6v0mIYZJ0OQRXTmXZ3EmSiZ0m15AJoiZ/e4pro2tYy5fSXfuk7Wpgp7e2HY
KYknFkEO640cs9yPeV4kPczXvWL2/fQMlg7LPejNV5fHj2A2R94zXousxDJXwUT9y9haEmjeNJXu
Q+1jzlsdH9Itgm8ea+xd6Wk6yg1RTsYwY05eR29bZsnK1kRqUQJzr862QZdTyX9P7/SIUwrerXTo
y5aMfGXdGdv15kdiJBV6wnf1AG14hmRPmuwttjv9uEOEi7FQZ+VIZwuMpBWBPzkvo408++uraVbW
DbRxUuXcQad6V/p4o6F1APsCIts4ltOGKfVGp1uIc+zBZlfpf1o/0ukCfjrAXKphi0xQctzDrv9s
LXmN4/tTQaPuzLPlqp69QZVZ4ajtLMJbsvxfvWZL57woG+UR+vYqyia7E52ErQxr/b8KrN3MiCg/
5yk9/2FtiEiq6KFwkiUYUATvmZUiHnDVmyDX0a7cZgmnw6RrDrzojz5zoKVW+la83eAplj+twiKp
w1UiuF3kBQJzr1yQOkzIARyaOXEujHJIhfXBoCMJwcx8zoMGqGHS9gpx5iYpHgI2ClI1om6NYb3p
YDdEFDVG2Ido+UQAEmCNoXU9uyRs8hp0y+9lw+kKCHaWCNQmh5Jw9DSNH0NoV4IYklPiwSZNCtGG
qFGfrBqrQ082pOZJina4r3/aWfEXkh5xzQFTnx2qCVGQmh6XNmFRyB87a7D259U09RCrrfdJUlHd
CCTfQxUBCyf63qBimn9Mrwn2zBiS0yU0rAlI2dt5HM9gsXc9/HKdBiNlumW7HuFY+Bj4jDVRq7UV
cgICY15WvC22aiKQBswkQ2vZEKvZhcPI9MlRKR0vQ0qCURAcm4rPpmAh00OX/koIkGq64KJO3E76
aRmUB6+f/iD0UjtYu3XRFopd020AEQafHvk7OtFcMnxWTiDZqGWDQBVO3ZRehoQ8dMzg1G+C0pGv
b5ow2Np5HdslRues+jc7E/LlLTULaPLtBNSyhyXO2D5VNt1CbF5dafG/U41fNzfd5r2M7NJN5ViT
AUaA9RQGW7mHyz4JU597206bxDYtt8Arcpk6ip2k9rilpP1BYZUtgvX8EM9owwQxAoEZlB3F4cpl
Wh+qwlf+78ad1IYuqF9Xy1+Xf+HOgwr2npEWQ+sR39RcGwLYsNp/ZW6JW4Q9vK5h2hI/PqJy7Juc
57LY1EpNIWKXHFW6LoHSKDHBvsJuwXSAn38yi5njlv0aZJslJD1KdaPJ7TxuDJ7QrxxEER6DxmY8
C/KMGIbd+KrJ7u18Xw7oOHwLuMQ9sQ6LZTnTT90Pzk1cvNYwvCM3xhqGuNnKMcKzj+995x9pjbce
hOSD1B8YrnIMdP2jl+L4YgD050AR82fTvgS1j+GuXDBgImBVh4PTNqqqkevQbNP6I+bTclqlM518
LgZ8S4u2x8WEKXz2VcLMPNrQsd/E86ZShxMWRwsnFw4klznV7J9CJadIwHWXgkc5kfjoDEp9ho3w
DxBIx8hq1UX2FZrDBTSPdNTvO/JVvzmjJGN1qDrRe3+8djF8UFRXs7n+uEYJokA3AJQj+ZNmX35a
+FJf1lDFbGpwgVE7IQyyeG+IiPnLt+WjatTXi5p8W/KWZ0IUqaKcajjjfOFLQ4ps0yJdi3dKbd/+
BYMEXWgKFcfKSu2AJ1knxq3z+GZ2xZr7Q7yJMvSSTpXnr2MRgPHmul0oVczW95ohPmWCwwkUQvqY
2iCrK7ZgfRuDH+e9xIWvdBtJ9NJ6UA+R7Y3Xvjr1BhPBIJqKr2JLQDnwOmEVBmBfo0aD2fPJ3D6w
x5SmBt7U+Nf7xyxGzpOsQjwWfxaxCytX2OudVNGJoWxnzW7ukSK+/wX4g9UQ09K+52Kx5uEd6dqt
NAUsFzhNeJIuymG58NTsLjOKCV0+ipMKTvZDMzW8jPllYFwbtvSQPVdRQjU9/eMYQcyDrn/4LXqy
seqmRy/r6wQeGCSJVo+uFusQBbis03Xt9BPjqyPCt7ZGGZS5LNEDv5l9uDJV1aD7fJXhP3Wf4Cs4
uFomRt+NE1+sQbgwqZaQDJMSrD/od638ImvDpVauc6BzS0UhAUfc9jzrQpIfchkmschSDfmXnWHk
zXZp3ADh+TWIuPhp+H/QJdSRhn3xrxKScAmcnUPio+XOUFjLmhGWfdUHy03HI1eAavRG1GBgRu0h
yOUqmSAosskBQ7R2E3iTBiVdsZOJLXV8+Y+NxLzTChOOw4N3nKNr65AZ6q+Hi3v/tuz4oN5LffHT
L7+JZfChUqvmbDjVw/ziMeD9SkXWyePgAKKevXk6FOmFUhBtIhOk58Yuqq90Zs6v9zKpdRfU11+6
VNBSBwVRbtISExN1hwrdrcCybXxEtXVz8d00hWiUZ/kbS/2LgJvSoeekIh6kKt+1zRp3VKdu1TH+
8wPfM4xI5Fd14A32Fl/0aFoXqJm7emBVGMRudMdLtx0jwV9mCt2BZ/6doaOODI8BznLQb7SIIbcC
kWaySlJGt9/qpfZCGD1S7H8eRZiyrT6q3CjNEQGtEiFczDJVuBeHrZzX5izXdEruBzfH9AMLGaJC
bTH95JxhjvpvZjtZI5lacFmx/SOR67uBsDHq/GviE4XuEkgjMG6VOVSRDJngjSIwI4kJ0VzZiapI
2f2lHPbRtgZe2pBNkj9KAZafejVaD1RWOHSxoDehtE483VdhxlhclL0pCle9xHh7wGbCPrKIDIVP
uhyTtOGjNyyQQckCVQwKPm039Y9o9elKBhn0dF4F19oG2UA+fyNFSwdCcoTQ8NLOrr9mW4HS405F
LmSKswGyjD+cA3DmuZ7nnmGRndwkERGsrVJlGBS3zLuhYTC6M4HFH14Xc+6ZPUKcTWiyogvcwZth
igK4OPG5jE3dawEXQmXTHhdQ0if8BRVRhYQFFgaI8dmLgKVJzDeqjPQjkNxlkLbvrIoK+sd9QgV/
sHSCCVriHlMkQaCqT2ryBEx2zVMYLWdGOzAyXQ1ebw5gaL16Y7eJZJr/1Y76kXsax+Vg4FRdumLj
I+TbjjR4owcYKuLMn8LDsFocr0IGoa/jhhbXlAj2Df+NTt1OmbZJ0JUMrQG3AhTRnGijRpYnBEDQ
TwABk1XygKNYaZzQ/8rECgI9+kOcZfrDX/oh5O1G+jKM7zHRFkpxWfnqdTxU/UEIZ9NWhKrc/4zR
tikIU4oEXQ10fVJhkqw/QUZdeaSGjNT3KnNJauSgMqySBbAWDCkAclQ0uL3UHdpFgjV9mKZOLHE+
78MkEQ+lPIfl89qiOQmsrLWQtppyImzYeTEEXAkubgSKpQ95gx7O5uGOkf6Z4W/8WJDzkVeQzZyp
KwsJo/wydmQc8FlZXb6/M11BT2UO3dN8OXLDEYraLYC7o2DbKTIoPBl/wO4QnpgUO36QzVg+hRJX
BugBU+DY1IqFdHE11hWhmifpQaZxPJI45NnuP4V54rFkm2JH5fYW/WS+CIsiRQs+AIx3j9sQYR/C
qrM/KhXm1r70v9g+ua6yDKcgsKVJfqZsG9MOIu8SgITWogDUU1sVVg6IMY/Robhd2D8zyPII+Bn/
neJVKWk2tyhtQntq9Cvjk1FUd6YcfYFaPJBK8VzYJhyrEMlFzAuwUl+Q5jXb7JxajkVjzsMwZoUl
asuNAJB5pScQa6egEBPPQY8U20RoMBvO/4RewWtIN2s2NKonB6VqSU5H6YLzrQWtydoLJ7KaCSr9
k+WMhNGqP1n91aVY5tU0hwzxC7XFSdRh9vYR1DP2TVlVSECiU4t/vayMl7sS1Ns1cVHpRA4Q/6Mj
f+DmKQOjd4pztAb5DhYTdJ96AbmGCfa8r+Xvr+bIeNHtNyNu7eDcA/7YGtDRa8ncn9c+iD1Aog+j
gNXzJAygo8rC0U1q/jo8I9wXPhiti/4ms72FOJsU+7KauxN2lIGeyV54PU4VJamZkYnZy7747nrU
mVOemlUEhJFiaVgkFi1CFwNVgmGsJdGjWq06+w39Sw1v8fyzENmmcHx9e28c4owiMjyTcxpQS+Av
vdObDqwMoYXJArcOsMmtflHiBnKoN1NL5mnl826a79VhTVZ3aI2ZP8d/PnO70mNZTBlFor3rYUX4
zudBbycdQcdDu46qMSdT9GroJQASksZ+TdH2qr8XLIjATm7w7isu7+IG3VmrmY8MaFu8Ywsy5DUX
Lci10QLTV7GtFo/Uttj6EPRWpT6owWy7cUkMGorhRxhVne3AqqN5eWTfjbuKA4HHHDA2zQh/SvKX
+kFeC5QFDhiuqBvjkuGGIWSptQTbymn7Gu3mHM5Wg/6mUZLxsryCRGBu228Hz6r/tzpBhZJuViON
udyDT0S4CnfWRWFrD4HuCA8l783icDWoQiyodh0kYMeYGHXK97e2SSVuFJlrRRscRlAQo5ttMCr6
LklOncNu2VkQT30CYSuWvQTjnlki80ruq50O+Sl/22sHhjE0vl3jnL5pXG6mtPKHTateCwLu/gpW
Axumbrv0UlBFstNzdnPH45taQCg/JShg6HJvj0nhItboqHX0QeaX0h/5TMHS1tWEzKtDIqgXBmVE
BmaWqJ4ZhviYTQ87Q/BIgGviz1d3TyuQ+Ytcxo9ByMeC04PC4F8BIHLyq+eqFe4ejSSJat1a5Lf6
0McCh58+zSY80UDDAHgjZ0rwjtGWQs+Xh/eNVVv3cf/JTzV8mAvdNPffZ2uB/xqrNJFl8s/Wk9Un
WpZDJCs3jdXJSygvZFqvhWRecZEYJc783NIok0G6rLNWR7nqHeWEyEfjNTLktUr6qiEvvRXAaXDK
igyaRguladOF2/JFEFwlKqqS2/xNdF0vg/8vYYD5rj0Ov8r6p1jnbqL+lnVR8bNBSaZt7Fngelu6
NzeJwqvAIE7Hnjq8cLmTN586Lm4UK+XiUUOJfFScaNhvwOpMIfLODvO3yHYMv0y3RrzQNL9oCWtU
IO6aZ3L/l5AHEb4sLBRJ6BKO4ltqD4KiUSr3DWTbr59qRDPAMSbWrpFbiVbb/ckXXrGg/NNywezJ
oClAfOzLBk9SFB939igTVgLWWxyJk8RZvfzHqX4obgqw1mxs1aBC22zgwZXv9/cn61s4utncz5It
Be7MbmiEcOCkOEhjCYDJb/AfUogzdjgaXtIy0J84Sj8D+Kt8vdmBhoFv4PCeRqDvhiNxH+5qE8aW
9rMXytwBymoOrUl+32YXIcWx01KEBZMWBkkA6H4AXepgUaGk/6p71IRfyjz4BSIAlB22da5+0Tdu
MokEprmYHjdkik9Hz5+hBGAzkaBRgZNCXit6kRmoSlNKcISG3Ol+dIck7/yCSWMKKuZ6jUBVIL6/
3pnPdLh5C0vsfOkuVEUU/kwYHH0cZt8GCE8FRJ+iSAlRzxn+9EsxQvVN7wccw/oAaXkzEB6/AB5t
6U6zh6QhSy4u0NGsGB5spiVmUYXj3lrPB52Vhg1R6VeCA01m+WYsBfDhGqaOE4YSDPVY4+9N+GeA
cSayhRDyXV/U46Cl3TgCJeN9WmA8pZLlXJkX9UyUMKC9RqwzoXlsELMpjmyMUgoxEt4YMbCSA3Zh
mzfvSUhJ4hGRxIxM7nVudjfNVq1EwDtAr5pl4GRoAK9PicNHDfIou7a8ADFshrSxAx2LN92EBRWQ
zlKYcRngdi+9aSlgKi/010VWg7wSKDqML0eT+WBKbi+o0xUfi6ZywUDHw/zn38pcfBNzT+HpbdDw
2wgLyqkJm4vqiNT/ZjNX1IG/kF5dcNjgEuXqpi57KZzeqUYWWpdgLft5HumbYv2W1XBKaDMRHTOT
nNKm4tvLmkOlTPdtMiXWn7Bnsk5/ft0Tn8KLwONIcoGWVmTxLVYVKYfPbaVDhnYdsjnIemWEVtc/
9CpoPNCbGVV9LDpCPmCSVqYU99oIOlrEKMn8Sh9vcU/b3Q68xXoLt6UGE97n5XzgVTCWL1sFcwCs
HFpTTfxKkoPdIx6X/uIk/ttgptaOdAqAIE5OlOrdEfzg3IPwq/Vsg4KfcIhOw6JuzBWy7atg364+
KCV9UrnQ1VwzQ0XeA0Cs0G1BxOptTGSMpInJnaKvHlpjbZvujxao2vwz2nPrXSmwNHIdedhe9fIL
rt3iBTxWaXIGE+5Cn3PLYLKg90n5A2Fl+pC7mJ9ApEIxLj6mpgoNlrlHijJ/llGq9k112DvZL+QO
+dMa7rO+iZvo21N90tyrgrJvDUy+YimcmkooW44Fl2xnpJWsV47Ts3IXnKsYGONU171z0aD/7ZUt
fsIoSWhnpvyHF7KBJGhMZz+RMhr42k/FsN2OTMawsvW1zLMjAugtY2exlovUqgPEiWHhLBNw7pOL
ewVfuEN0vhax4DaxqS9kCNP88qQn0K//Bbz1PH/Fgq6LrJjF9T2mIIe9zgkNBaM/fHJgPHHSweQZ
St1NHbWh/pa8K/d+LJyCMOS8V0he7MAQB0K8Wm6ZFdgfcuSc92cK9L7fDONU7ZkMJYsI3ZT3LfLI
5pduiP0bqIMF0FUTfQh1nzfjYXth5t0W5u+qDxNpDgaxarecCw1iw0qIc8Mvo9Z5m7RiRjQCxZDo
H8ucyZ+cU3I+oM+OfnJb02GBtMPuhFSOgjC/ccj4vcDT85tBmzoUsCz+hhtHaQY/OGTw+BBDVF/2
E6ZfgvVhrGX52WWG7dlqkiocPPW7mL2SNYrVPwE+1HhUjss2KcvOGSprUwlgoc9MkAtUbLgCIZ1t
vV2PHNrjeNerzh+w61Xm2v4YOKYTo9SgXTj6nLXkpVeUpJ65yV3BFYpoZ9DCaZaLosVIu1XDyZqe
mRlywVN5T26DfQOLnrCR5nk3QwI7jq6CDtzO8b/o/Nz8OfepsETOSeixFeJtgViiP7/zdV96IqU8
HrsjedZgXLkSEkl0kkQHVx9Ba5H9SoCLgemoWtSRTy/kMj75T3xStpDnM7rBFSM8ccnbP0UjQ1A/
QJey+j8YCCnY/AMOTJQZwk2w/+hfhTX4S9PQT8+iL6xjuv+cwhkwiAVl93411+eLBNXzJ/LE6oje
FBv7GkdySbmaz6KUPAylkBdLia85jPKDd0DQ0l+tZrYL3RCVlbd5A13zBkJoKjaGOrUof9fZkPEU
jWVftvyl6zLk5MG7NQhSf5kEXyYzitbxlinqiOAqcPPEHajIa30qE0MG7+paGIfhQA23wknb2H5O
fDmTgUnfghqk31AcCOSyBhnH/Sz9T5PaVbl7am31nTjz3bfsDvdnV/F7vkn5adPG7U5HE5ET99Zl
76Z354WfhG3Mi3DSQyEzTweZ8it0vIk+Q/dhKwQUxY2B33eUBlqPmd4wWA82YYk6WB/Ilk7bahEc
6nSzMsIBQ3HKI+VqSdmSupNgryA3+NM/aCUEfyoyOv/99YjscOW2mkVauiumsJAWJjrZ8Sz2GjzU
HZtfrF4fTD/5uq33D31mWUDaOK94HaKKDLqWZs/D0al7MJkVUqaaAv6HrCRJn5eQ8cqTjik3SSly
ULANgGeBqLTNFzyodmsqhhrFMhK8928eq68QBPBTIG/bgqWty67dbWqJ0BNKrEov5n54AZSMfUEM
Ma3Fwxnw0GY5k6dPoiXJA7iMk6+vG3H7RAKbN4HrI4GawYO81fyTlI2K5OsaL8R6XVHt59lhWEZV
X9jmOJpeHVnezj4mJgJCwF1d1Z5p+tKSMXMWDz53KDBRlgqSiCA2C8snWvY3eFex98jK8oKav5F9
Oe6K1liN8gsUjWU/s3qW68ZuTn4PU2PWFNVoh9tZRMzB17BAKr9pYSU9mWzam38UyYIVT2FqNu/G
vdQldjvxu1TzymHwyEjiqPmN74w6T8lgKgdBHzDE1ysplHlcuUjyr3mMYGIK97rJaQxaj7kxJmQc
GavJ6aDWxsIZ2zLicovYjxsPuCLmIj0KkhVYRjnT/z/w4qJjsmUAp1Aa/ALi1rTGVC7WZ+Z28jJo
l34V41dFkQwSQgpRZm8VKzAKaVcFfBVewcg5zY+O2XcMjLsE80X/xqa3pWj0tFOp8IJu3wuoIXYb
AZwDxXSlH2tzyCcMRHyLVy/Oqexn7vCTF2vN+oJgyHe1BagtyTpVgKpdlYideaMaWNgRyaw/uX8S
CUhIDGCaLeAp6k+sf8PvmGjpzL/i+gSP3fZx4gvAOUvK5N5fhiYiFFK+5ID1wSkPEE7HMbz1sTQ2
iZ/4DuY1Ioatftf6HsKHal5Jef1O4uDIHpwF9sbVKMAlhPvYRX447y81acrVjb7NaT5I+iimBs+0
sASTcdWCfd1v+4CA0w9LtPZkwDf1sGnb7DVhoRSUoBbpUgMb0W5ex+tq5egxL1uivSmLgo5banEO
ASu+kFcmjLbFmbEI69naMDWDinQSrAidsSCL/aM0aivzcQIn+xhQ0bBASlnLGWrTm1Mox0zGPQYx
FwRegnJyIKLuT3TuSmmF4bLAUQt15d22hAIVM6Q5rXlH1rz6D7IEIwmGqFnY8wxjpYCP9t4cNNGE
c+3x0Sx3tsiOKgXT1nCiVPN11WMaIq2L2MN4kf3c/VovKsNL7Ykqz3np4ur9MjiBgzAOOtodG7zu
vUSOEeE8eEo6VwcLlfuLRf6TNqc5FG/X3fK8OkspreHGI+eHMl2ViYeVtXgJx/SvgKhA9R+rQ53v
LIe7dhZDXIAvyAUarF7kGsn3Vgi4gXSK1jwRzi7LCEYq4FPVihvqNvkLPsVyvButT4Uwxbtvu/4w
KN+94XPu08pC45mqAQU93ICb8pfTUOhlCY8BePSuZHzlwC8hP6RbWc3mtwpITOCsFc1zordTSmIp
CxfxL2sdjmI8LI/RVfyhgQdDyYiji3aDS+8FuP7Viiz03l9wIQLvTwCchyctlNHa2zUlQ1lXtg7q
1/YC/89CKi91qu7y2VH/8ajomRiY+sPbKKA62E1KQLQfAH83yD7HT2z6fVBcxtwU6yyOFPxqdJCu
+PYy7z3eK2ZO0j+gZpB8ZD5LskWBwwXEtyT28BtOdke2jSspJ6WD/clc+nuy1qg9WskUjiiKguoh
i/mY0HRjtU5xtScmYHy8B0FYapzoelUyg1c7Qqj2CLG+eslAbkwO/RgvF8QHdKw9YOFSynY0Cdhr
uPTFDrQABTfytYdDTbbElypYx/uVyOGoT5HMtPqdsyFP6vvBaTiwIJXOG08S0S8xLAJww7NoNQfw
5codKOJQE3uBjPSmJ5M2Hwp13ZX9q2gfLF/Mm40N6gZDayYkH9w2ub9bq9xWfHICmVjbCNYSSJqs
/MQfbCaJ89QHWFTzGrG5iT6QS9dMbbGPp8s8R7EYw+FkmwIfpNt0l2vFPjjcgH8mpgluL574TzjX
0xwHr8nQHgQyBgNX/Z3Uo14CdkgwminS93J2caGNSwoHCpVYeQSE4UqR6QON1XwUsHGUryCH6fTC
Xyg5OskgZk9UEhIqroEptMTMVmDkv31Ee8WEY5+fEz8BFVTbTp9E1TMdcbDp1vCK1t6UUJhndrMY
UMnyHoP5GY7m84JUiwW3U3GARhOw+R72iQT/+o2U/5+OPK7zMnMZMgM8Qn5PzmyCevPdtNeOII9B
V602tdKP5qXAtqTAWUvHftV0s4zLDNMocxMpeVsMPeEGVAWD2Dq98Bs1iI5lrHPHc6aZkIQKX5LQ
y+hsXSwmzX7PrhMu+9Y4mrqcf/XqQ8V+X/wqM93x28pZvHwJZ8LrsLCw9hGQ5xsMhSRVmtxmUuai
DFB+0AK1eNYYftni3LwZtc6EFgL688BqU8B3GLD/e9WEvmQKbHMvysaYyM0duivVnT2Nz12BPFLR
oYLttu9jS4crKA7bktpks2XDC8ar6Nv4aTSDZZ2DJi9uo5u6Smy8jPcshZbWtzO9ej8cuFqDvNHq
b+XL31ZPdX1R1hEPvAjV9sz+tNREnKKpibVzYcPghYIEf1S3WzqUKZ9R+JoRuRaYnVb3zlmgz4Wg
yEU6RpAlLq8jtDCrGybI5zGU5KNYWzXGUID1nyKOBeBo93SK4RrRlMxGUBTvAM8/jV0y2DJp+9vj
fnhlTYlc8PE8K1Hl8MgOwzzVky04iV//8FWjaqyx/fDj8A+b5NxV4HuUe8Iu3jvi2flf4ceLfa97
kZFAvKGHCKesc6ap8hW6zIbkEkGjjubX/gVjuDL2/7v4Sdfg2Tp9h9ol2ZtVJxhjb03iHxA9pxl/
xEAf0NPAyW/P/yGqY9Dd8IXIzDjsM0uU9VI/ABcl0bIoI8gTTbTrkBzg/gUlfYSpaGm5/4NHTrpZ
h/JxP2L42IBv4YjjcV8kGeTmcKsD81ydhlfUwQpIDXvtRVM2Nn8CBYiNin1NEPxgWzgfClSNnyjQ
jMM4n1PeXdxtqjMwC5bIQufXBWoj99TlKwyyzCNwoqupDpziZCnZaE0s+ynX7QBXqIdAqbb78Let
3tLacFaXO78/BL0izoYx5cNvDS3zXHHf4p9CXFL2JkqpzBuRrWqIhGFMC1eEifWuVytDLlYEJlWd
J9rRWaRA29TrxfzaWxuoBSKMuIOPhzdcU2PJBHee+ps7QN2m1mQS3UMtv8FevOTDC93ysjmfg8H9
YrhH8LgsFQiNGjYABo5E8UMUNp/Ugc1xgjqh67nlFB/+j125LEV5b09TGjCpLfBuWC85u+cpKE4Z
4zyJAaX8twERX2BFOcKJTS5E6oHuEWZLGWek+EocqsRl4Ii3WT5PojWmYTCZe0cqfG26xzZvY3HR
obuTtyi5nEy40YjShq2RU6dJQAG/dp7JmXnWQ2BC4oal/f3K0gdKtacmcLOKLqmaogbOqJpjxCcs
BXiBgCptygZa0sNTZFD+FwU/NOVWciJ5DG6vC/63ko4Y9PWn4NmFLHywlX/39yJOG1/cnM5yRnZ3
OEAhRIrUx+iV5k3Kt+u19Z7CvDWSuKRmpQHYniFDWhhVPwXhJD8vZZYAmSeeGbiGmRrwCU/HQZ3R
GcQLyBwAKwPcjymXCTPbv6hbDMzFjR1KhBjAHO5CicLy2YqmH9BCiLdFNYTy3NgeGI/+GwhmzohF
ALcqbUl9fDUcQWTkipYLd2SB0Wq1OK1P/3PF/DfAT0ZGLyXpI4JreyFpW2dwSd4u9JRwE5MTNWd9
5nHyjWYy7eNkpAo/XgbteSvCmuztS1wl8IFlv2WYVaismzoCxiInVXZXpjpK/3dxK6pFpeYjw/Mb
KDoxmbC6/Ck/o3eQlpJ9w5GbfbZT5qUgYzuq5g7SWkAgZCGZHKFKup7PPOGqNSLcuFUrX8DdUZ22
HN6qLFlrQOaAm9s6TH6n6LAaNHnRjimiJurlbYYHTL61inwvTGn24kcV/FaOh2H1Nnyh3JXXzXbw
38Fme/ZabRtPRDIXYnXlqNyjZ7c+Q7Aydt5pADS9XQCUi65Tf/izCXlmcBzNwrQfHJ9XW19qF/H2
8oftMuqtgZMqCihKRul/bfPmgp3qqmShvI2uoPrya0oKh4dHM1MxaT1AtWiD038LuiXVUuBQ6ktA
2GMVAX+OjwoYF4agbYtRKdzeezNnrgEHyM55ri94muSDaq9imQyu8axw0rREXAb69xhLZvAY+Lzc
Y6DZPfinXulo62yef3BCwtanNwzGguTATriM6X9mZFPXJjbhhR7U3hWLltHh2Av+ztULk/33h6Kd
STS6C4DXR0/RGZ9ikWtM+3Ffnx1vzoLActsSZe1QZtZBH/a6WM3tXm2nxrEZTqsZlvWY6ElWnyWr
jf7IYVxaPMnoebWoyoUWcZ2o7AvPr+31nzdxApgI1E/A2DcxFiL/Iak4U7dY533NJQtVM/U3WuBM
0mUfUxfwxRxWkKBRf/EQXqWeAgfDtlSaJQpm38MPcgbo4LxhkwO1cBnvme6W7M6Cg6m3P9ak2kxj
1fCZEYaVCTLDgDgy1u+SSUBsK62M03jsAP7Pvkxq1oMiNiW3ZXUkNmAhwKgGIr8s2in7Y7sCnWMm
ou3866UA7jZIvSAd46naJKJuBE5PvdmGZ8Qe47C78dP5Jk/+9WtCv97T+lb5xz1m+HFRTi0YncWw
E9VKsr51320qZSv2vbq+n4gUBQuY4/ADmXiRXlowB6B+vzV0IHael4ab0Yn5JL80G3v5sPGhcEZU
bkytU6290TrLAep2GsE5wS2jA8m7XwtHPGF5Lx6XnAdXSBcvKntnPzJ7bophV21GZosaTiSdzFC+
IQgtedaQ3h0WwmrabZa+7aI5fd60P/9dJISeQJPjbh1msnaXoay/4C7ZXruK/dOMy3HQC/0TOlF3
ubsUKU3ruDXxuiTOiiYygv1djEWc15cPsFa3zMZcyOJRSsyUScQK3O1lBrxxvySpYOVMS5Wfpe4r
clbQ7Nj72bIFQ4gRwUGSv5i2fSNo7kB8r6bt4PghkVtT1oahQATl9jQo+UMrPZiddF0DAgWxLA/V
+xkWgil04vfHpC9iEzlG3pguN/YySsHogEfJi+IugTKmGscStf52bxoN5sSsi3XDpo5V0wlizYtw
eXC3G1KO3vWwOo7WJ3FSFgfZoafbtE3iWphT139qwEDKcalHPL7Jp4VRHNUf6tfCBzaFiLtt3ZZA
s6B/EMZ1qT3WngvcFdY7eR+e86edGHZEMuPO1APOapMbjDOLxYY23NE7M71K3usMFO+lKd4ohBkF
OQ4kUOsDVSZ3CrX5f6jKUkBF5YwEihnzNraRrOXlMOGYXIERYJayZ575K3KGKfwRzdfDlk9fBXym
WtY1TKlYNGgykqphwwMFCmdJeNHOkTUFkBzXwiOgYe0sSoCDEbDMvW2AZQzw3NoPPn2s8WUIlGcI
8OPXomqsi23g2VOe8lM8z+kzvFxUN5gbNiCYF9hBglVT5MvY8lJSQ1mim/6PsyM+RxbPWxMH9/Rz
Vizc9pP5X6UxjuB2oC98b5fAfGEw840nfmLrETm+LiEh+GBKOerR7l/8Xd87uHPrgE9kPI6ciFMs
7k6xmstcN8/a3gPm9YTnL/EuH9ozoW8a7RD39zIzTQTLp9y3i67l3BSSmq0S0mcGZmyTyPkNHBgy
oH3Lw3IcQEAxSJuG+thSYuZ9NPTfxCG+LMMjKQgF0g18RW218MXHg4GZr+PdsWg0+gYjw6tbEIS/
gpmXtKZ4Vhys9qiCy38W1g6HC4bByFuotPF8Ct/gT0Wtfim4WiXRx39TtzrkXNTGSP2wQB33CAe1
i7FLgSjl6Yo30pkDvO8UsbcwXXN0oZbWvIInxNaofVt8OU/vbrkNR6p2W7EJ/gPTf1ti0EjgGVSl
kHX/0bmUq6Sf0hRrHMzfr+8r1td2werdifpIaunXaL2jHFcYV0p3QwYm+NgL/TFYkkkoZEf9YKj1
TJhfpOIgdDRwhehUkDZfUEcMvJce4kmgz3bA3LiUFzMf5+IY8bAfhAXgyBtMC5ER0VU7/qTG1Yr/
HIshQ642v4wSbCGK/XCJ101td8OXj2rBrG+T9K52ycf87D8ZT9SXHyDESIBKh7kqIUmmYDTjyibQ
UACqrFb96MSjpQK/bT+Kj8kV8BEKdluAgovBZYOu0tPSOgu0IcmZsBfrFjZl06uyhWrQuPWTQak+
Ve/ipj43sKRWMFZzzMhG4u4ktz/ZMpfHdmymaUtZq2sUZ+rFLEXAElzLQz/Et6F1PhKcxztJzdfo
bEkDcQnebTZ0Cu6Qg6Y3w91KNidFoC/xeTDrClPjVFoni5R23Yd45gEX5G+EjwhQOqshg7Kc1rjs
wTLKHZvuyRgIIh9PavBvaK5pUpijy9SKJ4mKNAsZga4rrUITC3PVcvz3GpVMmj8AIst+rNCnj+NR
KwDq66wzcrRG1gNeJMfZr4c/PDSzS0g0Slz/UyzPB+k3DNs/sx+d+s89Att3a/WpaEbTzhgchQUQ
SlqO4j3b3FDpWKR5IOQOCLskf4/Sb1G8lww17e1ySBABz8MP3Woz8EZxCWNNbGyabh+pmb2MX3oa
MK0lXwR/pe4rJOqsovfTPeahGdVxWf9b93yLJLk5fha0fT+fMd7MczXd8EI1+4kzO274rtueT9uK
7OLpMnohjGgeKtHlbH4FLtNI0qlQjzbaw+XPuE8tRvYZj6zU9mSDId/D9qFQVhh25ioXJO7phNpp
qIRAZPIUWHLv/yiEdjg6GJahuytBTGd6P0S1tnQJAYIllouTGEbV4PHHnJJ4oo3d92Z2rxI3yWaw
4jnWXP/higD0wCG11HrNF4mVdEDRZHpowsmCflo5mCyR/YoHaLP4RP2aQ9oahctG2p9ZS8+DRgPv
xfA4HPE16oQ4RYsmvmpVX4ySkXZwHAh195t+mFeEe2DLJI64OvxSONjcftPy7CTH2W4Ih5XtAqAg
79iKiokmxDakpWOBmaeVkuar2EMvFgdkS6Sg9cRT1bXMB0Rh+1FU+d4jMoEqmbAJ7nplWx3/ek/o
N1GLPCVNbkpeCa00urzywr9LyLm4a6VUWDzzOuaTMNEIz3QYFszYcI5gClDyAJmDl8iRhgLGALET
C9Yh10k6nUTMI5bgUbMdFyj1b4+/TeVxDDBCshFEkXcHfwcX86KHv54lffLrf0TM+adCBXw2R+cp
9b6i/2Z7RAFf8wy+1r02pYl16vieAzmp5TFRT1I3yZfPlm0RLZ4CBqzGp/uUhEEwQ7OJI6uvXA0w
Bf04asv7tpDpolLSpGBNYb/QCt8G+5oaLyA8Tw9KZ0rvwmWA4pUCN8Dbt1sUMvbVmd8zlgBVu0Vr
C9i4EzyBE6wnIVB2gNCx87Par60sf6qCjOlB93hLXIAZ3L1G6qsWw05rlMoWNu3brq03Vn5DZvjX
Xt6U2iQXA/jVBgUdlhR1bcs04e3rF0rgjTylyt0tB3LFono0Tmc4GHAgfFT9k/jBvP380nZt3zAA
oStGXcR/oQXA28sQT16oytUnU7zhfyQ8u7aslDLU8or2qLLBx44laQNQf6wj1DkrBY+48LtFJvO2
i93LeYA648SY7i2HSoOr57G1NXK0DZ2HS1pWVqavakRRCuZNgMHRrk6vTPRQx+7KhkMcztz7gwzE
eGgFTgcQLBYzf+4JvSKq5ereKEg7e12fAAhRVTLEPs0S11zeda7i9I505OADidY7OO4ldohgYqTt
Aqb9RXDykj5DobFu8yZuy/Alr5soi+rzTBTvjYVNM/CcTD+cxBY+2pkv72eGJQD4Uyygqnw/pZhe
Gqp79tQn0x29oVjGe1W6c+bbb+JSfCN0JzIlpCdT8GqJCfwAo/bjj3uVw1tf1up4O5UAcfChaP0R
PYro4eA2Z2hmTMPA6ErEcpvglnBV5Cw0Nwr2oa0GXIcFdtp89Wn7IQX2dBi8C5jeYCwjAUbaQirY
lS0KX5gC2ZgnPeV8Yqe5JzQxG55k+hORyxlOPjBz2CYpJkCNhevOVCcTd8RZaR3Xk2txHPtdJK34
ByMwzi0AeCupJJ/D+prqykHVGuuHA0YMqme+fui+IWGZfay33dn+WbgCYmiZos1zTY3dX9utKZoi
3zzE4fCjb8b0M4poYa7OL9LnBWIDorAg+vQhVdXRGHs+H8mmv4OIS6WbIJqp14qGbrz7vpuWfbV0
LVKuOcr7hResO6oJnpYRkm8UzCmdWUINPkiDo/6TA6azjZe+Vk1PboUS6MmM01BAnnsoz/yDAVvW
Kwx5mj3QcmA2QV1tPhswepaGbjijoLUGoP5Z0Na2mC+JPAdsVRZX7s9Nf7oKBhcVozzlpBsnPbMx
Tl4YB2hP9rvQYrXzFJeUVCob6nLR9QdfZEyu7jSqIdQZvsEX4V/OOmg1wcykme/pr91bTAPPDOtV
Z3g5ReLVAAnW3lmeLt0nuMw+NF2SupqE2avz0nDCareqgGRNrEIYpIT71/bFMaRaoJ95TDZslnGm
0lBLtmC4uWyxHc4If/E0+i7c8KQHtCqHtAgdw/ue9huB3pemEHZLEQv0teBoqz3svYMBo1a89YLh
BjATejb+mAtnxZjZN+mOw2MPcKQnrwuO3746++KIlKTmQuwwkG14dRumEjWw5TyM5RSi8eN8u/AE
Y+2PDhDC9cq1to46A1QWSv3TEgvdq+OMRtmaQGrf2NlCxBxvNdyDNkjmXMBIJ9wwxeZU6sxe8Y+6
McQ5JvtNG3xbTpa24hoWgZzHiYg2hzipPMa9oM0HoPl5/AuJ5UxrbcKBayJPeK7u6UOgxKwVlRFU
OT+I41dwi6x011Vzxcir9idbM3UQKczycfAYChJyrGnxks5KgtyVKi1o8HXkIxDtqWCKyi3c27fl
gf2z8ZzA9etTO1Iz6ZF5ivjdRXq9kS0MheSXVSvGyn4L5hk7JUKwi3AHXASxVo/c14LdMVcTYubI
K+K3gRlJZhTBMcchhPQEnyGB1IjJCubmy3lTfTK8jj7gqvKCFJNb0qZIb7mVjh5O3rA+274ns77T
hZoGusL8lQkCy5DpzfiiXX74o0ilO2E7Do8KsSG5U6UBmDnyG+/Wkc48MvZWyU9v/ZhpFyUP9D3g
4K/gNJo0BYt9q506EbOVkHyZE/AF1KMgfZVOYyIgRzkiWIfr+aNQe5+T3kOi+s8s9aMgnDUBzFrr
FF5dUkX83Me90qpXtqNqFaw0ywRBvZHuXSv8HVgaZ6ftvEgvaRlE3MfAGLFdX2YOlKF7ZTfhneyT
ZgEixuXHTOC6NmOC/Banf7YvKOFIf36FIb00l06Jc4MB0dBtooPO98N40UPQ+BYt9LODcmc1JDjS
RYXEtbYn81eeCvmrM9cYd3CD/Xr+T6yS2LS7+mhMZgw3YlKViX42H8H19tC35vUpokigW9tFJJur
PYPSlmIsoRLNa6zd+jcDZ9BFda6fp/dq4r4TxS/vojJHoEU7/+Njo4XhPvdre4VwKjtooIt1GrLk
jUIsiXvkZBvVmkbTCrGO0LZk9Tjjkv8UUi7s6z31q6rtscWwdXWzk1zCGkktGADsQUV0OKoyg3HM
vfwWOx1A4/OomV9e2dbB6Xgv082aULdGIP1ODnG5tcKd4+7ZrGztkfcT4iPvfR43J/7idhTawXRQ
iVZhsWeiRlWZzSr2DUwhTBZY06ldQlFWbVw73pHn+IJleS2e8IRiL3c8K2K0PJOIB3NimLtYjBCW
KQwioU4bDccM5mpJPjsdPeHrk8/aJmqaK4WmulhZNJlzBQtPuqCjP44byPQYMFdRPNOhpYByOxD6
kFj+0WEBbPwHnJDYK8g1nbvkym8o172PeK5EGopnmZSpG1P8QJhF4fZA5kSfR0p7dqWqrwX/t1ty
yA3xDX0vn37ciMKdsFGDzvRaMVYN+Wb4xMSX+yCi4sWO9SXcFc2TbTiNF7BkcPxNQxjLhjmAw26x
MKyH0kMABNIa4bDMH72vtx18Atv+VfTLJ/a9YdqJpM7v6Zs3TpznfiVXXnvraWWyFF6d3KIszSmv
mUNfWCfbzt1VGnwB8xt+VzFEM+RHLvW1m81MAZttxfWrl9nMflP4jPa+LQ7tkZeW2XjINZn6nkTw
Q38qwsK58BiDmE0DlZtjij+IRliqeu6ZdyYvgaETlNGPcVZeaJ7y8DVOcPBXldrUXJ3mU46DCMaD
rldV4tJ7nHbG1v6jjn8xsCU1/0BLMyeU/IY088/YoSfnv3vijtTkXoSFvDz9gzqOZsCDJ3RHMAv4
Pe1XvEc4WFO6BYjtKMEYPMSxUgjYP1Oa+iUJ0PBhkMrxLXdA6mOcv0Jr8kZLnDF21GFCTYtY8Hen
2BM+tINl+9/mVm6aQbl3GdXFBoxllVceyNIeXZJu3JJrfVXnxWrkaWyY09Nh3OjE+bqSEZ5gzEQN
LDHzrtuJvTuIMZCbqmiDKjtEks8+thjdlNFORKpP+Y7W6VP+y65V9JYawtYsLJBXFBJlc20QJkwo
3W4vOUd5QXo5fhUrT2tZADTsgduFyM3q5L8zY6z0kHGyQJFipSARpgBxwX1x1spIznHcprUWmgaU
duOZv2iN0NS+2/2votZsnLWgRLqbuFbGGpr7KX+S18prQsbaC5DsxBzzPOet8CUn+Oa7Z+XVurCC
axz/1Pmz2K+W2AozKgjOrBdn9lIgJV6vKeNqYLuip2QVir2ea/sxFFthkA9IeSA/wliSdzwMJnzm
QoKqT9TM8woi1F2ezYjWCOMnW86+YhxWl3qilUO2bCUnv81nxk6LfHfpDnBCz21pQdcMFND/jPVu
cBegysnr+YXDcQx1Fes8wPkt9GppmSkE8PnvwSYr27oWQjhj/BtKY6CfI7BNlE9jNUHv+XEK4i+1
LI3cO8TyGoHlm43hyCp6JF3P+RpOobPPBJKF7pbztCxymjzEmrLk6KN8Op2+WQvX4bHs9k/IdF+N
znU7HWbEISF60S9I9jaJP7/RekzNBQN9kqnBPgY7ppnUo+AnWM5SuPDxNPju9G615U/mexUl2odT
zSsL7QhGi9i5yVPOYILt+UgYeWVlUb/7cKWiL9XYcWBowgp1qMNGSdT5l+v1X//BORSwY1bkFdEN
ywZogG1R12lWua8WA+nM3+VNyVFdN23lG7Xk4Ei/IZVemqTNEIgqdYQ5TCsTR7dnE6bS9Hu/cjDE
PGFyBA8Qfb/++WHCwHrc31l0KkE6GCZvcJ0vnxb8aFdaKuZ9bWEA4hwwgZQrd8vizotFJhcIN9+c
yygKtlRyOQp0N9jv/xjkbjoee//W3OBv/PTIlQvYfU8Qycw9E6snrblmRMhKfDHsjFs/gHp+Qq5S
xn3XmKlG75oZzWohpIR0ZGXouW7aY0BDnm7zGrN8Be7NtiHQ6IqPCnd7VAmlKYKK3Hk0caQZ/GNT
XHFvs+1ef1uPDmWtzrD7VtR4demzTuszvv3LCESnUHSU/HqizA62zPUiVLdsKy0qByp5AEjEU72c
Hgr5GzPI9FWLOTo5TxCuqkEBaD7GO888J8MZT6yVo+6kxWs2+jspQT5tGL2jcR7YQiavMVLcuGIp
8uMEnpWersyIKB6niBdOBDTiYuV9aEw4AQlEndEAVLr08UCVVsUCSvIbgxYuFQcH3RHDzD1SpW71
9wyl7hRMymvsx2WK5Z/8X27nt9AizZKS/cYuAaMHy9ZK4IwnH8l9qUglBEQ7LyL3ak9nOhOId9Uy
Knl0wHL0k387auRlY9nffoFgAVyFF7I04K/uBkm8KqgOtTlcvR1yQEBNF4kZ7Q59vI0WP1n/ecxY
VQWrcemjqJXijNjInauOkD3f3sjrN03oPYrw7gPNeP0BsyWgmV9bbuLf9HtsHinoQCWdvf+Oeca2
5CmVhYYkxbGDbmdY/zdOALdVEpun8LHyaLyrTFqt+eP+7Nxd+FMz9UbKuajMyBJV89XlPTYJ7wm8
w6iCD7xzAfVYEPIYY3X+GiWnKIzG+79f9HRXlQSrNR6Yxqbebgizt/Vp08nH/n8yV3F+pUgmC+zW
cQGUOlskkqL264om6uSc1iZJ/KPjYeSbWruf3zW971SjkargGscP7x0JbcLFiIxWw4oENCofiUtI
F3ve5Mjl1fZ2vj35cCaAJcHnFSfF5s2qF58EGIoSieIjXCaX4LLUaLNbzQX+l5bhog46sYSIpk7F
yFa4YDGpLQ2QmvMHr7vbQHDn/oyRs1YZ3m0mMljgS0fWve3z9JWTEp9l4Am+492x/LBilKhANfah
0rxFAQJGbNLIJVhWRsW88j5SLxfM8AYLEuVL8+VTISg+sb8yO/dbvPvlJ9WZgbUk4UAuACJCeNwp
X98vC+m4LtNckNA+UpVNeloiVvOFXJCZcHrq5tjHVlmoCeejJqv867eTFjZNykaE0bkhhkEvO7CW
eIxBhF4U9ZioeoANePQOa2JDuDhGE4B2qOoTL8lNSnN52YoGdxXxI84MvqIXKGXCp5eAYD9A3008
rr3dkDolDQEw6j9D8OvbSyQB1FXb8Arks3qQmGZFYPg+9eSPnpkpRwGgqDuuSJ9m13sXzjLJeEcc
O057Wh6fY1gBz0U8bJEY86yHJMv+4fqTt7nmP8IhUctjrriked6c6Y6hJK6fmoDBQgEPohVtu0aK
CPp/Yv5VS99q0nNuk5Onr7cNmFtqZSjqJbrVT+tbeI1BO9gYzqZoF1Cka/nje4hxzVI7lHjTZn51
N/ek0o/CHbQC79NMIzn6Bsv6pH8btWR5oogc6hJXVMg8gK22xq998zXLDL8BJRZ37Llr+Xj27NP2
41k9Sl3AcJmYbas6pfVrxi+Uhq+QkoVH7XLgbGv3NokA7bbPFsvcQzsDfP7iWzwPtqwdzS0JdeHl
5rcR9QbgZ8KeZJ9OMY1ICIQbWUpyDqCMmAmLTHTq4DvDA5x83wcqoJzcETGFKgV8YQ6QONdmugQY
tZpFTQvTWYP00DVfKO4WZmipjr9x7i4mCM8tyidpa6X7TdE+M5j1odVhLZxAYLqqhXpyEmwhLanq
rQhWiI31dq2nAXMbQjguKBSU/5cjnfLdh/Ob+DUehLxOIN4NbkPi0cr/hhZKVqKhv+UTAbkgNpQQ
MGweiluA1h0/UuelpfQjKGtnYWnIUNFdkzsqSRUwjmRQ5X548jZSn3+CM0Q1yPrZ9mZ+SHqhDEyh
6NaXj5/9JQEwz9Nfoy8Uxu5jqt5BqchaABkU7jg+hYRmxSRnbPWgfX4xS3wToJzXuxjohQ5muVge
JIiLWXXPiqBW7/WvL/dhe+y0qgfMNBTvKUnVsER1r0BUQkrGyU1YR8NQQOLRmmtsfY2XgH6Ea6A0
2+/rnsNSgUdhC5zz/U3kzViT91t6B/iKZxbb35l012kHEWPxBHE+0v63OGxNNN3y83eeLIbDLsnX
pCgeqsGfw8KMAbXvRNja2TKd3OqCkp8KDljLCX1BwO77O03U++pdKKKcUXAWboVL5Qqf/l6UQYU6
z7FV4BcesZbnQKUMrLcfLuF2oT2fgwZUF8CRmfVmhC+KxEyfIJxBT+QQmFtwA7wmKfcHqRS4m028
Esdp7IvAdkhMdQmWurBdB6HKDtBuouDn70y90QOJirvHSpTui8gDC4mOKNjb1f0YlwMdqSiwHkM8
grvWFtz/sX4TNZ1uvcj/aQnffZhbdQkQCYZ37LAyZjmgk/Fpc/9gKAStL2XtnUpg8bylQw1DXiiX
pPBtH8fe3ReYWjFYtjbh4y1jcZ0q9XM5wqyAX2OuLVRhCtQqjdfNBqWyx74dmyC7H8U5+FhMyGRy
Stq1J4RYr6RqMMVENcPjCXnD2IC+a2tBbG8ixKj4sGq7DpsxcfY1axWJMijfjOTjaRw+LdESLLIQ
TLrnK0qygJr+4ed/h8qcZGsfapINHVZoyHQlqUGj1J9tQp1jor5C56W/sCLaM2dmlj2FT6jLxi1c
izkDa3dmkWEogLJTBvydh9AY3LTniF7semzkT+rt/jyeWkgMXTcOc/6e17qGMr93mT/liTDXE/sI
u/RGAY82cbqzsv3lu+rC37M2gJhlanufRpfAJeWmG3AAXLAj3UxeTgSTs6dFVmO0/ZfAGnlWxMQN
lsnoEyaMrUEnlkEHBMzrnjB1yCXqdGwQYSmzxlHafEPWVLRO+Jesna3Rc8Dw1HGqFIpdxRmN+S1B
3DIxVRaiB+NTVM8DGwD9+3sNshp+O0HgfPILRAw4gyYby8Tk7YEqOEmhe/juCnGumXyidZtgI01g
lDo7ivBJgqsGkTxXN+gsgxcBEhFDoCtsDj3oKI9J7fPLL8lWE5NBOA77g3Wkkb5lgT9IlrgZcoHu
sSmSSQQJaOb4g+Gh7RDguVybsBnojrOkEY8IPbkHKJC29MXgnTFm3NpkRrht5cblynwSx9Cfu6hh
eR85gaODGBJZ9l4Ftp9Xv1yD6MRdlT+DvReJv1/Ik1xT5SkTntCdpN+d4hxToJ5OtMHeL71qW0UV
IJ/HK4FSUVtpbXw0vMBTqtuevLE2ieSxvdA4vTQ8Fei4kAh9jQHWMbaIazsR9mZc6VDexD1oAEse
R6mFSZ9MmOQqlN3twHwuOy4zLKHiC+v/x3bRffuSS2BBTVOqW69U7qf7rl6UdQXZHf653FkxRK6N
b0BPl3RqUvOCKMJERl92LkMhyuptevUzPoW+8u1fS+eo2XYuXhDw46zKyFCGd25wNSS5Y2pyeVLb
Jlfgfasc885xQyeYxRMKscWFSQ5RUHAiU7QBrLljM2GAr3eDDM+In/wlv7lsO5ce5kLh2V3qJ5ki
KmmFdxOwoAa8/0W1xMYurQ0a3DrtDhS8jaWIbmbFZZsfDaMf8R9+cMKpArtYOH4kQ0vTR4xb8rtV
9IJ0gfLwiDomDTdJNOz4y0bE0qmrichS6YpW+Px9R881LrKk6I+iEHYHxF3NZzOAAy6fCUpaLY5q
9LCcyaH1FnbBLuBJORJpa4/Bb+vb4jFPUTOyMsr/fw4mOtvvxbZP6tpivUkpqP9OCoQMclegvZJ3
K/RBALCkcuJKinvHJX3BOnxYxHBBDufqEeSgjP7eT8r0KBFFA8ofGRXLV4QXEtLhp81+dwsrY0HW
EFj1Zo3EnsT3IpqC3DTBp/FoeNCluTuBN914xfk91qim43L2kS0IwtXXKUpYw0OB4n+ofZql4uIO
cehU02GZxzI7E4Bnm5lW0FYfS6duBB4ZnhrgOEtILe8MEd69QLboBDrliVvL3cny06gSWwAxQuh+
VIaQTPXT9uHVXB9i8VnLYTFZWXw4aB/VtM3tqN2UKgkT+mR+9bZGuLACzVhy01fPEPj1kkG5v8bK
8yxlDidolJomFGh3WC5JbdIxWt0wuyZbyuw6Gmz/i7imzjqnignv4LtIigmXXJ1oZMBiqF7s+CV0
4aVpF8tp37ZOS5foHyVe85+5mCbEH7xmHwkU5DuVlPeOCYf2/MPkG6X3VFaxULsJgF95PdA2oNpq
8NCEiZ4YQ/bIH4EDGtK8V3arvelXHEgJlqYZhQ3i6iXYlEeEC/mnMHspajaAk3x45KT3YULQsfs1
po9Vy/gxG01mNOt9jsjSSCyDL+jaPxF7UOQmoKRfP+16O1z1C8VCXZm3Gp0p64obYFzYTSYa8x6M
eIlKgD8jp8gDtl1eRgo0NxaW7jw3RiOjvFoySyKjfEKg6mOCnUE+saE5FB0rqef/wLt7pcrO8UZb
kfhkz0FJ0kMOAXsnPG0bGoAzpWY6KKcX6SYF+6PlSC/pBt+o3prfKH0cNDrXSBzrO/YUqKquuMoU
SvJD69Sj+gISDabNADdqKHhJ5mdRczKjC4qzmQw1Rn4uLEeSob9btLZOGOsBPPm8WFYatlq4rG9x
HoWSchwdCPRtoG+bZ18LW5b6vSncUOa7VenYVaqd4tzbLomTbXQChY4WZzcOHOQMXJiBlqyRZ5AW
UrpvWRQQRAJo+TCidfEQcGVmJpr6f1kDDCz7t3aOuV0qVnVJev2qYgOor79WiCQ8lDUqRUiIU5Q6
cNFZFBR9uLK5vr8U8tuzOW4EcLRI6nMJluu/4o02zASuOsPu/nuQlt9vZyuYRa/XpNB3BKIWOmKM
M0Q9Z5pZsbyWsbCvZOta+XGhAWgt+l8/zm3yq+qiF4amHzC5Z2NrXTl7en1wd+cpxBx4Dz3ZXimO
M4bkjciKpAlOpomnOIGsFp76LcxbvlN7XZzXi8EVHrBjMuhfpoEX80O8rCB6rD0NzuXS9vXkZNIb
PE5uv0jWz4kUGogMKH0Ibrb4L2ODyRTksfUSABYvmkARJMDkb9RgPSwjxEvuGG9MR/bOkTIftPAt
45yNE5midAGTTqMjwamwPNN2HQwZIeu6n1kSdHuSQxYM+HCdqoCGCb6NxlOBaQ/xQ+pmlKBq7/m7
ZIstwhECwLumxOpWy8tdJciwDoEAh6rK1oANAKtrgW50ZhC4gxEG6B7sTZ31wr+aQ9q5r6XNtbSQ
ZP1dOwOTZBZj9ouMKaBrj5PxFsca4etGHS6M+7CseaJiJcj7gutCeir8gRrurGjtSdqiQPgtixj2
gHDcapZgu43BlGrBbEnExR8itRA15M0c88B5fDtNlX/KQ1n9cJtLq1fmeFrraiWCXntTjnKlsCLd
qOrBKtfo+UOXHvQB9JxmjSnL9janK4zdSCOhO+GE29Qotd8xr9bphUT9DnR8/1CPnNATdpRt3V6t
PN0HLVLr7mOEHs2LYlRoA0bTLQpn6VB655MmottFUAdRXMZlozSov3NC/mwQZCTjt2YIo/bqYEAt
8MT28oVA6bKYtx824b7YgqcKJYb7pTNwpyzSvuDp+DFm7/bxzjrvXyvSHgK/SiquNh0lIVE+7Nl9
SDSdYnu1Cd1RZF28O+AGZuY9GVdp9WcmdtGUdmPPBlzlOM7hbLlL4coMoL5YFDjPkL22OuO6qkbD
PbDtDG00EGSOZ06JDIRx5RWq223YIqSVWgHlw0biKMqz5Wyi4fkkjNojvl9eS1/fUeWdTrby/CIn
PZEfm7M5kWO8pwPuLPfqgt/ikKzLjEwis17CEDIEbT4/XUxl9WZ+veL7AmpM0p6qjiAp93CpsXGh
nX2Lx1T4amqvuuac8qmTwiyhbGLmfKGUT6HCQ6J5D4A4u/mJ7faU9Gjb65bVS2UIMtT6Fhgwz+ke
1lUYsHP3rSM/vsdNAgFf5O2zznTdCOF+sHmnsQnm4wqpatYiDBJYvb79Gj8BM73JeuZHnEWnHUqi
3Re/4O/fIpqWcyFfv0tp3R0+kcBYIOP3/S149zFhbSvV4mdfM6zUyJ2SC7m8ZlvDvitGjSfe49rC
itwU1A8p/WznDAGJRQavvxkV3Ai3AJhvJuLIZi60B9w7Yjv3jWaEXfyQUbbzNXpSBdLUC9QJAqil
yGNOYZaQ99/OF5NaOu/nIWz1I89Cg+NrbkunTy5Vq0AC5EzpoH3LgcEu3BTWwmX9ndxifGyaN92+
q7FgO81I6inK7ou6VYj2D1tMaXpFBKonzMGeohxTASlUw2cuU2uX9+D5dpUarQQviX4NV844vxp2
88O59QX1le7PKRxQApLYlAsJ6xwJ48mWc0ue3qGE1ezTtSX3xWairZTZHKylGCVIUwWCqTQOUsV4
fWkSGumrds0Cmhnk9uk2pwk650jnsB9tlaFsjO0vbR4t1mpZe029JQMonUEmKYtMRQ46TRQAhlfg
+QZb9HagwNfZbjvbx1MJIeUtQrKnikAq6kHkw3AJc6YKPVFKNXMbP/gNoJNqmROFkKKkuEMW+j6B
AJdQa8ahZMUgqaFJ4JT8rfyYQe64Ki42nrSMX6EgElCOtN3BiovYlYZ50ZmgAwUgGb9vH4Qp0v/1
RL26O9XAgfe9MNAj9SoTRaOR9n0howK36JrwplAQ0o31r7B0XBM24S9a5N3ybrSstgrbHQb8sOC+
Cx56dVXGZyXbD3H1mUiqYsbjE2RG2ZWoEC5om+XJ0IzOiyg3cys/yO62k7slCEEcpZGwaYq34o2J
hajZnAQABEExfbXMU59MZ4NfGmL5UN3lQDPUottp1e0PgrwFrLWW1BydpgtX2+gZ/7BaRg+3+Fra
DcnarKAudeYUNGDXnQ7M0DnQ+QZ6X2V7iNElGfX1iXsuiMDgom/kxRQuGhO77/9zDRb40KibNq47
9iOVW8eqnuINuXuaAPzlYlz+77qwjnIy2P8/Iq8DbksmxhB0FQtHxci8Wty1sD8xYC3fCIFk7t2H
jGy2y7leZT62xtBBXU3x6XjtyNInSRlGykUbvCw7CdajobCqkHz0zks5+Mww69xvURXxvrgtzFzP
kmIkCtf04pJ9abhgLA+bo/C8kkH2frQQddBQZ6Kmql9ZxZ3u1JXNhp12iW200t0gxD+t9BqYIioL
aqZTgUrdG1BTfBkxse0nM506V3jkBq9oUvtaOXuZ975Kdw+7K8yYtXhppCQQTRTZ6U/9PCuFnWTi
S3X7gNKJeN1yDW64KazH6H4EHjtDoIeV/+mK0glKkRG3KMjmQdA78R0lBSg+eLaaRYQScgbWdvZ3
331b/eEdl9zvE6MW7cR0WsrjUEZED5zLVy21MwfACw3heBEGThgdH+BUOjo0ZVm/N8z12KocTMjp
RrQ+KwG4j7kuqB+/L2Nb7pSf/o+kBAmH5b6R4+51Jf/E7uxACfpOMKj5AvtzhygTwdrEdRkpWStR
mywOEzZ37VqWYvb/RRjphUA5JB8eMWYTn5LJHBZXthaldknwVP4uWf9P/agsQ8QVtb8lxr+0kiuh
bsf1rrP1cKVKHx6vi4E6FHBP9tSFIE6BhcxCg4Nd1IFAD9iqyvbbtULt62Xu7EruWqwybuaTl7C8
ahWu1L4+CsDIUBzuXXwguNaFHqLjMfYAZgoN/jMHYYd+715C+E8lFlRu7vt9/AvThs27wcl9rOGx
Nb2zdcDVudTx2UNXsV3TfABEQG54Tjdq49DFYvA3B1YbtuWs8d2kzLhLbfHXXjNctv4YiUjfMeA5
39/jzO1HVx/6Pg8swyF9N4sUIAGF4bh/SQxm8aOPUnAZdIv8oGiPuDahljvM9540YLPD6qpJ9Eny
yYjsd0BhcGCb5mMTiGRsEx9dFfEc6yxtLHxtxoju4wT2wmzhZjyeLbWczjg3WIM2iYjZFDVmH1yC
SozJq107fhTLp3VOvFAlGKU7dCunbl7BdSq5PrhFcQFPpGKEW3CYRxABEh3fbVjUpfbzuKVjjBJl
GLv6AY5Bl8Whf8r42dwkqdlxPULeT0Nu4vR8LKY3qLqqL0EVaQa59JWqZKPFwoaKBWeOFg+dX69K
tkmWSiht/EaFdiLs7YxHHyThH4uqce+5keG2dRWtgcqt4bZlVZQhjKIKnvVIUW1MkScwSv75tZH9
8GhSnMvsu1RCkUXOk/rEIniQanwQCjLNpUILRIKFZw7acLyXktfFFziv5qSVosAu2OWEuLP8BgIY
FDGV8rT60ypJfshxhp2W18ytwzMmp6xnUJSdPR93UQBCgtZuil2Lv+S3/YADtcJGwsiW7TkxaWG0
7PTX0ZjgmhFUWierH+6LtaV6mycsSd59ozdYQbMhNAxbNxiPTP8gwf6jJCIUJnbiUIFf70RG7xDw
OrSEEyy8XF4NEf9RqZPE19x8opYhpleU375Yvsyzy5Tm/Bj98UcnhpyksDXgyjQ19Eopb54zlDIB
Ays/+Eq29rIibWZZ+UsSWOrPY290gDMDBp5+3InJ0If/x/wScpsAz+n9FptNgyhv1CXwg5kGvskn
lXfPMGcHEtjWDV9t8tFjPIDDKod49AF68BqbG9LuPSTl9afRW/PKSkjyF9qDDAU/syEIl0skTvN8
tkY0dC6YwXc/rXX99doNM82QNpHn3WKFx4sF/5oywvX5VwVb113qvvTFSJnhUbYd7z3dl24ngFw9
yPSq/YKB2cd5IG5wxmZMRaOtI+YLD7vHZaVHaqQ1Xj4wYO0tDPLhRU8wS0G9Ee3YW7t+zKQVn0vr
Wnx69BuL8YqhNyfgOmg/1twzoRtqpdONANNp41TQRN5W+2eATr0WI4fLzQXBXoh9zdTpXaHMRRvA
jhho/H/Srjq6bev8vLn10uwFcwHSzWYq0Idb4YPEdfrajrchdTTPRYpOew5coczn+QDAkAKfBUKH
4tWW8D2oS/CGgcSrjyHgRlBOCQbPG5oT8p+oVZzF6EFgl+GVCsjVBcJVB6LrI7JSyGU2fq6RxKXv
fN6kuF3fDD28QQmVg8KIf+H4bEJG/0hQnAEjab4IydjlcyBt+ohdDwBUwUH+1+lMGJ0P59eQtoKa
tQlHZKrIlg+CV1+a6fU/QgYwNO2C1/JKoZqYQ4Vh+aupWxe9nBonOu+zgM9qDHxdZxbhNrCgK1H2
R3Ww0gAWK8/+gLkW4TTgj3GMVNGah3AABD6jN6TrEOf5hykhX6KAAgMb0D0ZVwvyWGMDc2ED0fx7
r5uVvr8SS1IYHyi63SSlTHvqiMRDsMoIWaq06Jsva39LCzarCH7ZidlytLiO9rJLnmu7oq1S6uLD
+C/7VTFwh0RNdzi9HlbEYABaRv/TzsgZCR8pRtXXChMAg4IlX/tSqVrvlBCmk1+gNw2f+5DmW+Vv
JlR0n0skipx8FiSD15XMj5QkBYPkG0bs721ZP0k8m1qBu1o/SBFSKe4HknhRuCWywxE5nulFOvg1
MM1jc5ByNd7pLG4NQ15sYXLdqpS3dmHUPy7YQhIktq0oH6VNqU7f+BjOe/IbE5L5xrXrmKOa/V4K
TcyKBg3qSMQPejM+a6YovpJBrOEo+5fCMJPtMqJWefnBHqyXtFRczB5E84I6OvnciDvcOadzJLWp
TZzxhSWfWGA0EKuhpDUy8DCwsxmeC53NvE3RaQbKIY8d2/eIKaYBaeESU5SJjlIzK2cSSOqFhc0Q
qRZoYmSIaB1cp8PFkj79ewz5aehQBwWbrrs81ZjnwYLNTfiVapt6rNHsCeii8mey85/AovD2sTM5
9BW/9jfoaAPU6W13QbcC81LrlFPG7p3luqeYNPYmNwppqNPP2OLsGXRjioxZaXGDUTCsjxt8ZH20
h0uPlEPMHkrwMXP2rpSEstRCk5uiWRd2tkw9qniFq6voYCx7U9RWKhEHadowI2ln1wbWXOjzKJqi
VQxZ1Y/SQs7Ykt0nfeTmB2Kg+H6x7aFOBbaHwhFdSplLjFtpAdRcn2bJooImohzLouCmHMSCNztz
FWjHbDa9zGfjYk2C4HRFpr+cENzjh2Yiv2Q2WyVidOREAekdsELEK1zmveQPf9l5OVV8fRF8ZU3L
DtkDpHEg0spRxJm46jhn4u2epDZvPCtHItK4hzu80WYbWr1P/g7SEpyWk7LnuOR/7UCm4pj/+mYB
kHoq2FHv6n1aDXNx5GsIZVBhRKK60cGQbnTBKgy13NK7yJmMYOMvnliKpgAHYN8fPGFH/vBw6YPk
K2MyL9wXQvTdu6kKF4shVKRyCGpGnof/r0uOUsQQridtJSYFpyYMWQQS24vAkgbZOjDlwJhqueIT
H/brfyiM8z3QvPwIK9QtLVuwW4DgswqSqHGrUEPhVh80Hd/hJ3cQsW5iPHsDJiiD5K+CIwop2vgK
t6XdbCZTj24UcYcY90waxdxKqnX97HIoox9VMAnYjIOw06Jhv/HdkydNrkDtjyowHClEIf/ccCOH
SGh4CEbcMQqMhvfEFF3EGxbcOzEOE7C88ZTxtuaIT/cVzkt5ZzGXgnLedAeCbm9zY7JrLvcAEp7Y
9AdTczBOZ+VdIgde1VPy9+KHnzr4krRb2gRJqLxg4210Ssrae0+LTvi9sMrBL438Rcb/jvTIE2x6
lGlmzhpKk5SFUmvu+ocnuwPZqfSu5pvmUdz69XwIuI7JBDeTbNA8pYqQu8oe03X8xKM8hur+J3qO
2h4Tm3epC8Sm0txPH0BmS48D8xWDZPWD2m58VR7osxxs/SlFJKZ+vZ5DzxZmoZtC/BKNJ1kIrpKH
Q6CdHhX5V2IdDoIIFsh5nXR7DeXfqkwKpON3HN6JnoPdml0Gl+DOFriJbM3wIGVflfIb50XH5YUc
7HkXO3aGK74FGeoIryr970QzB16OItYWtcK/JBC+uEXrGm4BVA2wdEBXvzxbjV9U1H0Xnp3LBqZs
5Iz05LKmPkHB4aLeqmnRa/N4PiJ7ZZDg7i2i++okSHGRYB7KE+G1Ca9Lw3U4Dkz3WC31CmCjQQRQ
kIgSMEq6MXvWP16n07z2SOIkk2zO3E2Hp964yehR6B+Z3voM8r2s9hv+M1y9XNuCRx50iqbG03Bd
nUVDK2ZwjC6QfNoSIxgFrq+6Txa+liP4148mxfdgU7GyR+No4UNZgqrkIdVHmjky1oJmGdig1dPj
1aNyyP6FEswpkbITvaCYKzIvPkxkiPyfjcJTY0ZX9FocxG+DufXGkg1p0v97ANKpMevA6RiFpVpd
EFkAv4a9vxlHEUuHjiLA1mVnAfC52cjv0G5H/d6FN+5R7I1dCGmKx/M9XaZ2a+p9k8+dbN/5Up0S
DJCLS3ECcbHTwGcVO4WHFtMJsWJ47ZMeCOZ0r0El7IdSxJgQ7DPPPN1+hvYYr8QN4EXuTNIoRo8s
o8LLtQL3FrfnwSjJEE+j89NBZn5MHSLSOVljmjCEoPrcrKMF8Y/caqqpGpMPxM9gnUzLJu0PyGXJ
7frj3cxvwo4aSSsVFB/4USReC9OV2qvKKpC4F9WRMl9DtmbnEnuFe0A7643rO+fPdgzncfcANcrG
HcEHXF2cIAVGhm0R1q3eq6kj6v4E/7jfISkYEP1lxeG+RuXYOZrpGoNdbgUl1+a8BF9QudIPZpU6
MGvYndFj1sBDP5N2Zz6HUpsJ5Kz1lGcQLtH5O/FvjA1Nidi6RSXLY5aRsfvPqqkJI9lcmBWhPg/4
XNrILqAd6ck5YDZcKTSP/W/3A1ppsjiZhw8wZM9MnwBGDvLooqVkK/klKub1vdgwUhNLUEk1vLme
iNIb3NHjDlsEeeSfaEZ9RoDt//vKuqm6ltWWsI+K2EXGPPAZlZtFSrq0KVOxrjTmMuq2TsiVoaM0
e5FJ4Oi/xxWhfg8EgMbbaUjR+6TWH5q3/wB+sxaEMtVrYT9b79SEyEpsnOcRmCEJBrh/vJ7Oj4Bv
uJDNX8hBLEPeHwsZVgyU9gO906gW1FXc7uXlAVYPbeA5kiax9QGvfAycRWLnwyGDdaJjEQnNydN5
jQtwhxJ8WE5Zs/sVcrhxytoUoth84Q0FocXWvfxNXgmy+jj74ROZYADB/l76hlUttPkhZn4Yq+gZ
eGhvY1cZlmANy7MX1MeFIwe7EjEs283sEBBa+dHtPpvVvngfXjPtd/1Jx1PJ9A3n49miqZXsBMiI
3wo1WbbflGqURF2euFcFv0ys1FdkmFsmfRxT6pomH0oiy9bdJgc/3+TzsWBc2+br/OoDGHrQGbun
npw+1SFrbKLb6qpmcwkRw9sUJVq5aHDrGE9SNV+3rt9XmmC12YXmm3rOH5zDiC+sXrnCSK0FoDOH
olsU1mostcIgc+uWxNEhUFvXG8l/kUIBUTfXLHy6UQ7k/mRzRghpGzwNmiSVhXTyhAin2Sa3hjlI
t8XWEn50QYPeSkF5We8xmjLjrlXPbDnHMiOIi7kIKwAs5nuYiV6Zm/VQJZ7TLB121529qQpmL2Lr
NSWBUVloW/IXSWDCYhCmaksxpCM9B+y17kR0WWONXaAjmv80Blcwu7FtoDCnAYI35ipwJ+tZpBk4
VqXG76X/0Lz4ALup1c9wIPxMW4BeaS9fYvRw4tb7DAgBE/o8h/kKk5XZV/UWFH2S38F9x0cVfLQY
QLHc/jYsc168oh1wIVPQddb6yQCmnwUsWvGuNK0R5y7H74Uv1RY5MHPu3sz+E5dhc52Pg0L4DjlW
GnssigXJHclx/EWV7u+vk6RU+jUrbwn1iyBuadG5L+g89zRC8Fl7I5pHI86mj3ZN7MLejLFDPbht
Yy+PV/sgNjlcr6+TBxvaGsT9mFwa9y4suL3qs8CSo2kzPQHY0myYayKixYeR5SKVMm8vOqATEaIl
37XFPOGt0w4HjTQqSYmWYGd5gB//RLNX0cAvy3/mio0fHoULadp9Qe0sqqMQdDug6bGH1K592F9Y
zrcqvu89v6nspUR9XKTbf7aDPZ/2MOOSQHpbPXGYmU5GWReHX3t3u+gLEM14ybwO8R9ryoBFItlq
MuFrZMyLSmQ2gSS7/HAg+eKrjOeLYqazj93LuAfQDyhsGc49jIhBcE/t+Iaoy3xDWn/iwahtWmC+
fv8oL4RDXI1Txi7QT19TC1sBNoxSIzT0nGXbP3etdgJihXMohb8UoHFzQhVPXTGZSrvmgUl+6QTE
IX+2Irn6BtAGv9phqmn0hOtkIepfrzK0w0fAv0ENSOYzcTTMvR/w5Efrd1dK0XxqXrGlpyZ/mpaL
ySlG9tYg7GmgD8aJGmv+1iKoJNJrTcVOJY6dOhot0YEmD8Ft7uFQ7gqYQvVwLQgjJXVE/vFNwe4Q
irUYgXOfHcXv1xyTqeh6/4E6+YzLPeXvmLOQZo2OyGALa50TSQU+Iw+d0cLN0k8tykMvibdzdjxh
pdfp63GHz/o0FMewQXbKp7jXCYPm4tUGf4w70oxtFU1QBOtje8fHCNTSsXcntPSKl/YT6fDjVPyz
Qmga46kTzFo40nfK5vP/8c3kXzQ1OxmYSe+TV/AOIPWxB+0XPNl3s+F8wEYksbGOBc7yJ+wh5X9L
5uM6rw9Tmag0/7ZD1RNaa0uQHlPJ42K67QRwgJboftta1IIlQjMkOk4XQR/lP8E/f+I+LDQKaxKV
pF/D0SlPxrOdsRNSW2gWumDe8juV15gL3pJJ2s/K/XAx5Qc2ju8w1QMh7Nmk0d0RIBIG4wf74Q/P
aVTuo6CwmotRacvtHf0IeRmIIUVgtEpCYlSnih3sZjJRyKYHvWhhCGbbvmWszLVH9YpMYoVdURSt
6acWZZs7uhEJjqV9JYgykA+GUrB2IzhBGkBgXHConQRvTZ02YpQ1mMq4RSlyqmDiONdGopfwDRHA
aaBQ2tMFfKCpYuU8RvpduhrtO+6aFitr8W9lgcLGICpkbCbHN5d/5rFm9VmiDEwQq3bL2lJ60zE8
L721aJ8vp2B0tc0WUFcA+vix5Cf1NAzQ++DIM/lztFVtQSEO3EfAfbyMV98NFzw0KaVPe/hKTIsS
wjDkRIke4pIZZY9xKCs9MTSh4QdBAYfoehikp26pglN8cqgngNDqfv8kuje1+6FPwik05e8/Ofy+
6yaIKfNLduzDuUxRrb8NkK5MZ2tLDZIeTjC/S+vPAzV/DLpNlnY4yaWg4wMuUmbgb6GX4N8do3tu
jISy8dxVAsAiNtIAuNgOlDLQBEkDE8U6lyS78+vn3SfUaN22upspcdQTItdF3NrkIMk2ZoUloV/1
nZDDjyj3h3oXXWj3j/9htxHpxOcXrYfgpVDDbssFb9yd//eUoILqsJF4quknZNP1iMfjLhZH8Wj3
psayRH97VtqWj7TSCepCf9wXyvoY30TTlod4ofQrjDy5ROoQNnbdtFi30dC8AGP7pZbSRwcCGDtO
QG3OdP8p6yCbRFTbMPwcv3olgsHfa54mSdowetyXFpzfZ23VnZPHtgF0APAFIk1d0z/cSzV1mShF
A89ANCEoqNUkzFUl88mrvYMOL3hGFqcXGnUque/WLV8g9mogTEX3+PNa2/5TiWffyAaI/Fa5lUvR
5wX64bWwunQO0a3dUDnBPkY59Py6V71juRoTK8122Hdoc/MBDPXOpucpqTy6YpMv1JxIbTEZX+S6
sW5Bqs/n2OWo/Po76sUVaYmKlFwLNSEyIf8q3IHkjlNs6S3lz8B9b6IsdIAtlV29dy8ytvX7ESL4
QJ0G+BRJpt3k7YkPoIcfDpbG8qDYuDEbFIJO7C7lpebW3BGB2n7FRZrRLpb1urkggE/TAdhE7bky
Go9D6bPGAZBEUcYutRGrSz0dDNC9Co1eUDv8jnQAseYznMmePHehuToOwjq3dLYxRtlwNk2ttAWU
9p34YJ8XdUV5bwQ3db67V9venj8oRmDsombK3NPGbZmv2CuS6pDrgxseNxaZhf0NBz7lQXT1fBET
2od8W/1scvfCe6yqM9TU++uvLVNm5cZTyh2vGVB+XIptKC8Eu/eH3CzH5cxQ9XR6aZsxezNM6vAM
uKVxGc/3et6BZKkgD6EsED+s4dbhsddVbVJcO55wQ5KwTld2YF8EeU1V7fWP/IIfgJ0SN6Fy0ldm
jABympcateUWLKga+BlL8WFZR07PwxR3jYE36NsJSbRZDzZkOJUTIoD8s/EBTlJEYZzQdtkWymGM
GeYPK+Su1hcXZkS1wA0p1nsZjJnYWQBVBcy2upIP834Frg7AdAk0Z/qY+iCrFMZgd/gIQp+QcaRV
uAEfkAz9nCkuxpu6dwo7lOHU/J8jMbfx3pxL6Msw5UwROT6GPHWTZ8N/u27wF62ZLPHst1rvoVVU
pRaH/4bp8O4HRQA3zfVaDXG9uOL86fG2swnC2/UKPocxfRcg/x/pbgJh/Ie2TFobXQQEI54QAHDD
HvxoteXgMClWPE2mqWSOfK9JmIYSW8s2Sqwxt2uMKAF/a140CIl2Taxeaew1xAkubRqwKVjPmoqf
9o5LZtf+q+CjBqxdKcZz2UVcVwCRH0tOr0rrYJ6e/Utb+VinQ9+o3/m41/CCyX2FWpEp5+z0OSXU
K4cW27v4wkkzZw7LMxTMPMXtbMXbO2DnpJFpLbasEsSmUSo6TMIUYmH01OhdowyfSLiE0s9psz5y
0b+6RvQ1lEu3vFV7Iv5dLde5NwhxsjwtKzxNFPqper6/enaX8LDGbSH57ud9RY/Ja9mQjNUEsEco
9y2siQQzKkW79Xz71EgAVYRtdIHNmWpHoErg6x2y1Zc2FZjNVqD18toj+QLF6qeQO/UB8zSFiu2C
hB0iekGWVrMtR2U76/WS6LR4xASstjBXBe03EcZm1Yzshu+lSwmSBnfloF1fZpHIG8HZXfkYEtMA
oYC9Iy47TH0J9Wh72KeRCiKCCClkmavXu7mi6i7kjrT4X+kbpDhJPq6M08g45BwBrfp0PDduRq3d
6iq9D49gW+Mef8cON0d3N854KD5MGh/sbjmIvaka2c2bp5Lrs544Agk2Hf3cI50kNdXWqhWKNaDl
BOKKzzpqeaVC54VJdPUt1AyEHYy8fFEYuh+4TD4iCLfkWpNcJCEqNSwywuaRyjFMPZp/xW5GrLbY
Z6QrpF4xWRVWDE6my62fuTf3TVb88HQalib7k/Jl7JYwLAkxK5X4xjwzwLWNygInbd48DJS/BHL1
Z6Vj6+xulys6Lt/YwAK7DmXF5P/JG+tsRLCP6ShZxqithw42eIEVdtiO9eGfhc/4jBgbOlad88VJ
E7BE40nsOyF0LBvex7fsOcSydhkYFa+PnhF9blqdpw2PBfamHABd03ITPnAo628IzW7/yrPLgDNT
qxm9ZaEbU/R5HF/zdRRyhYSFAfsv7GWJGIj7vgAGr7S+mB4RBqTw5HRM0enXMX5LuKx6oEIKsBxh
ZythiWohwN9B7zkMcQiztMP4/kHWBGSPdkFvKiUmz67uar3pLKctzwsRewqaefvX/H+9tja0oTQF
IunXs+ops0nF+T7tsKT5XFeXLC/ddbBuMnVF4dH2oz6jO4LTvNZWRBVSSfEuBwtg94LanoAixpsL
733TIZbzpZn3Xncc1o5QiLS8wXHa91XKdo9+D3OVSAHmJMErjUMjZIUIQ7V9wNvSv05y7j/xtN/0
zd0fDpfQodk0TDPoNwNjXd/SNr4TXyh9nvorBuVnkPRgnyAx+JGSeoN0N6NQ2dHGga7KBnPhHCV3
nrbGKjk8u9z9g+oJwmEXz1KXuXRRDJ+0um3S+VbtjrvgQx5xBfBDUS4dQNjjfg6IJNQd97EgFFu2
lYVQfAKRSHRF5aadCBlTyeVYIcqjWPmIMtWm2gcBiODkMFRhW75QbYvspS5ERgVzj8xUChlZPLrZ
P3AxG8VE5SFZ0+rKfjmL4QnS5JhcPFbL02ihgk8IjO/Ft4Fi8fjyqHvUWVV0XbdBiRGarR11A/Je
1e9v4NThKz6zglWpBKl3je9Y1V10vaPSETYP6/CKcO59q2/Rkt+U2+0wdxdnEUOm+AZpLjG6/GLA
3epAVn5IGpnlmDHwDNw/BfD2N7dd252hQoptpdIOPVJxXoQVMdLiX7W/RDcqcOVW9T8y67euaR67
SH5fo5OHx5uCAcr3HYqJ9mh+sYte5neJhq5k5Hsf0PMohfiuJzdkuJPGweZNxrz37s+Lx0zsz0mq
/Pm5w4qdYeQJhZsP/xBGN3qDRZMIjm/z8/oCWeZsPZCLJIHrEesZOOkvVmY53TpXOloDvI/ImU3L
KuD2y3L1Etzc6YqnIqRrAFhSAOQqHbzxrRCVbjTRB3f+Vm7hqbrltijMhlRV/YMEy6iPms24/Sk1
git9yKfEesWoGrBH127xnv8qrPULB82RWhHxYh0C5qCvLRHVwr4lY75dYI1lAceDuRvdKK28Fo/2
0tHVAauFv82TH9FjJWx9AwRSP/1N40nK9fSwqUexO++/v0N3mdtzltJxngRZ7lbvu9G6T6sQllib
OtIudAuL6QYaF/ZKJ5xLdQmkzNG1qFbLLX4mGOw13exxlE7b0hwaJaucoNjHLoSGOUDaK46KskV6
SBiJqix7JMR1nvz+GUXjOjds2Sh+Y70w4tiYkH3QKQ7AUx/E9aMpaXQ7rOsga8Uxmzbup8YAknGY
TB2y+wfqUACdrUkU4PJL9IfUN3WTYSJ0pNOmUx0QeLSXTGr4jQTDekRiVukfM+z8IJOTOu13y3Rs
PBZKWECZNILeACXnQOX3ofdEL7ddnkm9UUuHgvxLri3NHm3zpyuFRd7nfNhrA0/t0Ok1Ve70g2F5
XIhPU4mUXXsG7uLVYYoJPre6aLFJPIhAmTjtPZO/iFl/RydVwfyPP5sDc5jvEsglcjZ3XltC2jAf
otRs/E5Ym4/Hfd/Z6/NjJYVoFpLUdqmu4A+LETLanGMzdBumlwCcUbvmHtw5avTaWTBCk+MvlpNI
Zryi5J29PA5ZzKCsz2GHQ8ruTu+kyojNGOwZ3iDDVCvch0YlyzK04WiY5bqzr/n5ctKQPRgosqLh
QDKddZe5jAk+IWUEcYyTw9Ucm/dB3fpYvrHH/B24+uLdhyeCltoelImE5G+R4gRRLZwCDK0yYRje
D9tJpE1alhBNopusS2Z6swftBFSQ+zjFAXcAh5HY45SxpiPQhXMExvkJaY8yTfYf8iSwhUmATkfQ
NshndCOeq8A5VdFCYXfPDO0gAYNGvImVtwpnK0Fh/2PdortS3eKTaA4Hd3q+4Lx6bdHsO8kWXgTl
KQBQha3sfE6Td85hdOScdp0JoJusVz1wfR+jn8aP41qVQt5S9uenTwOx21zLRwZZU43WDtq7edZ/
bSWKtlp7NnfwwKy7p89fKYWSnMtK4GfI7azU0oIPOsco8GhM9zreO9gWEq1Z+2vsGxAvrStSLbA5
IdbR8LBar/bYEaCtlwb0UFycbcM6cdPOh+w3QnBvOk3Oaf+ttsfXc2mq2p4HnlnODXfr5025+Wvv
KbEtXO1D6n+4GOAimbhPCbLirCizGeLgZkEcSBc3qd9au+vyUb6+GrijEsfe4uWGrpRRG4MWFwqe
pFDwhMbw4psmbYcbi5q7lBZDQCDxqEh1DDbFTlqRmBDEvl+cS6KW8T1Io8iwNp3bz0gmvgiKk7dC
NasxADlUkzJeduIhO8bQQzMDESZrXapMX+TZ5C/1LH7iHDKmr6u6q8+idS1mUpM+6O6jFOcDelhC
RlWWgozuHilQ+jOLUzwdAbU1LnZuEE+8sdNuE2N3NefUsSpiUaZGN7sWcm1uR4FCS0QqlcjP8cUY
0wnu9ZBIYBAJV4f8ghggIfEcWDc3moPskmnRzRGp2CyDRGkqivL9/QVvRKj/DUaeo1bLvLpG1sYo
+h5AK3/MDEM798LI/bHL6u3KakiAh8TDq0VT/Y8hdMifPkRzIxZ2vPWlU2Ns3LV4W2zj22f0R6BQ
NavtIZohkRB3dB1pKMQglmOd0IorHCXYrVQs0XPm9FFfgNMeXTzkqb/LqTS71+vcjrDgcSWW63s4
ntMRYmV7MEnszBmdXoWshseCgxR015rO4xSf14PfffOCfuzh16qXapuGInvr2LlMlFK8hdRbdiKi
WA54rKbAJ/7KijcEDkGwcsp/7Glmh175IgQR7gyiSDUV28ogHIii3ZnenxX+YQXCEhcOpcjVd72+
kykk4pk+jqxuDdD/0KG7atYLoPZ0H1ImAE7wPUyxxcQbVOvjoly/vW3So5bHmwiS+T3FA0d7C1rT
SxisyjrSWhppC/yIezEAh6UFfr2+ZkIUc+RFKLgN7OGJzpkS8sWr52qkeop05AufgXxhYRVBbCx9
7qOzH/H3ZYOJuHTFc2J9Cf7e7ZZPft3/AF5dT326uPQE7f9cTROL7WRtEN7J8gPVF3UvSyendxIU
i8JM/FJVBq/f40Z8YvIBN7wx0IvuTrCM5SJEPSC69C3oRhazmN2bT8CO/srwchqADFjCmEOQ+R1o
Zgz9GQ8p1zwBQ2X3kiAkUZpqpSr25Z+svHDAoLt1KWf305jpzopKPPuPtc6C4wo/oECVnH005Ptw
7ufjFjqqUcDGBZUuRdFcBNcs+c96RQLBYsW5wH4kPtj6Uv2aJmX9i74LJWnxH8SYHAVyyvZXwYhA
2aE9mZb+dLopf2HTYx3IyoJ98PzVc3oHHFCQRjvfoAxDSJFAX0nDP7JVT+4AShzk/ec1//7BlW6D
FpgygkquDN59YJBlfcpO/uNYHyHPUOoS/FprFgv33WYbKkVzNWbVdZm6dQjCeOj8Mwzo33/jAO9n
72+eXQi00M99M9v/dC55lUWxW4FdOpouYfvsuLqqmhHuXOgof9cyLpTzWq2RvQnuyXI8wZOorcDW
tCZ+Y//MSmr6sTTcrW4LlPAr6gwTs7aIq6QGhoY9TuQpPseNqF+AvnQyVqa6lncP8gi0onbn9b28
KQOi8OVx0JZxPSepcXwPXtSpT48p6V3Ed8B1QaGlcgkdb4TN5yMimVir2VJTMtTXRVBMDjiob6oi
4HFVh2eDzMdO0+5J0TsgLamU/LZzxTWwwtql2mGTOWK1H3g7x7/ZiT9kGb1WO2ul+EoF5D0PUqmg
+4+907L2I927X5VOARwBVA37xz8uzwiAwU6aP99wk9N3u6LfflEm2dUFdp3BQMWCSFFN5uze1AXt
asEdNHmtOw6txAsHcBFLA862KUrLH3JYp7Qzk8Vjwrg40OLwuQt7epjw6jGPH/SqBNurNv19Vtca
Sj14OIPBzBgJ7a8SPMefy5U7djB0pwKmf7aGJ4spJthYHQ72Oj4tj6K47ULkO7GTVxquhAUyvjii
/AHsVziOZcsJYx3iI5cl1oSM5RJZHhSdpml+VKM00ByRalYX0FRPe75LFLAwOIX8iSPIDruwT1Pc
cvJAzkXhlBPMPuOkFQ9U5r1poSrCLfT+0NA2OZwLOP93gaSTAXWahacY9t1sfv6K/msMPQs3+u8o
rwjpPf6ofDjxURK1zVUs9u4KeevKqCLlw3ivb+3KaNhv51mIqEqYCHOJDMXWOyBw2E9RAaUOAJHE
WHm/WfHSL3C6OLZDRssxGvtrGB0fjcm4QG4S3MdlfCZ+jAeMT9Y/nPBkXYv58k4CQ0GTYQC533i5
eOodjOtfbA7EayfGOWfQK8TL9SJsj4r/MYkpuGturLqXNds9yIeYIoyX/4QPHt0utTKw9HjSZsXZ
H/Ng6ygIsZ6zlXJXB2JQkfYMByLifj4bvdpA7He/ImX7BBH3HX/I3ESGwMm/xtSqBPfBVzUvQE0A
9lj1uPJ4M1knWBHTw3GJGu5OrOYvj1X0/6kq+BwiRrFEr3c8xmGs1o8pVg1TBpMrkoUa+x1QStYx
Q3ITGAvY+IktPh++ZtC3zkwly5mKkCxlB/erRf5vwuJCkmjtubU9GHhU7Kt1RgGROBQcho/p+nJk
hE5l51PZs99z8SAsdIgS8AWkcgwFVf/PSqPSDSL9sM/For5f+Qo8ykLHzTWa+F0TRnAtkBYxz/e6
AxMX4uvKc1RwK9iyL8pszSNB3/5ioqNvFPYvCVPs/ySFh/Bc0LOGgXsDbtDufBufLklrmfVR+GMX
oPSvfnOKb+5oDtmjtBsVxgURYzYBcb12wYJ14q9oJHkmmtkenicHol/tC37w+agdqGo5uBW7P3JZ
6M06YPRTucaYco6Nf9daCr+cEmbOhtGWjDz9M4AIcE2tErH7VU5pYVBFeA/TAZd6kp9RoLw1bWKc
FLHwKqNT0vegQriO5WHcNVjG4KOMgufKELTd5/h0xviBQbRN/gJFv9HjAJ0lfVgmPeNCzfDxnnvD
/iLTDLFj2urSn3ZTP/klifMSRZIF5cNjyZpRVCDn2ICow7Cr2y32iqZ9N5gq08bpxF362KgrREAp
H/n5CAWB6Vm6/A+FfDlikMUPMwMSUU4ZRB2JWCPcHe67oMHapWNvfby44Ky997OMRE9Civl36Siq
6krNm+3RnYgTTZuvz2j5P5GaXY7HsnU2wFaeAA5X8njYtouLvv8o+cxZE2Gvw91oC92gWAMz5iIm
XgjwpZaC8nEZcCw6jbFk81YUJlznl64UZTaaf1cVRtQKpdIlttX/6nuvuVYwnorLMTQ4KATGLTh8
YiQrZqlYXNVmvJp/B7K09VohTq40cAGWbFKNiUKwIuIj1O+hL0SZ0ftAVMBvQZ4CEtzJyJGwCybG
YOM1Lwx7AHvbwofRBi0h01RIBO9ax7yzvvMmmE3T7E42RVMsHXCkarnigp1XRuWh0o84eKnXMswK
NZE8c3SHkphOQBOgifcU60W7FVEJvRrdlVPrxNECdVuZcisGMeRLnqHozui6ZQOgXaqAhx00zFc7
vc0CZVPFfjuZ5LnTmj0MfqIEtDvi5g3Mydeb+K5PlMM3fcLfD9LoqztJM+cWKHwFCRSHEENQQD5B
HByZsS/VSXRFXNtELtjcBe3W8E7b0PccVZuOgZd0r67+U4OM1zKO8OT11tVSubAmoT3BIddtCiTI
j66W4DWKtGUn4BK0q1xZ/2p+2Ee3fnMCvUej/hqFccSFJwSWot7i8wo+pvXa2VFdZvC24IDw0l0q
QBrTzQMOX7zUrZPGA8FVg5A8n0O/vVHeTdjpPR+l+uCIfqYZTmaepKSs5M5KTRxFpRFDHNCbwllo
M2pu3cjSCAEXkUkZ6rwcVy+PdmhJFpHcP1lUgtF1nvXe+EXgURnpWZdlNmfw1rSnN7ALm+Ept7Yh
no88yFbLfNltQMptoRgIDQuxDxl9ilIrcugyIfUIrjSynFWTkZVqanFW4lnB1J0hPkIlBlghPWGv
vf6g3z8sFO98tU5f41trShEK2QGVgvUIs1Qbmh8ZNjPp1+SdbIgc9v/zchVSz9Y29uOV3q45lpTB
5Qm9XJH6/IfQGRmFLC39xNwxDBKgKmN1ffe016T0tXIf2Y6uWAChpBV8leExFOfHBknESL2XqnYr
tOMVzihZiILuxUKuFkJhHzR0t4lTHjP+FnDWSNLP8Bb6MKLUofKutK1r83SVu1g2HtOHFV6Nepvq
lYMLA6E4OHrGXouxwrQDf9s1bgz7MiAY7G4ORr9p/vcTQ1wZ+7U+0yBaTqDkx1bXnCg/5JlIGiJp
qdna/VGJm0fG74gpHIjhGel7BLsUWm1T8klLBh05PIztftSa1j+09b0IErGr3S4aZcvIKMx5Yk35
H4vVH4N7rYrQGWrijdDMMQ6MKiQYBTIP8JdA1SGzAUd0BSbaZmbSszkbA57vAJsD3OCaDhN9d4Xt
C5p9dgzButpGBGtFP3rd5IrSk5M6ajSih9nieBWUHsEA/nePSaLj6IPLV/rQRUeZb6lgakQ558Ow
vafzGpoElr7cu/xwJlffBH0M1Vl1o1htnsSoH22XRXSHaeduT70jyE1SeTonwHycB5pgDBAo/qQq
0+357ws5Yiwat3XJc114sYaS97DULa/w4LDVxCKG0exrbxDo+IjQd4eVrjYhuOiA2Jj3fo9QZrpZ
lwxNwt5vcPtpsy1G+I4VBis8Rd1PBLbr4gVJTxb2hN44CtT0NFYEEQiJ7MjMi1FUR2yaV25c6QXO
SYMvGqig0HKMoyTGfVpzpDzPlPSXVTiIX0c4Umz6NddSCY2r238I0L4jSxL7hi9pTRxqVdewyX10
7mppm4eIcFXSPhIcIwoyhaRUNfGcy/gYiwsKyO9p/INYjVqHw/i0RaCRCjqmCgKksEiZ/veD+f+S
t8Xjw6/rcHQqWQx28erFQcbdf5Jqo3IfsKlDiB6eIRQAtDhScz0rQn+i68Tokn83PkW1JuXE+5DE
5OGOpACGpWYTJcU1mA27GpNWnXZtA7AZskypF1cwuzIZVgGlOTsYwCZunF/GN6HPYe3RghgTw0O1
3Brf6poLF1r1xN+N5V6J/FqR95Wuxp/rRU0Jm+xef1sIJb/PMFVynYzhDVqBPQBbHQ6aKz3wTL/H
pMec0ieWv1PcLYj3hIwRhR51MhzL/6SXc1NNRUrPkEExkf2Cihvrl+8tuHo/KlKYwV0JL97che1U
mrEhyZjMPf8BcE/Zqr7QmU0FsPESAfLfANxzTLYrlIqQXXnwFRpJZH4lIcCvb1jo+GP/uK0M3I3b
BOXp+98KHkYJFZXZ4E5CGNgQ6rpcyZRBiYp/RsX36Ld2J9on5LgZeifkdTt7VKnOf/f2rjrYTIBG
heZ+7Z+kcBLLsBnPZaSlF+OcAQ8cnB7InimHeAFYFZCVEklx1qxxaQqNMr6zY0INdJvWt9uS1d/B
9rnRJzsn2XyURmLKB043ZonpAE9bIv9gzafZpKtGLowzXRjQaRcJxGVJs00VabyFL56QAdsjKkDT
mcbpPf/pQIc5M18FGM2MGWZHBn3ApnHlsNL3JsRpOVVz2E3IsflEALHXLqS8qj2EgJJzZIfneoNn
2e2RSVmiYcwl5byXsVwqoL673FTQEdBWIx9Sz59sjzAJL1ANrKiQ2ghEoqW1nSgYtZtX2w4Hg1CF
ag8WsLgZiKNX3FCHYRNFnzV/v2ZPf4rEo2j79rlVz1upayxBSMAbKMUlWpHXnxVHwvfSDSvfLGZy
ebEXzCj9aC95TpNBvvEf8Y5EEKQijRoBSsXTF9vzl2ipnKKJIuovH6DNGXDxhovgBqhuSEyctXjf
CHDsxdqYuqksm4f+U2ZNrkUNGD+ZoqkR2Z2gbKLxXju4fIZDZ8fTp87Y3z+iJ5AGfFkveUkXSn4g
bt9BabSKknz/e2pJkM91YAhGWbH1u/FEKOm5VD3/iyEMwyZwu0HdYH+dL3jpu1EO/EGKrLM3CK6q
ethKaw0qF1l9/xUr0WxKXYJXResPcxDpdIcag8Y8SPr5c/3+K0cFkusvwgWuD06Ume6fAry+YQqp
Vzgt1XGyeGhV06Mt9uJc6XfBjSb1sy3LIwe1/8B0WZsiayeXTy9VZ0jy9hxDm7BBje3YLtj21VWA
I3F/z/NHkKX5RMJdUthNv0A3rgqrfk+3Rs9XmiFkuGWqvoKtvVNRzfFlN0HMdFvbCumPQRUkYzfy
Sggn1z8qIXGY6hs1Kamo++6TJ8dX494hvKRMZhFPYu/Qj/xQraRNbGPS+0ltVvFl8ARGXyW3Viqy
CF3hzdeMv3TCZCJ4i5LnkPCd66QJaUDeEoIsKa+Wbx4p+L4IzJZmYzeiDz3//7aMCQHK7jKM6cgs
InWc3Ju9/oRDdJKn0zkO1oCFaP7YUeRss/lf0HjrAX9xn+LksE2JQg+mfWBhn3GQz1XGqFFn4fY5
shZ70h0cqUAhqE3dRrKlKEIdKQhFx/ddeFS12Q2XsUw4LZWVgd6ATI11HckitSdOyaO5q6pByfqr
FHJuts3snsirmF+bxbB9pPFQ8i8DhBFjfbadrYEUTKzFaX8i56u9mvSLi1hJdLtxgTO8+ynkaBAe
GVwRkWSFLiWZZnXvnK9UlQK6guEdWQTeMy9NRRWZAu0iPOH2KJ0NoxoJdMSs+U/cC89BI7dCfQC0
PJ7h+ZcM+IcdSieic2uERyxTkhVnih2gVeNBYtgWttmV/Uiq0rRUCYwSVDUty4D80lrKTFroNXTu
CJkCldBe5KW6fRvk9rkLJkxsRwyxstAMoIlnLVhCtqGaZYb1FYbKo1zckTP/PzIcazdVn1J6gdtY
Yc2GUs22sKu8HJ242FSY2gTsb6p5Pa43BEWIcr54rLLRWyS7yPN/U05w55iKfP9DNiSA8rqsDjMW
FNDxaM+xC3PvunI83+JkrTY3/Tb2auP6UowHcpXBSD/t1u+Yl8AR97iovGtvAL8uI4WqZBk8y6d2
bZdTIGiwDPZlpYhPfJZ/AomTDRgR9r4sixl6xETVnMnVhb1/J7gNSev3XonlPFsGM9BuYeHOAqpt
qbPMf532y0vpVtstXaRXR2bku2/g8XWE4xfTj21VtRzqPkTm2AqhRHqXxLgsHEdDKYjRZK4ekBhq
fzraxl5QH5HO5Vta7Z/vhqxI7SON77sOsMlFvLnsluq3H2lDljPi0nwu6kZt7zV9cOIz35H1tqIc
sIceLQ0PQrPZYDytfMlImuFUdjanWL4UEvtDQ5l9ito9RhA7ex9oOGWZz7laih2umFWQ4iWWunRe
6HoUwDNSoOTdyckp/yJu1ISkXVG0UgvnaYtdaP0nrO+is8i9342rLnHkWZlHfOkA4igGjTG5LiU0
NScy8zl66JhKVXOpzcLh78nYvMZzTPiiw43XArwyjOQxbJZq7buvAS+M6ydaZZiEpS55HbMQX0MS
5egHJFlSmDyW/CGFT2lDbG6FHLo3eX6ItKScJjCmPH14OepGwz5n7vZ2tkEHyzGiCnFiKOrVP/jh
t1Xy88c9yB65SdowoxD+Dv85nRGbjO+4yybh6ip/8YQ8/YNjjxNKp8nzvNv7lY+kiltbTNOJ4P5C
Rx2xvI8yg0zkrDJWcYSZ+Bzewfk8TfC18ohT/03eAzP4m9koimfP0cINUWvMUcp4maF5xxRUhzeV
z9gNw46wq8R7yesUc0eJuNcBBZrlSiJrf+GdxBB1mNgLYzAvo2AY66q/COTvt4iRS0zf9z4Z6n64
Lc+3bWNIPX0SkWvUpe4a0cwO8GmIMOg3Aj45BT1YNj7eF1MjqWVAAj5TjgDDB8AHxexT65y5LA16
bpKwiH2fOI0aj0OQDn7Eb/wDX9HgzG5sPafSjpuH4S6wKOQxQN8m58WfCcR2ctArM0gYefIp6Lzo
NMZnq8ipyMRCzgiYmZ5cyyXuwOyFJmavQD/XYkcoXL5L0yogsVpyxVBPq/A1xheY5FZmpdIVi+YU
g1YN5jOJ0KCsvkuk9BzmRAwR5wra9NafBrUgLLhK+MUp+JeLoSDq8YjbDcRscShlJTv2/YY/poMa
vJMcRgU7lnscxsgxAftKOTQc7q5csFBl0kGD1rxDnQAAcXkywOyQ4sop7/oeV/BsoGOn+lPX7rSj
2zV1miT7SVXKJ4uHElFfMEvQNyo8liRp69J7D0jPW7cKHtAqStzoRjPT7D5wJBNThQ5bOUr44YQF
HC9UFI8bEKo1LgXAkSZt+z2kytFRkvpx4VHx/v9GbY2joA2nT+kXTWdqMmJWTpWe8cbmZlLsd4tc
BTnLUBS1midP5GMC07IAwLnOgk/tK4uj/MR2OlhU2RmC+6rNa0IeSrbfPENo3dEQ0UGsJnT1nndN
J/tjxY8vxnP3a5frvG6Wu2NZZOqwio10UkX6WkUtSD1FvrOJEstkiLgxyQHPyrRtbhHgiVPKPEN/
SoKH0vXoR+DMAgQDz3l6Wrd+DoYNv6JoZLyb0pRA4d1TernUmo0k6A3Ns9jDH/n6zE6WXixCLBkP
iwx+1N5EZXxGqInBkSCMpDuq747Ty2W8RR8HLfg5q544asygK3DeNDNfUzXsZzRIlTacYxPtHoZx
wVTcB/Bvn50Ep5KCmjdLWr/c3ynt7sQVugdpAEK/any0NGZd4FVsb85YhLKV7Up5IYrL1a4L4r/v
F8oRQDwWZoLNliPjdWcb1VPygZQVcCCfSxhLJ7I5AaNVDbFcI3UrrjW13fP/4jXlfeZwbx72m0IG
CjkQsGYAMtmlYgRvKHED4AoWft/J1BR1TEayXNfP51AU+M7lXmXIcokzkA/houXSUyRH4VL7opyd
I43M6R9qwPTmhIC3qCv7e7YWW3RkUDo90xcVmxP862kQZwwk6Hn8/o3iBXbjAC0DGcVVGqq0UIcN
bwTU50qbik/ClVmYkz+X63SczGRLSVIebugbJnASjWGvSBK97gotNPBUKTbomLK9Ap4mi0oWoFtW
YvYhQG6mYp+YddfAANTGcjY+/J2EORQsL033Pe4ZBUn9PUtHPtAuHrGr7rFZUrYZV04DCOPkpjQX
QYe96K/tKuqdHKiiEFun4fKZ6VlzcspL05gzSfP8ErnXchv8QusJXReAYwb7giCSuSD6yuvgD6ni
N3X5WtR1Ok8phfYOf2CHlOTFtiaoQHswKxb2kfIYBRG2MAt2hYyvHBHmcCjz9sgYjqrYfeJ3LmhA
HL2Jy0HjAOceJHO8rq1u7CPYtY0lONC2MnbaxEJm4RlubgDv9slaNempgLGg/Fqv4o8Xv+ROYJfQ
kRF9bsNYVyEsG5XF9/afnlfRJKZh2QqIOaF5O8IYef1bexu27oJba6W7KxJhWJ0gEbgumju6AwKO
o2ny4shoUTojJLPxp4a+RW/CKOVzl8g3WBkfRQ7iXKwY2xJ2KlehSD3RqSJXniZXTi7urljUcc+i
N1cF3M/DVBxb496mzTrPfREyAoHqjj9UA5ei2ccYXuSsGViJiTdjqZVTWllBEST3f2CpVXlJ9Ckm
hUi8cdzI5umE819VVb1n12SLYpyTj/QD3f1SdLfPyeVegkVQTb0QBG0X1qNxfUIP/QWPa0buY9tL
V7xfTp2HB6A9RVBu0jmgMeEVSNErqFYsez0BdA0G64moX84uTEBfokNIZJyIeUcUnkwYGhH4v6ql
6BdgVQO0r2PeZAuoEIiS2JU/BYcxaV5NdUdBmKZMd9Njn+ecOOJBtLzOYZ34qK8m1gg0FiJC8iJ5
+pzK4iDPpDWUm9hVDWkjI+qSDf4JnNsKQXORGXAtOY/+4Pil1BzYdB3ZxG8+25B6yG7EiojbfPOF
3VxbNmj2DMEPndCxLgjSr5bW3+LrtKkcPLhkuWyiTidqXW3ZxqfuK940r9LxUD9rpK4iYHE9kw49
oKojvNLTQRJdlZ6OixNPKJgyrjdeXplggq36MXj9KazDCeHKtyDRxdLIOOKI7I24BJ8flWrV0ZOR
VGlk8Jx9Aj84M7qNhqR2ykWJDPXxhvwu5tPjGVIU3KM0f5AvS/imE41SDWQ4F46Ijxk2kMg8NKgg
Qyiol1aQFRCNdCQPXiQTBxKVTEFPUoCyCBYaMz9Ss9FDH/1juYh/h+ggAzYs2MkKT28/nT6UmNyo
ISFfz3BQkA8UxEidFxqHUVhtFe3I9ZAsDGkAfhV41y9Q44MRLC4aryEElOE6yh88kg5pPOHkHP/A
pNaC/wfa2giQ/3Kt4zaabu6Pd3fV2hnzI6RXvgmTkH+Qme8jsg7oH/fArrkWRxtk9a+KGtYTPjFC
VWIxpf1gFT9R8GSs7YiFgP3/3KED/+thsMQPyTiKrRazaoWfzWNjeVyi2aoSlroelLxxs0oGJBNm
9RltRODEPZoca5MPVFsIaaNgKq08AxqgpomB2OyozN6VF1bhspiLL0Ufqi6aU4D5uQXHWvGaOutr
sfOm7YKz0CbMYUYsZeUwkQb0F5DN8dDFMaj76qVOy5YCOU+dKmab8I5xMs9xfqNv+TGkRsZ3Bx4J
eiBotKm0V2YoB7lkUO+lrEhlU9TNJPUcuTeT9wXM63CAweepopRDzR5ZndZyZgIv/rpOd+H03Dlu
v/fqdEAmSFXRxBvOkIIUZyHTVKb6vj9wZaBkUMt+X3kaBHt9geXa+nIed0ZgG16wGHbA/9AIXHG1
UR+87+Gl7efBpAPoVcXCWK4/0A4O3YzNfbdr0E/ugXlA49TGINjxGovz25uLZAacK/R4Mg2GZmUV
lYBcbpNcn7UVGTfDn8dw+xmfOBFSHuRNBw3L670JNCC7W9aQZoGT+Jq6242eF7TXdc0/1QDJ/NXS
Wgq3zg3PY1fuQJbf/k+ZZikV6n/a1cFZAAh4orqCJ0TULXxqMEbvCp2l4j7Yp6+DKQGa5XyBJ5zT
VsINdG4tsNBXJmPrvUMrnOZEW4+4acDl3gfE2cU6M35lH2+gkuCte5Ha4lK9ddj8z1mhPDxq274E
S5neRthtlWUPVqfm0qDtSPW5qGaQSj00eNz/LV34QjsKh45oQBtKMaGOL/18UWcNYawRjiNi9IDs
xJK2wyY7qUuRydJ6KMSnsFF1W/7QLUAq/6opR9EB0Irm0FaxdSRWO7W1eeKUxHB95feK+GY8aqFT
qSs2izIRDn58vh/UbWRI5IkAX043FhXBflmLSSdLrgVU/OphfEnmBJSk+JXp7rDGxssMJKnarrw1
BG713NP0WXWTKDRzMc3JtlY4BcoHsuYXuOB4TqTgMgiRxqIMTH97gi6lWeqUC8BLi5hzJCJNro+V
0So9ibAARJU4GvyyfPHVZJWT8Yin+ibqJ4oDEh2wMX65lATI/PMxBhSQb1/uqBQtcXidzHic2P6b
vN0TA72zOF3b70JJI+zRF4KyrxVnQYjk7L/7qS6wgFu6/qBpwaDYHAC1fOzpn7+KWSakQi1Qjt29
8LWQ+6inr+6QJurpl6Fnx/6HXXfwSzMMbO7DGLOH46VPhuLmA0rlanuGmGiCXnqbG5zAmAyk52Ak
RN73S8gD+RBqXei60rhaXJWUn8uPxg8iQQYfBNamZ+jBOOqWMKwYUJpZ/owd5KpJTKlKcGvjIypy
dEKiAWQa+JqIbQpiht/IJBav0kdcx1+FuPs7/cnjBt1W/wtzjJB184Yfa3NvIubbKxRr9XrxxW9M
HWRPph2j19jFJPi4Iph4lcEoN+5s9S+5BwK1Gt6nEL61AbUx9Ywh2T40kg/C/wsAzwsvgSXtUTaR
kB3CDhIw9AYbIxIWl5daltMciya+FD3b2IOeexdBHVDzvs8cXtlxrQrYdc5GS1E+DWpDnnMccYn3
ItqqVtRfwKVlDsDuq+yQOKdf+5DpURzzJq8PEjV86eCGN+uByfnh9IWPLa83jSEgtF5+pzH0b6dQ
a7aUv6mYWVE5uAVaVbj7rZHCmFGW3HsUODcaF0WkZyZymqp01O+ZCXs3+A8zW8JEaO/Et/EWk+6F
ych4O3mY6xM4W0Wzvz1Ql9pONYOhJLODqLQGEQiOHcY4QbzeI5s0mGO4bqFESjZjrDvItace4Hu4
q5GqvlxeO+HlqrpGghzjzW8zxVRU9brsCcl41hdjVNqPADMlWSMq40Sjckw7L8eIlLbcj9Mzo+QG
HN4q3w+bDETqIb74tK9FyfB2dZ6ePKYVdfhdd0L4ikBTuGPR2zlJ0x3iVjXXKHyaJEiZUXNLZ58u
17UPKX01dV1aDJhnPPtMwK8X2iAr0Y6x1/J+v2r1rNisu7yo/Uc86h3e11rmNwAY1kaEPebfbwmf
RwxsONuXJ5AED8zpB26mNGvZwk/q0GoOLtYxmsAbnxfLS6RfzL9+fIvUgk/s8C8nYxnM6LPEhIAI
oanxOEpliU6Ji5sd/TY4pyK+Pj8JuaksNGwuze8VWfx1SF4VgVthTwQOn2lOgAAFgkLWFgRxf8Nu
W3tNMLWCAaJDt9bacQpNb/dzZbBO8wh2Xa73bjC39vB0RowM7c0jxadwGoDpjm1BaWO2MkaYPpP3
TsBwcqyeQETCmFKNHpLS1DhkpsRO8v66H3oo6lUE6IJbgDQ8el3/HgYR+0LxE1uHSEnKKrqBGSvt
xCZMC7iJt4RmpSgx6D0RspUPjqLp9r4EmVmwm28BvF50rAA1UZcXqe1WaWDbNwkBRBtlaRN+lAtk
9E9XsXCnRZFAK7s4iOEd9HqvBF1ifbwGF/fCQEgZxXiL7MMOLr90KI4fb0JD+F1+Qrtl6eQhJbgI
C9b13nuBVT0gMGSiwcUhW0OZ7nTxuCFhICJWZFq2z4EDDF9q91qh/Dz9Lurt6/Tt/9FQ8CgY6Ofh
vOxbm63uG+IKziOourvsclnGQEbKBKNO9tT442bSjgFhFjyX62eHmnYvpi1uT27zR4nfTJVTbDXw
1PP8JYiD+ISh/MxAKjzaTeKNELH2wT8Cfze25PNSQAcNMxXR5WLUhpQJNO7/aB9vnJQ/DzYshHxb
2Yra83gpLAPdBoUk2uix4C0SgL7oWtIAjXiYJ6nbjcc6lK1v6lETedaOIE4scsGiwmTLppUZP/7T
GiQ2oqkRKw4wn346GM5Jvibmo53K3RJQNON4GbTc09VVXo/IBABntuFHsVf/Ji0yh1mLx2xRSsXd
kEePZVtaJ16GNFBakWj5KS9DAGDF+Sr3c8hN0950QDvrEPJs9x3DI3CVYSKngvHvD64d5zme6+Ve
n7d0QFEX5WMsYVH4kslmbL7v8xUefeAtueGzWCNbQBkaL7NVC1r4xa1FKsfbPcZXQcFRqsAeWQ8a
4v08tTmaiHYrY3PcULbHfHpf+m/0CJ5yj40cRPIYcbqIXGHofbRuHH4bc7+uHxOFls/rddTRh4WX
1sm8NaVOqp9EPSpM13C8vVmaDlp9jnwA9TZmwJ9ZQrZ6r9RTl2Ddp/IrolGzq2hpvJosVi9tWch/
qUb0HcvRe+xTcYKI9DIrrVhhIH+ZUskao210Zlbmx7VftBV/vOg7aElx/AhQWTY9ud3MGDmlq5er
ICweJCDuYNNP5Y7p7vEVydO2w8tMcoHGdCUKr/BBA7W81NT0ZAVRpdMtiBfvyOOu/Ot4EatHo/H1
D36NeiRlbQxysJOa1zEN+xhrBMYFvJQ8NDCd9VJlutwdsk6u6N+8iL1UYgM+H/dnlZ/XFZ0ejLQQ
MT+XKKC9OI7NMX5tuoV3iCD1htnSNLUADdyVN+vkU4Pt4gPd5xm8HeNfQCvBupFAqu9cZxY3X2BX
z9TNkCc4tUTidDtSJ/zXnAZMqgBFvmNEuPuhIWxccuIEJEj0KqO9Gwj06/nCTjLEp5oskH2kvmhp
vJ/Lbfox6f4CksPu+4QMXqJj9fTYcvh7muPySYjHni40sXWCCF0snAA6SlbGb2TSCf9WVsxZbG04
T/cjFl+7AcrIxajhoAjYyfdmrVL1iqkt5/0roXdLfRtc7p7qsxAeOWKui7vnpOWZM2hn15WGaNlq
UmAOlXDbAWkC0Dt60OO/y12aN4toSU/47Fg9P4mlouZun0qy+oo2ueS9rvYUICl3qI4pfD7ElNOf
bfT5z2uTqVz+236D8kqDSmJhSJSURbMN3gQ+aM0LDNMG7rjSE2jTWjM3KcpmdrBHRG+aMLIRn++F
ZuCKcsWfkW5Xz5H/zaYjY87D+BugNqR//tyaaaLRCG0uBsorl7WSZOj7ryKM6eV4EOuVd7a7sD9G
C9rl8b+OLZqjr88Y8t4ThebLofG86jXgjR5L/6a94AgwfKGTkAaxXBS6YKSKcZpr/5wIz7yzxjNK
LwxxiFOWsDCH22pHeGSrWXJu3jP4eBYiGfmyRP2t8VT2Lbd1/B/GkKchxnkXKhmZRrNO+YTafM9Q
uOrpz/fE12dl+qru+UMMar8GDBkKgdcvlvYFJYxlWa6jYVdDnXDM/VxpbJE0Req6exaWsvAkYi5D
s+afVFfIaGg5wt3PbNMz4xF6N6j8+LNG40WhVrkKNZ6XRYaP73H+mE3kwzfcs3PrjepcjqxX6jgq
CxAYMCo5co1s8B1yT3c+Xik7OZ+KUc21P9gqnlnGkXvmghfEGdS4bTebWnb1xHS1d7GXpwBFOP7U
P5eddtwjUUA4HyDNehzg3B3+JvXm9apASGX5q91oVXeU1CdsfsPQuf57nbYME/4N5D/dvd+ueZxg
lCIY4vCKiAigwfhpaMO8LML8TT/v2xDRYKO878tliqNLq2anLa38SgYAMClHZ+EJTLLS4A0eQJou
TCKkEA3MMgknqf50rm9W8FmuQoPRJ9atuGrqPotnf5Hieis0iTXP4uXPOuiuXGVqdEId1HiPvVd7
EciGv8Y7g45WmIlAem9/8w8DgJVvtCI02FZRT61DxLK7O2A3fcJTm79FsdSaS3ttG7/KIuPXJH7V
5vO5wVYKGqSnnQx6aC529O5QB2ikos/NCCaKjCuztsV2Q+whog3fM5fUncchqk3U6+IAl5/bxpnn
vhP+I/+UCHJ3ZvaiHZhTTy8kOAHL6GAiFyUQiDrv4JlRWDOkjT0pgsxQgQO157fdGEldVWmIzq4a
sK52pnsfWbjJHyj0th2GqJhOqVH0iZ0XVHAKeFowLOHRKeBJYDjYg1JIAJugJIA7GNbz/R3U1NXd
Dp1+hBbXvTEJeWAdymvzFp4DJUA4drNjueJX5yCF5DZlEhWgZWkmM3QoHtTU86Hj+TVhUhR2fR91
xnPy0lw96jdNrPPE8B0zT+z7/JGcF1HzTR+E9AgPdVVELjwHyfTkXwlCBlJRIjsd1tVSRktKvPQU
1NHgjrSKtCm3PQKIFKtViFd+3IdlGvf4aZSPM6HKheQqo7ial/1drAG/EKrOvXc07gPqp4nJPsTR
UBWqcaQoA4zcrhfQrtWbp4AddpZDynyTxqaRmlGY+gQmOMfn8/J8Ga44ECfitKDulpIKjUX8ivSp
SdMXr4QedFJOgtrGQju5msMv0jXjjV2Jz+p7aaW2OyHk9InQPDQd+olD7Q6iaj+0u+xYU3lAK8+h
Hpeg++ID71ZaN0SSx8p79v5vWpVZ9MYJmXUVv6pBy05MzxGca5UgzoV9QEF4/ccDDNkGEcUcY4iW
/CMh98rq8dcu8feOnnZ++AvFatoLAGhlgDPprm2rB8MR2erthtMNpHGI6v8Zk5/Plbi+aeSI3O9n
7ldJDgi/xRamcQ/GRqWHYRnw0in0Vw84P2Pk7UGEv/gVm2G3KRpsvrQQ4CxWkeSRHXYttUX1ftE8
0TqDxkub54kS+qe5ZMEqYp9wPRkPg87S/QrYH+Pn2cXJpg2kJc6seI1xaJFSSLZfpUL+KBVLBReQ
O8m5lqKtZ0mwIb8N5sz3AT3IgVyIdjMn3gZVEjBSSYXTTZ8/BuaeScWkX6ZsKIQD+tcsiOLZ48ml
Xhm2GiVA2iso4fPM7bwrOEZLhERD7pJGRLptZVqmR8qoHZ6uuEk9kfrlh7shgdaD7ESfslfjT+M/
epFf9qsQ+PjcxOP3yVsGSlk1H+Wzb5DPmBbNocT4Mv83eicozU8jbl+aEMU1vPsYdUI0zjknSRWf
BSHqUk/UmKMQkXNiTdVCdQdGdkXgt4Dw7iQC2bltYPLbs5pNyD6w1GMOJUF3ZjpU6EYxsUHMPCaV
Kwe3bPTzr4mVcIfTmj/tNYYU89+HD6XaF0pPicNZ/Yp3jUB7TgGlUG6CsPJbyBepLBEKixoWzTOK
KrlUe5rUDCaPnF+/4nJqhc7qM7a+kK+JixMOKeh7WNDqUA6J7s64PZltcBR/2NKoZcEPkZoqrLx1
YEomxBM/IBk0poyQZIw60jJkkgaK8xHslK0JMVksntlxUdkNXNLvAMVIGZPox2/3QOo18YvhdeJj
2lXOThC0RJ7jW+9WKNYSr6nG+dDJ++sK4g3JTVJTcV/qraO0PWoUy8t7C3TPLa2hxs9O+D0flUFV
6oPe3mXQIn+P7EZCk1bYASFGNz/0ODkj55iMR71Fuegx35fRTBpwQkpsM8z5h9F0oDFblhMg2gFL
KI5OKeXqDV7PBSawAjcv4NUV87dtFoRuz4xWbepP6WKx1/H2aonzSdWBHChjTz6IrLZP7zLrTu2o
3OnL7ORDexMp1VBBOSmoT+vPWCkz3av/aPM1x5g1791QNgx+ILuX+8WOQ6h9AwUpuon07ti6QrLk
j8PTbaxDobgJ4R2tIHK8QS4FwqKLu01t9atrSe2ndADB8q6yfPPOW9dP1M8EMnJERwZE/QffW5YL
pVk+ZEtCuAMiDGYbBAuS9etEw/OS/nZf/rVMHnOsCEVEFYce4GinK0Wwk/UDegAvt87QcpWIOtWG
yFgu+LgoBcWErzB+546BsYvN1Fv9ePq9Jz/+yLnmgOVe/uOHHJpQC5d2mEgXEapRmHFAuIEwASpS
zNn6gmoirB2gjRSnWc7aLOZFlHPZnQAWkIZ1j+pHTRLNMeh5A33oKXu6dWQyj00fraacHDkGaiSZ
xg4Ybprh0wWnNw9KPJ1K6jg9qJbfFtmMGuhCQClm4WNCE6ODImj0p4O6qjxqIphFPUGDpj8thu7m
lO5mfFy91lfHegr91SlMX/lrOgKEPfYVPVdVU/qDxomko1SLAr0Bt2sfteTqd4DuHWUDoE1QL+p/
dvX8MkV7/IPH0zk2G5XiipXagELAwAA8UoC1uroiW23I84HNdiRShAt+HKK+EKRWjC01xKpJOZav
vzXn2yBDQxbi8OrX5OaJWd2jvONiIK6iXrHUUAzuDrqLvOw7zG63XKghxW8vMg5QxPOmAZHEX5gQ
rmYAgTxYddD2AJ3cnmCvhx0JDqWojMh6wXEosAcOpJ567zXEe1HdjXIRuSWXIptDY1Bf2uDCREBV
PHguY8TBwp0tLKR1EXLRBqQWXK8HQ7CZMav8ApHZfBVVlqrdtEBdIzJMXJY6BBx5gTzQSOPTUgRk
MqUy6J9V8g8loUqXztudCAlJY/6oYEGlorAj+4EwE2deeD4ahbiQYNsR1uh/iqRZYvkdc0kTh0ie
QhoJaaMRqLvZIGzIfru6Lwz+AC2ouwWeZA31Tibjjn2SjJVB2gBle25VrDeq8ZskZdKtx9ul0XcA
+DBzaI3acAtEHF0cvJSG68A3xkw4ANpCYomTxF0HN8XW8SorH/XacKUvISegGyUUJuhLFa71CpUL
ZVj5P8biLgnnB2wzYm7oNkQdMwbKTbj9NogG23SiUfI3J1pjm5imOt6/34W2ZqZPYpSXZBWJGTDy
zrhfcoNob1RVxHZH7a9TtB3CDswhZr0/q4n7bIqTTCCjT11fTOFJjgrjLTAbZc4gto9eVcD5PYZc
3D8UTxLXOlfk2LSAKS4q6mTEyLgKIa0aAE+7N4sRL3ajZh/eFB3uAMdV3BIvoloulX4sw+ti3wp4
ZHYrXAf6iIc8vOP55KePG64eZwffQyPacOLs+4myQeueGdFjQ0N3JVhAKRAzkPYHtk5t6mN/6yiO
BofpnwPX7/x9r+nvCfjl7yx2LV/pgwEMolgoWf8dKxAqdnsA2HDHpIW0x+vJWq1T19oyaSuF7g2a
0MtXxZh2KFafMxwMOpZ6/lwiehTn6DBLBTBfL/Bgwefwvnl9RqhOWZOcVwLktezvl/9uqdDldoAp
B312rZ+dUJjrm1mM26uQvYhH2tyCVOBC8fbV/eohWUjILqVltimzZvn3b6cLIoa/vpV5qsAjjyM5
ad5LlBTb59+HM2iK+SblSy47jYvour9ob/+HXkY3CIN7XYIm48mOnaMJFRCQSppirMtyY0/eR1JF
f1cecijrgICws4w7jOKQDxf/YUGEjGgmvZ9scIWyf5RIK33pl5nbnJrikqk+5r6Fy0v7hF7s/Im9
+MP7mt30BuiuohM/czCaGG41+3tD23KaBv9bdnuobhgJw7AdMRYl5x/CK882LkM/BIeTQ7snENZS
xKkpIBV0nXGj4YSEkJxFzhheOL8p2HW9+C5CRLNVlV4XMbl3wcnjtIf0Y8gWDh5QtJE6Th5myNG+
Yd5XmmNze+YIVI/UxbJR5S4qe97UvPzS94O6fNa3JDmMA+pHmvdQMFRPYYQc+kS0d8Cqqu7W9/IH
zrGzPIa/SR16aRk1U8YhpygtbLuQVLJFpwGxffXuiAoDejCy/xiYh5wONeL8DnZ/7QfhmcqHiP9Y
hKBWdRd9mACCHKMN1gp0Oti6wE2G/FOuq+zg/P0oTDqzzLlX8BON3a38A/AUgtwX+HS/jOLp1Jk4
S+29ubz3nGnJDmQLYGdXrTakU+6ku6SfMuph3IA5zUQh9mgdwT6csz47iaOh4Y05pvodPL2sdukd
xVBiW9YOBUHE+mAtvg564G0fa5nhsvamOHERE6wvCwVn2xSxfSo74zRjNbyhiJ9Ma+WGyf4t4dJu
dQFck++o1lK48ikMpeSbwDY1BNw7BnWfTSEernrQ7DzQgAzL833MS5+WE95dEXAyl9e5kF28ZjEH
9Q+Ok83wck98G6kTesL+cduXQ0ooxfa+YemPHh0GjAjsE/J1JtjggDmqdma26BAoyS9s5CEiFRK8
I/gdQsS8TMqQHhq+2AWQ5X5FbyTJAIJvucVmzLGl7pKl+SaETZN5qBMKLbJIpHyrnBKmjXcA1Ls3
xLCAwlGLGhyXRzxhNJk82pUvohrn41eMWcI5ry19VavDia7+m+Swrwu/zoLLgoScjnLsACZ6VoPo
iSfG89ejnl8uAirUeAr5b0/POqUCwUDKcpyoNwnCUT90DZiIP228ssTGUEkZqvDzZ6l/Mm3+W9mh
Qr4ssBs4CuUAx7uqCOQduOKZLIAgDfG2O8KE5BrNeLFxVMQvwpR4/i8K88GeayBdgRBfM+NWdVfg
7kyWZTe8G/4PI8kNrRxOXbUnWH7EXU7aK5BsO45nKe/Bq8NYDHUpr5E1a8Sx23us9zHqeWRY+1XX
CbhtbkE6lQSxD5wL8Ewl32f9gRCXJk8gv5NeW64W4+8G4tYVZDY87tO+ArpS2mv/mEDljivuf8k8
aynfDH1GmjzVBW4e8CpdMmYoAOPO4wU7dH9je4sESuybUukMWzv7AuTfI2KbwFuNb+mnnzXsQ5Uz
M6N1vXR8sACUfjPcsQng1nsozPsPEFTeQHB57YgBYb18b7dkhazX7PwHAl+0sqr0+fSsbf1qo1bp
OwmbErpR+d+PCwA48VRE0i9q9jrheuw6bjc1v0YEQshNY7IObOg8bNX7B+xRf/65d13x/K2RA/vA
TZFlb2LmWAr/8m5DbK6iGVufGQ2UIkqzTX+K028C2ErD3+gIvHsu1ZtDKVQH5alXUFnDwCCWT9FU
Zmt0CYNpGKiHHeTxxldr4dZD+MuVXgn8IiwTR1bvrMBoyour9dnBpzmMag/u5nKVViBrp22iHEpe
rosWLp6xYuyYFuTZOW+Q9pZtgDo+4Qq/9MV1UqqpO77A8irD19ORvgD+9Tlb+tUYEluD3c8P5PyH
epcek0rnU1HNU5kKzwZpUOXNjQaw8oHWRcOiJnzNvPCLYBR/h9GO8Gu0Jp1uxmMlx09BWCaEfykk
bm5nRhWjMSOT7fZFyKDpDx2F3B4oEs2xb2TVZwQ+2w/YCzZuunB6uPcG+v0SV225q15+v+gxPL7A
7SJ85hzMHYYb9xXZRhRdM77aeWwmpSnyKKw4lj1knUzqpXi8yskeMOLOFHiwrEohBSKM8qIazyqx
seyO5Y932fSEuG2tAGjSfkrgBpKuVhonYXgLweRKwf8ANcSUc2cuWst5xkUaS7KEjSfvlx4+5W2w
wLVBbnq+rKBzRMRi8udhYJnKouFtK1qktSPoNcGrkgfmP9QCuA8sZv/x2WhhdiSOGQkzWQtYQyJX
6dF1dFzu/WRT7HlxyZkjeS+dXFgSiSAGYHxK6KYsKrXvm+7ZFskhakkB0uxV/U2q7dBxGAMp21+R
TBf5kCTdZ1WsRdbytUMOzb0sAxLiK25go3mjmCDayIJaiOLekuZWNCxjrxopJ5u5S0vFjCSjzSBx
fQqlLdCG5pRD+1EpdULzz1d6xwE4/x13c2vqCb3KbyzID3nIFdi2/Z8CXGaHBPXfLYu7ZYmsXkJC
dCsdDvkBTHJakDyi+W2NJLLq8MuLvQOvaFdCeuI76xM3VF7xWIqV/S+4ru5Z93Eq4Z8thUxtjqOG
cxmaNinQsJrIqMtoBaNBiMB4V+C/qFdPZPJ0YWSUzaoDX335fnP4PIDXeiitCdz80//Uu+c8qoxB
RE5IlvYSv9gdnt9jhvqqNTtEMU1KRk4gEm1A1rY8GwjGq3Gw1kZYMLgH9IcQU20wcPAP3GY1Qd+V
j28VQAnb5lxtD+j/UJsrC280zwpqYgKL7fAQ/Ae1By8RSpkdBkJBykKG0k05CnyhnL5BwbCHR+Y4
qrPnnyzCJhlgK4Gsw0GZIIF+0GU1df6WYcCV50T1Y17Y6qtvqPbIf9w07kJvCyGnB5LIViwCTQUz
7t0K/a+a6oP9WIvAYRTJ5L1MU32i7CI1puUsk8PoN/Iwnej0GOt0PQFID0zRM+2MZEx+gq1jfA5c
hoRABvXkMdTc/aa+N/ewf4x6f4VBB/oMfpUIOY/wmdp88uBeqf2+2ZaBox8mG76ZATLI2Oi6/oVm
QX5weLfLdmn4zr0Zxu0Xs7UxclV4HPoN4vP5lAswPHR3wc6+AwLrUphfxjUudZFJWN2UY7tVzikn
CElc32FCZmWHl5dPY6VIs+eXYX7TB8lQwIf/NDvXvnZI966zDhJRpA0B7orD0NjF/XBz7BPICj1w
xYvvtE70cLKpSswRXqhAAzfkdtcgtRXNRZy8h7lmth+ArBXdduc7zL026sEl2T3yIjpKHonwRLfm
feM++gLeAkR5WJ2GzAS1uF6XjMVqBXvGWSQUR48Wa4DSfgFwi4EPkIC7lcnFLpEzQTouCqFtcH9P
dRDnzFgaqw7S3r+BO+geMoOWmCvZu6O4XToBE1/1AYZytkYAnv1I5y1dBjNGg55G1SbpYfToogH4
TowbwBwu1p6CUe4E/6Kk6BjhWNT66gU5JZ9J0iDrnFoYs7Oi93rQBCzNBwNg6QsSWhWgrVFBoLqg
KDX6wQ+CeL51sWzez3Mjl85vMMB9GE0CZ+t7JqdLz0MndegXogF05WeG22XL9jK1QGUKK2g5Dqi/
siJiixquKBv3pbsAA/FzWMtDqBlbk00U+X8BqvlkCPshFuOyDiZCXKijZDBO80H3W7w3o1X2Fbxi
nvLU2fsaza0LG9/Po51xI69e6+amwby8UsG73rjh7RaLx94RNY+2seI/4xhb0Vld9VkmByOWy0Qv
R4frtEM4gsN8f3xzxCvyNFKVPjVG/aF7ExGOmolEKyHrMGSvedK+vpg5im/vq6TWQ2p3wbW9uC8H
AbdM0D+6CQgr8uMxsxbbHcorQXip6UyEf5zHT7VEMoS6pBMWEhD7iDV2oWc8Ssu5lWB/O/BEytSw
EJGSSjV1FOAUcKcuDyxKnUhDKABLfG8bKkBxML6IiWhRBAYAH4PxzLN/4rxqCSdEA67itHGxwhEZ
W0WHjB6McT85QRWptXlU4ppek9k/GLc6xW4ItwYyFM6v9l7Vlt/8pfNjA2ZioQNug09PlRmhJ2mQ
VloeDZFe17k1OJkTbC4PIIbuXmoLSt/dva8zj+UsUnv2kgjZ99TRUFG+qHViCNykoxyGgfEqp0sm
uaBE2nHbnCL6+FOk7jXHB6CdCQ+tpKNzQVsS4vi6J9wu6IL2c4ByKhxraLOp78hUF2u+q8HXYf+F
1vI0LrfqYyDDXAwrvnhb/P0Q8Y9m9wZRsbJGU21jQX3iLQ4EcIoLa2tSnY7g7eWPd4MMNR3bML/F
ozngeeoPh20bQZzLlHxW0LFeNrrE26/RP+IOg932tr1F/N81SJMCBjE9M2En92hfQ0k2fOJF8pWj
MZMCcISRM+CIcz1ZUxdBMcLhmcFJiMSr5pDnDGdV1h5o+S5oppZEnXZhS241+uYrGDJ7SMB/Efd5
nnRw3g1PTbhma8cQgU1R866Rp9I3PyylkUWDO7CKAzJqkV42QATC4c6T3bq642W79LZQ/HTLYvBD
BBMvm6ICEH8Cv1BNzpLeGvWb/knIH4R80e7tCK7WXv/h+A6iS8GDbHljmnPFeOLukwQ+upQTS3lo
l9vNgW7VLN4dFz5UNbyGqGISOqYS2aK9yUBJV3lPw/VhaACEIr9fVxhrvb00uSlPKYHsjJGj6yUn
rPozXDZJk0X5QQXfAbX6X0ailgBzqqU+KYCH+kCZqaPN2NGAuYaphToikUbDuGUMqmsE9aVl4ZmD
GJ93nHs9tuohMmN9JV+jFr2K+2sd6MMAkpKnDG/mWnUdYRJqmhafCInc6GzyiEkM8mShrkZRqbl8
e+UlogmWUW4tldp29L2XI8LmvANqV7oslklMnnpQaTavFf8jmMuyJ6ZMpxgz/iFv2zF4loERSd/U
I7nfFT+kOorHxPK9NlorZOlSHVP1Fi6K+l34CeVs759MVtD228EyWpQ7+rbzPJP0aUuMCFEu3e0G
OvUM6EHsqhmaz+d4/yU2gT9WtnmZ23bmUxxyyGvbKA0mTX/IO+5wl+z67MoxoGZpgj9VU5sOE/X5
2fL+7y5HY9sj057uQGLjpadVs7/3VrFwQpZPxF3D/+mwRfp+07Ktz79UlFPda83wEuXze/85Hi8C
eI9QQOHNuaCrGoOjhCsXJUwd3m1THoATVxq0/pRUxarODipfBOzGMIh5M0/oxltE7Mbd/wGLnSdL
DyOpqIJdllw/RtkQz0qq7MSp3O1uxxPy7lM2kZapTHuuxPcIiHnREWT9MlTbAes4tSX/aWIBGF93
RKtUS6Q4FKNTO1cQMaWI+MjReXeYoiIFEFQjA39KrMz5gfpel4OgH5Dbgrwgnz31HgizPJsi50GB
PShZXHxzIqTcDxnJtFXX3PCsohkDNoRiDwyNR8qbjy4HMQDPzpgWBgasuGomzCC2t0NWrzc7+Pn3
3EX1w9jxhLOrCyyoR04ndWT39VzA5nhtb47lbmDZd3R2gVHHuhy/Q2A6BmCuuAl9+ZXzMhuV9VNv
/Q81X7knxfMcchbelhhhAIR0isqyz1ANHAa4ZlFG3oGYN9mZSPJRjWPekCTTB72aXVnEVWRcxKKJ
of665p9tVVNa13SboBYXwS6SA4ba6NmPcZ/zmBNfuYTwYaxeOBc9aSq4TCti2EzLPTekfLyNKwWf
1T/l3xlceS4hBN8EteGz4OjIMwV0zdOelPKs9TeAzqQoj1nqTUno8PxxGtrdwhXbC5I2ookl5f27
o8TgzkduIfPd3y7kDz7SyZC1SxDDYTzcnCqAvvKXIKoz+DG6XWITrUyDKFvp/Tq2RQtKebCMsq+D
vOwUCsw6aD7QadNnJG5cSR8b8x6PF2Y2ZnKbj+5tVJ2noZ3obWKz2vW3gEYBsbklX8Au4ahY8Wy7
6ILVsSvCv42dAKA7gpK4DlKAc8g+FeU7SuMDHmHNY0lHwcBv9GCvn4/mSViwbe+8+/+0ID+QqQML
Oads1qErHsLMmYK5vMZ+UgESbpYbazo1N5o4Lq4XHScbJwKL1pqeFZCeX7iv0pPMR7kkSj7AphvX
OxVKBYcgZ5sPb1kWqiaFu4oWif7Iyy4tYTBr5jmD1OEOvjPMARe3rIoCjZ/gxZVDvReVb2YqRd4s
JYaNkcGmbrtT8l3UCHTxFkc6dfLOcZOcf6ohW9KcalN/bvKwtYJcSOUjyrQKNecPJz1P6wPb0LTy
vwSXEDotxN1mCqolCwBS+erp8Dv/9B5oCEEUGvRAF+fH6Yaeg5h4Dzu9ZqgDYGm1/M9QlYGdqoD0
fLbEjMuQ4bB8cFdbj4CWeGA1jha3nbyhCtOD1AExjE6SjMs/QYM+AvuJB3mN/OD6hfPOTrSTffxA
XevE1WFF5IocyNhQihWPDJyYmh0y91/h1f5UFYvYjCnTebrpDWU2okopVwe+0IyuRM+ol2diEkTJ
uk7rNqJdfSIllI2ZDufrL3617WDj6ds16d0ZYYjvBZ1lrbetfWiU9S02nNfplA4zUCNyOpOuVPfG
BrX1dSyPAgW79Rclx9n+IsIcs8GH8p2LaIPzHGX/QVENP/3IWETj2OYtJ7avC889+FhM4rilJTKo
9MrL6QWS3cMBPdjDelAJRteE9kezSF496CDmdrd3d0B7bEY8GOES5Df+LwETr7pi+sANts8rqS6r
qv1M8Zzf7a3Oo8nFYn+20FWvocxhRWO5+0nwEMmeLHKMxmebqPizy7kh0O2oRnNZMdiAFc2azyY0
an76QE+jU1h3hHzyKsE21wk0RudIcI2DBE1c1C9/ClEKgixZv/28ajMBD072UxtRYIXdXKyxgDum
sJncghjR5Pu2LmlfmY9Ujg4ij/JgkGBmLiR2s1G8hmavK5WraTCLEP2xiMQUsDXDcrDBL7swBKE5
NTUVOEWVpBAVmQqkubnkkErwNuBbHsK5AgGslk9+l+X/z5pB5CVsXmnlhG3PWeYZFFsV+FbFF3vw
cBVr5BlJR356IUYXd8cj/KqmXBo3vZ8AEVzibwsn+n6m3lgxAD2/M50R+xDujt4V0u6cKRvShQW6
E4MBmP3hwExjnwgEfNOTO9SBFYwQb1T7sDfnrXORt4i7rtlTCa+3mNdpd5FYe4k9ZEjf+/dQyVRL
n9c+S+tVZBeYjIsO4YENe4guepQjpywqfVvWwmBIc85pYFpHh9a2ijzBO3koCMNE6FQI3NYqjd/W
cNqSCbQcfpjnfhzUV/251WDY3IxR14k4tiW4+eXeSUda6LLciMRZM96TwuHVdbytEyFqPmFGfzYh
lBZTalbDrZYjZCYskx7zOWRnib8jRZ2MXqo1IQ5Q6rk0TFUHKL6Fgv9MZSkAzb7P78t7u3zwd96m
SMWkLrV4feX2VJXCxqpqHXQ5SohgSBYZkEgz6oAPppwvlWtGw4Knsjev8wOx93IcCh4gC78XSbXv
E8O2XzaCbjfrDBmB8N373zbgpOx5QwQ/FY7N3X07d8ONoyg7k7N4Zx1Kahf6+JRchlmCvKEltir/
RH3SGmnV79+HCa+OG+gUL7LkD6E3YbtJtwWgy1zpkpIg3bQG6q9gDcw2AQUE3u41AcKyRRaGInyf
xuegWH29uTCrh7cKeDTXB6KoTjdJVh2aRoLrXFoE+u8YvMoxpwWDRDQkWzuGaS9FDaqXglrRxFQI
JSXkQBvwtXQOevsir8Cx5uhBLMsBTbz/0RgaaMq/pPNAufhWkj4+0sSlZxE3PmsgizAQh3mW/aNO
oKOVdJ4hKdK4cI0rUm+WZlc0ETy1l/0r30SJidcBG1hhH0kwtaRTdrxPAbZPKU8YAk30rvcsZUa9
eSNPJQIeBVtRETF7rtUNGvT900sEwoymxvpOYU5eHg9joh9RrDQqzO1OwNFqxZOOIebTZ+3xH9lo
KRDr8pUQi1GEEHp8Uk0mDVIOdWw1Y/sjxjoDuBdw7eF58XaBFM3wtBTJnBW7OWHdQN3Hh4fTrEOv
/70eeXk0WXhx/PS7ZU6vSv28cS/EaGu3dd+O95DGWL+5k19zjNs4OTLhPkIozpHRBhIo5mjWF/rq
/a/iQFPPNdp4M8BYa0Z0OIjpUiw4qbpgXwYHZemk8RZHqNqCek9aHXfd6GcXhmoa1Z5tCpp+h/lh
ndimWAEWWHDL302nWo254oyBqnUE43mm+aMe+OyCTt9nVEvsH2WmLaK4M2GiH/ToCm7ku4/aTaM/
qrCMBGbH3tO8TkCcmnfXc8puMM2zx/o/shZOT5uDuvZ00NWJVDsI0gHq6irjAgeEvF+1sLa0P0z8
eRwX/Pr2bXnnXC63KGqeyjpARbQi0tAIpX8oRS1azgh7DAy3b4Y6EwiSZd+K08XCTqxt+tv8SN8a
uZ2QKvJ0eaWG/4gsAgqIR3uZCct4NhH8DvHIycLsjM7fGLEVYibKYCSTWDnBA/wwGKsFJ7JhmWOj
l5g4wcoMWa1e1H2YsOirVxaJA0aFi2ItPGhTq5Wm5k/ICpu6oEu/j7c/nxtA4EWIKv786uh5vYQe
hUCTgN+IWwEJV1+dOk0qFnHc5/R4ceOCQo33l56dM9reNF5GinZIjGN4nwcvhZqUEVdnTqKV8cqh
00SucFOQ7kduW2TTxCRxF/tg7/1WokDlgQI6Ryf/DXrSWtKWTwgszeS5Bf/7yKTlNyC0W8FA7FX2
yE4EdiaobVAI40xAGVgbvO1yoDBhc9pNIO29tw9q7zL/C1IG9sNfbSbyoLMi1po5YQmxsojWvFu3
gprQIK4or78cpzs+uYuxa4B/vhNKUn6pQVKVQZsyGoGHwRSn5lPK9NtTyHLoGX858mlk98WJx3em
Ue6GR/EHujcH80JaZeqolwmJ7iCprJ4SUEKAr33grpWF8n3dVqbI7gblxSbrDqyZXUGO7TF+3YrD
IbRJKHNyMyEBSPErpiDVVlXqb1z9QVypLhAWGzvgiv8ZBSTOI0IaX7xD4rDMuOm+NsYa804xdWr8
r/2Z/w6Tew8NPsrzzOHtRhPAe+xVxHHT1FCAmbG8oYmbOfUxThFySlUH6csC05a3pLKs+IuYX9dd
ysaH3iGrb0n4eDnwTyHEUhXa0w/rsD0pVphudn5DHWJh1Ft9/fCOHz/sNSZCu/Haomm8AEN/PEy2
xJjsULPoUVsQKURJwosXA3YwDOV0GNknyeyOzwwynOxYFS83WFktHtRARsw5RGkZ0eXSKoGVsdkr
PpLZRjbvH2p80PJo342TrDlpvfRS5Hheh89sQNZhO7eHN0oGZl3k/Lnc8xrcFqign3ulVMcBuNvN
GKNFbNh5nBY5HqllaemfBw1QEW8t6QqvIHgso5C/3N7Ez+Xf5sx4ZoUO+TNTrC+Uzt9JVOQ2sTVZ
nacyxfKuLx4NLsr2NVDbP5Z6V4vaOXwyf3tS/oj7h9DV7MDRUBi3dhwVsihp5ZF0ZfEWnVM7tbnW
PVITHZsO53ywX/8FI/Mk6O0uUFtOsPExbu2hHzp9JbjMAwufp8JSzRdiug2x+uc55S+IDRhcO2D7
FMsE38OrFMlK7CFRAh8Z1cbw/bTObvOxG3195HVK0O/DNhtf30DHWYVBUcM9uJFqiFlXDdBMtkFP
hwodiNISerfHJXfhyZAVPPJrZl5yaIL01yOC8Q/c6wJl9TmuIJUSsR0Iu0NJ/1OqThBWkK9LJzj1
R1mXDZXkpB9EuxphoPEYcMb1yvOT/r62Yj8i+O5QkMRlJvSrLQza6N8VLEhdjI09TUPwdswznF6W
Cf4eCmaNVL/z8InJAo6mqikyJeok5WDDohKKBgLPWuQsCIG8M3j9VcqlpU7zQPRVAFfv6i457vc8
4EMdfnmmTQKA87bXbqEwjtO4Jq8qPiEvGBJXSA+y0v6xQ39dmXNXolDWwZ0gbTZOk3pSKmzSrwhw
TvG4lrZyi0sbL2SS0A7vSBxpS4sRf64f+5OGiHtMT4GY+sQZfu7t2WN4cQbCbX3MpuIgUw3pZRAX
KvUvjO1Mj99/+070cC3TF4WizF6a24Anc7NPSV5nOou++w7q9fMIokam6XUuPVbW3IE+5YXiJgiw
+1aSTmbG5hkDbwpVr5356W4Yd/F9Oesg9b/6LCFyY1LJIUCYb3FFSgJfvKbBpVGGZM32XLe3BlxQ
ts6h37avxxkP85VZ3WmBlDkYj6X9JBQOEZznvo+NLte5iuNuytPkwF0UMSKATWJLqiT38g8UaVd3
bmNJe6t8KnepOm0QqVYaKVERxLy0Vms6nyKM8mNnxZ4H62ZxKhvHlu/eZ1wXYa4CXlCRfvM6RNsX
N50X4BqrXXS6VsmS2QkI/GYMSMRrBU2l0b/LgsaXHjRZ/PbL+wnJQTbVirFJBzkJa8MUJx4zBCO+
nUF/yRKyCLZWVr9IKDokFr+rRTy8F3FgQXmGOUXVZViA11kI/hWp4Qhi8QtVjkacgn73Z6CNpNWd
xi3KL9sQuifeJOBJAH5xVLMlQIiqDdJ/6/fRxsmwwGg7m6k9batqMdhcGuKfTvcMifOqla1AIoNs
yPK+I706iCiAWfCP5K0fzc462nMxqDB/Y/Yznl6yYKOWGkTiswgyRAUYjMubahAxsJjSvcwxnF7K
s4c1rkI/FhzdBuF7g5paQWYaloe6KSlr65jE2QcIRC0pCfzZOTtTl5e7J0biHpVcibBEzBTqUrd1
CRePtWPDTehhJ0GzCeFNTzlgMN8K5f/TnTtNxE07tkWveZd+4c8GzrH7/8OEEU5oFSbeJTRsphxK
InPCGLLyNG8Ujt4a15E7Il0kFLM5xrh+HIalxTt2SKYbKYvZOFEBexim5H1pRfr5gc8HBajQnz3S
rO0DJh7tfytxpbuXGU5Cc77pdb7VmLl+EdI3rySOeQr6GEgOqqK7yInxsDAqsU90ciV7N9I8EzEA
3bTWOJdiQt7P1cvbcye56x/EDVxcWWGiYJM5Ja/MNJemGX/wTT24X6SHUUU0dkh7tBXIoaPDKdYk
SotyI4YvgHTOzW2Y6PcWE1fYUqB2iDQQiXTSdcJiGQjm0/YwJn8xAkjb8KlGTlFgE2u5BK6g0NT2
+vI+4sMJeC+Cxies+oFzPmR366MfdOAJB3Yi9oEqVEFAJKI8pk8ZRKAVgQy+c4o/acMD22+2+X0s
eYou7IDKTzmal8DZvsztiwUwVQwDmxIzvDXrzlWh2OHy3/ZZIylVyasxs1EQS2SDPKEVDHy5RpOk
OKQ2uQEh+7cCOD5xPXdRbJbBncMCupavI0UhwBiO91+4JR6iT6yQCsm7fLFlAvccSiG0qkabtrIv
6lffiU4w9LumeCaZlDb3vf1iU8TXKep0gq6v/vcYtgukVMy17zfvSgr54ThvDee9iRZXfyKWTYUG
0DMvqdZzRDDBiEQ9Lw7kjqSgkVSbfsLVN7KAZ1uu64PTjiF0R/8M3cvoz/HYOe4kbsHVMQTgNTBR
FclL3HcbRpJJ4gZXkLYquCf+jSj2BSGLXMpygiDS9bPoTo3eRGpDEMREUh8egwOWgd7t+JgtEpcD
d92wH+J83/YLRHq+Xz3eF2wSU/LmSrZLP0axc5b1/T8WR7s9tAseEdFWRJy6LQXYAgmlcCoEYKvW
7PyU8gT3avhDHujHfy2toDz4FwaFKpdXYiqw8uTfhDz5b/9ct0YpLSBy/lWGns7Gsq3eZrw4xk/z
oDNjkLmKUaBofGW8KZdX8sIDOMaHJAXhnDq150ynfJ3fSVXr9/fZ7fbJVtotHrULvCV+Hbfw5bVN
owSgccdh57vl46M4daG/mlBSco2yqLCvVFQVUImYnVBhT9ulda8mhDlqhUMNp5U12mREExu+cU4K
2hOb6KWPAsOezTGCZYpTdSxVau1+GwzLNZI9QyyxkdHT5TlXK8MWybK7n7PlPyb9scXExujpQEGr
5mpc6sGkClpov8sx4gGv/jOieV/QxfbXoQDH/7kb209Nmw8xJ3yVz/KLR6qRiUQJfs17YyBMOyRY
SM5Ion93+dqwA0CsZdDRQk9l6OTA/tYRhmBhrb0MCVamUmPfqJbF64AZ7HRU77yON+IT+aR1e0xK
WQ0EFquj+yrvbT0WjE9GchOojJz44UAlCcJEGgSRprZERIKcE1ITGFxRx+CCB3x7NKe4SftuYbZI
7dMjEfB/+n0C97L8AaIAS2s/aOPFe/V7KGwSk8tNi54Zqo1pQ0lAO/fCue9uWpH8N7cdBIP9LGoI
wwq7Zz9m/AXo6eBr9KZNbjjcw/azEcFqkqlUATd8yfPe9XaPnYXzdrBe4OW+EZ7f1l8rmp/WYVE6
r1F3c62agF1lbAjpJixrT6EgpzdBiIVAlUFrqJ/5VvYWrlbJm15G61WsrNrFdLLFhDxqIp442guR
pVC0wgjiHptey/F4IJS//PO3hj71m93NmINGKalQMhCuJUVWtRrF8O1hGQecGUqXsMDaBOpq3Bvu
tKVwiL0toJYF9HWxgWTfD+KN1h3PEFk1qG4jGBYrojKguSTS0Af/Pf2JtrVSm4M6qqi3qiVmiwvt
KjNEVApfff7JwD2gONfybL1N25k87We1y0qwkOOxsNWA/k4lo0XbGG2AJkfcRYgC9aeK1KiLbxWh
uQXTID7sJb9vV+f3GmC3c89yVXb4hhNpNWFgumPGRss4qZ0fOSsio60xYyha3YJEKpCkgx0XLU2o
IK5+suztI5I/Bt4ohKRolsLCa6f4y/uLeEmRV60H8g8kAeiUmvaeXUfg4mdIsesRrytxTe02fi8b
jgtWGd7Q9hB+ENM1BlgLL7/BYmcZYt0hNzDDkT2u6GN/SvV/bo/K1qCKy/OVU2s78+JJ8NnowZLJ
mvYyFAU+vd9peLJ7mh2sY3rcxvtqmJDR6/SUf+OVDAJ3W8KQ/o3dX78QYJ/0CrcX+EBaoiT22K71
b7ud8MnueJcXJl0n4VIDlclrx7qjlJFT8jbiYZKFPr5cwLuPkk5E5FHC45IUvpZBFCYYNuiwMlih
S3gcjJtN7XIAQkvGq5Gel2Wy7g0HGDoCHeaPqXkv7sypinkC7CrUm+AHQPvZY0gGuxMrPHq71jn0
55AueRfSUAGoMxUJvf1TA7rh9dOSHTgNXrjQAtk6KX84/vyODUVg9KyZloxmPW4obqXKsgcelqiq
VcA04jhhpXiKpvXLCB136IPp2hrs/EqqxUpJsjLnajmNavzreAJbkFTvzym8HVrtW4dthh5qAsVD
VtGFja0e80KCePkenJ3G9qFxjWMXfPkcMIDp1DEWW3nIBUo2UMVXQVLZUMZjfXu+K7kwx8tbJpkq
76l8BEV9aFSybMzQ96zoEcgMlqyaWLJuj9ad3sneCZu29tJFdKlv5SF2TvwVuk/5JEjmw6qss5P7
VX5FvXkrELOs7lqeq87wGYlAmmIDwOr5+Nym4DkusH+PGhH/N37abLcwCY9gMYoB6772vGgZ66Dq
wV1hJtpfvUEpS/MdmhcwoLpgEFjsyVhZU5avUd+NVznP30utxUuSzhuKr9Vvi9F0T/6aBlJMkFxz
24LsRPnhre3oR2L4kQuzNcEtbr/Ky6c/TfPqZTw1AVBe7Hl6enhIPobAdnbotrtRW6RGTk2CLVxW
2kt7G+x06sR/GwtkGAEZ20gIBCqXIDObWq47V1iKm8wyC9haALtXweoj0t1Nc9KP7mDRaf1n9OVF
x0Fp8K8CpP0kxm08Gzx+qBoFH3fQomTATBntB5f167OKVs9jTlWtNz1UE4nNBgdo/7L//l0zAEn1
ZzKdz6EB7A7PAVa75KZWJTpQ7ZUlpp6dUcJ9tXe8HSAX7e0u1I+sh1jJRbU+W5Wi3rxkZyHPU0Qd
4tCQV5CdDR5LjvNKsXQLOR1fNZrIyQ6fhI/ciM39f4EuNE+EnpWo3b3Mntxgmok1eYlmVaDV+ioF
h8yxH/trOrbFi+Gj95Wadv6hcDwgXcAon3Lbv4SgV0UvSm3dVfCt2HPNI9Rkms+se5knxz8PhTN4
FnRkMT/6KPB1VgF0nDqNF7doBln+2BNY0oJC/n6apXKK+UqewtJLInGs3LYv8DLIpbpxl/Naq1wp
ELbfLm7X0+DWeXqWOvps25BSRR2FFA8CHjieLgbkQM3eV4S/pD1xiJH00dUVM6B4ZKs+5LnEtg9f
HPZUjt/PUvdQescZmPo2sTbBs3doZzRr/M8WchjxpPohMzUGNKOnyQb873Uk6xd/EENgEQGXCaGO
U1ETvbfi9/DlsSQKYDjKhBLwS4og2RftpcDwTk6LmlZ7mYNtCXOf4wNfQi5MLLEXekj0OUX6AKe4
D11XrcfbgvCJ53Zst1pXt8jk6WN8x/tpSTmS1YqNntOeuGOTC/+VGEFAtUL0BASMdROup2gMZJkf
caFIvsY17B+Z9OZ/6Xq62V4cgwhSoSdxN/5ieDV/ZlICuFkHl8ejFy0CeYO8au/qBf0V87WGGM6D
w3/CmiQAS7E0JmPppFFO08PIm+XR5xRrqGgMG+XfHoR47s0/l56Xoo7qfGlxS4KqQLlNbuXa3OfR
RkffE0pRqGfzXWWzyguLBrkSfPvyypSBFz05wbMghWfDztjoTcX1hHwyl+IlLEobBwlaS7WxdCor
bDOFsObm+isM3yUzJ8Ia/u2XwsJ7rQk1XHG6qkYjk620lbQKghaDsa8/rc1N+NGFwiEjcLNJmIZ7
/a4JQqQWLfjAZwl7UP9KwUCpVphHvf9LNfg5IM9qDG7gK201eFAafc9LV4or22zFwJ62vg+wYFNo
2lBJy/lPNEA3M807mQnw1yDh27OryT/ZFfTpp6HQcFO9g2oOaEaPyTC1obFaOdvVS2WoDgMuWALn
1IkvkyJP0ONsAXj/DI7PffW74KIyd0KmEmBdblK5fop8cOvzwlEeSxdvbKxgU94IQgNHb5rttKFB
JlMxW7MBFeMTPLq1By56ty4CXbYjfcoyEx7ORf+kOC/fc+klClD/4CY/L7D1DLvcnez9FrJghv+R
EBmNRadtH6gxXI6x6lNn2wcsLAjAe5S/X5yif8xYtna5joYydGD7VNtsTABi4+LEHGaDhjCMisT+
9C15v//m6Al16yHaMLTRdytwsr7OwKod7hVRtP4l4fpjVNDnLVjb+kIWNzBKkaxz3jdUd/23ushG
BWHKF4RibQ8dYI0jln7MrB1bLGvjklfLzwqOc25vAFrZnEIcwWdDN1EPZGgkLpi7gVpDdStS89E3
f1517Sdp9s5infFnMK8S+zYhxy6EVP2ojUPZibLuA7QDhKbWWHyWpPtSxgbbK6faODdh0KejJwQN
8tXVkGO7fwxw3py/z4oa1NzNswYma+irq2qKmCOhNeL0Lb2BkMK3LtNQ9Vmidj20w/vcyc+W+/KO
jBmAQTBsjpSKo4/vRmbXpfZXcoEn1GZ5YIah1PPP79ZyCWTQ4NM7lyDWPTrh70SGmzu4DCphQ4bR
sg5LldNKV5wk00B5UqncM3gASiqcoJlBjFXGK3x7gwDfXdsm+Na6hRR6di9plefYON4S8zF4eXaS
t4sG9VQlPPovt7tWelrQzytqnbgLz1r6ZjfVqPxDzaXIRHQYF7o5kZdLjyx78GvhpNCY01GI3LP+
cFMf84ec0btxh8bzpCqj4IWEpj4QjYEN/jMo1Ga0PMa1C8dPbyuOdiEOEnWibc/5Pbcwma6ny2PT
JnZ2uiK1JQzLYgh15MIg2wvTPbuch6ouc60hpa2fhLSIZ7i2RWcK3B2MBA2NFn8mnjqMhdkdTADB
62l16Mu+oOFzJ7ofwoBo0s+We1cmhB3acRUAJB/jOX5iK9jiIU3Op7T0/mjG5zBvfHLIlWZw/v4b
ekeH9JZQ+WkGw19wwln8BCZ/t6w7h13kY1Y9W6uS5ZFX8oA35RCkEt4plNuMTLIfkCPPpmAQILNs
GR4OjIryWrh2iCT2BUYqfpzIlUOwax0KubpJ4teH/ECGKZQ8NQa1A10zEMEeo/yb/tLXGNA4jSnZ
ww+Hmd+NWxMWRnU705diINeieLRXR8S2WOfd6Ve8HWWa6fZgsPHw3PTpGZbzoL9LlysLDj2ypZGZ
/dZZt9R/fVtXW32UzQZER8YM90v8nvhxFFgadcS0CKRiou9mtbACpNJnwWwfeuskzwpwPclc8K0M
yknXhrI5vY0oldVO1j3OfmnYnz7+JQkqGLvOv7sTerHeyCgyKFnt/3O/at1wOvZBmaZHIILrR11l
AOutL4HYubUNTvSQXYjnG2piQsLXjZpNu0O/g0IAq0TsAL4qzs7EfqwwQkQbSm13LUJF4ZIs27Qe
25mvUxqK9LbEfjrotNz5OulW5y5hMEeR4WwUye2RKIr6/3QYUBnS79hcum0foznXySb4k2acx7Ze
aU1fJ/jbbXukqg0m9NkCWOeXzh6nC9CtuM0+xLKlVOJfoP9Qb3ZLkHy3ANXaT1cbo2vSsWko4/xv
HXFIIyzUZIfHSqYAgTR8M2QzLN7avfI3FeIVc5AuGGVkfgblDLOTMVvWBFAFVxSgNMJ94QMfQFrh
Be/DXa0mzPEhpRX342ea4xPyXXlfrQrsitnX9EGPKqap6j95Ct3OyQlneishj9sJhunp8+HP1qjh
NQh0tftUJmPWioiKCWOUfIoIWxG1uAvPdUSvAodR8Qt6uN9WmLpRyU3SAjKbnOhxuSGd/5psqObF
0BXkf5JJIgYj+ZxPE6wasTOJ/bSyPTvNgPPygaLvY/HhMDCUcxZsp7mEw2/qT5t/0h8F+QO+VeW1
5HmoI90s9jY2NsQg7ocOdx5RCIl8bCNJV2ba5fCp0br+DRqO4XJ2x1iEqOO+JdDADg7FkBwAXTKm
iSbG+r6WDGJT17ro1j2RyWGAIGeKvLe4pxDbWZX16nrCT5omjkqeDW7/2a0FGymbljL/X0ov53Yp
YdSfMNhPLsrSXTuKWCWwnpFzkcEqPzS4uwohS087bnNS5V1MFBSET4oeXNbwgRdnqL7f6c87gU/n
juFwaEptsW1UZVMhz9Teb8CZhSyFmikyosdLyTbKuHNm/eczNHGkBBXdWVMyVLyWXiHTV8Jlz6h6
/8M29j/IKg190ZfwdiJdRT3d3QsRhpqMGY2BNOZzewxgveaU6bef2Dfhop0XScow5BQ79f7mB1np
eyYmL+xdiupmQ/YY8n78JgO6oRGOHEekRA8JD/oeiqa4VHfKKipzEID+SiYCWZxNGos6fC64g+Jd
jOBFYAHmTZO+hj95itLEEnXC5QnlBju5WOUifDKgSU+iCiyiAl8D3EM3YKAd/GhM2Ai0kqNW+2NU
c3+Xp5d0hgN41Bvw3rgIkA+JyRRwGq/4eO2jnnVRakSkPJYaaJKf6YOEzoGqOiy1sAwCh+pB3I1B
cRKlmwSAhv7RGlbh9P3EQEi57OnvdHS1OdCM8fh8vRTKkg9Yjv9g17yA7HDbL5hTiEFRX56LAjzI
9mcL1gEUvLYc9Ac51BJMBijrMf7DzjEPhcxUur2lo6a9N0XHS6wrLjgo0G7BSk4NNSCIywM22FXg
0t/H+afYrEaWgK0YomxdUpWswTxx8lSg/Z0HRbS1xx2t7/83zvtHhAsfEYyDY53SE/Ytyd1W64qG
apJjwHF8XdkGVvH2D8yRsCqeKkGY6oGySp8NLUXPs393KCYoCrc2aSn4ydGHmdgOuQu1XMfxVaJw
ZSzrqSgSShq+8VBYYT17KKJHKRwjobkIEF+qq5MlaUcm4kpjiZ7TB0j2b8vqExBzBMj2ntx0D187
cvLP8ouIBM/W/vye7UzXpjUYNpkdw3EXI9+SIxwbymI3Yka172k/DetFWCtECP9jPQcMEGacjA1P
lg6N2Iqyf+bti5WSe2T7jtCjdy1AmxhNbCHPBtf/0DgWX6U+hEvEfBgXGhgSxxgsdMva4k0NDezM
oOepvlvVt2OSeEIe/XQW5zkA8xZNwkooETX94+pAhCrNyLZ8SrXDv+0fkqlYobDTTMj1ZwVSzLm7
KqYHD0WwYyjJ3fepkOu7MYYU7t+ItkDANUqDbfX0e+4P3FnxnKh35eupWA2tZDWTU14UWa8ig2dZ
7fmgw81CmTmvxyIa9NwYg4o7WM6Y8pFHHyXxMhwrSgoWgFA6tF/NdUeXKTaicY4Blybb4bVcaog/
oocJ/UQpx6vqyGBHHfR7WR54NhARhqFYjHnesrXtVD5S+JrR9RJlIosWgP+IEN4AqT2BZcYsqIhL
t5Rxx082CyNNJzeeJCxEId4FYPlWETfN3rQPLQl7Cyr/q1yBNX04SVBnCLqPgm0XsIDicvR2fwsZ
SUqk8mtZnqdt73b1DYYnE94FJO9kcqV3CrAusTfTsyWk/sUWzgLWwfdWTgMUwRrR30b5pzKR1LQP
AyCWgAnsots8oV5DCukO949aC0Wqy9IldOd95q3tbN3n2YZNq7xckpnT6vU3G63bRT8ICHdW75GJ
PTYC1nP4Mcfuhb15HcnuXTZP0mZluWCx/RLkMQP59zleQeg+QgVVmY9iVGe3bQWP1gaxJXZX5aYt
8uvmPKK75NXsiv3HVhgQCr6+q3Q5p8s7mGmNBiR9fA8yvNRvd3Wm4BCgiWivC9keeriH9QVLXat0
oZrVmilExiyLLFZOFa2g4IxWz1ycG3nMklIXy+krjpLJjZXCZoyJ+xYAjVg0MhlCXrKA0vIXGqwn
C0+dsakGuPf9RnWxgB+DLuestgDIgiYw5Eu172dGdwBq4MqiliJMHTqWybRA52Tx6I9nA8C0dHb1
V1Wufc2QtDtIavl5ZbYSzfz7iJdL9ymO68kVbiPYwJtGwLTVjsi9wqHLi1/cavCo1ZLDUGv+YegN
gn/Qmu6PBsbstaC9Od74A3z5Ye0rNT4VrzzofpULePC3MlGL0zNKJPbC6CVpeKGUEQkYdc5C+zC6
5ILVg2hJMEAgaJf5IKiG1MafhPgfIjOVzouPlCRMf9h0uq8l/RgQWcsUY+OXLD/HsCfYAosiWOsc
mqbQGr0rX/HIzNBW+Ri/2HviMebUfsF+mXfTir7/fP/3aCwYlk5P0BOyCLncBqX2xNsVa9tfLjdu
WnHp8Bb6BWH5eQ/6RJOsMG7AGD82IPGJ0zBIJt6xm8Y7vyAO1+KnNqE+Jqsi5hsdTzqyBijDPmNl
wS++lF0Uf56nrHnDOWOCcJHvwgS2GxVbWxQ5yhSftxuh7wrgVpOs4IzBX65EGVOV2xluulIh3kNM
LlO/WTZXUbV0ERtkwyRpnAjO9qlF78TLaYhZhBNqUIQfGLN29GmDASHrIDuXFy6mSQiowaASssea
BviuPiIjzs2LxKohlUcsgAOzeO8PgSGUvNuAM6hbhDPcHYkJbfjxp3eClOHVjHvVTRd1rGVOpWxU
7Gxsv9lCql9EounWYV/HrnEV+1PKAUcj7e8MRaNB2MTE6OtD+fFtwg9U0Pn+VrGG00frlMAUB/Fw
whIW82fnBcKwYYOq/1VeHqon/xJwZbSisT40YEay8P6hmYgVzqzmu57HDePnz+s/+J4HNYcp2mB8
/pRbNDndPsmEm5aQUg0FYFePScnI/rq9rtyM4K9FoGF4+uBIrrXHPjx/kCH3Vy6Pds6YxK/fpQRb
v16nF6IFuwzzE98Tth43fsCHXc1TV7dPlo06+WowamqzPR4qWwIxEQKdgSQNs3hEnnIaA4KSwu2t
eBrXRAmKwH1QUguhMmtsGUAvPYlN4GsWvLVBJmjTbW1RfG2eDUuvSw59fKD003DbnVgwsyzQazsz
81bvlpmFT2dXDYYhp2qRNbQMYuciE4w7Urj/lvqLrtc7iDF21g8HRePEif6+DS0hMqThYKkpFLUW
kcESfEZuNaJUhUFbcxrkat6Duj3d5FiIndeOdtm0HtyUEUsM9Y68O4iNhzHPzWPM4meDigFL2dfG
JJ9AniCFJl6dvWQwwTkvMlatQHlIScnHLejI5/xhCL04QT3OJayx3wnPtnSaefZGSeGB9JYIGP8m
LJGQ3tC4nCTxL+OT/ar4xHORQeIJ3/d1qW93+2Evn4HQLjoVojUXKtMeD/8r2EvJ4gLaFqZ9v8g8
TC6GVHA7BIfbSa+7fdlH0HfY8Wt4lNYRbT47wuJXn9dI7Gt9IuPZG2otcfLaIewm3Vw1ih+NjdW1
WFaCLVE/lQiwdMcdVhI68AiYL3egTh5jqlb/HTQ9OKJ1JGV5fQBIB8dnvIYjTMcEtI9vkq3Fw6m4
oFQXLtRNxCTKJONEkjLi29l66+Y+jUiKUF6dFoNE1xvknSsXzQ9TpyhGHtN/mVbVd2n9ZdA2fBDj
lYEmIJUk4RpL7f4Kcrzo4SKcBAZZbv923GzQJUS7uRzDTJ+EmRsyE9VRvX1SoPnkYwBw/LThWyGO
xi9auJ0AiZceaD7YurcfRlj6xjvAKnfe5Dol5K0zbhi5PwfrHh8BrU8rnBkX9AGNjt6huI3oixrQ
KkYFQN5NzA7vwd1JrPSB/MCPJn0spgorGj0aVqDEEjD80D7doTSRLawvLqYXSfdXXVyLnlELzIl9
IJhOocmoC9pW+gDwTm7y41jt5afFM3vl+7vN2UOu/ZnntufMODxap7TLH1cB/9/IZDCFe8Xd1iz+
37E+/aUVHrsoOTLOTaIcIu0M9AtkFL3FB0ncfQLLbzq+lUFlrgYnL9rtxBPKoYJAHFlLX7szSWNN
r7354Iph5hkEp2HZdMtB5MiBArkHLPEooQ8Uop3DXrJdkY9a2X5hjNXy6EzWfjDgqq3tgP2QKvx3
PiXGi+DyPNeXPpwTgusph77GvP3qBYzEfhRlW1W4VrpcvHu0llo5SWNxXnS9QWz3hNtAd4jCy8ua
FhgI6DkJqY6CExGNPXvRWKHUS3ELlTHyobgzbkm3ft8BRbzHX/Q1nhn1qWghlWvrXJSsqxvwmbFi
KdRniH3auQfh2e5+iEPDaWorQVk2AngoC539scehlfc/VPOJV/AV9xHOKBy9Psz/zSSRVwfnNuA1
xYGiNoRukwjN1pUSUP3aZdSHKofZr3WnD3d6xvlufI/1nZBmz2y2WJiMJ+6h45MJfIiucrQcnqdE
AHuOxPilSMHjaYjcaFJKwa8v27rQyjDVbQmzcqIukN3O4KoyaA/RhbALps+1/wABkwecw/5upvgi
h6VGpMo+VhnyhlMEhI1DLxB3y7ScD15LA4uFz7sXT8sF6HI7lzMSkESnz2rPXorF/NdpjwYuxEyd
2uLfoYF0283jnqIpEjQCBAuxK2JbrNMDIZMGcUEghGdySxo2OyuyeKCVJJEZZ9LgMYvWG+7xdbVg
3eapMHAV/FaMDYewHifQaLT2I57vRYLdcP7zuRFCkHfFn70tngPpM8H8Z/CNpxCghx8NOEQiJpmF
GbQwpwgF0UN9/cMrkJd2ax8jypUWWPpR/dN+iPEr/wtU9j8UYy83JP3sX8n4gak9KWam/Xg3769R
SuTitWqmOrgNPFG+4vDpEWvOXkLfEljM6O6fqzkaLc8Rwk3mukU4JymLQX2PEegJrsyrsxnUSXcD
M8HmhMquL/98LLgAFYs7Z/9xVpUxM2y2D2ZvYrP7bEp5km+CAKT02mvJdrjzhqoOwbqfmJOnTZDu
aj0ZZ9HesOOFU2yF3R4Ek4iRKpd8yeObIe00+7qvtZN7hvvvMk+GEzTu9kzeYnhBgWO5c+C4Mvx7
+WBRdRhELbq+n55NOx/xPUbVgNNYlqVGVilh/iDuSOuhijJRFTXS3q2qbmKxFtX09nF70r0H3C5P
AgV2gXReAGN5w1GoV6othTcV6SlvCGaCVA4N+ftKogSuFJZ8jjG3eoD7K6FjCsk+nkzyiCF+VBvq
plkO9nzK25daYZbe0eFRe10ghkpfsFQcCOlM8OcsWfCpi6aZx+ZXwubm7y/UiffXukUWPLo4v+Wa
oWEgDnKG1b/x0/qHOTpj5OoOzgDlGyfq41qTun9n/0No3z5zkmyKTBI4NN1KAVM6s2DcVd00UkiW
10oAtJmihPk81dzWiB7f3Nzo+k4e2J/LuGKz1lllRfGDeiCrqEXT6z9umOBF0QB9yFz/Apt/3U3L
NZfb5mce7OPW/vW3de9GHmYPj2B+m1pr32Lwm2GEFsj9oScyprALBjaz2I+51YXvhFOD8grEodRC
+Si7+xUbJUXMJru1IZDozDEgHe3cr+Hjh6QbTG2F9WFrEd9vpWj2Dd4M0hI8CU97KaKUwn+ANjRg
8pGVHpJjB1GP+Y/yFksBvEnI0ly3sCffjTk3jVhQ9c40MTX4b9lzM35fiw9OShoGg/MC/Q6bTftp
NTG+ucieMPswJKOWNwTMBy3fSyRR9pXbgVZBmp+RwTG2VN41TDx+BEkUHwaNynxy3f7BeSFVg3VW
sasts31awnJLnNtxYZLjs3GLJZgQ9PN813Cmzb5wLGqpVslanQmDI/fjblWrU90sSzMZJQzg9MUh
zOiAq8eraO+tXOApF4ih/NxOlEbzWELIsSPjk8ihJSyqShx0QHRTfY0yOFV556bzTncmrb+JRm0q
FvImxicwH+CHDvuPVQ7wF3JftK14nXoBVDE6N2wRg2vy1VSnQNLKbgmYEwV9RJX7RtEbBdBiPMDp
JqV+8Xr60OnTMSg6RtEgpib0Pp9MtpJqRwNIAv9SHt39hVqTN7PF2RU7hkG4SuHYsxjG/ro5oJrx
HX4S4/W2c1vbpxQB2UUWSz413iwy1+SUhYU2N1IhSSeJ9ioVBVUnr8qg2ALxZvc2JTZvRN952PZl
Mpw/pu4PJX+yXIX+VQzyzvmrP/O5DBeDtjDZ0TpUKT83MZx4Buez6V0gAkfR09op8Na1J13jfzTq
P1fSOOF5fyNquHUpA00FF6+hkrj6C2Vx3Egr0pRZ6gWvMa0lHblMhgINaqe9TXkFcW4F5RMJXLVk
FfDNAE7C/T1ZMk6CznCqJaKABbn/y3vtQWc9gM3FlNJh7c6+1hjCnWDcTkdERTiVrc8ZBJrxzflt
Z9nwXielYXRJONSV1YBrGyMACtor9sgZ9b0wXd/OfNDXNj9Z19RR+CdSco17oQPPJvnYL0EjKsBK
VKAxFxcj8rTB9qdxsIT7eSlSS0wiZoQjB3dpfJk4udkpDRw+XUvRrciuQgBqlwlmsJLW9ORnN7vM
YA4uAAEv9IWhqJbDaO3JsPULqb5GYFcdtsYMMDJdJEEcmPPsaf0p/InQdSnyeG5ReDYnniCpWEQF
wLZcavfwSSlNfmI+7hGdy4KUR1k+kLysi+r/nbDRLKoQjLLZ+W0DBxCscGX98mVNQWSDwvmFbZOd
6MzLGINYd4SpScjDEPoAPGkpa1L/HDCCtoKRav/PP7uRdclISLsaWAPtZxXw4SC0abpUxigDV86d
LUBS5WuETm9+MoRcKXMApRNRr5e43hG2fN1mofG0mK559MYmGsGE6//IuZ2FggcYLv0FBhmQvjDh
3RV98fN7Vb4G4KGRwSFk6ACzLr1sIfr1Fs/KB+bV4SmBP/49pw3Z/CkhdDRYI9GBNEXjp3+oLvW0
XHZXmybPY+tPsz/rrnm7/t5h0kDlhxjUId059P0TbOZlsaZ3vJGnTiHXbr/LzO3DI5uGK8mNG5aM
OkmhVPKmFd4/n7EsL1JKNV8pKCu1/PgzZcKOtB4XJCvDTaLPap/yX9fpSizqPYFW+yRQd8P3Nt7f
4GUD25R9mbSPSAqbC+/jDp3O/38wHqq4NwBOmu8bpvHhhghTd6rmA/2wv1yJxY/jmObPEm2Ef2No
LNtueoNAL0GyOrE5dhZc5TYCo9bydZkk+kkwAKPihq9Aiz4sbblc7E97fmRGKvyYoWKVVShL8u0M
sZ3lOAVCDVpYcX58h/zUf21kB6c7WunbaHaCd8NyWlJWHCWu57/azrw4xEB4uLOFPcsRbvEx677Y
CS2eXD8f7VoTlAD4V8VU5oC0uqySlIZJ0iXArhI5KPzEo7HrAsK211nFACt1UYmF/9Y/iRYqZ7NV
fHGVkQe8tpzRdlt5GJqVYS9RkxTievVIJfOk+Skxkb1ZTYGPmjBXIjdVHMGZbMrYnvconI+IaGRO
JRuQI2kNSQcZ+gkR8LZXbw6lRZWGW7hu5vC6CN9f+5dukXthSnOV8H7qNOMCbzEj7O2Nn3uPfY+s
pPktwleN3sOGnhu4XJ0kj0ZEoQVlVZV9qkNismnwzdKikX69eZ9au4ajiwQba6/0ihIdQZXgEB8s
xMyzRKEAA7LwCH44gra0/g7wtB5wgfTzsjMHsEWphiUDYD+aBxQEDS953FJ5tGT7Lz6Cv/lmBr5y
idZ5XkH1rUhfEkV97qHUH0ZLuO1xAucYo6KrSBEQyCmTM3kQDxat2KtwybkWxsdThNwp0OaTWEz0
1ByEH1a4q9lI1/+4nZtdtaHnbhi4aafQmD4t/H+E72MMeHT0g/xXbJoRMpbNPm8LO2Rr5GxOjfUn
a8eCxqBbGLskN/Ry/kVMMYSRDPLbu37zn7DrKk0JzB/j420EOoNsjuBth9zkvSMN+jDSuZTs/05m
erhEaQS1jgEL9Dk35OQ7Y4k3divpcJCgKIXjsXeuFMSC6RfzhWQKQoGqK18STRVOsGWzAE03u4lo
ob2gNfcqBj0pZI2k9mfA96JmwmUft3mM90OoKypM7XBmm64AUeu7AtGhQqoloUHCXCNB+KYvOEi9
F1sCSzbZQJ04LxPT4IWsD09/IMcZYXpd4CBbM7HTXeAyACdfRwAIbGmV+SUgntO4n2/tAE4LhbvN
Y91LQz9ZjQgOOqaO2RXCPPDbhQlZYMXUb/mO83TEM5N4wTMFyqtWtoZzCrCpG9ooU9myvRs1S51o
WaFH/sABOr3N0S3aT5CucpxlVx/behfssLdUKbML7n8pQivn053030GhDYD/G8tqMQaDe8W3UE5e
BJ+roU28dBaWsLUIt8QZhXd57mhA3YZjnC6zUAD0S0ylrzBzEuLc8YWrDg4VHIEy5qGPEFrT52Ji
v+vpa6Kat5W4Wg7KRDAEjYBi+GUIk24Yy6KiMmeugbHGFRXCJeDXhrEVCRLVAs56iF6kj+QLjaKV
Z6hLQkXJYFnnuQzMS9uIraaE8TetshZKDV8E9VIOXQB1MRIwgsMieZcM0DkOK/YPcBj6RP5zLDQ1
bmwDyWMfJSVk9/L57OynU5VU4fCvjyDGqX8DHvJ6dgf97Au+Znl3mUWTUgBWof56GgQ1+vkt51WV
uN9bUBeN5j6bm/22J91TSPGUq5dpVVLQJbqMOgM34rD2COf/Ns8vZKNISx66C0Mo1rzk9ROj/aP+
zaAtZipOZO/KkLoCa7Z3hthb59LqrQclKtQ0f0t4Y7WHjMeaQYBO2HUavsIrVuwLkkOa2/nm4L6B
xQesWdQGBoiCvwoOIqWgzsdPqbS4RRtfSVTSZMuQ3JjyxUrVHhUzS88zVTAKYGivvrW4W35yumDX
hN/dPr07t+xa0O4UrQp/Cc7YvK2dmGtxP38qiNnLYvLfdrqSdaxLADFV5Kwzro6KEpUG0CI/H82Y
YPcrrlAuig2YHu/c+gbU2Q29veO2l0JU6rUzBebmCfUVTVL7u3I9C7A8jGeeIX7JQ0aP/6/8DziE
X+dH5UY84GzSzyy+BXyHFJutg3fxxcRnNeY/hs0gMdB9wSI5DcELvhcZUmSo87ve/O85bHLcwJ+5
mjAEIJZG6IhOSB2+3N+539km51FQj7XiI5dIIngqqVUCtcQtx9l3suiE9EIq77Ut1K2oOztULnMw
N9/aEUrXWFqN+rwWyFzOOPGh5vKzT/RkgaoJGrD2+T2h9DZjma91339PmmtAtqev456L4FqpllHr
wi5/lY2co5+Dm2PZ16ZHUTnFZWH/7yBcLmPNyNU3oMY3EYHU7G9dHi40uSGMQkitMHmS+BNy7oD+
LpY+rAErAD7VYOV4cLrrtYc1QgW6hMBq7nCF6Qif+PFRjj7bvYdeah51xZmMhpFPGvFwivgEqqUY
8xPVZqRjOSWGLf1Ne/p0YJlD0Gu9TeWnK0FPnRPlDsTi18jKzcQToqvBQCclTJKAwK6oAiDKfxID
I/qDFyUPc9JYWhRywpIXxGhRy0G+CQmEYykalWX201FmiYtcKzwDLiru2Nl6fLjE3Vq4+j7txjsk
Z7oLK/DMPPtaTZGNGEoKUmiChQdZUm1MAGzB1437cFaDlIGluBwig3MRCNZuV/1aEJWcNhWnWUNZ
6cfanmA4ZhP9qfoh0UKL4tb0ltMrvUjibM2euTRbkuTnHbmP6oOeGF+tTDez5LCE93LgHu29sfey
3MA484lumsUoX9BynARMeixziFEZwMVXR/M15IepgiZ1PD5g9EmaaRlcl5pvJXmWYqEPOqBxlNpQ
rpaQANBpBBH1vlDwbLlnGOvuD787FgfEwXJZjmd0TId+5cLMeoP1aiY/KzUsxwmeC/ELz0pg2MXS
lZ2gx1TLWIppoO9en54quxr0MMz//uiSgoP2OQQx/VaN+49sYUDewf6PDq4WyXY5vfq+gXWISzSG
A1kwK1bY6D9p4Ro1B77NiebW5md2rGef7wn3Eu0wUUti2BxUhI7aC5gHqqGjwGJS1/7+AOom9d9k
cYA0w4lq5EiaLbzAmRlc0by1uASDMulToWfnUcGoeLjfshT31TZHbodlTYA7dfT+9kJ3GKHcn8Rk
vx0BzxhwgNjIYfv5FMJ7d7rgmSr/cLwAaUQbf3gFdHibgp2clqYSmJRfV2fiER3EMpwNxAdz0iXn
7U3LCALgPr8VxIM60fOxe/g8ulHUPUCw7SawfUcdCyOUNLL58B15LNgjPXor2gTqk+M+4Na4IPqR
Tx+7fUyhSmy3eXWrNj2gThx7BhJc4CrVJB/CdVbeAYYy3zzI4t+Vlo/QYB7sC8vgcQIOu6C4WyFg
1JTmlW1+MIx96h+ZZlasTAPe0Tf54qDeSzG4LFjyHhbUYryio+qidj6+XMyyWw13ArqvA+d4A0i4
mwQVOqelz0/1vugthU1ljoE8ktfWnqQnt7B+k+sGcJXX0PRvtFht8wpNK3eJmNT2+YqO6Mn+Rbum
peRZFA+HC4Jsnw+oxPcuSDMfQ9oA2mwdnLsHm/PQVjIervE3GcBi9NJQmAzL4oTvoOo/lPH9jGiw
7wlk7toYkwj+Pv/vvlhz96GdCtvT5eqH+lzp5iG0WLAyQoldIKHyTbFTbmF/u1qX519uxyHGy/So
tmmvGb4yz0b0IT/Zt5Rj8GQ1HYucTB2IiIewsSAJzZAuQr1k2NFc9jjHEsrf9xW8me3CZqYQkf0F
dMQJIB/aGfPobhDZpnRIpgQl0S06WlSJg5RlpngZcAOLQeTzu5M7SOMuyG/D0I3GrS/WvDaEpPvp
vU4sSD1tnDJe9YQGaMLc5Dgb6Faex59D14vja+a/pnjJF/xM1iTZ7zqngCiKI3+DC1v533pdSGo8
RkubVRITGKpUT981hVl7y+4FovoAzVKnLJJbyokfrgtnijNM28gft0QYzdeOrs4mTBTNm9QqjEx5
uLlAy0HK5P/HBaG+15jUIUMxIbJu/GV1Ghx3em3/LKLDA58o76oyB6onqNww73OA8JJVJcPBgs2p
gjBnbxjHs1u7O+zbzxHvFfEia3idbnwNAIeOu0OdPdbDceDzBVFEXoYGiIoegW6g8BT9ADKeetLG
x9kn3ZARdXUCtLUFfzUbIRKCu42ApghJvd9HaJz071oM2nbCJ+TCEnm/L9WdEiz13Mq6g/jKgp2X
qa3Dkpl0gVdfkbROMaCR2MjK8t/q6fqtrP7g5Pdj6TmAZjiZG8x84wBDGYy8pElKykboFygxSwA7
kri1IURbasmlgtF0uo5t5uzh0oqrPxV9wjn0ittiEdEL2lLbwdzfr+5NE8b+8w6QjP3CHQHNa8YV
ci0EL46UVGyJfPY3MYjZvMKMX3R4sNsLasBYxMj2ADshcxlEYHZL82+7XSjXitDN6My0UzRV9tLW
z9vha76Sqy7ccog5pdYRdxIHatlXB1jMmqXKIDk67fxxWxm5sBdLnNkuwgaLcRxaiV4VHQVvSN4Z
PvDcJspdj9dPpQNkFFIpzGAxWH+qYMuE9dpX+NKNRcWFmAy6Wpac80qiueR+Zb+ysSdGM8Sft3/h
1Tn0ifFtzYIdQuH169FSEJEfYPc2Gvc3+hZsFQq7o1AvXTOOBPw1trVcuY3Hx0F5qS/J7+j28/0S
a3P0643qZz6VROxW3WUq2rfex760xJNYerPGFsjgaOFxBeRZMs/0zwZW7QsXA6h2HtxNGRhF5WiW
m5qoTP35LFP+h/H0JXE4qoZ7yL39c7FfoSVBiL1RXEKyVMSrSnoUGfLPRLn9xQhiOUvNQAMcrcT7
UhmxnireDhXtmrc8sFJkIHF880UFZW7FZn4LQcmirBlAjueWPGRWNjuQl2GIVHDNAaLp2zr8vYHJ
/aqieo1KGfPDZ0z2p8j8ETJtdckAeENAImNTQ+oTy03PzVDyrR5cDdsy7HSF62T8T1OTLdISud26
ns/FIdPXBk4pD4Tlo0mRfKrR9+ClDs7eYjTgg0P16iRAbCW4hXcunTDdvFIviP4tgLRj20SLbR+U
euXYz4acHha/V0lh1/udO+WKziDetJ1ZSHpHXaeDbNHl0kOkZZlQizE8g6uSXn0tbYr5qLlBQsiX
eI25RA5gHuOZevV3ldk65KD6P5AWY1FVdek6k5bVBykHHEKKtH/m4bYZ9HCGOA7BH6lZZggGpqj4
fUwz8AuZbst4A5cQd1LnQ6B1tdL4jcumUNW0WgaTW2ksHRNd4vGwxBIPuJk40Xmtrz45jJ1dN1Le
MTx/hd7iDZADBH2qyB7FjbFw3claqeq58JuoCfuFOv4gxXk5E5ccZ/lTA4byhTfE/jYYkCVRUM11
g266W0VSi99VwUkqwXyWAObdMT/F1TfdazYDgjSXXBK4x+amWT8IVB2KqHohAQ9i9El+HbJFqBCc
WCpXdtqPxLAKuByexsVzKtBzFpv68ntuc6KYWSJG3awf4iD5Rfviv19BmJOwqXZy9aOCXfwgvnnj
XIRYQ0n9Z6odSGqTh/fAaWGm53yAc5yF4EWKQm9kIPhcGGCeRdz5xcV9Ai8dly1pVPCsMwNf39Ma
0IUo9IMx7uoFcwYXVXYF915uf8CYrYecsqRI8Y2N9Iqv1+Hb4U2TCE/PV34ZyjrZ2LBPmmftC7LF
WiN0hb2ffj7aEUIKHjmpKQGveFqWw8aG7bN5ZAxtizkIjaIE6WnuARC2prNVI83wX3LrjFQs9Fbe
f2a+HZ8iVrYNeoudUTuE/em5BkkspCZxVGLZe9asdRac4fgTug3L83Kx8gBa2kdDJBS3T6vYx5Dg
IwfxtSyUdEmnmUNsu8jMLAeH8XNrjOhX6lLi5Nx8RTY63kl70wL+zJQacJakSwCg7cdqPFsD60v1
PXkpzKUyw9ZauovxlSJtO/VolgLdrnUBx1WtXYq2RvmJbdU48CKCx1xv32IWUvcwDe+ks4V2xXk5
YZZ8pZ4eudwnn1LPACNaGSkE/FoQKoDDNadxe3SMoX379VsnLc5zbEvnDHFL1af8r6dQpwqKhFZp
CFR7VVRM73ZkPUM6cowvBxkjyqPavIffaHR3ZsqGhDZtj8p0hmIWo4ZNzGvsGTOKD+iarqPOb/SH
/ekNZPctKXBpzuenQXljGPljrDDODHfclTi/J1oTAN9zd1TzpXxy2iQTWxoGNyHA6wT3zO9byH4b
g52ZNfReCqmaJdGyl7jogD40AB0zS6/GICCu0ChSaCumCfuGt44fx6JcsItw+DKwprYWRAGD8K4u
F31tI10cONUB6Otq1KG4ySbxsWrPCnZu7zLMkZpeblKKnBM/S12fZsLgpfLFdO5/9+yEX2a4iHgf
2+/s0AtrAds0c35kxd3wns0H3usn4iSv2Hfy/0Ofi6nxSyxcDHV8n6PZxfWzwc/vRG7xu8hm1G2S
5y5KhYImX0xfd3eKBNgeauwrtT6NzkHnDmSirUvNyN75mWvRv1r1o8zUo34lcYI4fyvL0U0VmwE8
pQqEztnrNzR+lRMZPmqWy4pnspB6weytICjuMoxYryoVtYUCfk5KRM8CRaUWM+NNKRNCLR6KgkvU
VJoPgkz63D1vdeersRTy4Gqs3LSWj5mDIrObmHV/dOqiTuQPPtBsXT/Xle+BwDlHowAG5nAN/pG7
Lm4wcYT3OkV2iAPh4bU19Thqi/GXJdSIi580ayE5nj7VMccOVFkdo7A4uyL994Ohu/6gkYHTQjDA
/sHR8zMFziz2G6GOLHsjQRX4XRlE/Lh6F/CD3qLbDVOyvAbzTVWwAl02WXp7NOLy6F9hi8xmfGUF
BOKJixbrfRoRGJjNEqHtV7/c2DhH6ZaABU8JBaMDLP8fdszp9sLUfa6hpVISYapHTUhaiJ/g+S31
L3DtQRVdzOXZkxtyBqkVIDBUbuWR5fZAymWKDOm3jpbBmH5tNc670RYXEXzaUSSaFjyi45Suwo7z
/gYR6I5I57wg2/DlQOqWa9+vL6ONXYtvT7ZP/wGwgTI9ArKR0eOcl1WFR/7LWe82XGxmyjxGeIil
mIw9mV1YeZcTOGBhK2FHCGfRqM1aPrqjAWzo56ZAu83yXNRjnnkhOO4LIVxAo5Y6Ft3Mz06hE0mZ
CkDmkhs1Tebng6vDPXdRJqVDkmi3vcDYH57v7ZBXOYYEU4ODDahPzo7ZRkumgaUxIRE/RjDasGWA
vbfQibDbpQsWWvt1V0wW80JhsMQjBispDG1CT/ikVOthlPMFhh8Ub484GfEQV76Jj8cBGlGcb6eq
y9Qomdw6uvi8lzfIUmkIWj64FeKNKYSnxJf9aonzuItoHq71LmRwX72x6IUoO0znwPvbr8JIQJ3/
T8Yk/Xqu7eWqwUIL7Gc976Z3+qwKID5vJ1crF8RkV9ekCmTNq3VQUGB8OUEusY3mD54dTX+RkOs0
9FJOswdtEQZNNX9fPsOFQavv03j3iyYMVk69Hah9KSxZwDZKfs43qCTwDGxeEOjc45zQCilqrkFK
V+dbW+jGdxbRrJG+gnPi7QnNn7XwHXNWagzuolJMCui8ePiX8U/2aEplIOf6E7BvCrL3gKKtRZ61
YGs12d1I72MSPpC9aye7+BzcSoX5kA7vQlmBeqsk5U+STNf/kZGIzyiKuXmqPfCtPxu62LDaoCWd
1bH/U4ExXNi4GFgHN1dP3V08Mg2OAIcmdqpUZwcIX2Wlsj4tKJFQLVFThk4a8D1epfemRJ04zMaF
GsD8O518pBL2OAScyk2lSW1fZYGF2IiYVWwGV/sLIfWwGV1DSuCi01izj9ZkgrDd30HR7T1dik61
1j/ed2FEyymCKXIbeHwY4zNDXyr9W2KbEi8Wv8xE2jU0zWy+BVlT8CXjobvHRCrcnYPDryL0up28
REP9kJKxKAYfqkDNX9M6JyctvBGqgKM2/EIw2WSFw0MrI2OMf3QOgCvTk9Y5s6G8Hg3+yeih8MBt
yLn0a/rZq2UPqRE6R7td46ruIpGcOrV9Z7CPhn41x3aixptDVZqYhbl7pQS2mLo22tyztn1y0w/c
hFdRTsc4usYAJOUUNGTteqxc4rgEWTZe+U3Y7fZQsebA2/3xrSCke+G+9quJxQ1shan/rhDP4eyA
ALCJionJILUO7bDN71SyVK0A6EMtuC70dz3QctmZi56VRZVMwqGkB2juSv9dsGk3QiIV/dc9Trya
OSGGRk9TT4mCEI3NFlXaD42fPo2limgiJEdPrmp/aH9/RCy7KTOHWQ/Z5A3BqoRbRLrPZG6eyux8
QC+zMQBqxRkCoTPD/XMEFn6d8Aas+Cp0CLJsYE0jYbFQ8JFMkcnlTFhN3stcR6SMuM/67Wm0ZgY7
g+FPYwzNf9x3qgd/QKgq8+aqUtJTgZBfK9SybmF5gSVeKnmrtPCWQV+HHbe6ymWRynKWUAt26zNK
YepYsxoGnKmD7XQkSyN46CIg71xZGKO1Nduj8HgvvI1Q1JkIqzDk1xAi6x9MRlzK6lSMpFJT0W7h
+aUawIXKJC7ZZrnJXU0eS3146GORlmMFbGBIJhS3zic0QZ5k4L6mOBaS+t50HCwCJo/a4snHM7V6
ITfqHdW+26vdMfyeuklJ1E/427qFjAmsCrTaGkq+q/Q5w5cEfO1ud5UB59AsIO+0oYxnLcSM5JD+
gJkTiHm9mOXfGq7ncJfchXAmgJUoPYyqtFSHOHVwVs1EeVynmgmxaggpp9LIHVEncrlLTurVUQDu
IZtKCr7lBDcYjrw0vIY/QZNRv4pG9aZ8XRqfgOFe5/rYmzeEJZisiOmCDer+1sIKknJ6y/2TvQ4n
tP4bxdAx6cxVdecGDGyplwWJItQT2jl6ZGuXY/4FtA95pb1OP4bQy5HhCfK7msG6heMqoFR0Wxc8
ORatZU6aajkdujXCxXgSj9Dj+y7O3KdGr+LIrDpPyszOmbOATftosslvD+55IgGFTxQmlOud42RM
GN+fZYEsWIHB+IMjBLJOY5nmG3ww+3sTuXX649aocCpBETTiklKdyqOTDSP4WVbvon79WV0Nu4iP
/XGvSsHwYF1vsdfZwwScejTYFJgORsipXAXGhqwq1dLOsNqrM+p8nUiCRJFhmLMIzLDT8S5JLsh7
gOc5+x2Z0zT4CS7LNDjgxxZDJmED+ENejkAJR/3IlGMQyh3ie+sW2Q4s7Nqqqd9rnIscHRNieT9/
PlPQQK7KykGzIP6sBwpHuR9w0Myt6YxFwuhGFhX6OTc+2dicSs7F+5M1v7neBB/UPeZ1gbcs/1AA
EIWCDaCxYT8tGyJC1ZNw/Hv+bn/karomPTdjbjquzOIkZ0YbjtfeZjxu304q55QIMiwokmunbN9o
iiS7hytGFnq0gOJv9OToQqaLnI5Fqgkl3RGe8Kwfsberxqw+EbXNSsrFmjlvrcT5tH36JO8XU1Rw
NqhCUVBzyzxducymhxOwGOsZhXGd56ufrVTgdNdOUvGuLg0W1H0bBKFp7kEHJw9yeny7mHJhYuOj
BJ8RIEqzYcOYgQ9eChdGxkCFBhWxo4qKLFrDiZxZ2wNAO5DeT/OIusBytPVa/Wm1Y/a3SRRbn895
Y97x2qfhvYH7rTYj4PNkYrXvLgV7v7i6umOwm/YYchMIXQ6XeetcZv0y8kTY3F52cFxoBYuHxVD7
nDdr3NE2TztqGxcSiiBSyUMfWqC/TN0O4xBTrQcLLLQ2uFWLqSy6eC/duGnDnn2X9Y4OSN45jncC
KU2DCjxrMVy7orzMKc2Ad+y2M6JtZHESe/ZlgKeedQVpWqSN1gr9Y/TBzEcHeEbr2Yg2HZ52PDBo
R64X5ZmMHAff7kipD8rYiyZMpkop2yY1woAc1KIkp7NXpoUvVZfUV7gTjPFfnylF0jdfqtGGDQub
IOM1gxEiNxWtKWTdfRPaDdBC8on9vfhW5BiFBsRjaKC+uWG0EjI3uvuH48Vkj33WU03EB1RnNZpe
UW7gVWL6c5ggP8auyA4NQaT4jRAE4BKC915VRCPKHJqpYLPpHb383D7/hOqZe0fzmvQDXXbVAotn
2w0cQgC97jcwuQY4EBhlZNz0rhC0IXPnjDgSA/keds/u0KXzQExtGR+dtSDmlAsT3D8imLbQPGX5
z5reE5n2MpZ/mgnv7f7R94Nmaqij7e6ofVrJPoD6NKSA8W5va3V8iqzxPlO8TqHbUIHUQYkD5cqM
fXAc2rgZoDNq7bOqMEOqmuYmNOnR/CxY0KfGNh+/p3CeD/Z8MSeDISVR8NG2rpgVwl72RFfvX1Yu
v+xQ5kxRTrC2mQN9j3j8PVPhEvrUjCi6EF7PMiTZvEwejtc45ibffebkf6sWvSA1ru0F72EzzCeX
TtjDiIDttisLgX0MajbvXiNuVABBqz3FjKjU+kQIOs9SqWHRUE72/cpN/b+Lb7vy/AX6HFe+XWLc
aCLr5sZetiOtDXV6egVx7QRajzQgZ5oza2eMuSFoofA0brNtSOkoKm49moDIiyP1fWO8C45MxiCr
8bE2nInQ9Nt0dh0TRX8TMKAk1m9KvYOe6yOtTZipP7uJAm0X04v5CcyppwWgpzD+zo90ahftpmrd
UC1c1jH50Hxho0e4lO4De5xedwMOdMsQ0MS8b1IsYJ+AtuRI96JYqoBYF9F0/8lhmaBpRCb+jhoX
4It73YC35amGMaeNFLdA7KkTSMIXNnMHHIPzJ2dD++GY1aF3KIqixZSGROLbr3yTztjJhy6r2ZX6
UJSl0u/sggd8j+BjkX0CPlv92LQ64taiPGfvUDNxfyVOf2puGfVoD4jgzv73aMRjPfpPFKMVn84g
nUnL8hehjHPwXQGhHiKLj6qtHnjnqZKsVbD2dnjLRdlKKSuVTXFOQYX4XdadA3kqq8GPltXduJ7a
cMxGkeyhffbP0DhQZTwFYUxqVQsAFFppCpKmDTD04s8FUyb/y2eRbS7uOo620wukc6/khf69VeNO
yXJNYDVJ/Sc53VBSwSq0QDuNJiZrGN9TcXFUGnsen1dw/SyMkLX7G2V84HgaKXiIkrAihJ7HEs3g
i/+9dzfvJHEVRy1HHEKri3ZHz0HxvL0IZVjtW1ncLN5T8KZOqsm7IZTYHIh0L7HY6oioRLe+17CZ
KAPyGlgQJarMi52CbcJelmuvzs9AAt5H7U5ZMTVEC89hUhKDqeJ1McFFjj32tSBeFXhztuVkzcqg
IeJwUeF9zosPqnk8F+609crUJUiIJcvNS8hmCuJJWzvGHObqhCb08Ss93p3eLAQXPUDBvIN/H1/A
t+GRd2PQ+MPXoJAu0p2RFL1X5hHuOOdwpPphhUhpvzdPgDoo0hBkyYIPmGc55QArGFN2MkXiWrDN
dps9AwNx592H6TnmmJ21RbUgr1jOBidOY/BsaHExJmeK6sx3/NGaZ3NuV117Yx3yaQVLx8dkV2gg
s5WR9M0GO71uOIrIU7MQBV9tM6U2ilr5caHvjHwBuOH8cc6Zt1FvG5BAiDTl7GHfgFPXi2HDdByq
wyzp1OKXCczbpEAPQyNnwlqlJ6YyOFy6qlKR07UAw+sJN/KE9nD3knvywqv1eUeo6byCt/lhUf6e
nfggPE/QzH/LfP7w1j47jfN2cTPCbGE17XKVNtqsfjbzIHy8MvrICN57vs1U5dBTihetBjltk97P
drdlZVrS03yUl1C6t48Tyb6XQyu0iMTK52RgnyvnctRmYT6zyvtR+bJxeHcSGz2z/10HSqt5XpBL
PW+AnDZHpQb2jq0VY/bW1ZPSRxBSTP9dfMGAHyI7d322Oapc0CdcLq8QPPxbzgLs/dVDgNhh8BBO
PDCeevxvd5njRtLFywXSHfp832YGE2BPwevFYQM3nmtUgebpRFkxO3l0RIpg750PegK8ODwQIkd5
VL75taNmhAH9Hg/zgTDFJPk3P/cS4lMSAtEN6SyS3cBO/Fi1HzdGDGCcoBmvGtLLaQpJGxW9M/A/
H6te4KnvrNk5pI0S9a8xftbEx5fV3ARNBUtex07wx/pAeZazwh+opxpDXJLYwxPLyKF9B5glrD3P
9mjgP73dULmVQGnaQQPiKgDDhsZhpDGVeEzbz3EmjaGoyGF2xoyAczmKSOczqfia3SuyPpjiySp/
8hLc6cTHf7fJF5xGle16922hD2+s69dzavt9G0HX8kF8R6wPjKjm2StoxUcdxMj8jv+Y2DZAqWvE
ILO/3uktGtKor1HZ/yrSUqWCERlFlmDIekhzgD5VqFqmBwBGK/VYvkoIooNqaLv8+PyF+ICMg+me
99260rV9H1YVJyEwtzZdVGLgx/iE3Di94I+ivT2sOtSZgqpTPnpFSvSVJRRFBUbBvEDKctpE4mYD
+up2DmdQaWD+3kSQdSgv/xsLn3zuZ0vx+Eoxoa0nbolO+wzaI2XGh2SOkbFuJwthw4imo56jic47
YVLBgtZW05HOalwQomFlm09jpdOSJt6KZvD/9IRdM4gV+Q9GQmnOrFPbVe7r18Us2QLRMEp1Fj75
7JDbc37As3SRyZWxvBK8lxXyNNc6LnDlGmuCaePIFoXS6wC3mU72j7mQraeM9x8qOis/utCHLYJ+
oetLk1xGnql4/4UURITNhfW3p5Ltq8o/4ilYC/uNQ+EoMLerTxatUl30JzY9/TY4R6LiJRbnp/F+
nUqQVU3EqU4izjlAg2hqpUwO/m/Nx/ClmFKcX4dOyFCtEhIw3uFuNfDIxQwbYhRWLrGyz3dNzZde
h/rTKySFKyfr4/223WdkT5+QmMmRRc0VScYKYunoTAhL5AHYjWH4VzHhSth5nKx33BSua4LprJjg
H2C9s8uu73EnMmf8eoAe0AKUUheITCD6ce8FyqmVgmQ1ZGQZtNZpV5USo17EXv70dNRozYXOdxNU
BIOpKrLfb6w6FTogaLDu8kZ8N/KX+o/aLxgchxTKQueL5lmsqcBsyWOVRUPFWVcTuBGf0GlM6Pwp
A+ls/Qd+9JqTIqTcBGyCi81kdvj9YzrD5bVsKDxRzpYPyrY1IKeMzsSvO13Za1H6hUpv1/EqtQfJ
nNCVrSWrdzL3DQvFh/gcqWWejQ9RhJ2Uf81ILuengioFYK0lrs8utgUZhgLgnDpWuGcyEkH1qJ0a
p8/s89uozuf6eoQ8wXntQRu7wYljwrK2lYMYtyeJBNDswoVgPM2eJuGqBv768nGGXkUBBuiBFD4I
lrTu/BVz45Uw4TaWtysl5tF5xG4kvqUdQbQvdFGqLXqLFOOjTBETn9K/FCA3P0OWyCZyygp+m223
iv+ebRo1Y/Dws1UUgF4wklmq2udwMdY0iaPIduLyFxMVT4jHD/u8fwVjDrKlegkUWgs4k/6chMK/
35mOpu2bKHiqtEQwByMVzwAGZa8ywOskOOuzUZh9RtErTrR7I1kyxJAFJpqFoMnR6dZ8juXlW/T7
o5250yNpUElp6o/b2ZLc/dPuh/YKVt5MyVOvsW7ov9VaE9uO63ef8IKzNsuhZVk63BB9T2YDYwgL
0DVXzVVEmuKfNq9DjLxVEZ6Yj6Nxgqt9Y/k5kPe60jaydSM7JclycEktcHY+lyo+dL601phGYERR
vr5Q+vv7TxbZiPNkl7hQ6r9rL7yrahCnkE6nKNSLdnNWkbvsXORzvtzmsvw8EWUMjFGcu54xCfjc
P20UbuKhA4EMhLVRJfh5OauZj7PqqqOQxmdyOhtOtzBViZBJq659ISjK63YjvfLQPwY70E2IhZ1l
vCHlU5IdRxcwx3ykmIfV1wCf7v/205bhykS55aUWXtgwakJ7gu/RV7KLbqWg6c5JaVsDRkqmc6OB
Eny1abQSE6K++hnHKP1UEMTFl/eX9pwY03zEjv/USeYUp/Eq7ZzirD3SmvQ5f9ZMiHltz2kW4VVv
f45IbH/es6XT706ului3k38afrR5v5hY+KXP1p0MEOAtmiY/6rK1231VySYzYaSZclR70v7n6GsH
/eau8F93rDK2FZWvwkFvnMcOPWjYcsu+IZL7P6QyF2Hqw+Djzveca3dYgE2VxcNV0NcFk0QYH0OV
/RjWqPcuEgGOO0FbenYwjGGsWs6NJxRDYYcRkK8C7cRwW7mt8wogpWnPZlRKA308eFN7lI0h1pdd
A4TG/UvCshp0ppZlKcb4M5MCbn77uTj5RJCD/bWFjjezNRdyIPuM4ejA5Vk1EtxvaAMGJaowkl5J
au0G0zjSDg/2alcGHJdg45r1w89IasJ3iyUz/TSIdiq1kOCqDLEx9hKqXRRN4AWO1URxLxrAvYBe
0nnZJgtPLc2tref+qlDbZ306h0lCBQmqc6bZ/dtqYxWTQ2lpvp4DiYxUBJ3m3GSAd/3CZHBsatr8
iegXzkDtMLHmXr1ajhAzdG8MyjsWyhgv58DifDbuuJ9dYOjbzsyKOhbMCofT6jVeINoJBwvqYKnC
GUTZdoEGM+ex+M5L2MM8sfuVeX9TISwxVfqowpmzscabvqpM5LLyz3JbPmqYVguOON2GL4wz00UD
VAt6lsNvS+aa0nrQ64DMXfHZKrK8jXZfTyipBW+MjPORwBP7NIkAlKjI+tsIrn+kjnP/WzpbsXeC
dkbqdLmSM43r+2a70wJOVsVKmQaeXmIi1rTIWia0WsSqNI938BY/7NN0fBU+gCgM5iDbOz+VXYLO
u6mu8+7wOqqnJF1nFC6NdTNum9XfNcofrA7jUzn+Cnaxa/CB/gH5LEzaU4iA9Z9QaDQnHCO9tqgk
yH00cwpOqNG27QfffKv6EJ1sprlbZJcGGTIpbGwsBt+jpFtB1eLee1Q/hSALZWQO72v3BYX9cKMj
1aYAzGfB6SRuKSSzP3NLci5fywMwLdnZ+XFUT3v5MdkxtlAxU125rwdc38FuYASGIB2KCLOR/QIS
oqGe+nVk6muhO5iBpVqCOXNjDi8KYqr3j77HNr552ueQ3bIpWG+7K9BL6q2txEu76ZtbsTioLpBp
5sGMLSJN2xVoA3QN1szmUX1CI4NEzw06YOI8Gsg7Qhm0KZejpo99M0WkUMGk9KWfU6eo481pRyks
YMR1D1CalN/v289vUTtMC+X5rAynJAUHUJHL0gVsAz1XVOpuxingrl7ykVv4g/Rtygk3deOGjmU5
2/kcNSUF0dwKlkCGVNJu6TYAw4RirThnqJNtGhFmNr/wIfnAp319zTYui0j2CyjP6EoMFr16FU0b
1BqYCNy2+STbKqRaqBU7SLSzMrY4jLj2tjVdMksMHe38Rarq5s/5BP5/siJrW97wc/hRt9HLVaRO
0UAvxzAPz4M0eYJBRtEQtLtD/jazQ4pyDiJKG+zMRKbpAft4TTvtLMveuiukxQGOtEv+FcBoK8U/
lUw8Q69xZ9ejj5fx+kIc4wSAEjNMn0aQt0eBWQ+HjwGsrx5AS7MoGXWuM1Z//ct83bhKZvm14fdw
gmrzhzlkHHfSk4cf2SfWVrAsDFwjyVJzu7CZOBiVsnx5nA5Z5UiVaWX7doUbx/haM09Dmx2XsBkI
HE6MJJSnTTR9YtNTLo3haoonX+zE9Pcu5cP4AEd/1XmCHB+ql+LgOUKXMdwFJ6zvkPWhZ9SqziFE
VpOfZQ7Qkk5b5eUOAfaCI+SFYfTY0t0CYpWy6UMlsU+ltg9MVvqeH3gHtuA5zQEp2fm3Y84s8rtn
tGGQnnZcPaQyjswEmHL0k6ogYg2kBC1x6VBRCmo+OIzRQuPdPe2iOS0a1zxWFiEJze+7ZwHQRXPj
1P5L/ROMB8UBwlBSTyj+xvm25Z+0imAm0z1fPq7J6hEvmVolazyOHWH5J5BSM7tLQGjMr9mGpX1h
gwQtQyQnjp0FlD6DJkF35DzthJZNIMPmZP5fz8jgXSfDhW/78E8Ft6mRBvO6LGEI2cBguzMr90Iu
EjADPIyoGAIeVwGMKf9ipKCTfGjWFaynLI7CpGnXMO43IEvnKqDHj9r3BBly7ohWPbw8uTg4yKnl
ipBSerwVXgfiDqkMotv/7JJ1LRtq5rRwlI23csTp9bH7Xka8Lq5K6xwT/5/DjSr7D6oS/INYgkku
chfXZJsVJj9LUHx7R1varOrFceylknkQm/3Zrd3lehL2egOHwuqkU3sRl30fKYnJH1FBVSTrvRuM
IwwUtuLwnp9I6F+iI61kKikxnd6HwqZNHr86q+2Hw95tWZgtfqyutRIXRdxH8vhT8uhXCBkJbYSi
q44DLwgJXBh6EjcuwKKcjLoRQi3+f1g5+fsfRwHlqUln9kECbq6yetVg1j+QJ3eZ66CzV6GoARIJ
mIKarGTOWVeEMbof2L/dy2mD2XgUaLZJFIuVomC738YcbwVwFv9lcd6LqY8TFz0Vy8wNUMyu5NXV
Zs2bjikk5o+a8NX8c1yPr3voL06OrSz+oomqaL+QU7pUcPovJWSvJqqq6O7/i1lew/36DJoGBghT
YvnhY2VZ8KGN0kRcEnIMul12cFLA/zp5088xYtGZo4j1ofpoTiSFPceVy2rAp4sI3ov4/h177v+b
dmxoKDcecYSQNHEqgtZOZIwx0a9Kst3PlfHjxe3F9G7a9xEqWHp56zCeUImD+wC4yZQk9Byl2eiD
KrJMj7yjuknb86cd9rGcCgsY7Bd/Z9D2GDa/DY14L0xfn+qzBAq97vVlFXLwTsrckXPe4IZtKbeh
bPXWAwN1jAoCpNepmzA2jmqS8+Mg2w0P97tsjECR/Qwplv4nFjdlrh5tAFQ8nay6kZ/hYALLMbRg
H2aTb88cP6eFnWAXo9gQd1wF5X0ywnc4lnRJpYDis2mPGLBYwUBNmZtXy/S5ehSinhhZeD63XPpa
MqDU7fIrl6EgoQ7qLgvybvk0PBOPcKGsnng2LAA3snxnImUw56N+U8YznBJUWso+PaT9db7wiWZP
tmWhKvEw/wDR6Vz9HbOjBpYfoxAqbuWkAhNvrNTQGmnukr/4ES9KsNjIuJwdoNligl8QW5F6W+U4
f/XutyNvJMHar+pG6BYxA/cVGSULqz7Tm0kzl7BOBjn20fF868039A4FDomsrprlpzc2r8xfo2eW
QVy+5kP2pr4r0L5RnyWIriAY0Z1T9k1d7TFZS2wG/49Ofi45FdaMYA2dCzVTGg6l0q2dGV7xL5eB
4pD4U+njIljHuPOyBZAkLXy6y+I8k4ohtXiM8R8Z/jPSjfpkrEB+tmx70LN5Lvc0HM5WHhbMY1dq
rYIyt7JgQHIka+BAesnrtj7OJdm/9UsnxXnuTO+5Sw/n97rETJIL1fSVrxRmwnp0N/wiaecPgVqN
xUE1FKeD+8kmLk9spx/PhI2W03IFd6oXJHX86tj4CZC7o+AT2/YwWH812eyM0KGVxFmhBexfHgn/
DD5W8VVBuiGZ7eapkYNf42rl6/hf7TqzXbuHZg5pNRAcs1TbNEdqVqSGeKsAlq5Tocnzg7BrqVD/
wu+Bz/bV9ZVf6DS7ERqHdIVuOBholLdhT/fUl+fyJtirBqrWcxSCgLYHqUXg2KJ/yQHcSkn/jB2T
NAmDfJ08tA0PqsC1BsOF5gtFu314IJBAOHrZxZ18VMU5nJF1Ny1vhgN8i7tSOK3PZaY9TgmtrBPs
W0AEZBKNo4fxESTjbpgPXARtr2Uhx2Wy2rZzRRv2Ot2MG0AZhY6JLn7jR1k/EhTWOrcmGUN0aH9D
taCBj+h+vb8SAByqIv/fZ56fgBKAFDIwOzDjJjNQyRqucHMm6vuvBsjwmTA3NRZnVlYB2Z8UI/K2
vx5asO8iOGr88Wx/74D6T3+8UvxQgpEEfviTSfeb2S14sD/sVYJJCmXnWR+NsNgfP2ybDyJomqlf
npVz2351PwNUDBcePQ0Ptt2mRUCXtrLUfSf9sCPH54tXM/zMKf0PlWvgMVshTLHqCTboaplRG83r
21dntQavQLm1zR30cFq2+CkkdWxugDqh0VyLqn1yeKcRgvZ+YwlGGsnzvW5QGZuob6qomfRGeu61
6bSqZb159qTwG0IYkIBoStWOIjQfLV2yJnrtS81rJESO8SOxnRR3JIUXd78AjdkOV1w2MeoIeisT
dL96E+5WsQzsieKMmlA7D9G5QQcAWnL0hRAQKKM7F6JulO/FlEDivbpfes32jcZb0bdqyW/BsMkr
fgcIefe/WS5PkDr7CYtwVA3ePPQZir4eKibc0XUlL58AdxK4fUh1y/6Hh4ikHac8huO0nUA9bJA1
+itebkqG/6yfkLsLv2SZg4iq8Kd4rwtoIDv2d7H9/Pxmx80kyMZDHNqwj9RZyMJXveRY3Qncm9Zn
37Ao6ehTXoZBVgWwtTe3e3rE1JcJfRXYFXUpjQ4DN8JtR8VXFHpjbrO/mUYVHnCHXJC9ACsJwavq
jUJgYTBOame2g0Xhi7gofmN/pMGMvhxo2NiV2evAotZUsXp3DD85t3B2pe1RDsGOIZjcHngQnZ/E
JqNsgqCpFykXgGmyGXP/yPN9eGS2CeDONBPnh4f/lnlwoAK2o8c7MRRnPfAb1qGDW9EPCZm5dkSE
/CD6rdW72RpfPLpYDDYJK8AhkyfkR5C2ANyzUtt+0KVhsSzEv1oNfTvN6w8l7f/V2mn9l9ntNplA
l7Y8twghZi/3jMgLWhhLF0SuPrJKT7GQEPlRaEVqkLF2xe4+mxF+lJuPOxBS5XDHh6JE9kRrKeId
Zj8kCyDw1wXU+fGZyQMFYbSvC5DT1hlvSiTjgLQv/BwH8kDJOU7N0k+YW44Szw9t/BZ/ZGefI6Tj
1XaH3y/fgWZSHJDgeGuk0J1j7tsZBbPMF0V3E0wqXWiYdnrmADwhgHEV8HhxptTiReIR6ZUq/fiP
7vrZRR2D/4t73iLF3O+Sq/jnZ0TBKnqa/F6gyLTw31x9EFOlevxrtX8rbA4V7YKiQM7XpEbtVKvx
QwBP+fMxWlXpEcRQU+d6+TgV6aEeGsK1B3QXMnZ8uUlsMz0j2kwhKco7j1EWccimWGDW9i/mo4MS
NVgA0UQkOoG21MsnK3op2UVmK8heWw9U7ghCD02BThisWAvpEgCr30+L8zYStWyOoJr1q6Q9rnxf
NAvsNrn7yITkVSlC71cDD7WBqD9BGtRzOcWHZXJgQ5Lu1T3ltaEmNqBpkbWh4SO/GsiEaQHEAwuk
5GVXiRzoiSnbDhRcZaOH6KO+6lxYnSRCNH4UaRX44ZeISa1Hmk+n5ww5ljI0PyGGO4JbcY59Td2U
jTE9fcM7guYHmQyqu41EXQGrhqesU6f4vbJUv1vInoVThFM+Ja2XWEP5BE4ZlaorhYMuz6SNZBlR
Zqqz6rjRYeE/WyZd1MTaRxYSoqSNInl/CbqJ9hHM8wZIrAijHuVW5xMSuAupqWicJN3bgHKc+jG0
HjPWD4Y/qkICJgvzIhtPKnxvUKnt/yLD+F1TSKE5kxXz76ClD4voBR8HZJzZZUdBtVHtEmi4sr7G
9molwU44DhQEgaBr9A+sOGK5L3g8BZTi/JCXYxKvMBCaGgookVoryKT4/e+lGuw0bwSslcsR72cb
+JxSBWPhN89dbTxh8jtJsS8kcgIZePaY6/O5sX8AI2RilbpEv2JLYdT59WhB1TozUDCrOXm4FhLm
1N6dbKesRSKbFj3qgkYLeI1aS8rh76om2UXptBLCSJIVtxaSgH2sV1OAkfgDvcdaGH2O8XzrrkDI
6K3eayxivctB4j/nVL3bzypIh/7sS4B5gkGbufVUXcse1JFNcUzwxf5OM66TDfbMZlY+NULy8Sfm
GshnDpkqCwDD3YSFKD6MDZE5mhODjz+LGS0nqyYqUPQsxxTuQAD7BpdjYywWnQWqtdf6w6n+Ywoy
U4aZxtKw2FM/0kMO++aU5W9FihNiwUD7Dkr+0j+M1DEUaluTpzBhQu685l2JpnvSGf8Vxar2sqkI
eR5YHgWwKapvGd9yK4utQGizd7cjAWjoqoF/5kUsyLVoetpfBsQUCpdi/s9ThJSNIawt5wTTRM8m
sBKhpE8Zup1cWrRKYuczbJ+ux72OMk/q61lee8DaB3UcfaYD71F5jeaBVnkpedFkn+7BxyVo+As5
ZaaxI1cc9CYcFpeCMt3uskQygI3NkpaLJeGzVMyhWiW33p0hIDexkL1BjT5e2HQY47+M7lNbCwVW
ySdwmMfZydkPdYLr7hoGgC/3zaXwsQ6ufQ3Jw5HjslkbF4y/wXNxOIC3sgcxmN9AV5BKUQ0XFdJE
VZPDM5AKmzRy0tGGaqByaH5+M9wbqwlNV50SBRnVh86fBjDsR9Bd6FIk/raCLIxzi24AWck4GFoP
Uk9+mQtu6NLqw3t1nTwDQ3vaon3Re6L2+dNw1NVZrVI3Uamcb/4V6YLvhG750OIA5XYkaB65qad2
c67FqAODpS4u3/Xf2TTVvNiMN5Kb/wVqtRD6o2U5g7skP9pDEdqPaB9heiHodCg/bkYnwC0nto28
n2Ib0eN1bGA/qIX1bkVsUXEl5XbnmswHm9D0rwQuwt0Y7fKt9ntbFb5G5vS7nl7ZrhQc9Lz+VbCr
UtF75hCLWbAV8WfeB/TJzm9OukbDqjo6sMq9QMj9KjDZY6tD6yBYM50F7kD4wnDUsPjU/9u5gpMk
jjfe6zQJqB72Hfc+dmiTFK2nYO4MAi3SMS9WiQgZWsmMN09k6WRe/CGIxqWnp/EY2HTo0uh4k6LB
wo+5N98NwNLtcyQHsC7cCEGLwT2gfvn45Z2v3LVAHeVaGSqz44QRAH820DEELzLBZG4j0lj2zp+o
FTLOt3GNRNhrtTmu/ZtUyBr8DoHlWqo2BWidE/WBrbTFACgB9syxaG20kt36YwvsTtCkuMWmOGnW
2HDMNVClIU/8TSWIlabzJzdi30j7304pBRRv6fzVG2AdkhiVMbHsK89rrfkyCS0xu11lTtn2kGLm
ObzlIu+xez6kArFo/N/brv4jA//L0CB+AxR6hZ3ofNKOna4fclsnPb0y4m0DiMupI6ehCzmwj9y+
RBhWGFK3Y7sbZiGghn+LSceLlhYkeh4NcB8DkAXO058/i8PHH6Th9vNOcDNUc5xwk0dSGo7jWSNk
USh5c12T0JS09jGUFvMcXdL6YEdEOVTazt9WVDH5Vb+JBOtYmvXIkdC8SvuX4GSCRXPu/h2SvUld
LJN5BQHjcSzeXD0wZO1XG4UpDACKBIngH0olKMQ68T75m+hnQgfWQGnfaNHFNWmzKQu3hQzk3y1K
yTlP+xxgbsBc1VyC42Rxc/J8eAUpQTfY77McuNhGQgU7rHAxGuwUvr5hgQD/55BogeWe8M17p5og
/ktYTDqsH+KPUOvuKh+0QMlEBwMvyprqUIXCoY4LYKedEP24GpPyGsMY3utxpls4aBhD00UdLaBi
uxA+xxhfNl6bvSEZB2hAr2fLB4nSkMg+2dPXZSJ6stMsmP1VIU7qHCWLZmCOindxCk5npiWfzLV5
AWb4FEk8oIMClMHgOmrNcf9lHUkDQLWkXXxmkwoBVX+ROGyUyKF7FCsYkUm5lfI/F27Ew/+sObVR
K2Y65C4MXJgzWaW8e5OtOV2SQpBSz5/KqlqT3GpJSNP72TXuuwTl14MsqgOSXqlpsI691FG2gfqi
+Eyu3M4/UctQBD0pZ98lR+gIvjeTXpw4bJ5TWKskEScPeYTu6oXet4AAyjIiI3Ua9HDcix36lNVY
bacidTk1sE1p/rarQ8sT9qjkbRvmJf5jDtGXP+73U+EzHcGbhN1+ezz1X6lLb3yfYhju5D9OJMXM
TslmUuqguCpQpLmQ6tD9ZwWVVDkN2SUJeIuoJVG4YrARi9IJQOIDi8XRIAuXfJ9SWPfuiECwO6v/
qvAdpZLLKEqZH4v8IT6AUhTSFuAyrc0IVeVF74geFjlb0YSW67M3wsz2DVuRLLvzubS917MoHlpt
Py45K63kvdo5csn4hLlmLdu7hX2/KfZLJAAZIgWMFQLSN5HKMyKewK5RltPE05Ha0iG+P4tlxUL3
kT9/Pmw7P+I8jDO4Qka5aa/oYvGp6+QA4XY0fOtw4nhTZ+0oEgMYGiE1/9StRq1ZUmbuCRvGHvuQ
bNOI0HmuZVqm0T2AeDpzCqxBWFoAWybOMOgOnaoFAnW5PFJ3ZA9n1lP//gZnzF37YY1EvwRpJu/5
XYteghV+JXRYZbibEQDwU1Mq8dG17gGJ4uWA8Gzd1EiyqIl4ui/B7eWC9Htn6sqEXhou5zO6/WQ+
+Xm4B9fz1HZimH7Kw0RZBIzf4Rs5QnqbD2sWd8EYuV93pr3hpuWfCUgJaXBBBBroBoPYNh/MGUwD
5zPb0IA5d75AnbmofeCFi6e/KuwkV050n4fE996iIjSpSbGrtpnGfESjCivse/oTSrHK6DKUyBKI
hyyO6CFdXJYMFMSn6jm+B4evBkIrpsKZ/eeFQaGZSfd4hAq2+ILRET4UisWE8KqAbVml5XxYS6Or
bLhUUDmyi3WCwfAeO+dkMkG68QMwdiBtZku8WfaTG6RVKDrJckGYzTYoAz2xqtT4tknfQ87TFfT6
0hE3ExV7FA1CbVcT1lZ0+rNyvuTAWIAxfkLDv/kQ8jndh0XQW7nIvhkFogeCesLhKdlF1v8kjbVx
/6r1vBBGyn1qc72fu9vX8KnugFYDZrhAMu7Zn00EsF1T/9rVODpql1YY7vQamm9d+mxEsfWJ9otJ
CuN4wTqzSFokLUJIhorQVCVBIEWB/dUv8JZBtssVtokmLHvPNoIJJ31Z4bfWNE1zHYF2DOYQtkMX
HrRAJ699+fbyX0Sn3fUfkZLOjWw/DFpDV+mv/1dfMluQcFBYGQcadT6IS2ASPfFiZjlpe8c8ZYVg
SEtVGvwBEM0PIw2UTnF9J33aaPHPsUnsmoLEmAtuUjV/+/OjMtKYU14mZzWltPY38ahf9H4OP3Qq
jyF71urb+MENH5nAuMppPUlxILn9WKflZyJTObCowFMMLPVUfm7b3FF8d20ZCEgkG6qzRJ3grHoE
vPhVthixvGq/FgYWOYZK8Gi5qRZvtIMxCsaoWRDMKnVoD118PFmoUNt802N6zTUMffjrM9MsV2K+
zVbeDI7eHbvV0UucM3m4G/EwAUFwBRco3ATzI7Fe8JHkuNWbTYMWkAmFP+gXNSk73sL+Mn68V2kE
IYlq3pxdNFzlpRB3inJZsusW4K9M6jr4Ng+wT3HLLdWemP+7YLyCulPpLfW0FwGXLuyXfF0socjJ
r17lY/N0pcDYfWBW6rGu3Qfde3B3X2DN5dYBx4JPZpz/woYlW+psHDpUGAm6MpsiX+93u4SiwznG
e+s2euDvuQnfIHjpr701Agpx9uEHHLzs06nPmLQI6pNThNe3UiCyMuUqIQmOuwXvQsxTL3NIozIE
ns9eyl61idyqt36WZcwsLUFCMQvPBPMyh+ox5oniQNdPCtwjuRBjTf2b2cTRDliSjdxrYFOquya2
fDGFaTsltQ+U0I2ElO1VrdEmPCTSC8LQRbfDX7gzqJNvG89MwaqI0ycoj2L7xQxboawJ9OpV2jRY
sZo0ofRwknjy1NkqXBz/TH4eajZyqWO4XQuxA0SVN8pfxnVmDumaKgP/cq7FZ0H6tEHXmFV2ZK5Z
ok+VU8dKzg5fGNXQYi3a7XHtmQyJgLAZqfzUg/R3xIFrat+Tri+VW0ajBxh7FL0sZGCg5M2ncIki
MDKVM+LyRcU+pYD7AN9xAHFmMfw2UCCHDNFbwmQYn/q95S/NiPEhXUA6d4JuwywnrBCbbUgOq9R+
BDMgOK/KXZr1o3dzwD623V/nmtxyG/l/CbUq8BxK3FvNjqrZ3IROmr+U+wZjPEZ9PzfOC8eYCqMQ
YIa21KLvDH1vLXXlEBYtdAjG7UwSDuYi5r5CU0W7gtLCTPBQrrEbwOk9ZiunHr/GN7VmTcvDhEui
u8Im5Xgz3nWx0IXBg1iRZpQOWks+jCDwXNTV5AlVkqjKurQSlhKwHGxRmpTNL7zFiFC2OiY3+oyh
XdSV++pO1o9uQk+yf/gsnQdJ72lS0rUV4sQkJrWMEGZqxDgMPAqXwknUQg2llgEQ0VBGTd+RYWeK
zwqT1QLJntqEpJEFgBDgLYzBt2cbFQ3kCBcWbsb4L+sKshXKnC5wl/0XY6P2yIjjTnXMnyoOlb6W
hEUuUveOfU45urgLZR+wf9f/zy54prktXmC8NiNLMmwf5WDFsUa3w2ObzP3++dkVamjvcX1m6Dms
zyTD4G0kr+tW7MigNpnwyYCoCMb6AdJ2ydsXv/g2Q8nUwSC0I9SBVJ+PQexAbwR8lfJ1rcXQKjCW
X5WWtFgDCOpB/MVl+E/UJV6HfusEtcyMAWONvUMFCdP6+FrPErkwyn0cKUpNjLlYVAcTszhNl9nu
4Q2oZNdAYCVQHMmDm/Dywm6PpqSvSNIWoo4JIhXrYuTNSMlPGrvvJpNnH57zdZPz01haZ7WlVbp5
6yau2iIjapW/VOEML3j/8VG0JmzR6GjdfiplDvdzx9SGrnn6FVOGfq28Q7JqqbZaqUpCq0QFmuV8
7O3czexaoyPFIIzaOAQoYra8gruAWLwQFOXZ+ab0x6QzstbBDNEE4Kyce7RI2upfB8aBRd2fxjtS
dIKezm+vmtgRjFUzoltkEaScBT9xS8WuYPUAvHw7T3Sw9MjD8+SVjxjO3A5SqtegxxvSS0LpDIgb
gswS4IvonzqEHUoJJH+7sB0VzgnF9qsaljikKjh8XaWlUlG60BX0LGxoipW81bwo39s3lUparGYa
7UcoeGjGRo/+Zf0Ph4vKXDZpQMIRGRzQBKYtM7BU1XiiFZpX7FhteGH64AH05pehZUD05Bjq3bpf
9mtOgM7EFqbb8hhiB7RIaczebiR4Kae199UI0UxrDB6zWnrxoxGfZU87EmUq0HDfMWdSq66vz2K3
Hh2fr8ZtWQ8OiJ+qgXODF2Pqb+4kj27vum50hyoOd0inzdUOh89uobyzIb8Sb0CCyOllMsEhaN73
M00MYM4VgTMnZdtGUU5pnJcWme9wGF3g+pCXidMzBfQLoALd8lrQ0O/sy0wm1QUQsSuVQLBv9S17
uCNs3nchEgAdlG+WCLDPR8SpxG5RCBNZV1OrOJe1BUxycMvG5S9oX+0HUG0Q7U9D8NUYDSdjYANE
kJ4kBfjexGaOYnCg++SveC373xvl7z6HvVTWa4bEIwLT8dQ/P1ERXJkHeh943Eah+2EoHhI918jb
HonaBSNUsQAnnmnARNaejDmzowTCCtBgZSj+y918nFw5KBAA7HQ3Q1qJAjcStu4sZr45pngePkF5
lJ5Tkk1m+xK+nxh7vo/g7vBlx4nHtu9By7BMUwJ/tvzdUEGbMywXDZ9+NYWO1FgdwheQexCxvCbe
DkiuU0sv0b3+lL0nsQhdauct3QnTZ4szZHSUSOm97wOVyPvE264xTcL9Kpti9VOgUQ9I25H8hT0F
MiVkhEUwGD4L7actBd40nw2dsuzGSRQTNl9cR5W1Uu1oxlEIxtHjSLiS4YGlpC3FlbsVz8Maeq8w
Ehe2RySNXo9ClTKHpTkQLg0gLOn9DJJS/wQQrcZBAfrlm+nydMmk5uMbrCsbZgmnm0oShrtu+fCm
8OnlJsQKenVahvu71iOhF1yD99aOyh4ee0gcnfUd8hBuJoiKb/80+iERjKkXp2Y21EccrLEmAy8R
WORnjAqz8mWFEQO/r2an2gc3OX3tzdM8+Ep0Dbzqfnzh3WHFoLXzvshbxwBbfwYSQLZBwhobH+ZP
AU72mx8kApZQN8rgpNCgsOiaVq+VAiX+FVnjF0IlfFmXbt7I22r8sONo0pd5zajKcN0if4CCECA4
7sKPnNP4PdQrfBspTDMlNqkMBHRe/R0ifA0pss1aH5EltHWtchBsFUS0KdMMJfUEQUrr7QIajakP
JqUuQFq8xPZBLM1QUei//E72412l7I2ZYITxtTzFZS5DadEZcFyq2zW7d2GR2BQ5wjmxeLY/XD8K
RiaUai3J8gCPiV803DCJE6vM6DC/nyUKyEE3Z29kqhMjWjtAiYrgK+qaiqn5hZjnuMdbzB/ryg85
9xiGx1GeZmDBj+Bvm0OhdaWBmXxwibK37AfSk4Jh3K0XHOKVpKqCyUJK+51+TYGRbHvIL1J1cDkx
74dVmjQoyQ51KJ5Fu45LafxbywnbrX/SIkbXHYbI4bXpSrrIbW7c3qaPKTsrCSWkKfWNAIH1H0g7
Bj7lcK6uCvzcqfJv8kS2Qabbf7bsZb3z3TI/w7WYqwUnP2b8bFVgPV5FaF2Apt9vjm/VjN9TxS+W
7/ovLQhSq7p4qJt+7qAQaoLYfWeAoXj8E/y5cY8gnwz3W8Ce43Ct5X1S73zrvYA5wTU5Z16hKZuv
eSG/6XyH03i6DeMNZWDgOX3LRPVV3ZbNuMo1wSaB8jEsov9YGk3/DwJ4OOw9cwcxJ3JOLx60PQbq
xCssNJualYdIiCP5Bp+aq4RMJYcj+FG8KtR/pXbswfDMm+TInUyh7JdQiEMYYfklKkWsDlWOXQ47
KYTJ1ointAJyUp+4rOueQjU2HhIRcAM1SEIajNlEzBuaehpWxaAbADJjwATllWyc2thNxfQTWOM3
VwmPVSZhOhRsj++05J5HnhUiAQiL6yWOFwwQMnlbx5EcGDx9ODnPMjUeEimHmesQlyTgdJfoKjF4
oEIhhYs5U2juigwZvs+Fwrf2yE2R87aGFTq723Tr7dGyYzQIrpKOyr3y6l4W2oghtKlwdmYCm9tV
wM4xjU6BnPre99PH9ctWIEv3CIIdcu5V0O1gxubg1YEEmlSfu1RxUy4AhtoiYflxyU8Za8HgwOMS
hzhOJx+Z910Rp2uZpC2yG/4KevvES1SDZxN8EXr+HcFoPlVo+n9iJKVTkoNzrQbFa4TQuw6wqCeA
qdv+uQxQuM1VSDFSsjpYkxTkaiCP9zx5WsPGAYWdIkRKHO1Kv+PFUL7t8gVqoEwnswJTd3LuV84W
Y7gWF6YtzOhTRdbK5W9MvF6ntYYLvA4sLoJdRr5RAz/9kH3PB/k8a/UM7SIGccStfDeO7qpZRSWR
qWADjilazjXWpFvbEFjohUo6fakq2d1uByDVoSTCJMvVQab50/mI77tAd6nU72nk+LUHPMoWNOny
8wWFCKa+TFZ0HXYHyRoO+50ucklRQ/ktcs+PgjXqWFjmp81OHwIPBTXKImiuVpfQNa4UGai26PQq
KUc79OMGZf3k+V0hdBhvCq/XR92vLrfmNm3gR7vUKtKBFhnOj7gbxAL1N7/UUO5uMSptYMltYp1t
6yhoNh6laBwBkRBa4FJw20B1rOtRmZnNG4E3MK44qIo6XyGRHuczrmsqzWQaGgXlSeVSvqUvCLX1
BOIn27iTSFPa4GiHKQRJUAs2b9FJGwvEQzzUXMyJILBj+cdtNX6EnO59ZQWulyqENj43+HueLL7Y
Zk72ToXgZfnerXodTbpqokFuVVrIV8pH7A1OUiOFoLS90lXDzUptAXocB2GccH3bMJ2Q1lRweda/
wncUBtNJkl81Q2FpaQ2M3gTY+cUPniv/8StdnnC5J27q942pt0vXll+Eg+vIKrmZ8iKV/OIN+d/X
Cq9LcYGRdiLMWzpOCz3Jt2bC6gOGmtp0Or44Z0Zvxa4EI+6jB9vSURfDIYwotq/0QccE5NbzXd5+
b0UcYm4+yfP5YglrKsGkcVt4lGtk01LLHokS4LZIwx8eXuwYzANhsiRizfOegOZWD6lsMFzjCX/q
pwyIVj94Z8aGwP7ZdXZjQe+VqwgVDY17vZWD8c8jJtECArS/hwWFaJU1EZoNeKXjC5fl05QEDyor
kFsgNORBUcWlJRbVwpgnoLwHsjbvPbP6On2LsXypI412aoTZQqDuNwUn5/MHCKTNRKVRuyaxXCSU
25IWHKOfJaPpF55E+5fi0zi+a/vqSbHh61UehPjaLS0J+eT7BtYZ4x1qmzxYNGqjADgOxg9j8ooq
IUD+3N+F2nweChS9ZpW8TeBB50gj+Ke/m7SYoRmSenTQ5LI7zoJrB6NwglWBuZ6JdCHvnEmx0jHK
uw/2xByTPOA+50Wm/oNf2fsc8lXu0cbHjGAk/BTJC1vZm0m13y9j0hRB7zyFTITI26GY7ogCWeoL
KYMQnS0h28b6uBUJaMP0Welk0/jCU0XgQGoSsdcH9tIjpajVuO5TFd5EuTKifTqIpTHibssugAYZ
sGwx0Rpw8CTl2/6gYdR8gMvGM+eQ5xFqD9nvTu06B+A9hTNVvXqhnn+mwTXgNXg9QIcqmqKssaWB
qnFzOXFzsWs+BpgX5HTXr5eu20NnG1E1jlYHexTmUugjXdCAcggQuz9ZBR24h3rhnh0DrkZ9oA+L
STWS4TxaqsbCpdB9rxPUESwIHD2tTU4lSw8ec075fT9ZfROJnQgHyKBeQUdtw65Ph8GOLrvvPdHn
OGmvMiNUbl6qWeYDoU2KTAGWtiBOsWzBN8bI9zPiaebkjTYHPuLZXBV6CoBxE7Y2HDdrPA64VMRy
Y3U0Fp723ZgcJJWItUWLwK/voe63rUC00quMuvzGjIuzYf/KI6YvcCA18fsmC45C3UYpaoSIiU1Z
LZwpTHWZ98C2P+M9ZnqFhhWjY1PPj79NKMOiaCnUovHB9/seyiF9ye5w2BU6F1oXHBQ2KRvttGki
iddpAKqQwOO3CRdfYc2GKFS9paNX4cBzhXogzjIR9Y5aWB2eWNkp77Zjx+kZWyoHA8eXBAZ3oR8n
lojp/eSd9AseLhNMj5SBO87FHwJEoVdYWVol1rH+UWtW3rEPiVytzTVcQFxwnqL2EWSn5EhHA784
5Q9GTYO5yElpGzh+z5rYKHwbK8jGeAUafgAzvC+Ix5LenMtQnDGbSArXJtKOiGzyGcgJvFIMdcyl
1y1FemJJ4F8hnXNgTrbEmM6SBqdqqcaAe18mEbTje5es/57vS0wauyh37LyR+PjF00iznQHqPV6M
/37sggQZXBl1Gd+lx+U1IC/7RwyURwIXitTfRp0b1o+J+8B5zDnkadLrZ3XrS1CE6a4vgOJuL8yk
Q/7DkPH71IElImxa8qzF03ekNIeJ6jb4zUuut9kAahLFZohUGP4jfmEZC9KHfQlAAUg4QtydFwCp
+dR1ZPURYsUcPquM3iSS1iXzga3zdCC9olBr4XX5+99UWV1g7MdS6lTw52/MjsIbEt1qswcjMkn2
98DvVoJHj8HRqqNgg8NbAeP1xMNG0uKSx4WEdzV7Dk2M6BbTkILCrJa3LNW7/ocdwCQDvD8WMpB4
hbqWADjXHeB4Ck5vVotdYQH7r/ppg8EArK9NQZZZsFhqIimQOeMDhkxjRCtnNeDG2+JDmFnOwWSZ
neqIFPdEPn3sIIf97pq1P0HjExbBz59vVBY1ycojb59KpUaN/zhM0RpSlu6x7paw5u0GZ5Irnimg
mYq7gxpMCnyBU2jCPZL2tFbr+xkR/c29yuF0DqQuR00ZZlvh6BdhL/m6EAV8hpkOyIatLnIkccnj
0BsqjHQZndA3wac25eFczpraUyj6rjsD4zh8utQ7Y7SkpvXFeu3ji7I77aZ3Coa12iyFC8qrkJtE
IQuncnHiFJME7nDB9YTdNSujbK3O/wdLMFbYBm1Vh0nlph/stXBa7MpHPNfD/1T+DAi0W6QxJKex
5foOzxnKESPH3a90skCuFhrniAMYrJtIdjfa3ECjpiJuPKJmO5filU9aOrIXpvD6V7XXV6HW9LbS
kt69a3wDKfuLWoFdC4NR1q5FzEilZ3eODeAGMoh+g7fk7cLUtkBfKR1A9Z+EPJk2ekpu0fuZBWYd
zp6/zXKfBC2MVvutI+1TAnQ8u73sTAVoFkkAFIMKO1DPiTf/pS0ydQOmFB7T6DZ2kBVoEZO8QPUk
853b9RTqoDnvvYdhpLYArrNRInM0x9gb65E5Ffzk/DiOMCRN6hsrrqFv65jkv5gVymU5HIIXeE06
npU25avoJEbwE/N7RJT+qwwjQsoujIffToqAvUYiqxdZmWPymuAb4s/G4cxj1A1BGxUomBU+SIp5
p1ldLBU3UMv4CXnQdAVojDYC6o+P9kcvO1FVQd+mdB9P79JgAvxRMhjnkXrm0j36aAcpgb3K9O5u
8+3q0bBErKvGLaQASzS2ZlxXl9dpjiG0YtQWiwQKTQga9Bsc7qJd9fSCtBOJqkT8SmjkzxKWaO/Z
L7y/9HscDk1qqxxgfUeHkdXaKpsOE+7+aSVCmRRhof77Th8fpMzaotfCUZpfFsGt/9tmtZQSyhai
Uc3MlkqUk2fKOOpOWhty0NQUCXA2HbBtyprGHf1jtu2RbIpnekyD1ITbOaP7yJIq88dGZRfV1cDc
vg0X8T5oFCfp5fIfiqSzLUcraWv8o7JGbbPK/3DSIUEby9diKQNwuUD8nvP/OqJCHGxQFzPAgGAu
WClB2vkTL1SH1/jDa2fdFP+xhGje9dNzx/Gb9gmbt26xWxrjbBybHyLLQwfffQqDOGYZSgc1tlts
+Btq1QdpECvhyqPllOPJzEFssrJDqNgqt4UXX7N4HfAKwvP4NcTiHh1hXhgQWsqcgwnSP34blDtE
PM4uwW4jVxqFb/npAQG4ZsfEK5ILRY6TfqaVsIMeYieGLd8xrYs3A1npSiisth35WEojaA7tKg4i
LaDPZlAzhPLryrdiG+LaQi70yQyKyXZA3XJXgm7bgZCwyiMBv6Y7wIJDNRkhY3p3J9gF0iY0fnXa
mIi5EQdvOjzJ27LZt54BD+1p7dSi5YPPKQcEqaJDyp3+bVqtREFNVh6iSRLvdVDbMCaPho9KpfNc
FiAd7sDGE7qYZpPcQrm8KnWqN19HsSRiY3ugWzTMXv330AC77HXEI0AmtbNcqdZdwxbIgPmw/xrK
aqT7QklHy21CaKNUtwg7gzKZUbM0ADxhi4DewcIHhQ507w6dlCSEoia+cAB31zrnvKQUGVCGF4K5
hdgi9WvjtVOUya7vQG8mxqcYuVGcL/MkZR+SMVhdPVieZg4hEZ2LUDsXvI6/pBmjw0Mv3I0NhJod
CQCpiJxE+9hUDE071EIQ3cJzGg0CTa3IFTtR2uj04HyU9LJh7gJrx0DNPPhk8pr0S7Ez27Oq0AJC
KKt8Vq2Er2TJJQBXrn9kH0XCAg6HkO8WO/dFoqsFC1cMmewAmNpJyM0V6csdt7Zfg+6JMYmoq/PN
ZFxNhj6565CKWsjHavVpOjMXEmqxb0QNz3K8b4pUU9QujzsKAlnbGDY0YDR49FNkWk7DGFAvJ1aY
R7X6RlIgw2SEdOi1ANOhut/tQS9m5FlO1XobKpeU+swhIHHyQpPOAmI5HjYednk8OZaXTU6VXknH
QIXWBR2DODkVD6Q+pRR+Sp9QDFetjfckEcQZ119kaPzGXieE8MMUfRZ47Dp/qTkrsvXs0YgO7eoT
D5clNab8lIpwxEQFnWceFlo+gf5PL21GKBHRnPpqMBKAMOa80xJsVwQT+NG1fah4tqvGZTuhLynN
HzuGwNBLoqoZ0lHKzR6gsCpCLBaWlbMkJWS/xEOjg3qEX/2lU9e9HMU/BU5Z9exAfgbOHEZrqQMY
867UMV3c5xlQewWvNtE9xnSeB+G2Po8s1h6FX1xmc4ov7BffAdVjOXvbk6H0gb3vDQ1K7m0xauK9
6zMLGevH+F4r2HWQEcxfcrsiEtxsh0uyCPGkCjH8p4Du2zI2ZTS7wJQMaT0PZx0nV8I4v0nVInx+
IVRMLKxdIos2+yYgXjsPSr03ZmhYf34QMOKIAJKJEqW/zjVLMTz7HpcymGMar1PKD1XrJ9TtlUVh
+UUWWzADmsmdYmGNKCPIfAFnf9sLKBYsM7zfnli8FBPwIUAwJfaCIgRZ9e0sy/7JDiDm1wV4Gi7g
mKY56y6ogsN4RLRw8kBm8SHR/8/5HgUXmodsGLKa5U2SiJnINfQpCb2p9gC6p+wOa9o4T2kNa+C7
f10c1MwYdsKzUMy4mgBxJXZ3U4UptiPXOzruFS1vz0tAzgI0L30LJ+FPEguS18P8cByklJoDAGBg
vyCPYEyomkgtiS0klx8hNXuwUsRLrMX9Ua/A0Z595yBkQsWT+uOLpMx2SLxQNX6DqEMsTI2UtGP2
CunbJVXoovVC8rtHLxFE+Ji4oFVtfNkCwLKIJwm4Ldx4Sfs2F32WbapcHDBGf6ZCmOVcm0Fkpho8
GU+1FdhiwQUEIwwf79Q8tpZ0Rvx9paAdP4jdIOOpg6bLlxEZsW40l/WKtsXqKomaJqQiHyNMpnto
yAJ/sBxhe26TfgduqBxybHhSFf6zV+pB+nR//DxOmM6C573UmFTyNAuoPyv/ffXe7r18C+4UyNyZ
rgZSuwMx2LcZxWNQWvvQR42x7PgURMrvc9alxt0B4wT5V15dkbxtvonI5TkEWOQjuuAg51wgC6uE
YpTTZIjQGIHZtBEO00wlSsp/DmmwKdtWsrRVlpGoG7wjv1LsvHYibGTb5t365aJe1H4Oy6Jgk6sI
kvsGwOVdkNOW7glHrxny/z5aMk53S9ud6yyboJM+N4/UPTluQoL9nR010wdsBJlV62eUnG+t6sBG
q27Yy2QYOHQiJPH6ONLZVdhryVrdZh+pky1uP76ajcW1M8PkS4bHzvmheuDCbv8e+JaojGtb2NCa
kj8v++BCnP9sGny3h7bIt8VIgMs+1xl6FqnY7zfrFETCdJ8hPlyO08EV002ys/AK15+E7+ktEoU+
TKdI/+a3ex0Cj8TkDNdYN6kxWVe7U8JTMKI5FvmW2FqY4Eu3xglW5OedQ93R3Vu2+x4nv17OJU7a
jXhME8jILUgYsx1Ork37ttlqYJ5Pps06/Ii1M2hkHNqg3UEVxjx14aGfWuZiQXYnNXVnR4g6RCli
Jug2qZ12Vmdl2UBEadSLtlNDzc5qIQh42e8j7xUFAbHsCx3gDGLu98dWAU/yWrHo3KiwuVZSwK2O
eQIGX15yLNdaPHtoXIUtsSbbjUPnWqYAYW8hbNmhrUUksqmJPoopQ3rbFUhVpD8vNAl3JKe7Q7G4
aiQGgJ6IgoK53VkToosAe3P9S0blFhOr2bIkKboW+bbfLArTC4nZkcMefKDYvXy0M/Y4hM5xzMA/
xvdEq+7ly0RUs9QvuOARcLWmENG7ziT0hSxbqH+AoEB/UGwXkWxczUhomCSLo1myzayUjJHCabjo
mYlhpJbIn6gd0L8Wa6fwJ5HC19RwCsnwaUwTymU6+40VzzPSByDJvS5YReHfeEbfYoH8NvKnwIHX
9Nf01PQZpOCPGV5c5N1V6yjC25P5OuT9ZF14pnuMvDcMEYhs5QyT9EfZc72AW/rMxUfoPIdDH7Tg
F2t12Ht+3Ag1Sto8vIdHvjMo3qlWE2lJJ5HIXjxbbsX0H/pqWZ62Yopy4LXMXlhxmhmI+8bv4SFo
vKg5mAjOQLRQ6WraIrPqR3yZhaPyNVs/c573KZ1D1aZ27WZtnqONeRNI9nM1VdInqd/qqwlO8ZKm
mqgvvcQr3njhCR/oVAm+3U6P7mm64xHgNzWs7V/U7BuxFkjakSF4kXZZzZ+EWCkS/PMOP2S29Gsm
RcUSlNTB80XCYQs0xq1RqYfp2wpO34liAj0k5XKXrjn1TCTjmY/L/BK5/HYpriWFEkH58srRvA2E
5D9pdvgb/ceKk3w0SroE1JnARWf3PlGIYZKviF1JUjGs7RaOAUM9QVJEu+sOW4QVrm+0O1UMBjRZ
tDJ6vp/8fQx6vnM5+TtYjanWugx3O6LlHuG1Ba+2pt+b/9OI0WikQ1nWFHo+CwuwNNRhQNl9SMeQ
QYmojhUkFN70KV+EwDCEYvngdJ5ZNKOho2SG7n64eIsickJs67MxwZ0yJvNzzGPeIBryKsNKTdUC
V2D2guHUm2vXP8y+2N0RRwOv5xLveS4HdQ0WOLXjbmKIhovccsGtXq49DYjfGvcfdrYcIA9MgqAt
VRIyAZugSoyxDdAmNqUM5ovNqniAHfRHdVBDRzgiUDmyRGe0s7cVwFFy9a6BRPAQ16UUuQgBu488
7PnMmeaJRYnbEt/uGLVEjNPBwkI05oyvENUXfEiP+QDvsxrQsbFgQDlJSXg5EjfQ5oBqJG32pTbI
yeE591yhIm90Wb3g1v4zDi2+nHjIg0KUmluxRpq7aGlPhyQSAZPRsibsPOEI6DkDe8DX98KjAUC/
OqcWv50RX0jdVsxTsIG/OJWB30wfcIWvn0BPnSLWUzyWVNso3ZE2vuGduk2SCd0/N9oXfm9cG2j/
RYFbyNCeVUepdx1jAI/ZrtHcioyI1GiXtKCJDk3yo6G9LofMvz44oKyxtm8xZCqXMQRvrmuq0pqS
xZtcflORcDD3ih4eGCgNvqtB2r656XPuWRrlR9ISHh6TuzSipnxvn4+A8RnMJrEjWDcZbmF9Ryt/
XOwOCs2shPZTFCIl/l94kGlXIH8p1JjRjxNyRwRJ5sqle4xmhhfxIjmns12cSMicsG7NCcFnjQqD
/e/SIrnWG6BhliubysvkArjlvsE03Fux+VLtEzKgZ28qxuwuPj7dQIxUhNM7gRQQ0kwp+3xO0CKV
8wfguKuyDD/J5tqJmRvaHkZ/BHJlwnNjfpXJx+DdORniRUa3HRJ8bfOwI1ZF2IBjljgmdNZPFLRN
bo2hMuWjJ4bvyTaw0XbyH/VwnirKxXItngYjv9D1ZNZ5PHfEwAfjttOzYLOKWJYkZTQtxEIYic6m
+jcGQXh9EpttBEcBTJiU9O4JAXPciRt4jSEiqLJ1tIUEbRhjm2nO61jQTNOqZnZnYUFEO5ODZHOY
+8JFwn+GehNk4kSEjblyXzy7vgfmOz9rLmpgHVzBFVYnvUaShTnB2DFa1RdxpRfNq3M/mEMIXH+3
fUrKt5F95ZCOxoJzmRz8iNtCvC/gyj/RL4DI0jCVy0ouHaCVF5dnRvUfThXyLUosljAI+SuEaPPo
a0iFWUMqaBn4zR78nNJmoQMg7JMOjLa5OCID7TKdmrkwJPN+0H6+woSsw24xFMKMlfh/4nkvGVdp
+9qubO7c9iORT2ynI+kyf1mcL1ePzktcOU0O8rKu3zmUSLq95SdbW8wuqgVlzd4o7iEhg2zEcIew
noaV271n8/0NG/XD8MRjv98ltUf7xEXzsgDTZuLT+0fD8N0nDzcq628AvfatI/CX9QdOSot+nF7G
B4VvcotdaMyU9fWyVvAn1U0jRfvtB0zA/4Vig0/n8TIiq8UvFDY0qahnDRNlx9TNQ3DoW/NzyBop
/wjOZwfm+mzGeBrwqQh7So3skDeJs6PyLF9MhcqYVw5isCXI4Ljr1MRAqHadcaozVUy3PyzRnra+
hmPxiI3uvACIwLq2NWKsk6XBLv7hQPW8ax8aRr7NgFmjR7/r38H+EA9LCyJGAHWX/9CntsDMXvmr
LrZqPohq8lGKzgnRdgBlOPMyB8Or9DFp2/Vlyy2HswkhB6NH0OW1JRyD3KXBywrj4awaMUgicW7e
8mSoQ+9sXeSWZMMcPIlWLUsUA44z9YBxIZWK4rmy0RbRktj0C0GutG9GsTtkCRS5TqUFQat6ShgQ
XmqOhExF6ckJZ2Y1eeMrTd2Lp//iF8YacaJv8nJ7dZ3k/ifT+O2eNECs/JHp7e/o9mZ+ZQ+CYNIf
Il0sjxtB7q805EfqHxlXNQOqfMl+qASWkOMnXPESOVkbmX6MULqvTTL6PdpW0KcivxYyk1b7FV5g
VfRj8Pz8Emz5Av2SaXb5zZmeL0nG2JMslkCWzRtQAMFk/N3EhIbnwHYV0MWOmEjqnAeoMIaLQFcW
QIO226ATXg3sSz52+vUKjDULbeMzYizGZj1Zd8KVffHWD5xI3n/fq5m6N4WdeoqDbjw8lXQ4xl+E
sHVKi5HDKBAbhPNoPH9mWbQtI9Q7efZ1Sypgr8ME61bh+O+fxdVvayMQ+idaUKNCpMb+6AEwTri7
V+StSLhqUF27naDAuv62z+EvfnBQ941JBqs0v73e3PiBuSVqPRy8sbPPSzEtbtim+HHRTH+UltD/
uDBZX8EHQG27QEyQ0fuJIiAh1SNpvnFwrIKkYcOH1h/N98ZNlsfrsFt7ArXPX9uLiYjUMAT2+Ulr
JVWU3H+FbYRsZ3B3ze4Kpa3rZYP0T/w0XRBjjAblmOBIeQIUTqyilOwtFcn1vJSJntDODv3KV1QM
uMPSMq6twnw+Hq2zQmVms84kNYUY97cENppD4ECdWuINJTXmavlS/w5h0YQsELoqW55dC7H5Jylh
fAIiNLer2vU8wg2wP9o74J1lZinVujgYduCo9BRQfLCYRO5OBmFcUqzh+BkmA3sq9zUC4KicpNJp
dZmfa7FMbKeuuU3YWgFSNaEB8XDaGtEIjP6BN+cbsC6J15d8MuGYnspc+llqQ3ano6ZdNmcRmlbT
ao9dU7jx6IGY2vJq1ZViiM/Wpy7oJFuHDl99a2u1PLMo0oi9W7UuQrKBjL9NXjKNRAril+FRo04D
H9tVIQdsOwistN/O1qMGzp3Uoi8GCUHs0oOYajqaymvn/GuutUxDk7C9zX99w1WjzqhqKphmY66u
a5fo8i3HvB+LFFQSJCFmkj5PsNB+sPozWdi9qqJJecOFFKjZCXustEfnpQfQnfmB7OZVI/rFBFZQ
cFex3XRbAx4bQUNv3EXX9hDjwnMxO8LJKVxnrRJc/4EuT1y2pqCd+QR1Qf3aQruB6xMVqRnIGVSy
yGRxI4toxWCWup2MLKfHYkanHyhZE/JfEkLFZ8qUEWExnzadnjZ8zaQDG3/F8HU5YPPlFhr6lpvi
faz++lboLP62dZ1hj+geXB5S2t2EgYV1WIYCCWWVl34vTcaHi1mIUJF5mP7cMZ9nAFZauq9IWu/8
osu/f9GgrSF8lgbz8v9myy0m05F5U/r/5ubYiIPwT8uaRqIm08TOioq11tPnLXD+H6rdrCOqdWsV
4NH6MAgMLiOaYJqdR9jfX7dlpMN+7bjUEo2a/1U24T2EfwovvflcbKPKBiwxS3V2qhWaPJ/MCJRU
ZT4WXLf1/L0EcHDYjMGjtekLNeIZgiW3kx/zWOJVMqurapl/imdjciYkw/B98OEAqD0y6UuBZNL7
2yfbV5/UJfq/Cij19Q3zLEJi1SdwnXK4zrRi9nA0X1foHiRVMBKPHzXjQwA7ILtfxjuUFIAImjkz
aBG4OYzeghyYtkUDpv6YwC0BF23oX+sKRxpdGCOeXPgjWYk/a/fPKlmcY+wJQfvX7nc874SEq/Re
ReyIEGw+G8Iitks9NC798RifH8+PD7elct6tWPMlDxCzYFyT9oRtvKr1zQTltCaWA9NZ+pNx9cLP
yRwni4BWBIqEnxlJBzkZPMZoNdVx78NnWFAXtoRgPFU1bKqiYbUg4XP20LZqqyEwhYFXBwPU0rxy
mgeC0QnGQFqz6uEpZZZc528vSMxyjBhhtPFb2x2Q6Nu+dOQY7zdc86yRlUOY/yHLEWv3Yri9EBGT
zpKlXvHJSqYhJ93wSAYqo9k4JH1pM1jIjqIu9ywW5o6J0Xp90dA7lTmcL1+UXNcpuBDKctRnkDVQ
ffLRarEiJXKWdi7kc19OfKG0Gfa1Pof5NKbUzBQ5Wfyb12YuSjIyUD1Rr0DGgPtrR/i6RYrDLqNJ
fXi4zOS77hGM/kb74SAuLhjIMDW4EvipxM1akvy/oB4Z7Vo2ni1a9VM+Dnrqo0Wa7f1LWpSmN4l9
/6JAbM6PGVDGlheKxko33uxVJqdyoVCYuFNNkT1nwef3wGjHCfNKNVK5yypGFrJCKzyXzUkq1Yk1
HcCxzL9lnxgX28pDiuYLgMsMT0/uwNKzzvXXDI9gzgCJjgLaX01NlNI/9VAGGcHb0zT1ithyiNcj
zxzqkQHYXsx/gz552xH4nOI94mUDFAIeqI7T7OLf2Q6US+IFXZ3Mb33XR70bH8w8XSqkglDmhAF1
hYWZkxd2x42MZM9saGEOtr397dYe8Lq4LxvDMIjBjBlpHrtfXNNq7k4x/lzyc5un4xl//dJHh0Be
gf4Qn668FosLDDkyj3FqKfSGNjnfVgzROUPXoS6fQKUIahM/eDUVr7hLnQbqNf9/7BlW5b9Yv8Bq
pjXcDsAT9mF3WNFhXjcZjg8hTa/TtIROWknYfNlzVATNYWU+XmdgRNETluSCsy4VuWqLZXj385Tf
iMxerkmMeGnu71ArZPuOR8uxnsL2bqHbg0zMUL9pnAVSbCBo8wn1l95NtM9A6RQMGP0Wx8pZOqrD
ZAj/Y4TH/Wd6y3UZO1agfNhnfN7yLgHVCFMm6yYldq02E3LHij4DYariXFB+mw61447Zpsl8P9rI
MSqXuL0bnkmNVOPKJOUrTnBv0gDv+e01bsBEWCrctFUHgLfAnvvTzXmyRnCA3ddfe6q1+G+rtjAf
vry3VBymj3QTyqLJieZfYYTBEKLOjL2LYg5eTlc+EnZ6As6Bvcsi1o05b8q5YRzQg/DdI0/S7hl4
b5y7nbneb0Kyv2Wj99ZU6VHLCRzDnqrAycCiS+hT+eidt5/l+Lgs3imHELLWyy/vAa5XKOO++Hqq
QC1FuAF4K95dUe+PiFHIBoXk5qvlkqdkiAm7z7ObPwv96uMphHbjOqv+p+wBxNNEjo8Y364xoxnb
RGZ3cwyDhN4IiFcq1Y9a49LgfdFS/NbOuhnQ8Qzj5VWRL3otq0PbMuLtJ9/jJ1+0X6iNBUpvgtO/
YbJgOM4GG1LA8LC/GASh4seRA+FIGplmWSW/OCH1q51dLKaqyPVtz0woJLWkh0p8kd3k4RgytJcR
ee4j+hTslaHqPh1HOBWRZWpIOgDVQ/0z3uOAMCf5Bo2nI1LQyFbRC+WOrY9fcDLrN+hSO0XZ2zbE
3iMyvjViHL+E5MMPtTQZrAqtq+Uy8fLs+3o8FmEenDmfJArU5n+ysm5a56xl8fmZBE+NJXBvOhOr
gZIw4BAyxfaxaR+oywZXgfHfew/PtqK3gdQ8PuvFeEY6lpl+/1zoqwM6Pgv7oiZfOGIBpR2BJ+QO
7wN2m3xsk1IntB1s9jO3I6JLcSShzvttnlhQzBs6gQwiQT/fmsWupAeJxS3CJWRzRnVfZIqm0r4m
0q2r9QAU9fFinnVYUGlrgoHigIv+Y/qANflhUJ5jH+DtCL7A8qUkRlfx1kn5m1z9u9BAcFmSMLy/
ICpw7FWTYlV7eqsVMGqurNf8ojxgp32rbvdX2d8LRtDhAXk0uZkAoRMKveV9GQtLyiY6m4BjReZP
RuLICT52ZirIko30cYtg55g6Iq7nfbLFWxu0MDrYQSgGeZdBbBCs4ZO43kio/XhYTpaPCXYNRNux
kmOtGMUeuk6SDROeYf/4rk/Jhv1FlxikTCv7VPMw4qqDRBMVWVb9BF8EB6Hy+eiC5l3y7gNCacxb
yz9X/ciJQfORNiPxu7OhpdMmHJk6tLYRrlcouXUXUt7xquKX7xhC6ugweAmK5UlNMd0xx3NswYul
WSWd7e0aEgm5PNwTUvKLfyGjWJdjHr81bO7SsNQV0lO/T3pwKdbT0gp+iwlIRyI0PpBEKBmlweV5
jKQfSV52K1bZZW8L0/Z4NFUNbfD6519woKuXzcWC1fJbOQvQjw/+ESpetQQdGU8NYX5nl8JjwGt2
L04oLm17PbP5RHjdNE+TQm7MR2x8uXrkk3jElJS5T6JheUkt5bvCgbXyXYMAPmIZ7c3H+iigx9+e
wt22TcI7cKoSLWtmO1Scyt3GaFNNi8Oh3BYnt0X2ZEpM93xgaxFKxwTFgW/ipAVVETs0hgDvJ5Qm
oQ7AbY2nR4o04qsvdHm1uJwAvJwT552L4pc0RdsIg7b6ah/neaq/OyHIjHIGbRC7ufnN9rURgX4a
XwM+I1T3TXqxw7B4ZN+Xg5adXl5y+pmbjU8KWXfLs1imp9KNfLg43k/hFHmcuN2cqOe6kGckA+g7
MiIu1jJA1oLSEQ8J+stXBye7Vco168WxqIxHZb4bcv5WqT50OFGcCt4q/yGtL7RUKIZsSR9BeE/V
HW8P++A6nvFdkDwprImomfLWDJBoN/V3/P8MABPtBwI3hqCk59/zKV2S+yaaVtyvEaOmTw5AYRjG
4qyikmquZqrfKLvXCUaDqxEjjL4QPpBE71NW7Kh0WWhfzkXzjC5PZh0qlop+UGff9/hI2GqcFdH6
pNvbb4O1EuvhY1am8ryKn/US1F/K8bc4ZWSXg8J8TX4hMOoA+OPzPm6PFEbdr+5qDA24N+ZtiYxL
o8pgcZY/q40OmCqmPu84tJwwJqdYG3QEE8ZwBHoS2LvSV1F2pTLxseAXeWDzPgtCZ78mYvCHlr3k
JUdoSxvwu2Y8xEeufWmq/XF5o2kVeYsebjM51IvblfKRWZCmLT3U/0OG+bD2TjfvlPreyMwH7YKk
KY0MOkBhu+LGmPxClMDnvHBQlXpiC3PK8c7oTISfwqbzovg2yAd+YDrI7URKwgVIbwRZXz7NB8C9
FX9A0vYUopqDbQ0XKxdBO7RQWxa6k0g3Go6zNqlc7F/fVHk+vjqo9HTpz7lbLChcJe0/qjyaAGar
Lo5hl8OgK0kycfZwIHNh5YCp0Q9i62/OeJXs+BbLy6+cYeChe0v4CKP0seuYv0wIKVtNe2/C6585
gku28v8kRfnu9BIMepmuf9/+GCEH74HQ0gVayJYQOfcFtmW7NigRgS0dOvTDnWjPYNnOZltdm37a
BL4YVmYrXApbbbQGk16qTyP5QIkfIPTHw6vEMfFitqP8gy0TjoCJy8REUnq/PVdb4UULNtSm5phA
sIFOXD5ye7+WpwvG1ZdlFLoU96Tvm6Afn91N2yzUVUYlpXyfdOq0NVz0m5TFmrFoG4CjVedS+VXt
mr8k7VsNlrSsPnJA/hHXAHhFW3M6IFH0O2PdbEwD154mnjYl9lB6XhWznQtwblQNLqwKHjCL/mCq
RoT+kStmjcNJOFYwOdSWphvVCSqm7mBk8YmDuxAs9Sq10Fd8Se/8+rImI347sQT6kB2H1pe7sZ9B
jsH3uKLUHjLjmk/aNSTnVL3fl+YQQ0cRwubyaLkWzHoTXsuYjMKz/OsWT39ooVTdnZICtMrmlw1+
A6VqZ7z1PZz1tKeI91/n48FH8frGE2aVcX9LIlRwwVKKkZMvK1oZ1jpTliB1jXSJuP7lCUfuTtm2
E7mqoZLkq/Hk3liyvwWBaPMaTr6Gh80/LYK4Ud9HDRA+ExcOO3pp4TfKpJnEaXXpCD1SxiG1qOAU
IB5jgq04pFXubOaiD9zW01iwU7tBsUK/iy7cDZruCG+pcVzeGtOcMhd1/Gzd2IAg00Oai1eTV5Zb
Fk1zqYnCaidVznH5ECUqdGKV5cYAQBLdLe2T00oWnLWABwnE5e9a3nS6U4su88jeIoNtLHofmGmQ
Kg5A9bcUV7fcsgV6RiIG4iw0mB5OEk2AAXjprJf9CAAsHZpfpSj/PzFvRWRy7N2qlc/NsBAjpZzW
eIKRg/99PbHks550bD7OVRXwbe4IJFRXsVFhbnUQJcHpNh7edUTtX+ienePhGRRBL84x9dBM8LZD
NZDNsFi+/IXqQBQpGfkRJsGyUrYDgrdmrAJe9BEqlQVujeDkxd4EkAU+0ixSyOQzVmr7d8exbT2T
KgZ62kl7QKvKx/l/dtnmOZ6tcOAIEevLj2fQS96vuYvYu5ACnJ8Q9UvmJ0Uh/QMtdEnMRYhhCL3M
ah2Hae9+xVOOmy6WBavNYB/VCZUATkH9YsLqgHm5X0FqCWSI1MB5nT+XAHLiRAc9auPkDxlWi5SB
knoHWawMJpOb/rvOxr1jQGOLpbLlR/EdTQaFxR/PBWYXDtmozSapShOJ2EsS4QsfqpbFmtjSfog5
G6ZC3R5EgYhnjDa5fDY06u8in23NYNbo3bvI3DQ4+KpHDghj7VHXMIxr9FhZj2sTKVk71n7pG8+K
6w/10bA1/nVpImezj6sROeViMbU2/HFlUuFuCus9lq2g6Dyc2f8aFEWIBdNq2uPL2XZDgxreVmIR
BfceTGrsdKRJ/d1BeTGhET/aqiS0f71G9TL/CeTBj8cvEFTtPBmwmTF6sgHmHo5dueFgLC/rB/d3
NBMH/42EhVYiq2soXFn8ddudnEf+dA1oiHCwBWosKrIGSoJ20UASWjr4RQRfVJGNqrLSlaCo6kIr
GupG3YaX3tPVgQ5OEi05RWFAAxmP+A/LUQvY4Ecm1UBYWrqzl8hMctyCQbcVHcDKUqySEKbppxpS
Pm/8miIB9WXP+tlnhafOJS8079IEb6MO9Ewf88YMcu0hnV+hO74UW0kOmsLBq02ObsV//WedIiOd
38SEwFe4wvv6+qdUzPLz2do9nJJ0b2uyaM6/Ky/2V5O0lhYrQs4MYpmaKab9Xqw0O4eQNiNj30f3
r3butdmU5vWhTgtVLu4V+NUr0yfspGGxhqZRrm/PusufIuIqUkyaXJGIKV/0w6TddWhBTjS3EwoS
2e1eN2Jf4YXW1y2+2zuTSBWZHrujy+kj/SMRrSsnnnJJN9FFD5HrL9tu4E6XFVrLk3nwYo5JzDzC
g9+hPnnSOz1tRDtaHJ6P1r5QAx0jV4CxOilRRGyQvURpAARc5t28olShGqwGVzs6JEnaf/brya1x
g3ihlyt0fCyNK7P2GKbYsKYijaAyQ6HA+LY0U5yD1jSPOzv2VQs8gZFYdUPeoi68CkDZ0opL+TIX
oJSdGPEhhhgo3lftOhUGhiE4T59iRZYQXd0tRIImuTNtqS837eGqcwAASupHaS0KG4zoaAwETIpr
0WH3EBVe68SI1pxvlInUw+6eW1VwuoA2FxBxf6oU6ddpy3cErn25GovTfFkDtuBcM1f5Zqpjcwlo
jhc0lj4T1NHYj9zD0Ohc3yhFFqc9sAcv5HM/DxS3mL8Zw2dKreOFu8k2Ww5yTio8kqq/x4nqpeMP
BKVhSQoGO2hu2M8Qb1qpIVW9EaAVFiF5o5U8x7U6/s5oRkgMI8ady0IpZOu7o/XT58ds2B0FQVac
3RGv6Cs8HGZHLaF5Z3gSKvn40Rep/XOh5GtyqwKphxgtboFzM0ZsGg73giQpIalm4+2hZBj9etI+
vN2BB1pFWmxlY0iEJJcQApSHmjKst4KHYB9lMe20E5ZWCHurWCblXIgpeQ3DZb9ZsOPYQ2R3M0DK
RaKez9Yws0ucGPem2q/EukuI80lwRspIcZ5gjhPK5UG7C1i8hISDnrLTF+X6f4K2KqXjLDPjdKrp
J6M8mWygXSCeKmvEUmASMazPDqMhDjSJYITWtdhOoSUJ2wMdc5VLYWwYalhHzufvWq+NBXawTjBJ
KH5N6WNFaobXbS8wdL+fb2sNdwblJrz4aKl0493WXrTWEuCwmMyPGUUb7Nzxi4Hz4xC7prGElQ5Z
Dh/O/CJzb5tB1S6meknmxz17oKDMY01Xt7th5+4eDXipPASQspV2yl55kToFUaw20qBIKaOiwXKf
CyndpWWEw/bzXNeEYBX08T01khcteUdwjnUUwF53l2u4p2qvLTCLlM0k4URfBO4OvLDEbtiFa4Us
R4yNYxWpy6QQL26+UGE7E6NVIS/bwL1DaA+ksZFXSf9b8HqDKW6ImNTGSCQpAiWsLXUryfEvRiiS
A+blVXCaYH0/EOTmUl+Tq7eEy+ygpcby/eJ2+fi5WiS5J3Q3WjwvP1L/fELDTqW+daFdfPn0zY6n
Ux1zjo/qLZP/hrFfXU3JfMLNclplfjvJHPFjluTvVIhXnsqfeWEPNJZB7RTlTBK9ybfwrF1EsLXC
M8NmqLjmpscv2SFox5rKNwyeENUNaiXSWLaQqeG3rJRq631wjIEt06kTitYzzIWXWB/Z1WlrQFzo
NcBoNJ9J2uBuQubgSBjaAi36dWjKREXcSXN/rCchNqNxAWli8E7+0ojxw9bUAdKD8phRix6TCUx6
ffHmb2vmSWW5T28p3gflcHHX016PgHhMzIR4MdKtfHH4JrUeRi1JQTv2vT5AIcNo04PI9jSViLu+
4dGSDPIL5jaHqz8OzE3zysGrgc8xSfqU4T5zp14hDGyS4ZUb19B+YyP875nu8DfbCPr4pVT4NTOW
PZaEYtS+1U6Ql3Nrki5VBEQTMuy9FRRBAQPtMIVefVXpiF8ZQPu2HvhfG3Yk8UMUO9WRn2P+2t7l
Om7XDbjgcvz6Lhs+/QuiUtlbt04aOKX5E8tSMJBHZubOxlQRIODN669e5M69UNAgrFoEPYjiljlB
f4FH1WMBY5MtgIbvPcg4AjpHWXiYuxEczwHFS2PeZZ1KBmGnAbZqRzEdreZQAj6VX50KrGTZM4GH
gfmJB+slvTqSpasrPVSNLsDtRflKMthHZ1Ira8whHHQr8UCNHbzgmgLit7Ta1Yx5ooJzGwwxNkb+
lQCRR1F7Jyvw/WqrhA2gnXvyjztpK+q1BkVeiniBKOycNx8hmdR7v1vwg6PvFkMh41j+fn4AGced
Tcw3psy2Ikm3BBRKK7r6qc0R62wJrVL3tKaHUcGbulf8sZiGQdf2J0ns9th3pYIQvCwukNbUMxZK
LJNEM6uf6fJuXMN9K5+T4VXmfRzzSJNmjRbicvVLCGfJttIsO4PR7LVdcUvQ2veRftlkVhyXpjiy
PR7nFh6qWGhal6cZNV7/PsqU5STQqe+aVXo5HxqYaHSabyRdKww2H4bpeQYyDCNqBC7rhv+jtRfy
/EGhCb5tVrScg/27gJEYflW+wbfFe534VsclSU0ShuQ45LsD3KELVf+1I10tzTUAmepHabtLDrTr
paVXxWjdWwLJ5rmqKnLIBo9pgdkfTXO7lNYpH8Dl2phO3UuN+60lc0w74pmlq/0cw2Uu28dULRSf
YyEmtu4pY91s6+vnivxHOJf7dWqujHaIc2Gpg+6ENuLtY7BwJG9khVuj6dKemgY562WDS9VqLoDK
QbAMxiNRNHOCY8fsKBtYkZFnr6IzJDi0DF1QpUdYig+r3F7YeLlzjSP+vIWXx46d9lFANzTAHUEb
3+b9w3SdvE6TCwMyJtj9TkCcAlVDyMPxuU4gS+rSRktyByqNL/vDMRGF1jBcZyB7er3jadlN23On
AXqrAFwYEfxN87X1xi3aAqIe+6t8uErP1iBbLyQt17Ez+PCMqdRRkHy4katsY1UfJl3jg9YmZRrv
wO5dwHwYJZh3q9tX+KeFoxDp4SQeVKXGY2J48XzEfbIyjw9rkVW9RH/J/Z+t3D3zmHgF0eRBIGlZ
vWDCs1xBmccR61KillJzlK33QFADsEZUhX99/Z37uq7YM0ZxMLQcLYtvU2BurYKHuKcgc1/H7S6e
VY0+46349r8U5FRKc88yJ+1jdmPnaE5MTlvaXlsojCd5WREfGMMOMqaZwx7Zv5QJuus5Iw2A0Z2U
R2/UMxA+RWb5tRkWpmK0Rk8/FH/hZHzjebc5kbgoN7LCkFfnX1R4PdSCZX6i/UdQryH4ODQ3ZzPn
9S8YZRdodutMics2IMRVaJN9Y7YETbZCFPwvGwuc+CNuc2oIqNf7SUrRLrmJIZe3yoGwzIrvn2Qc
dUmf01Q5bxPABeX9xJhKtFB/hH4jcFyBZPaNRRa7Yg0yE66U0Uhf9PsoUjIYHnqnbkT+R3bf89p5
RDVVbyGbELpZIj/uH5+rVHjaz8ErK5s/fp3c+IORVhgJQFY53QkdfN7SvciSOtQNsb3ewKFoPwKN
Eu59O19PZx6z4kcU2l0jbJ6USBbPG1+ua93wp4FTyi55fwQbs4eUKZYdoAPMMoXX2o4miQYv/WA8
FQ7lQSkXzjkdFWHYsNe1ITVrIxuX1dFI1MX3GmoSr2kEVTxokzQ7N8gtsl/rngVH0r8gWJGbPeIb
UE0+wT3IiWzzc6YqJAaWkwLyKrKyaViq/VMb42n8hbspccO62SOVX2/75zm3N4pjftlXqVrESCt+
Y5FOKzFQxRNY/rgzSFVUBv40ehko0bRiZos0C57csH1kTVNh/6GQ9RgGOMlvj7z2LknSX33LyGQm
J+lByYsIuluczqyqWW1V4QHVJo6499Cs9FKlo6ZgZMZPdsENV3ujQfn76G4iYWEoQgmIgk2LgTx6
Xf3MJqgKdDSY7PIImiREQva2/txBluG+03z9dQiD2MXVo7Yl47/mMGwyDZhOl3DjzDz3nEAAG4b9
TRpQl/FeH/2mRLEtHHfJckSfkKuD7sWcezSrpHnuJJ38yaKCyAi1RNt0dQrQu9pEhTjxmApnWJWA
A29tH2Urc+scWQUYQuPjlci6eS1t2H4giK589hkprVsGZVoBT0GvHinSW33pqF1LyYGXSI7WvBnd
k+UgS5f8KU9LijkxIL77Ot+pipPJlavIzU0B0bvXkYwDYRt4xxEQ1Fn4YLBBgZLxul19hLdADx4y
ryiT8VxAmt0/KLxg1G+NSST0i/K00lj43/GyXTbzcCkYbT5xU33UHQGotM0KQ9QJ1WS3mSy/PeUM
0HiaAm9ZyVTaJHX5makkWGQ9+MfqA5xWVl9wyYpeFD5O2ddW9iKg6cCG8XEy0iqHdPuy0/TQ/Gyy
BfCxPYoxJ3mt2y2p9RDHbv+orisgDMhC1LH2AhsyD/hBA3W2dfqvC4wM7qNciP7PYdYJOiETx5u2
b3GsRtf7BwWrJmWmYefMLlxIZOoB5ZhS9oTlu6eguj034QsxAK2qLlbRe4eL75MHPwN3Y+v2jiMX
mJXHguviEq2/jjXxt3tCCDP2sIijxaqZ4nd8m2o+/mKMQWDaPlj85EPyUO++W6yt8JGMMqEjMFtw
n46/VsgYyvPSja9kvzIRLyd6eEndndBMFA0iD1KzVjaeqQkWbqLzZOcH7YBNk7tMNXtWZC3UTzCm
Z3b6+ClqWZkfcn2TUknQ8T+R47/8MqE8k6bNrkmbQ+kOSgZG7Nbg61Ex641FhEx9tv/RRnRD/s76
2ujCbgged5Zf/qaGnUZdACKfboSx2nHjyfLYkCtNpdrKiUyXwiem5Y57S1/UP7duFutnw0neVU6W
zrRKvayOfHTvlQRfTEznYLLG2kABu1jgpvKOTna6P1aCQ8Io1GyBTkk7w6E504sCCwPY3PlI1g/k
8Cd0UJDx1MI6AZ1v6XSYKWDtxBf/gsF/jF9vDgVBqflwoqAcdZybS5GxrPgx4fbtaRVPhdmwSl3k
r2voLGp4N/7XZ4QX5kEn+Q8WrZJXO4QkOo8giiFsdaGTJazTlOJ/zVcf3YKzqeHJrP3BVBp6YCNm
mRcxIxWPVxe4Gn96HXCtFUhvAmu2O456un/j3kChfkdPOOUtXluyW7Fos7hm7GyHfnzs5SaT5uoi
2Cvw38NjPhuFZ1mEz0LdHTp8QWApHUrY3Bb38GB8xBrspYCE7pAfnB9M02kNrBCE4fLyrJpqo/e6
GvNBw/b1dYwr9HP4StYO+ZfR1DVnJ53+bc34jE5VHWWx6bo2yC178ob9/bS50VLCm7wrPpbV25G3
nlzsYKfTiaXCuBMnfPCIRTa1b/D+1Jo57+c4wOtl76ovY9f2/KxL2jM8cCaOrUQZJuBHEfkGZL42
DtnoDsVuaILPKtGMdmZv90bKkrIXYCcC5GE9Sy4jTviI48JcjR7HFdwua0CtCJGyYFAgyEQwOWfg
nJeoaqtomkavWS+zPTpqyTAA/omyme/vuCyN/sMc/2HxY/UsKUH2moUK25ltf8e6qkrJahtl0me7
YD2KTtwygUx4yJM5mzmc4EsYJCqkWv4Z7Pldv/zmFDwwZh+dUCif5Yoe9rUot7GAKP/i/hW7G/vD
fkGEkC1PrmZNFUXBB3f1Dzs36v5YQEa+esZj05HsAqIKcfDYwluFUsu8ds30Lvt9Z2hk2+IzPThQ
00Qgj074hZzk1T1cdAxrneWJC38kP85CL2HWB2fA/R3y5al0zRRdc+7DXLnv1gmKqBz+j3pNyQZi
+pyfCJpzcntEknCBmrb7hoKIa1Wdf1ZnwnzTeShwf9N2FjO/YQWzWKOFiYRvUXKPJfxMNr7WaiAf
j7WFnFAl/N6W3Upq+JvfpkHZqXVzKSvBlUZCi8yuAwXaw4Jg1h++bpdVoH4VXstjWAfIUyfY56N5
//lNKXnaNuCnPSs5m+8VYiXdSs5EYuyYwYhH6xrZx7nmWkpvI4Dkw9FxNxN3FRucPHr6dmtku/k0
ATFJ2F00fDiSUq/g3W3Xbk6yNEGeoQS8dYeG55L2MSy0n+UAgIe+X+mBe1wOgGsnbt3DxM+QFdYh
bsRcSnPZXG39qpCO5eeYvZfOskHGkhikSUIukPZNQI77jtLaI42LCZOGKfk5a1Emb3VhMfc1bw6W
ZYecGXs65tSfZS/8VxHOWthgiaqPqpR/rrpCXlFud0BsMcqdYU9XfDuh8zcqmoI8JbCmgSnR/8eD
NDcHJ40g1htuCKKtjcTb7NxyyhvTIr4j8Lu5sHLBsIUREmMQeOZGPFzQh0bi4sacqHUljR4gd15b
qxn0uj25DLDE9O4oG2WfSU2QAfwvONalbgu7iJEk97wG+fmN22+IqDilaGIrGtoIWH34NB/sVW7W
TqRK//k6JPSrNTw0uPuU62r6JYsnJPFXGSRVury/hKVjvrTzJrAdcU48ghT9hFG3OsM+d9QqVfoh
Q46o8h/DLuDSliNaO7gvfRGx219secjhX2azZX8f+1uMh4Ss0uBBtRO+C6aBG4CNZcnBcDYM17Nh
EkwcmkgAx+GeglyRv1KslqhS0K/6/4pag9Cw7/Bq3LlUiP//sxUrRoOKj7AR2YAnVrRPtZw9O9Az
q8TW3IYUUZS1OrgMnbvajvuQz2cyFQ+fXBewARl/hZTWiPG+FUem2d8gasNsuGab24vBNGY0AbiO
CHkFhHlQcqkVxG1pTw6QM51H7KdE1Qhdz/Cmc0et1tvtioDy106DDmnyh1kWb4GEtZ1oMocfcsJP
iu2tHrcvMgLw0xqkLpvpSg/mSGvmCLN9KMCNwTm6ckIpggdpSl3V+ZCpi997PQR6IeUJfjd300E8
BoB9BFaTrMf9bciZ4nd+RnEcO5oHOuCnaNC39WBUAKSjxaeRF88RK8Sram0fgQsOzPiyyhXbyvbn
TNkhVz7h7w023Xhdy4A08I6mdD4LtiWByi4VGqvsMzSjdbf22kMonWBf+jDebZ+bG8kq3MkvsPpP
sUZvW0+qQ8Z2rppame80cGyfjQsYzfCWlu1cp0XCm0LCTWydEx9S63y3/aFKspsyxO3cxhWLvqu8
K2KLjf40iJ2IUdbjWtjmvTiHnef/VsWF7S98OWpUVWvGBOKW7VrZ7uyEojM3yF2u614pFL9RS4gr
vOKYHHv945WQ3UN+ioWMJZqhvXIDXFfiRWtuXMGcrposV25mPyossvqynuekvmjIBUGti/rX2V8n
BRZyMxJO8mWZpSP3K7QsIIa31SUbtl8LiGrMPJ0bfmLORtlyxzOjzwafXv+HZy6uKhL3VWjdw4Qs
GCjBkoVNmgDzZ6+dyO5QOHbpqHk+lM0TOjC9cdOhtmIuk6/r1z4wk/MJLB0bLLT44vRFZhyt8yIR
5Bo/fYoPCWzafVKpxK9LXOp0Tr4Ih5EJBDdJKD0RmIArXXNJbMbF71fPCr+AQ4BBFZfw2yXmXbHg
E26nHs8mfColrDxa8h4g2EPPzoyLkT3y5YqrHFuOqIUgjZL5OeyYaKBMrXba96hI8WzV1wUuzDS1
VUNQ0s1kDQVS+q4HThOiXpbnFDElIqJz3D0sA6QDrbFggGL6HW6JQoGRJ3sodcHcwZqOJBuiZb82
7VVpf8Dv2Eu9Bl5jj3qXTzhvt3TSR9xv5hqPpAuQKwVIh+v94nuwJkTBi7LVjXt9yR2goIz6IZQs
byGSnFGhoj3sA++cW178ypcslpqP2Nffn8dEEYhbyyWw+g6GFb++Z3Jys6oJ/USqP+eAigAK4cPe
UOBc8sQjBT9XKNy879QpBNhWzFywnq1JPnjBPUnU9cagX5FrbCBC9rvhAZjdibMmWgDGSdomRHMH
kgyMElaJgcl8PROGNJyFm96Ln9B8NhuDvaAiPYmbccx1i3UdGPmtxJHSkUT7WUMJwXZe6eYKlDwn
Na7dvfkwE1iV0KWlCIblly+lr7ssFz2FtAhH2ncfPAw3VMCFghkzLdmCCeNE6In9+HdKlorReSmI
W28SDGsNxeowRjV3GTn51KZcavC/OXFakruuHg7VgRWA11810pVkv9KYesoQ2wt+NjVjopxVAlE3
R+mo72zv8B+xc3i69Kdj08MeSFdNMZTJcScF0ARRKOOSN5wz6FPWBZHDyN5t0GZfQHeR1+mGb4R6
uFt2Ex1cwWofZ6nXbV+uRP1OTzI3KFV5nUmBHqnhxK+cncD1RYnJWyHDjz6Fli4lVR0BJGT56VUh
R9UUv47h/W0rjcT69zB3aUVtCZyvbKRx86/S8L6MW7TV1bqjC4JzP4QGHMQvDSDwkBh0omuaaWlM
w00DI1DfGvtd6IKzAZz2WD9UWGTReblBzla/j9kWQ0zyeks4wMOPmQ26qTB01Fc+mPNYTPFcFz9a
5H57fEGsZrAEs36J7oux1wet70ycKQHAH5jDelBPxEGoNes3MtRVSOY/szKGxhc9p7DdJrmJSy7U
YP2cYPy81tSjBm39T0c9ihrixniuxqSRKOSXwdCjJo0PbmujVljqQCH0jfT8lvsubp/EMjGb/tIA
F9IF/GZOQMeBQBdjhqq3oUX9ME8gq2Gevso9i3fpquUGioT06dUXim4GIHYBqp6jgd2//s1hyuc3
sBnOpV26tQDJvx9izqIUEJag5gYIBtos81LgLisG8VKyQWdGQX8q/dWr9zDuywvKPbkeCRQAD17i
m9eJ47J07NJfEg9mn3uTNnz/09T9FQUZ+KCYycunA6dQs4JvzQ9K3UCInO4HnmeU+aQYzfZCE4sc
ueBfod3jbVwBIpbmZYbs+NyGiEq0DS+bSNEGR/Z+7r/pnRmR7+fWF43MfadqWMu7fyLUpr+vQpKu
5sBItudVk9kgUXJdg4xYFeDX8A/huofukaOoZ7q7Q12LKoJTI1g9FngMEAxBpgX3aprp9cFPT8FM
8YssFHxqDIf1anysBz7Q8a6WrYxDtZOnPTU1jHI71QvyebmS+hfLVY0UjeWekV0zqyiz1DIBTY/P
ngGmNlDJ9G9oHnWb4uqjNiVl1CmvdiY8dPVPklTW6W76TOLDDu7L+t4aABkfeePQ2nfUVRvheb22
i2M+b3AvXsdO0jPs6eGWuqViZocDhm3MTBgOmiy7yCgJoNSThnxLmMrliWn5tXZtxqTOVH65BtcI
ar3DovESOhy39M2m9rwGMvGC87yaT7h2FcMcPlrIcQFm51USLBR6KVLKuxQdnCCWPedY+PUwuJ03
4tiOaWMrLmjlcGMQfMUdgJ0+/26OjoSW4CSrx6IeJZK8KqiF4iN2AwJrFq8rzqhKBdi63ydjzG+N
Z/aHb1OnxCdGuLArefCIv6GsXvT1ohVF5iOfDQWKnC2g0FfJnDUJQ4OYJZeW307/1xVv11BhFOwC
ZkPAC9Kohj89Oz2WMVEhZUWnTviZT2Ep9vqWA3RAGYUQKCt2yK+L16knF3QLIGOGGrztC6q+XuF3
FdApHo4IMUWQtZ/hn/SMxXaNLdkXHIVjdOmlkG2P0ha9kvndXxuEy2s7bYX0fEMDAWjlH6dWKe6M
OXcIR9n4JqadRU45cL4ivG3cJLs9vNgD5jYOjNsORtaLt1t+wPfsM99/V2aCjIfhED+LvRyFSYJ8
DRM15Nme9h0IE5Kcw+Vi1Cc26AVbQzpwk/pP3eLQpvUFscthDqcpx7wgOFJGHCimIHQr1x50aRSh
dYmD6kXr/WSJtSEf6GF0UFQGzYqk1PbiLHnWjHqaQi/BZpZeCCOFNOzK7xD9s98DTPlMPHzgutN8
cpr58v8Rj3DCMQtbJCImKBtcCcaxc+xwjfIRwsxL6TToKDCGgmCRLY7V1ERdmWMpNYunyt6k+iwP
k4uBx7NL5HkbEDEo/d9ox1lGYx+/adWyUhl93NkDjUzNXn1USEVJDrNTVxC4Alrv//DsqhpUtu0O
2xDLkwJuE0yVVIPHxu+/Fqrf2ge0cHXuxuV5uIaWWzG/EZkyXYbMKeuOoGIbNuFT5ArT4+SCfMn7
p+CCdaYY55mOHIDZ4ddefjiwjIrGZLwi2kiwT9QxSpI9i6dgtVxfgvHtSVaa5OB6oIx4RJmj74S+
9B/9Vtl23EZFDPCUqaRa9Opry4hvgRYDRANAJm2X/3U66c9ztV1Pb0NO9D0TxKOUGlQig5XqTc1H
7s9qqrN2oHZgTea9FTBW5d6Wo8JDaysvA8naitESoOubiBSmdn3zd0qVAYFT/j0FmP1vLfXBtrYx
+W7c+CmOvVBOduubg25sv+mY1p0Bom8V71tFtADIHQ2ACewJgYSI236m//zxqRb6adkYgu2vHwWG
jqAqfSlGEW6WyPDlSDxFeI//bCug8WUQLSJFODJxtGyZlVJx0cPdeKo1y3RvUvJw5ssUadCYImHH
iEjh2eeByVtOvyJBHe3mtTIZwywTsTwIW/86RCONENpTCHBOjpEvuVj5tdrn6A8mjU3jMQLtsh+0
ZgBdTCVY19opWBiu5dT5jAd1BWturaNq29+eNyP2Unu5pyiFKByxBy5te51tGewm/ImxiyAG0SZm
KEbzDNOjyRiK//aBqNcMjXdTdkCuYfc+6OVJU1HIJGR3RRAnki7OPbLXS4MGxhbQwT60uBLQxbI/
XEGCshNyGoVi1l//SSSDxZkGHCzULEYiLwZA3Xk8AB/Be2DM13toDCYoULJE1DMU8nYbW8qAyDIg
8Z6qdcgBllFldQyg7ubcXhrfPaekZU3ACuQ9tFfbRd5eH4ty3zeSrFEG5Cka7HsQn6476EogNLEM
gehGnqq+G2d5/Of2ge3/wIVrBvDozOpFeEJzPvm6QX8catsXaDFsDVVjhuh83jnbUOz7WGs0mTlQ
DgKQPqsWNvpOGALzgi7ba/6RUyzcYhTtTwtSDrwD80SgcgWYrXBNK1C+BoGkRwYuSVWekmwFOfFk
7ZR5lOwGJ1RrSbwHCX4HdggFubntMTUygpQBewCcaD1YEbLrw64CGuYBozPU+eDuFAvsaJd7CLpn
AD9QKoKZuA0T6SOb/xxW8IfdbwzJF4yNAuE1ubRtpJnnWoSw4KIitT9qbdlIj7743YQrrTv02QQ3
+WYyNrbz5XVyzo+h9b+gZBRYzYUXs+0fBzWVEsV6yj4KALoXeSSfLd/FBzeT9EDK3pGAjrzUrPap
dtP+dF0DsLiuu+jm6uFPKyxivfrCZI4l52ljcAb7hCygT1tkqga/h8jJ73quyMJm4aAprFPunEaJ
HxP/psiaHWXlkFQJI4wBH51BL5VToLaN66139iLi8+pCTQy8mLokHwwUV08xHY9adnxPEeHzuZ8w
v4h2OhOU3kCAx3AAQYLnpLp2Os2umDD/lw1CpGWy1Zi0q01Ayd3NJCTFILfWMMHkSH2tTxIa2ET5
Rrvmd7LgNdX0cuJLAmFdBUE9sdCGUqfASxX2o3JMOnR4Aggch0YRyYZPYLDM/Lilat8rxJC9FNuR
fRPdRYWJ2+EC/AHYHzgrG3mCHlAdnRxs322GK0xCED/F6troCytKQK9uBEIz9F3QfIT9gIz7XnpG
VCKnCUQKzSJuu3E43JcqfdNlAJBmB9kdFRi04p1JmMhM6N58JetT+MM/xkwwluB+k42uYl9qzAGG
uDSqMRKJjjafJwn0LcIk+gcHZpU3siUDFx0n22hLs40jfm8C7U6NBcpMiAuR+JhAMVfsXjjN9URj
hZnFH7pYqOARxopSzm8LVXooN+0tK4jJZm1uFwNU4H+seQT1TbTaRds42jNPGpvZctKJquUxsAqY
Ty3csPrppuCCMzgz6blkLvuhlNOlQCEJ0fSsdpRP+NA1/5G/nziGAqPR2jehx336JR1xv0hbuRR7
6Zl6mDHIorhoslxgsx6s4kQtSjt2ZrvbZ2VOWk2h+UM/zrvtCnEY8WdRuclhzQYhhqzEA593uSoz
PHwZY5K8wJwwy+f2eM9xtECVi39ljKyT/BWceGdMbCij7rASMF/3QdLkZd39IvUZ2yelXqcjXUbp
vugEP9VHHFLRsXMNcJUFrt2L9cjMmctmleDPu3mCpskbGjYJpT9XOMIfxXJMO9OrHN+/jPVC8wd2
Lp/uzVZ/U7DWnLrmd/SqbMWOpy14C8QZP0iX860gkJy5MjvQcy0MW/Gm5pfuP6yN22wT5Puzb4U4
KC6CMPdwpy29Jci8FqhmcPf8hYGkE1qAJ7VPZXIxH6QQFHkkvEM8f4IuO+4KvU/QwSgOJJPer0Vm
PaFTDQx2QYDY2vQ7eX0Wl6zM3At5/7aAGqQQMspPaAsx02RCdjoRKRVDqghEjJEgWHbiXjZZiRTQ
ExbJgDx+Pu7kTeXRPo6mhRTBsMOHfqvyxP8Z8l7Rkc+qCLs8sqDRmAh3l7CL6jyVmRqOEojH1v4e
1l1zosmFgv/eaZ3Msg2MwxGS3lFp9IiX1ujCaJgnDkGvPoXdL9jGM716fu/7NSSKNUy8m+k1gTwC
IYvFzVYwxtVaRIG4Gqqac0zH8q/pvu1DyRLUp+sLvL/x3pUzG08xHVaZOo0rSy6QjKVtGfuxIQd/
huqcoOeVPZIhUgKiyPU79Q32wh5e+dVfXsof2InRDTYzGCWfaroMCVVmAyClJwGzPeprDvgD0oiK
hRHTFXEm+IsUjhvYDtSggp1XpQcpFqecwrVsTvooOaFYgb/peAnTgsvGfCEaVv/+9yJNhw3lBX7t
VXj620N7A1TSkONueBqiJQbaUl5Mb45vHC8H7gWf6JfZEyC7bty+Xpk7EFHqkMOZhk4sdFyk/xy1
IC2Ohx79i8btiZ1sGqs4UGG658i+tt03mOYPcmaEmbs7gnO/CAeCXYtCyDf83gA6bCfQBRAQxB2G
mcyx9twfDk67p5Yumus/2SntfJsYOaMZbLcg3W6ECJFhuvjAduZDrNxEbFf8uON1Fu1g7RSthmge
W89vz9XJtreocFPPHIhitNYSiq/YrrRQNFy+oTJ8byJj+C+lRHuTeoxZg3xYoG8UeHs8shCO2nx1
ygNc//h9l5U7dts9gkdvSoHNlQU7c1RG99UNXCx4Uh+B3q5HTm9ANOGU4kcmvQWP+XaiG20LOqOh
+p+CIyLEuHEc7N2tkvzx4Qah07EbRwChUQ7vJu4VSArgsIjOkyM5A3kO8W9Y94oVFZg4gKDfGKh2
fpDsPFaiy6jPhhlRcEp7fzB1yhuukOH16z8zkyYUp1lgKEF4UCMDj2W/hGyl1huZl0GMKQ3mk0aO
cIOoPGuVUKmteWQ4L2lWnkqoRYuXkddE3o2XwWiFemSbVUfe8U7Z5hVsNf2qEUWtNUmTfbo70AgY
7CeizJLcv1MVnJcUKv8Bg7LtQOXvNkCLSAswNFt7wYh1qSCMQgEnbGuYgTy4tb5nYRmkcUBw964D
9R8lZrLadHIo+qizBskJGFnrC9wMBHjcd1R1UyaSN8uQNR3nHgaPki/mLzt2zfdlUxk76JN37XW8
3eWt2VbczyRgKxQbiFb6pEwNH+zQPqRx5fnn6jaBOuwz81NYDEQ0Pjv1cBx7iSgjpdvMIUflg1Oj
yvKGA5XWpeQwH/cUXDof+k5TRvCSDAJtydUmUnEIsgCX62fR/ITnsnLNSj6viGXnLFjGIq9mZYyJ
wNMpJhttkXLxtfQ1D9Cm6x47rwIXUENzzvfi+GUzu8faVFNNYJK8WDjAYvn7ZYHP49gJGzFnihEw
bBkKV8lJKcIxA9Z6nuv/iMdbC5Jk8+owv3Qykz3Mwzicf9WbpibAtvIB5GseLuyYUAcxKdSOWDzJ
dBrJxxWgieusjR1mNWERJ6RicW03gq/qOZW8NolCS54sCxLC3MTcfqxY8OamCeug6fBvg2g0zA2x
a1OcY2CH1BmX28tHT5gfthJagfcmSJy8bMQoHwW+7V/hSII/Ev4xdWK6cQWFEY9CvXc/SfMUjmha
whTM8bulnE8j8w7FdT1QKOue5bGTuyymz1wxg+TYF61Bi5IKgIMEyPn84ZHYH7iWExmXmW7MZ3yf
vLIo5tYE7PkVUKHbhJIKrqsD4LO1Jsuz9ifXY/CDEAfZR4aQvcpvR1UcsWKwBk+VYPNdsVq7BdFD
4K1TQiv4bD7EXKh52zLV9YqPIEjamdnKQTgl6yNBp6WUl6I4+jU+XXZ1Q2n0QfZXNb5lioSs8XAc
p3OeG2O3v8SLlOrQUCa3tePm2JcPfe31OwcSNkjs0zL0tO/tNPhSONuFNh9uq6y9Ki9vyL8LWVmJ
ROHi3aEMjGJiQySvW4TNeHyqjwEl1NSJHlYgz7nRLCk4+DotHwHOYxdntKooVRyj4jt5e9hqy9n2
W007QYOouMv2ZhKvffMmUBIV47t0x89omniqYX8jov7hbO/Yp3veQkhZk3r9aORcWyu618f+cAE/
16QMF9fAkfRyaM9oplutsqDKBxcHnVi7u2s6N3IoBo1+yt7Egm/KE9sLe1b3bLwxq82Cr1KefkX6
o+QefePwTVMWrswqAuthgFaguJ8bCLAIw0it70ROKsxAE4Hl7i43dtYl5iwWNbWUgeR/a28YUO8z
ovuLt2Z+j1Asvv7Bw+GzzATRUq97HYxFO5yOjbI8NqgMyQA2iUetfRATAZPE06NVcw23PJ51bmaK
2RpoUE0T1t5DHuz36QFNhW7gCs9bNvFbakd/UfV1Uj9BPCJROlpzeICDkN8kTCo386LppsFLmW8X
9i6JwxIyIgZDsCBUI7A8zrp2Lr1rxkUjYn5BeXZ/Lw8mh8B4AQHxx/zWwR6SJeVmL2i1Y8k0nDig
W4L8Z4wB7jVCAiN/AY/0HY3GRmfD3wMqAeWqQzsYZlxPKQl/UT41EG8mP3pwkzNTvRXLlAZmx8aN
c7+AxWZgSnH60tw3Y7M3NfMXScUeBZTQwUWdnOCNuBTBwXMMmr4qBre7TToS76wW3H9xAoEx4vfg
1nlo4e9c7VRAcQ9tugxq5dcn6r02pPQC5xUlrafxNkmCEoCrtuZ/3gMvI9E2W69FGW0WDrV5aeGb
EoEkPjBbYSwp838i1wiT2zhK70m5SELTCWXGpSmarqLjKEROPvjyX3CHbxh5T2nc7RKYoB/H4zc5
yag/0UWL3lcRVp2a7wchZGEplBItqXSK/60mH7OjGXuZR0DdwObVmWvIvw5QsuVEdIYI365bgyj8
U9X5Q0tDLBAkUHM8OmXjpdP5xCml+mLGxsPhQ20qK0JRTm0UeMCN6YXJN2SkVSJAdaiPybPdN0Kq
UIK6HOB7UFPo39BspNwAcGdexV2GjxBHMXs+47hWen/MwzB2nqddj/wKN8x1VPHnJ/b3AYSL6pBW
urKZmipayPwPEq3p4FZlmoch6in+Y+8FMlZ0sNv9ny+Cfanir8sgSTvG8R0M7j75CRzFxFIDr4Sd
ApVPSsEL4+GagahSqdmmGgOcGkTKpQhCkCXFboUe9ZqJIDCtYIIRURFnNXdmkMn6vowyPEHG1URd
dpAGsGQ5EYNLaOzw8U019uFHJFXh7DbW8ehFDCD8IrTFpsRtA4s4kK/FNSv5MQVmAv82BWKQKAwq
Ts6QdNP+0bxlh2qqDOVrRzbWO/sVFvEVXEzJvO2wFzBIlw28nc6DWUqE5lMjN8h6uZ+gIHtTXYtc
L32RMo2geHXgzyfFxQ8DFQTw4SFfFTJX6OhQEXhFvrMfj8KrNvVAvcwEGPFYwG0MdCF9S3SgL4m/
w6UOpFbflghbg79Xat/y/s2FyzzHExEe2JZty+yR/SNz+Y2rWvaJ2nU6DpcxBMiEMOkNO/jDpON1
GAryvnw921lWCzRR7kQuFknuboclLTLvLKi8eGnYHThvFac6WN6SgLavaOipP3N44/PIbcK5ZuPv
Oi+r3aUGnLONyN+wVVaHHxCePsJK5xFmA12SqGS4HxMnAK4+0+1ABGpBx72kzYavjfOvn5cLX0en
DxfEzqYnXIrKcSnVNNH3kFmSK+I0I1dlVyQ4YKkFuBXTm5LLwH25S+Dr1HRJREdGKT9ykjBjAok/
aXUTH2nUCvvivq27TZ7CB0zmHzCXgYbRc3iYMIBn3NLcwUOeC5jJkYodpCIwo+IL+tQAJ9BajgaU
0A3BBZK6uRAXu8qliJ+HePqB2AJca6+esq6ZJkZUJQPY7vkFkNBJ26TFhZHM1k7QQIbpU3BoD5/t
zvvSpU0sItIgvv4PMP0Ina2FNHckHiv0p/CTVmPF8JPvMW+wz7c0FpyC0v4JyDh2Gy+S26ILqnut
5bIStwgMUMVO58M8f+MhOgYLeKwqNbUu3z74BoZ0aPD4zXu1TDLOhIyfc9E5XtKc/m+ej+aDtQ5K
1Mjk6Yw0AtB77ZOyYP2lc3SaxcUxauO1dRpgfCkZDxvzmyIzrxjigLvVJcedViaZ29WdCdeOt31m
x5MjBX3PlOlY2pxdTin3Sq+OIIjgtMHLbeSwt22h0QtlHlC8bxlh+JXc2o+fhmYLqp6wnja60gx1
1bKLwFCUvvUj4dcQ57BkEYxt/4yfyetkMBC2v2JckqBZq9uXAx/iTC8R2fj4aeei8LKWJytf5HxK
qSrr6rpYww6bGvgQvek1Nw0mxk9zxHewCfmYdXaGpvttjp5zMqANmCtAhM5rKd2h0/1q33mNVssr
MryofoqC4AbQ2D5hTGRl0Odgw9NJlA85SZxAFIR6pOEF24Al6dMO3I5SSK5pSGa104Ow1YmXK32b
CzWk8oNYvbW4FKxqf0J+8MkJ85TduGCtaReeec31xuksPQjShlBIINgVXTA6VGNla8gPbexcaxIh
8SoHvUMIFHizQhczz0wop6nVzRXi2XD59eyX1d7EnvA4yEJf/3gIwa6HKsyWWItG5ohUJ9NVHW04
28JcX5cqkFfDoX0Az+TDgfmM8rRsu3ESBOQOSyK44t5Q1Z5Lrqh6bpYwBh0bfsmrObQddsz4gRTg
bdZN4jZXlN1RjUI8i2id0csEFkstYstU9oteVCNV17uMkYFdzlG6HFPgl1fwBm2suFOvngA7jNzv
OKOfrwb8JnIT72XkNIaQQ6FpXQQ2bb8IVc8ewu9t/GodsgZNqw7T0RpYw7vUeWbPjBukRFePk4uT
8dvtPu9g41ZRftWkwvI3pz+7apRwBNPiXsLEovII2mDyBJq1+MpI0Jc14/5fS7gxq//WzrtXpOUV
3eq3THheIFRTl6Ht1ueBBFuApJHDo115x6kJRKQUxP170NRoZNEhEfw9RbVHmPpSFXwBO81bZHEB
PTwzfP4n7VreSJkTTll9xNGo0AQWGxKrvdPMdyfRMHAusqCgqyb0C/bhZm8/R65IGsNwPOCE8bmD
JETCon5Xk6FGpG0272KEi8bhqNTveDrGUbSv39+lceAq6fAP8fs/DiUJmNcHeKhHwlgQ0AjmeJMv
huEH+Mmmhb9TpubCzZmOHfG10qqWjf7I5wUB3GU/c9+PZvTNjSq46WOgWJ/+6mvFvKA2YHTYFt99
dGNRCJ5njeCYgLLq8Zx001hHEkmxRN+/vBtwlACzdj/hM4ZBFyfBuo/8W6qCIZLpfV03JPytom4R
3Au/DVoGaRe7FnyjFCBKelTGkEzBzf0X1PmhG0AownZt5jSW/HX9CHJR6sOOX/PDtPNNgIB2EGdO
fFQHUhpF6to6RARbyw6T9vJ13tV2FpeNIHm0GrjwtRhCaa44XasdYunikyy2QTxD3jVRIyDZH5jP
KMbSlOI4osmuE8Gksfm9ZDH8g6Jfn3i4trw1a0pX3dV3kXaraCKUYQVZOf6hDtky68rm8KWZjRyQ
dZz2Igezn3A3cfo5u+2ctktHcgFOkkLEPBeqToGiHx8SilAsB6YtUmBd/ygewqxDJ0KCZI5r52XN
9KxgFvOlUca3Nja/bh2ecVKF9WVRdV4FlNifRdZvcNbaMz8nx3pXmUvErcl8y4QLpObn8LSfZzRA
DtPiTd1G0IsRukDWnEd0fiaAzlEiyZJThCgwID9CqTh9QYD6fvXxah3DQ2PiKZTeAt21/Pj8M4qm
XJm/tJKbP7R/OcIeRFbmVVbVifbcLsD9T6cnYHX/VDYpgSlttdTI0UV5JF3lf5xPs0V6CmPekBYW
VXaBZ24G/rJKI31RJqqMX7ibkuiCw8LYFmNhwMt47Iv5p/qO5DgRL+EfumLgvw3Sru/sXsJoGxND
7AvsJlc1OLndttWufzU3Ym1zZEAvMkQiuMdfMlRpNm3eHkaKKHQGZu2n7xDgNVoJko136DevFTq2
ysD77nlL1jJGZV0ptqXi0ekm1H3ZMg8IR2lxiu8MpyskgvdBFEtx8YgLPmWhKBm46DKbWc25rrbD
S5UkMZJLH34bbTI3i+i6u8z39+jVRdkqUVVsENWHyfLsC5w0KINZzkH4n4oy8R1GCOcx7J6cnOzt
c+LnOYKlbqr/F1bAiAsQl9ZeuRotYjmRU+k2Jd2aa+efZB9TpE+kIfpiezm8pwXh40A6TwYKKdMY
UEeJsurCSnEicshrQU9jXse6lldfu/b6IT9ECtGBXPjZYXl1W+jMZIHeHtqi01VoI7gdKIVdX+Go
xZHU7R9nLG9ScWUHfmJpkPpQLyOuacmNXIXPX/fUmdt/zE4Ga3DwGkckn3QePBiK889nMohJBXqn
DJyYIAjgWPW0BmxOlKL5en/C2ddiQ0vUjURqT/mQZ4DQByxBqQOlU5b7SaWrF0LzWqYnFQVWqel9
TngwASvCYW5X7UeX85ukWvG5sOZO5v3D9HFBUclzt9oVxEVQfa7xhCfLpc5yEm45fji+fA/+on9/
aNGp85yeokomlhte9/5JDO1cIWl5S5o3GEIXGfrTgQKE53QIiK+JasJIDOdna8tC646Clp0iVt00
tpEVBGkDTxOCD7e+/7mcxop3JJUxsM4g4PJ/3ICYsMMPelCUdlgakqoFiqNOKZDIYdJ1Xpcg6E7P
DbcID/ewvHQIyQTtpJx/bXFLRW4hYaYnHzkXmwudrhmLInVPOa1lA34uTHnYd0jH2wEF/CdcWdAM
2Irrv6TMIbJj9HgbYqyPlGPtGIg1rhHhN4awmD5qWC7+F7wC4vR3yYytaECfPhdubxQOAFtlhOvQ
bHejSJBFHXZXrxpEpzz21WovvTS2n5UQ9b3ENPzetgjm9sH4c0wlEwMQaq/Z4pVOn/8NpMgzbf7F
xiCZmCNEBhEvqvFZ8FJ5eezAtPId6FYm3Dw/raDf5HDCEjhEw2sIQIS/kP4I0uG4vrwNXn1Bgwlz
ylXU4uhtDXQ7MHArKXPpvzphaTQxzRQyEyT5KBC4yHUm0NE8Hcx8L7AuebxG/Q6XJkrKTjRw9bNS
z2NILjXFqxbwOUOjQXIA6GyMCnFBAcZ6r27ek6Pte6bQp+NfPWmRvyHVhrf5iFOGjnAD4e8Rl/yQ
Rz6NL6zGKgWqoiWxFyJGPpCPhAU/tc1eun1BQIPqnQH7Xdul5OOZux6yQJRRMQ81g3HcLNU+/PPW
EXT/JSlpykUC8BBRZlkL35eB2+gLX4aADkGFIwWmaQsa7vtj5mePmNrpo8TZkWTALmiQYY+bFi36
fvSSz9Tk2xoarftJq5BApyKTndfvLN/NM3PkivddKHEMP7aR+eLPiZuBzjziq8TDeaybfQys5D8f
FTOMzL2wDXK/LkGT0R4KHukMH+LzSaGBvF0vcuGulIJGihN6K0rkSE3BG+ajz8BcoThTQapqS2yL
ss1GfyyW79n1T8Pflq1zOrLhO5T+dWgItRHahMphS29oTMDmTWm6DcV0TGa+gxJK3zL9y0DS58fm
WXvddlEBzph3gtAJVyzcmniqDgOyXYXx9fD302mLdTM69A5Rec2ufz3s5mhUjap7glk+6qHXy8rC
wsrjHrCRW8sfjORzOYrpEqmjKpQHQXxqLhkcRTGVCSucpN9Xc2Wm0plEG36cVZ9+jhJWswtASeEy
/H97fL2dSKcbt7Rx+I51aK+j6S0Op1UidoeP89bEb38B/EUMF8K6ujK+X7Vym/ZdhofKrWY68/dR
A0Y0vrrjI5rGnfv1AHp4HOnucCOY5LR3qYQ1PjIpEHp10HlmccZ/y4NAS6BjOG5hBFjcJywKJfVo
UELXEpmqyyjD0XloQ9Z9EvMeBmTjahgQ/YdK8h5aTY51Vibc+nVroclv7DV1n8+yEnHBbPS1azqH
BXgHctyv61YRgRVIk9B7st4dJLmHveoC+93Q/TS0t52BTErbmvrWiE9vjL/jO9avLmNwJ53Aedp/
Gfe3L6grh8rdRmQcLIJ99fkLNZlxvrGWwQCAZwBiewCnSRV/spDLqJJaEdu6EGSKoczdytAZ1w48
t7XoD5Npxv/XLotLf7ndZb5qo+9IQwO6HjNIF9ZcBbpW/bV+PzZrl0VyZalkdJZ6VmLgSqb45ehH
wj9GQ/j1x4UgGKsLKBZc74Ze/+r82CnIdsWt64Ha19e1DI+tK7tp06T1SxLhPdGdpe95TRiJ2yzv
BTo7ljo7MMw8JF2N5i49vLX0BMtCWmMehkM5Qr2fHhesgWBlnX2QAige+HLNJLu9drNlhGaPOMuo
dwQUTlSlz2gU7VxgnoKxPU1xXVugkK1m8qM5m0NkCP5cnazipst5IqGa+nH4CeoKpH85Fu7EtU4+
3UvGeKl5nWAZlT49yObs7CIPFoXDoPIFbtYVu24F11581LZ8dt3mxCTX58aVMqPHct7ZND6pCudo
qsa48Upen7Do6M3JlKzOp0/f2YU70rhM/SkvDH6nbk/bFJaJYeJ4fHF3iN9GAZBmgCCW++5MNHyG
xGSmF+FkyiokmeDEBK3duwU9Z81Z+M8c98f4Z5GpB3gta1UrIAFnnU1oNVZ1mzhSlL4LGEJ6iBEB
Y6DkwKQibU52Vhy5UX5u1u+H/Y6jHTynDPPo+z5aqz8bTAXXgwFmZUys08CipQM1Ni24ATDvJLMX
gZBUsN4EQEMNPgLwSXigbglzHxN0pAnl6flktMkaSTKqJUovp8LlELRKnMJv84FPl24XGOLMuFmd
K19NAIbZ26JXCWrk9hKbACP83aiBvO2iL9X+tCAOLnpXdONFy0dgxVIZHJVZVhRMXpR0kI1JYQr4
WECtbr9sKwi5bXhF4NMnLjUjsnzg+2KEJs6zbTfty7hIshAwu1UBzQ2FqbrU1xpZqUFPE/Lat5Ce
GCCgp/AXLnUD47tH8RA4NaQWR+oR6SapI7Y/Yc2g2ubogJ3VOvPiuJPOxUCSxUW7peQgZn/DbFIs
y5d2U9eQju4/uDVMSC30/uX/kY4PObxI9wCKCwz8n3Uq0kpOjaeH/Z73/0UQNsXJvimDsNIZiQAx
K7hm2bxe9tB5GUt9CY/7AEZ2LDjA0DkLqW9EO51WQtfmbmiJL6QdZa8J5uxPmeb3DqcHbxyUrHG3
OpFb3d/rEm//GuS1PByLjFL7MTqkCkZZZSkMHxFSikKVzZ0/fSEA/9jDYF00bjxv06P4ewAoPYLC
JZkg12qnZck61iM6pbYT74uXKeb//zWyJM+GLOmvYp9bd433mm14u3Gs4hvWbkpC7CnX6fH9Pqt1
zjFPEuD2mabGQL8hLQnBi4BsfnZ8AAZomXWTZ6JlJRnt/v1nbSbqjhjRsGCwLXDC1iXx3EoChhg3
8k84H3mMeil38lKLPanPfly6vzEYFirG+TryJFQyMOV3STRFjvu7OMoc8Vjwr80NybIxG6tACcwc
tKRKE4S/IijQrHjtUHYwjD7+RDgEMKYJjjI2LhAj2CRJKcRd8kbt2/nIs2WLkX7HoCKRtuqQ38pC
zXaxQv+FS2s0zMZ4y2Hw0H2w8NXndVVuQv32S9N3imF/hfJC3KWwBN63SCL1GdPi4ysX8TbWsOTp
hAlYYP7UprqaxgY6Z8+LTBqs+ptDukHZw/QR8S0id4/7D40Ld7ZHPoZgtdX4UTUHK75pioB3MIvH
RPoLl7WSIWUYToFxfNHw9kXOPWXaPlQ/yXxyDakq6FyxraPgAPg2YLpNdo0BlK2DiuSxyVQ25UXH
wb5r2iqB9IEePNUtP7M/ncFWllQP3rEUpIuSeTbVylZki6NC+ATDpKcsSO/SALIJcmnpcZdby0Er
8CH5lmfvVhIZN/pO4h6q3Xiq7zHJ31G61kb5TDn2Vgshre6HhvdPkVpmQIGZkiAeGhdRXtCBTxFc
aDTK95iv5XHT7HSgZsMstVdIoYl1nMZMjmAbGLPGByRFCT77kQhklQmRo69iNAm94067j8mVjqE4
6+1+W4TK4L7LAiHRu5nnxqT1Kfr2YiEJ/MCCJ376Q3rPHW/Sq4mXFdXuzV+q+hzJKQgkj7pwg9P9
CLkQ5EUvAdNJhUN5rTq1OkuD2NCV0fG71I0XmFPB7Zgzkg+V4ioEYsQE2iOHyziUvAa3Vh/LiOpd
e0jCtNU/PnR+p0Cj4USJL8QYEEWkViyYk18QgMj0FWKFQ/wsQXkKIsIjqJaRqUAJdmmGPbNsb9/o
fwQI/i68cB2Ga2ANNuXrbZhN/+d2oV78qakzJabByX3+K+rK06vfbdan0N1cgZq6o53a/f6KDooy
tnr8en748GvRepLGMy7uWfkFpxMyqhx4GyPGhBq40zlaQwrOErI+SM7cPQWUlXUtlPtxeyUmDWbK
nBY8K+LYzq7j33zq3yXxNv8z7oWjo8525grSGoIm0d5BvBIQnHup7mhmFwQXSig+ArC+KwClWdNL
NNtMk2Teal9EdC8KYAsy3f3Wk6XxLSiKssnzK/YKVPeNdHc/sFpiJ5PIQXXbtb4uPcUaXV+Y9VeA
3TJ69gTcTHuARyVrCp+Luzrmg7QHOlNAdG/Z+mZilxRlyfyjFq2sqBFiizUEhWAZ2C77SxlJ7kiq
U/rzwwd1Hhhv67YoQKGwdui55Xn4uoF9kcxuu2Nooa5uXoJ5kUv8vz0R8GACoz6u5fnd4yGScHF5
upXWyKDDaZBE1HgqVBLZYHLDS+WaMvAFjpIX5JoOKfLsbVvv4oD5rSwIc1NIxMVM62I9clh7rq3V
NoBPATzpw+WW/mD1LrLuHceao9J88FKW7JPk4CKvZ1o6FpAQD0tm8MUlvH6RAZeGWHwjqsJGml9j
Tnjk++6UhHdqbXKSBWE1Zi5cykAvJ4JiszG+oMI8nMYLIaMLV8l8ValV5mMnfXxXLQ341BpIWuLb
ByQREy31uQGapGL6clAaCuhG24OYq4QMLepaMt4ireEU3tjz0bnZ5n0LTtTAALYsQXUgptTZPeGM
wOhMK2ytgvJrb0Pceuopd5UYQXLppjvScrNbIqjeygOC97rmK7TQpFsA21iMDmARDJ8yziIK0MoT
FLpKWhJM8hu06QpfBQFDZXpl/S3rHFDhZExhA7feX5e5qa3cKwiR7Dsu8ILgC/X9k9lIZNYiMODy
MPj4EUh7bQCN+J5rG8L1MZXa0j26Ksd+gmOAeP73mFeWgYEKRsXaFGyRThlWacWXDdvbQ7w0i7BJ
vncv08rcN2vLyiVwYLXXxIlORL40j0FVcb6kyFKUzp1keukprTzDb4f5+HXZ8G/iuNNYlupRtFC7
sD0MdPv+nHC+eqpIf2JsGXXSvSPbxzEYk08ZrmdNiXQauEE/aYUBbkdO8Esx1N4jgYr0I7D01zfg
gmc8zl+2c8G7T1K1Mm/yY3wl09bX9YHSPqJhJ4WkslcPj4Kd8VACkk5YCoGsZkbBijI/TBKABlXT
wC+zfojOb7wIY36tmUQwOqi7lNjo3MelFrWkq7EaYe+pf4OZzYm3yEUkpp5h/XHupUMD+ZNC0RI+
fceuQsvrui2pREjecRIHdZEiGAqVfb0RQuoM70O5bi7QJxoPcV2NglS29T07sAkMDgl8rlPePhgp
O5iu0p5iOY4Pwg9Y3qIob2d1KFsb8PRJyHVSNxtsXGPI/wAjNXWOAHG8qvLgkLRXcU3WXOr7BIYj
nRQT1LH2o9STpyZqy7uH/1ZKGq0m1Kp4urzAA6GinD28Q00NTO/kJFcR4DiE93Ap+VAtScbUDxvT
RadYT89YH6yPZpvOr4uVxBW9WigtUgYdQpnK+svpoMhawXetCj+j8U5wKdpIMuNR4a69CjaCzunE
fwNvo3r2f75KRmwbczfkhj3kEpAl7KPXHnFXHJrzLYmtxlwikBT3ccL4P59EC6MCmwkwx1MKz91R
n95TWfkRUVAAPQ6FeuBAMRG+2x6zvj7iEie/0HrT4bfXpPZNMmIqOay/XwYe1Fgqx0EAZZSIe8z1
byrvw7zF6L/tUUyaK/riMYPCJDFGdKCM5flDb71/rCn7hQVKkH6hHroF2no3V61sCkdvQvO0uRr4
YqH49sgYgrS19vJsPiQam/hWGTWun63RrdGIsaQ1ZdFOoWYAh+JWQL9QWz2PmvbxwVwRWpKjNZ3r
S0sFsdaC+rmfiXkktmc7z7R5IkSoVkkAkzJHSrdgF3dAi5fdJuRsEH6VZBWdLfOurogqCyM9UyoV
9r1f3z8u8a38ERbnRiwLqO7j1YI9UAvbLqKIvugYVnEOKms8HLwlhV/HKVpEHEaaA72oOKqt35gH
Ytp+jxx9DRYKIfnNakx1Fx9I+EGQIZBPasY5o+53o4qjeNRgH6UUsjvH4Ii86GxMcOpzSK2v8cID
+IH8mnecSr7DfIyys8heIyTC+Y+dXxsUjvJj33LeUa+ZzLS4VkKTqarxE/GgHH0/0qyoVPAi68tZ
mF4gKVACHt1XS4F+0+rOfjEgw0XKRlIVi07Au+Wwx2Ihc0lu/U/x8YrzgPuQtrXV1iuPxrrqqCVZ
scTzP4oVgMr/ZEXKaniJzygOs9QfvScBHtX01YdSvj/SoGd6JSKHdbyhDH9kyH70HZn/Xf/VYzDM
8uWhSEazB5PJCA2wlvqU4JRNw5rI9OBTFLX9KWjCdToAPF30lOh1EMLUGKdWxEpma8cOM2c+Yh0z
Ibh29Yw1yYg4eWP3vnlu4ZejwflVrw8jy02tb9htHxU/WyLWP4sP4P7s11oz4TXY9UYDusUXSza9
tF45uF5jwnDHkxkWoiKmnpYVAUchDhLF3zQhpfHXn5NNaC8tcETVeq8+V4fHavXhRAx82ip1uxB/
/bxk5DZhL8ja5amBKj5RBiGI012yh1ppNaeX/Qf4OwZeV3MIGrGx0ZDiMQrZ0bmLCAAytFb3Byw4
uIgOf+kZlbTRwHLqr7EF2keKXuzoPhfk+Vp97fW3k+QDxFYOVGC29ls8hLRTNNgXl6lTtmXft7s2
82SgiosMmGlFnCWO60OKHaXSAiNh0ks/WqNbi+eVMg7oebFw3RDrC7j1d+M0pjhUUontWekZxQVq
7loZBHodtAvNpWCQz08Lj0IJB4xfnkbvDodbV1RrsMNmTjCU7l0n4y2OuqMIXxef3aHeqS0ZbTji
fXjOnK2Qe1gIBZRIcfkj82/i3eVASxmIkPV+iQcWFuVEukX9rVWDv3cplnUPnQTa9TWFrfNFxKIB
ITeYBdUEHtTR5C+ajSGlYwoMzRtq0JtVVKFfQbTtz7DEo6M4oBR6GycAmHmieR2NyE7IHNHRii3U
sZmI5Fy++FFIwgvH3ZY1A/mlbl9i/RN3ohxAiOsXyy57WE0OsO88lCIWNZOFS20Y+FiG+vULKxL3
yAFKQy60pI7fIzAEQUb5MDWfnfKl2psfn3sn4J/+1U/3/bi7laYy+8YxxUJc9IOfidsjtUL4pnOW
tNBiy67GomrSOlipcM4wbgczAldJ6laSPkdo4lSVxTbeUxMP3MO69H9zCRIl19TP2WhoHxQoLXEw
UgVqbXRtV3k+SD39nNH6SpCUjzOOpWIfrr1UaUdwjBZ6NivWEQBV7VvIBMhl63P3bbAhccP2HPXT
8g+3rAYYPcAFs7q4sIC/NO92jlB5xboLU7XcoBq0FDUN4GBgNC0ddBH0PvcFF1UMulJxJUUtU1dh
ambAVwM0qiHxchG978sC9Yoqi09APq8rjcK3/9o5JVjh5LUuca7SdZq40H95iiBV9QqUoaaZoveE
LPrQuIUk7+EhlwK3KYW/QROcalfLLuPv+9E1sPvFEqMyjIrgVf6aN4hWmeLkL95SVMf7i7t1Yqpp
LhHEjyMrxGTXbeov+XwM4z2I3B08u5XmFXZC5qv5w5Va/6uisNUVuQfLMU/1SRwzbEDHucY9V0YS
qE1zjX//+ymPLaS9nOCCGIIUFGyFjOWX7TCfDrmpGWJE+gi4GIs2HkTFQrPAAWUjikUL8LzTGToN
epiX6wpUYcLcLXntG5NSAA9vklLi3snfhy1pqCEsI0nVvA4NZFlwAjdtFY59Iin3TZ2yXPFWc/2/
IkKrcEIocM0Eh+lk9Ul+Jmgh2TMzRT3wCSbT+Y9wiZ0cPFnPgoCpouKZP29vUdFut+iYYExZkMPY
PUuJGEtaZrdsn4gS/ZETqmAlPsVzpUinLf0r/aI7AIq3ilDE/RbjEOAV7Rp5GZC3BaG1Z/8Yq6f2
3szssB7qACqFdkEtDYKO95dU0g2aNLjNwC1sowwpiVp6MqJTIds3USi0gkuudDI316XsN76TAFal
84pmBKFrOxco4stG3yX+Y7/4NUeRod7dW9uaZ0QmyfbW8G2VNWFH6wV/fcnbmAxwyrTGP8Jjr64j
yQalDg8bpFPh9FkQV2jq2CjQ9s1UWYCLDubBrs34lch5BmvzdSetMEJqSp9eZjh0dyzi1ingaqXj
C3xp67JHfSL9ePgpI8ClcbSo1fiFcDVDqrbSBCnvOOLtX0RsIuL2amIWXYrc90MH2LXnDrwkis27
mrPWnY9Fez94EeGM1N7+30oYCgQTy/Sxzw+JsIxb9XhtwQEapkYTQdFIpYPF9mQufzn4j2F+STNJ
dLm/pDFjsIPycuepgU2J7QMkxQusikppmcLc3hjW7qQQlph3mN3AlHH2kSAs0rq67r1d4UWP2lhA
aoJCt/52iuzfevAr3AlGmGEDmSOY/p53jRN24RT7kXkJ7G+QSLvL2LoqD3i359WPSFBZD9T4cX1U
iU0F8jlN9FSLhGs6ZlzJzXRHpPpWXfV2bsyvBXJFP50pZX6FNHy1ZfJgtYee8/4SMz4K0jF9Fx+J
mU7j61JMYmD7fwcDCegtcb00CIOM3IXElcCm/PBsH4T8KMNvgr2nMfwES/5d7m8TTFuiL2GBNOod
IINPzqZkV63FjWd59vjdZe4IWUCK5rQa9JViP/jzMyhlbe8i5GgrfBbVZtU5BHl7zkWvu9agmsfe
3rQ8MRWkPDlsS70Ov7XjhbRxYjGATUOhtgppRFkbdJ5HuYcjUg2K+hZqa/XamXopX8CUIXCumuDT
OhzvPlcZcIDUd8N/GxNikD221Pz/5oMLfJjqEPs4OtgQf3G57QEGXiTob9yaysi1IgjolO4xKpZ2
MaLWmLEi9bSqLdqTZGQ5jdPw/XyFxyTgSjMKs2GPEXF6QAGFPW7bCrXkwd0LmlR3cAYJjVi6V6Eo
bOMW3rM9/tE6Mr7xlixqGjse4rcZRxuxK5ubc2067ZRMhpIMSPyKX4u8PNECJA3ezkv2R74UqoId
yXZPXriz7E4w59aVeesuN2EqYxor7iKCKoC7MWkhdArAOv0jdBZDAC0rWhZcdtd8q1rpCfOV5HZQ
OPQJhsQl9pcl/5p+HhVElSczu1KwS5xqjYEqeMYTkIAPG5whip2D354avFsp8kdezzu7tVQdT8Nv
LfeQzYHFuuqupfe+kfZVcyjMSxLDPY/PtCHtTTOYW0xGxyzDPpigOjkJIgW+Z3X1JRqSInn8ZjZQ
g8ASbTIpMBl2lwHr5BfEJrsAZClvSuKupIh2djQQOYQvQCMzdsXIvR4EtKaaWluzxBz10YNrxywo
vCaBiUndy6iPwuV1g5/H/Zzb7WBKGco7u0ZJvAW8xpnCOU5TLMUUmOmvsVG6QC0y5TYdehulWCO/
WcnP0al6uBQEm41fHZ0KiAqn9V3C61M3ZqcGp0PijBawbRSG6GAF2W//wm/7UUX1EiQv0nH6mKQw
3+hc5M4Fpf3DDWYRFAmhP+tNoWAOAceGz9jnAOsaggAgyKZARS2wOirIcWCuWuS9lL94s6iza4c/
by16fyH0b7SFQ6nscDnKtkTvZrF127Hwl3+wrJ01VsDDvWl7ZnZxSqFh5EWNPkR3qGMaKOcXNHtU
dXdgyN4x7dWtQJb8XcMAicnKe+oDJ0JsWYgeKInJxzaMspUka9OlqdDpWDHSW0PNLrkZFz4XYjkp
uUaNBOvbm8MWgz5tdbZkSetLLZsBF7pIwIR1hla/yL9uJ3RArHcjpELZehPRQpgZenD2QFsoG+mh
j+w41hoKUfRk0byasNtxxscUfLahg8+vRLAU25unlPMoB/NoBqXydHRW6q8BvRbUT9ZYQt23Tcrx
6NCwq1C3b7hd8cF0sArPhTC0d6uIFsWSrD4mz4S7bsyTXV4lY+u6YAgLEewo8zutn5rLXfzOu3jq
nrGH7lz5VHcEO9nereXwx4gw+xJF7B2nNcqDzkvequLSQkAmxaNdKNC4dmLpTcWU2QwC+lN/AaT+
OeazlSNdwHX74n+mf3COoZu8eHs1FRGQC3u8HdvcJs3Ik82FP+iyqjRSH7DDvY5b31aWxmbLRc2R
Vcs2hK/kRg7uLRYN80jGlTgtev3xPCaxQE0FroNEmqSGAUI/WwLE6NXHYULvbz4kB3BOY4HDAPjo
FzTgNmShOGAhuFB+/0m4sQM+c6cUBOB0uhQD3G3cKEn1yltIWRTI4Ihs2jBevHunUnjWe4uswkKV
Y0B7+1243VFBWqJI57wLFlO/7oaBuA+4F578xlp+Q6DqzO1BM1BBSw2bopTxOJYFSQc7DyAH5mMq
Bn5EMZquZiSIUcAJb4KDtopisvXY54ISsQPX7+7QML4ImfAUnk+x499IXlKJFDjpyBVaXjoqDQnd
F1kFWyeA6C5NsgzPXMApZPHAyeb4p/Dk8ehg2ni7KtE/Wm+0ZBCyyAV7gJlJUBQFwJ+S7xSvwCo6
4RH7OVlUPWDU7DqXkmENpSdtWmoXfo66eNyRo6bgrDiYaCdavy1jKbSZcISPANQ9k3r1GD1wOhwX
gfBioJEUH1T2CsTmV3Bua/pnHuo3bolnYQw8nr2q9Td4X+/umWeMyBFdkma+7PAO1hF8jB/6Tgfp
zeFfujF2j7re21zcT51KPVE3Ojd4jk/fqIk9SY/Kp0GPI+vOaOJBHWWdke8NlfMb5v80EvXDXDWX
9ACGd6jBuYoO5zAvxs7jcJ9TLn+24NEMId80uKNQWkOfC9UqvXicDRVe88Gtbfx6FosQ9Glk4Enq
7PyyZdRBflb4DDsCiLGzKRB2LTd+OMcbnS4fT+G0F2MugePNEditmJTAYn2jkIkeipnsQrj1CZP9
u8yUaLlgVfEIh0EZLISryCTnA0nd7Tn1yQJnupfjnF9/IIi+lPgO+QZIWz3L6BWJ9mMco5JnZI0g
sJ7mLBIUc7Phw9weaX1xNq6jJFtmsbPHjHyBA+xp64TSC9f7nQtEsbYk+5WXAOgSWSHjuGaXcJiE
4Kr8zyQyunNRbNV72gJfia3hInNNj6DzS+aV9QD3G8wGVS1LT4/tGExnR83Cwhcv6IgeRruJq8++
8eOcbATuHjfyB8MpLnjANffLwifqhPttWJHAxozYXUsyxthYhvOnP7B3+8fyDUUkXLVz9ihzX2t9
9Waskyg+W8dRFg3tTHrImJqd0D5rvmyqgs2HqMn4mB0BNEnZxU7DXgXP5QLyHKAFrLZNRn9ytpOo
KvIQzZdG97eAbijGwO4SSPqs8UU0sAhxtC8kyo65hYyk2KgaYABVrvnBdS8mw4dNNTTh9AJwke3M
txBDmXeExHw3/cSkndnoC7iCmQE5ECVmU5BrIQqNv6Z0szkOogdEFuR9JftOGkuLTKzSEheMX4kC
p2cArPxxrBilhXMG8u7ZugYaBZr0QjmvrAHAQTLueg430jxIw5o4mCvUR9t5UetOQkf+t0/APpmJ
+Aq9Pj6NyXBqdZy+2u3kRSSfwgjS1wtLPMsMb7AjGxZgV7Um6heYEB9JhIgwwlUtVmWb2eIgPAaj
MajCOupzix6yn4c7+Pq9HxMSQrpjeFoviEDlR674EcR7tm/IFRjK3XB+5S02mpH2McOIaj2W5pDl
17TRaxSKHwqtJUOXMeutQiKPn8fHv/dV9cm6aT/62eHeHtqQ5E/MJbkk/jVTgmawHzkSpqlTGa+K
G/6dxE5jdVxF0m8aePRLCvJC4v5xTXRHMWmaohWT6cxBopJr56p63fHS73AyaYib9tbaUBptNmnX
sMJ+MkAzd5o/PlWQMBq1voJ4d6d0q++zCCiV1jrrMUDnw3iISOinoFyl98FSYUxVO4o1J6zF3ktt
V71JTbY9xMv4e1+NAzZiH9qC3a5hP+T5RrVcET23CSq6Rggr7e1PvT4paAEN9pg11w95DpZGnGkX
LIipe/bnKR1+GmvzLKnh9l97VlEUSCS3yiXrDQHmpKRSTi2DaKz6usaBjVsD9Z2jG5qlGhcQPQPu
vvPx6Y7AKvjvWv2uVqLQHnLVJ/6hcxahZ+pwiD7X3Vb2GLun4rKRNnljc/hcudMT4sHLU6pQYdL9
1Jr4KsX17rXRT/Loe2TZvmItsgOmKtZYYBy/uBD6Jf05TIPkVIQA+atqD/nLQlTwKbRAGCCAlKMq
ZWgB6vnxrlWphnOVIWjvdTRiLDl5us7WYVBz7q2FSWfYmX8nxgxyrNNxoKhdw+5EH8UBxRt711dz
fQNqcIfVDiix8V1lwhBBZGDKqGmTH+14DjK8T3/Xb9hekSC2y55JZyD8RJrJRqj6+oOzhybt5/Ht
8ez/wI55GZzxRcfo6O3sYwKFKSe3LCR9LA/SA1/LAxjUnzg1hqHZCPkZBdaZkT4kYlj6rRz12kJL
RsFcAZNQqaYUUdJPryaItT6NnVCQi+wmzGtYXZ3t9TS74ZdUJ1iIzD1e0FUMP+7LVY76gwiGbnpI
ORvqOyhA5tBsC0nrzAyVVgCAyImgr3DD9/8mdtanfKLTacGWApR3xQOu4YO6i63Z21Q8kBakAfa1
4uM68LxPlCFIUAn/R3AlhjY9YQsrpHcEjcvAiITeJ9Pit1f4PapqFN8rv7KVEjE7tuqQZgDlA3m6
Ijtbkc4tiEI+rGoyEE/Nskn4CBih+G1wKZNbw0RL/gN+RBZwtfBfhgPd+7A9LK/9nkcy3vZ1Afr2
taNUa7HIxxxBNZ5xrjGBKH68lmTSJU08ioiXOoUFuwrDuxTEQG9H8fHYDmwuVP1/kiy/jibjqc27
UVse+UqBJAuXMLac0wCt8UTm9Xuh0wLnDsRmXjJBm5zYBSeubZqCtfS276hfD5dwKaRTvVsXfkMn
ZsWwbAXwobG73pXZW0Zqw+m0aZlo73RiZmxoUo5YmPNvFM1k54QW80IsJ5Fc3k4AfUTnmpBhzotL
Qy1D07PJ8FRUBb6L+tN0bufJypedqJaAazy/HQxzFDHOPTshEn6KrgWJR+gX9XJDdIKh0OjIMzKb
04NTjBB8BFDAf01xIH2hbiFemXwz2VqJ++WymT1MI72yNvicvVq2ClMSWYmD4ophuPdppPnr1QG7
YOwCag5sfS1Rk/Hn8uHeP8fU8PlQrRnrHseg54AXqAcXjxDJkkMlbhJup7rRwdzHYKs1v0lIPNzV
7Tv0yqASrjBF2Siu6N5Vz4pVCS8eF6/vUvLwNGiMJ3eXS7FhsXSuG6NyvqHldOpWtcdfX/t3EiN0
Ye9/QZJ8hWbU/0agDLhzP6EhYFEJQ8QYeyVuV1Q2SrYoLakZIjphFMWUAIrKNUrnujhuWoZzTgsF
UexnYT3+vSWGB/Q58dpZDPiEnM39ZXbTtBW0a37LLZjZjpl7UMBwYmGfDs0z6SknSGVcny28Aeq6
yjEAgEPKgWK5+rJPrCgS2OyBa6T99PQvGx6FlzXgAEnJTZXGxdWIaz/+t8QXymzvWLDOZzDKX3Sb
arh3tpPSljOgovXs3G+OuYzrY67fJejQlHMQC53Z1ZvJ3MUXTVs8V24MwG6Z4LkppTIfrPyISGah
2ZUp8p1XdEccE+jDGR1mr7OLlPorSbqx7sxVQRHdABo2VHOxPV2E4PBBrVptG5EGJKkwczKNX8il
KaSHk/SEC4nIWeVBs8enb7+6Itx3p/7dynD9TiiUGQFWbpw7mCExUiMO92PyHaaN5aaPcdOv6AjD
kUYG8RahlUNW5yCBPm3gg7CRFxjomfU2eKE/fjhGeJ+Wal8dLkQaUGfSay/D84hh7O0GKjJCq5UV
21gJfTGeT0elkTJJuzGhiYsSvEKf8zoKIB/d/0t+KaUTLUdLaSwhZpKQXVs4vQ0QSmFIf+Zzx/rp
w5XR7AEfZcmB7jDJVLlUXEKwQDn4jGfYBX7ZEhDOdHSvHOuCzdrNAshjvsbhzqW+5phf21+My4ns
rTIDqFLllWI0FZ1e0dfHx5IenF3TQyv8l7wEy9mjsvmvrZEepyUuGE8JJU/LYryLQtCh+JIkuPHy
9FWpgSgHwN5KTW5VXhTJX+LywV6FvZa+copn2d59onS9S0ul6DU/Owg8flOT+8QU61d+9uTXf2oB
4eePgHVMBSk9wW0WYmbq/9LBuRW+LeUyGhkYTkrGgBQxmw7O6AsWZ4Kut1SJqXQxRAdb7MTTdSjr
LBirzrl4SsczGLwsOB2kxsxDJ2WicSjgD6RmRdnZXldRQTRrtzXBzocRaAD4zG26CJpLeoRWkTun
WlsNwtP6ceY5d3g8pxnWcs8Pxt6Ye+qFYtfYAz1ME9IJ/BkLk1dKIB2MjOlnAHe0G9N48vQmCDy/
kAe69ZjueQyMqEZkSCHwJMFY3nWBPBwIFxuetDV9t2s9RqCS4BG78q8pZiWdYsmMB4tt9XN5duEK
ct6HtcKV/Tq2LGvWOgy7inSwW3LzUYCYZbyeh5EpVQyXm3Ehu/HcFy03RxMXjj9dcJ2a+Qt+W7I3
RyaIczfwiOBoSLuKzv1Uel6b6FV9ddZhAO2A+fZ6S6Mb9zlCgv2fZJnVsmG+0IVpqNk47rNVMOgL
tBL92uK53P04cbfSII5mvQ7bSSf4fsAUL64cG38y1r42sZ+cTDWFFiNUkf1cVQ7Tzt0TXRsU4Wq7
G6ipqtQCawZsRSM0HdR7ALlAictx8hVz4bXFIUkLOE0h7ESa/iJW33H7xTMwBNjbXX+rdJE6pcWw
fMa4XaTdwgRDZf3xsQidno4viX/5IrcmqohDyNPeKL7Ro3KAFZlo6OoTqW2czrBKO7z4FSMoVIlq
XPrr2sULpCufOVmssskeGMSwcG/SJ34g4SsEXRoP+5OSQDJ9iY7AO+zoOInEa8rMgbbO9olAYz8T
41inohcd0Wwz3xP8en7cY2zqBHOQfQaNMrV4rA/LZF1oykDpBugPqDs7FcwgnpBEkoLnwYlCNNQ6
yVL5rElYFUJ/5w7z4iX2H0xk3GE/ko40WAFGpiGAd5Uc7MwoUVlCoh6EG4cVKDNfNIjQBmthtFMp
IqDs9/JBdunc9tZFokZh5Rb8LuTTNf5koTbQmCWfYBg6TaE9M3PxX8tnW8DsAVktjrjtI1U2xcwM
qxhflGt1O4jFkTiRqtsuH8FmZWgXHiOK0xGHsIMv0DiD1t/HhNNShVqOuy3pgwDWyapBGiq9dL+1
QWcivPhXWXTwPIk+SmagSDBvguHCWThUt7+6pH8TvyJUvAtPZXii089rlEuwcqONxnvYa57227qn
7niXYwDTYqkNjZx36oj1MOyPa/qiXgcv5QNjYMU7liPtz4jx+iPw3zZjFtwrysZaN/2bFi0PewYJ
xb/RIs/LL40bEngvXqfSGQGGJvtIjoPU5QE1jsrd7dV23/tQSvV3Bb6yHDDTuoYT6jAlgq+4PILK
7UIQ2mE5Ievk1FC0cBxf+Fp1vC29AfTP8K/7xqi1n32TZhdyBM7lSJ35Kp1zM+4oaNkWJnKdMNdk
PYceH4HoO1R+fUJciHsJ40aeipBiLgr2CmTOg0IpuBen6GI2owmuLs8FSssgdOKfS0a+UL1P+jwy
R/Tk0mkdWDTzVmv3ULUc+fVUEMgeyBxN4k/EMNNk5RFS4Gq8iaVl6WNjwW86mhcpX6goZd0iUmrk
1LnJBqmREyYbl5Hm1Xsa8Ob8eYYbhG/oLeT2d306DxssTlwraT33YgCduXFmNMPZxGOTVPV80iKs
HEfK7wtvh7ZnIboHG6JfgWyyM+/PiilhKlJ/T8DQ9f8QkpKubOh9xmwTEQ3XoocepPuTQNaCFfy3
gTd/OHegl2z+X+sHk+UBMUdJ03a4KT6U6ZZd+sYM3FpGvBkNa+/9Mj2HXcagQOywUVcYZtYq/5H8
/9lCUmfNJBZwj2qD14mdsEu6XHvxHessH4gWArdOCOeCVGZa4d1dzVMOX1NB46TWnrAjcuM5qGX4
uyxPreFKHwNJdXnBJ1BbQUxzNPmQeN3v732+0VIulYVZOnARF0MD51yHaCdszhBSCEGkJDpEOy1v
piUBWv8rH/NL6Gg5IsO6RfDQP6vGmWF2iRTh6T85IQZf47cx/FeZsSVJtxBBKwDWCLVTFhdIV4Ms
Ds0KSZrOHsGy8wmJw63Rn9y4pMCvkaLk0nxPuFDhQd9vFtwSTfR6B5+mKZKCz4PFYYgD2g3YnBy7
yuBtvGwPNaZ2sEBfHMM+nXb7golXTkdKqm+FiIhl+kOyOfSBHxbmCXvMM58cS1ZOoZl08QlQudYj
U9wPXRXK1FMPBW4m/b6YZ3THYJdH16mgrXMLdTeIw10v8f8Bx0uoWzulVENBVWPNKg4Oz7AIkJ2f
CmprtQ1+0+qPKZmqHPfk5S8ssLxzqSXWnLnDhwah1nfJRA5krJLYT9bLRjLEYF4Hk1RdJTg8oF6l
L0GDROODq9QzStGDnZu8Qw0ruS3z0B7iJuR1aBbVTMx8Nu11b7Fc1uAK6eGFc72rz5zGCprL6tMu
f2zoloWiW5HS1to5x5GpjPcIF9CcIJ68jpeoRUu1dh0jFGE3KkaYmL/bYq4omKE7XR7c6KtXkdLv
qGVZEd9I9zSaSXCS7iM/DWKQA2EG/yZYb3FvPFO8gGLMVHa0tpiqYA4tfiHkh/G1dL100eAgmn4A
vpAioBXuLbmbR0bB/KM9c9JWH09ZFYrXTV68/I3NWVnuqDpURUh3dniA3T6yYjrPj+UtPGCe3bUi
6jPhMJSfAk+UvXRbh4qO8g/vrRuHFIOqPgxoM+opKCUt+GieZUX4Ubuul8uFCqFFHD3nEjW8FUm+
GAq9Zyf6wfHNTu5sdq2n1jUlcZHAFXYjrOUp7NNeSakAkrzt/xqMuHUlq96g+r3RLjtf1SIfruKc
khd8pFTeOPULoRXnKUe1JR0WElCPUmDKX6nN4zlem+y+3YwaeyTXzCLrBXEYChYdRGnu05IBhST5
uzBKIhMi7Qdug2nmzgiT7UMbq60FEVY/taxoQjVrwfdAeBYzsnOEt8tfkAmUzypmRN3FOjBEIu5b
FuzufjkrHmFfhrCrQTZSyDXUZQq1Il/3XledprFqXbd+f5LFLNfKVIOiFYRMDP8Lk54DrYqkIxwg
xNFnGnKFm+Ll2Q060VVrpT/Td1tfP6KEhydExq9BPpqjvkmC/JQnfe/H7fBX4ZHIk0dQ+xC6s6kb
zjGuNYyl2VFIoeH9XuKezXBMon2ZxQTJfqS1nWJ1EYNFkkkHSJQXlxCU1MyiarvqNVY+uLYkKycw
Q5hH8PoRv/CFT6eW4OXCoHDWB6TmReUG45TuS4wkjMV9zLikZAjGKoYluiCi3azB6kQrdKbKl0GE
QB+mdhrffqM1gQVnPhDIiW2Kav9sThNICDdZ0ByM9I/fu76PpOR8NQEG4RMPS3BCtkziVLY4tcHY
3QgHN2EC+L+F3MKNVvFnDxiOQb+96cf2CL2Wz8EXPDiNVr1Qg2cl2mAGT3Bkylur7Zc0d/r2G3FZ
MIJkyRvIw5UNg0AnR4t1vX4YkbdULpKRp0JgoClwPPXpS/Bf2vBy7jy6aFUoZK2XkDOGhcJsg52s
60SKgOLq9v649anduJTksflH98PiaR9v/aAvB7OP/41bhEyb/s3Jl8a3/Jj9JKjzw6g5NAaTTE5L
DasS88Wm7Yr2c8MqUIaAVvnekdG5UZLABm2fhsYstvYwDYn1+DRiCpzgzi9FBlxJDuiZgMGtxGWv
iSPftlQt4BJFMq2r/SOd49BN4FftssnkluI2Z+XtrE692mwyclmyV3W1QxdSUxl020O6n8pKWic8
STLcjCtaKDGlfutmnnszAnCcsGb5cSlOkWz1gg/uTJA8Ro1y2YgpCeLvL6zjooad2UbfIYhOuy43
1g+9O+RtP5wzQIIRpGnWByh/L2S/47iVJio5wklRBqm1m9aGyg8Kkglv0qmEoAg7LnOiv8GUNYry
uDJLW38UolRvRjaCOohaiI4jhn0Yg5ehZbqCza7Zu/oXOQn7FrxPYdQNYjnoRFkAMp1i9cL+dj82
l4pY+ldzT5oSUFeDsDS3kOUUQP89ip/cAZHQZeKQ9JG7iE+nl52yc29YVBToC6myrlSUIyLv8bQO
7gxugojnfk6+SFU5bmQTs1+QaY4YEp16GXrAzZe7KsJnTzih1KFmaScFodvIbIzTfO4aiUd95ZfW
x0MdoQ6zTApQRkBokjas6oisyGWaEEu0f4LdQjzOX3dGwT6E2e7ta1Raq/eGpwLCqP4uFquSUsok
UZC/vfSCc5kv68n9f46IrJh0G9x33P/14vcvKcuJkiex+mYYHqIrmQfbFNCGrovzyM4fJm26+iqK
oDl6MJZsBGg7IpfTjASXdu38om3sveXcj3s8Vvag9iJWvwfqbWyl4A9+1ARvMgpYpLJedCgElr5N
bAiNarx2170YsVZhqH/8wjj+l2QQ4d7UJi7I7YDVkPpiEXAD+O1c/1P+A/d1IWElFp001bpxR0lq
s347nA2DA971q7X525XjVDEyC4S4HfvAhPZ5v1nS47UdVmhqonGg4utDtd22wiHxNCHa3YuQ1mU7
vk+3IqQcMgy2DqR8+EaRTt7ZV+4GUv0FL99tTa/yVJ4Iy+To1qIfm3tTHGKcHoVWQFLHtCDGkTkd
HW5RlWuQz+aHaOxpaTiXoTK+Vsyxxtn35pXknjm/gkihypurvwcDz3hV6K0RhghRqOzEZdQZJ+v3
MylwXbJwdxHBCO3LNSChv9IKVnfBKivWwwjxSKL3JYpAJAUY3LijwQFz9NrgCW6LaPLeM0Q8pxcs
haykfduMrKZsaedK2Hjjf7DjsqcIERpC7uTX7wo7P4K3wn4AOhh4cTYkY788XYf+BciGfrLqhdN+
9mP6gLwPJUNaO9yeJuUaVrvwCXktLAxSTW9WUbg980sJLRMZmorr54SO4GokLmObo3rcEe4kdnBh
xeKcUnwWo/b+p5AlceRAooA1iPV7d1P66PnPOKwjuurbJY4OCK9OoSHaihgRhWtlml0HM29UAOYZ
2cDkp6PK3fNu1Zdv/AxzVjClC3k1ZMGj38YcWM3UD/WGZnGHFqWyCNrpYBJNoD3dSQYqXZGcqSED
l0XF0kL6AYj0vGjCBFqOwgngkYdvlxEIh3P5Xs8iZ6Fdr0sPfLfui7CrSdR/vWqe1Mdi6Oy1AZpD
j3YCTBw5YrvPUt5wVKyyfl+6Bh63UD7fNG0lUO7r1AzXv8b0AlZSNON5KXvqtRKSKse0FZzCWux/
o3LCLKTzo8tvCtNWFrc1ng/Q21xgWkbyzpAGbbSZ9GxDYatkm4S/yLjtupkK1zB6nfdy1VQof5q0
TINx5wTr91XyLCXd1+kMou+tnOS9R7cea8DywNBl3QjuatNYPLV56Te31U6dS8tuScTx1Ukxsv5C
pUEPdl/z93dhTQhtZoX7YWLsuWg9Z9vbBL2Yp+Ibvt4f1F4r2gWX8on3qo7oNyxVUK2VpujxTVi2
dzVXs3PK322H6qYiYBML7OYAkhyNxdNROPycsGblqS1c4rnfKrGXaOYzZn0JNCEyH9gSSv9R5+Nl
+4Q10sVW+1KFNNvql/9y3P+rom74zBXJf4sqjDsi8gWc+HfRQgP2dlXcE/migt65reMi5z5nNezq
ydqVWF450T6QoyxIbtd9dy5l4G3D9n3thKrVHoDtgx5LpSE4A342mJpC37wCUOwfqcvXFFcl8hbE
sJK1E1i6qkMfpvmrQgkStoOeuGrXH61DNSSRL+8j4dP2k3TG84KQOPlTDe4vFQDwKjWI4fmQHsEW
1SHSgZnjlzSRrJTt9AziqxpqGbam61EtbEXVOHNbyfQruDyYKcvS6k7sfZGbcfrtpivL1ml8eJat
ahG/SYpoZ6GdNYnGXDpyzwLBwK23b2pX+XGPIw8z6hz1dD9IenBDIJ6K70DtzCyhiSbpH4YcWapr
XESg0t4ouSKJr0XTZxn0NqWpbWOlRXKFeXVpx9mMo5ojV75/Y2ZDC1jPI5G15n0/ZiTyJMZGCO/Y
L38t/yd93e/VUC94UoHpfvlK0fLkjpOWNtuq9RogE9vgMM5YRwDfeDt640jXuLdtjQlOh8hZpGHF
V6E1pSuS/3VavdT+qsjVaMESzYX/C555FlGsO4xKP1x/1PfJcF2m6LA5ikjsR2kFafiPcDLBnKz/
i9o/CF7JoWR+RsZ8uYe4oXtbKafkyKBoUKWLjQcdaMBobGxtDMbEnIjWeyLQqhvCJuhCtsmWkyjf
ScAz5djRclGFVaLgG2upJ4W+3AxEfID92jY+Vh/mfaT8K9pDvxvjWWZRGUtRfQzNfpSIUQXXpZoS
K584zRMPnnPwt/RfVNU8n1x4IJ3nG+eb2dR+9NaM8PZsM7dBJc4lg8WTAHE1a3obJYzUT4n2whyA
POMdQ4dLhLpZ7n5axo9RBhBc//mAKGbhQdWm/P9nOR/HFGClOzxsmP3erK7dH+dRgzEucBHYhYXj
+1QQv6FJGuBcGKQHSa6qvHFJ621Q8jd3lZETT0gNtOgbA9HDKXqKia+OdOUwfYzvM8IAaItiVN4F
r15TrExoEfr7Otw7gh7RymF0hGGExJ+WRLCGBQMwyRYWClLSf4EXx8hub3EG/pjAgLcpDncagmHH
IE/i1yxLMu7lPRR/F8JeNhrN6ZdB9Ia1K7xQDjX6HPbD/ioYJflYKK2Co4v259FP6wHxMu4to24s
i+6FlCYe+01Ct+EyYSze0H66KNV06+IQh8flWHeoATo+buoxb9sjKFHwXdrpnGIimPROPujDKdw7
QSOLahtHifgZvIMPot+hlTbgkb410QmZ65f5pRMIYB3/Dngf7+hwy4tra5QqF7CgRdY9R6xAgkNR
Ho87dwsh8qfLYZdSQXNphyNt0TySnahiwYK3wGfAqSXg+rg5mJ0s08DjqluhaT0w375aD3VvqrMT
QgNhFrAkbEQFTddAVJk31cfEGL+Frj5DDcYbvCX/jbzdlR/LTTD8oca/+0YuXDAL1sbAU5El2W0S
bY40cLYR+ZAWF2h1vM3NWEucUZ4miz8INitXJ/uXQ9zF0MJzJZPIAutbaN9TiqHYUHXqxRyVu0Pc
BY+p/nDXK2wFt7MWhhyEnIGR+rcuCvwt9o3u/Fg2CZrDKE5JoOhxrIG7fW9nZlRnhnAJlXPIjUJ2
5O47gRgjmbqABg9lHh02+CtToYIeA/xQS+ODSN1MHTFj6Wu7TsXuz4jxmpAa634NlaVucfkkBZcX
v7DA+8MySXa+pQrBPk2o1cbvNhNvM0C6Cr8kpJ/rUYJmRr9RJh/rP9HeDUHeB/CWr7adYjVQ22rz
ZYkoMvikCNbBluLi354RdgvVmn3oih2iYbapr+8BBUES/AXwjJVIej6pxZIlvQReQ1QgNTf6/9Qw
FbHKJi/fERz2l5tttdUPdxWUn3lC5iPpWyl8b1IETRCuTXApYJL/+g0bjzS61fXwR92X55xQ6vzi
Zf24FJ7GotNfMoTYyyWdKtPJrX13ZzOCTXLkeRyWfdt0Nmz2elB9Df/CalDToyl9b20tWKc3jF3L
9lsw8VnqovYYWT8zQv+PSbA1J+KGFRXHPn2IVyyiJ8cfckbhKaxRG+vZR+C0wMjhoCZjdCfXMhCc
0l59EWFI8zR9QhH/a/WIQ4ktUJ6Q6x0ECa3vmYhC0rjuYMitrNX9YJXPvJGlhMBmp+Uu9SJfacdz
yno1BnLSSLRhHz61gytmIIeXowhlUawRvgxlJQqU/FMf8lnwaIdo/C2O1WN7d4iYHi7dXrQJvvsp
HAVym8v7Lt/rvy7jnTAOJGj30g8qpI28T5Ol7sHJ+AjzTzEvmyXFWM/sQSmJKaIw0jxBsJr/bkTz
kRbVI9he+ONAiWLQTlvbmpwHqn49y4wJ13XTlX5zQzuhJOyVLvBgPp57ARDnLaZojQEA39d3wgJG
VPxtI9jTxMjC7gUq5xnU7m7wlZyUc0mKY3Oks7T4j0uqz4IWxchXSI7rvT7uZB63LbStckUol9lk
nylqGdzYhw1XyzyYrvKKRf+kz/13giN+iY5/51ieLNKr1XsNUecbLDtntzipG6n7T40M+BABVoOi
JCxA5u5HR1RvDIpDcQg50rQjJpuZ0wjhm9OqpDXGBwlTBWlhjE1LavTeTYNeeH0rk3Nb3oXw0pUm
/ab7pwKes7qlIVMCfcTPK9F123sgo3lWcV0dbMAFcO8Ix6brIAdcNYBjcgKuSefB4NZbAenyxgVF
A9BKcmIsOQvcag5fdv0hiR2Ac+ghtIz1L3qo3GQM/LhcvPr7peV8zNNmvJItuaqEM7Z83DWrj+cN
XgZ9lQIDkk5N3kHu81aVsC7snv0U6GlP21lFc98GuZDssM0XIUzW8NarbdxbkP1F2Qt1X+bGHqli
NFsLwg9Nnlm7yRlGsuI1R+5HrolycJ8kA1FViHV47GxVBjqK220qxZLKaQxDIU1C10nLBnKbjR0b
36NK/2vYvDMCzH27Tj7ZOKDuVZBsKGtHR2NsIaTLuJS4K6Fkg723UUzh7KrGkrJzrEieai+ePpT+
qODRDxQS9y/t/OY6VHijwmkJm5C4oe9Aslf/fPA0KrmlXxUIwdZyRwZmrXd2OHLxhtqKCsQU9Ix+
2MjVeaOxO82DSoGbQsIRvo1CwzGrHwgXSCQS2rcDAngWRd+4Va/Xpb1WjTatWc24RqyLp34tjlom
WyjT9eUhqnktVgKqplyiJj+M2vgIFJ5rM6zy4hHRw3lBpRIUSKHM8kYi/fNDl9sNXYccWBPI0d5c
AzswGdDZFmjq/Xh+WNqWemkbfcfJ9xL24PNqJFFxmVkDg2l91x8qry6sMbrOey1fS5XJEz+lehL6
NJsZFk12QUAFQjHyEzk2OkBnUfDEtVX6vMHkIr8wESm9oCYFKEisv8JIY0VW9FTk/InPGCo6amNt
C/X7wUZDvkwoUEqqRighEeD6AVLPth4zZO5mIaaG75p7agz7WeCS3DzcY/5hKA8lzNWgbu7nBeeH
tTIkxoT41ukBM6OoiDN48d9s8e0ApqCCbUjdEHxRAN8WCvshZKEALSukSeYMsZMAU3RqXb552Nx2
POvPSb/rd+0rmBjd3STYSqiNMt4h7jY/7rwtEF1fuW12AlhrghA6XyPQDSoghSLjIFbz9qaNPpuH
TQMTUXH8WKrvx3P6E/g8x35UxGdN1ztxdmxKob4bpHMxxpUn3nOppI60LWmRS/fOX2wPP4OASOsQ
hkyhM/Tiockvvc+sF1dhSZrtZ6EMhW37nt0oW6dO4dp/sKH8lhJjMIFyK+N9UV0LYWbX993rZuDi
s25K2z/P1wdbfv4YU1Y2y738oABpnCdhBubUPta/XiUAMBCsWJpTrQql2Q54ZhQH42nhJUTyCqO9
QynYTApEUwZJ9k5JHPBHh4i1mPFjG1Jvb/uQbcg94EBK/yBNb3jXiK9WxWxvgsefsGMWy0XSBz4Y
WTcZ1ZR36nM3Eet9d41S4BdugS9uj/dVEF/0BXYuUyM/YPvyfF2yGB2JWRrzCG6rx3Nm1aLyrhxg
f6fVi01DOJVlRraLPoLm0HxFhnRQfZaSlhXkGSM2aPNPk8j7KO2KzAyyPrCU5D1wDUudvx/HZ3S/
G5mP8DUplPswBatf5poRKV8hrQ80tjWG1BnEv1DfAiyYqLA84jTqLvvNDTwDzhNC0lBQ8AFBJZQk
cxyrxXfR3Os9cv79lnyuHrONd2IpDFo2LukcYgqFWaDSkDKtE5kL/2Z1+xbJiaq+JgC/UQ9DC8P0
SNNvvr9vL/LYAB7kpZ34G7+FhSd+3ATuWpXjX4VEV4EfeDvt2yS7FNPt3igenEqUmnBhHO5HFKvj
T+vXpZtXC3Ryat9en8sq6FHqjclE5/cNmVCU7uND9nhFOiqu1CmugNaG0UJSENdv2mCoadPBbdyU
l6PPPO4yk//7R/ajHreqXhEhtXaNR6RQ31lbMlUrlE9ukYoTlqBRfN7LV3sPeRkDl9mQUQeq1r0N
ERe2pCqcFqjR4I138ket4UDBgXHr3X58VOV1ymDwKjvWluHVPvig8LikUq5SxLYUanfroZ5KTFbs
SBTVZbIRgxoYp86zUjt3rvd9Kg8kuVDO6xhBMaloYydhb/ZISYyX2m08U6giu1xr5fDbtm35KcjN
0A1PP34vrec/ulTzLkhsVYt975r1NgxmvGKsDBi/rjHTsDE0ADInfUE8F8Xnql6Oi/ZHbDEY2M8V
ZRSk/h0VkDewnnIvahWs+9R5T9rSETE0hAH1cNqNuk9Wu1Yn2q4h29XqsbmT1tTtnPXgAiIzz6Hv
CVNEYm5Yvhcg1wQ1O5y9yW3rxol0LuZ+1+FqZY9JTiSTA0sxDeZ/XKDVk8+7dnqhPeBGPSIeX72K
NUl/7daQE8djRcQu0Rx8Ep8CGgCnXfqI38wSw41F6FpIWq5Hc1pmtIWeyfuV6Ho8S4W6/aXcaY1o
NuEOC22t0ozjeS0ZpptxQYD4BC50vRtFsM3RsuYtRSu8DMiT5Nwxa8cdcD+UR8N/uFrxRPhYDh+s
F4lnv/wLfqKDaydM4Z+hAAug2bobwm1NkWd71Ob74mkUBuznhLELQYGF0S9Jx04jHlFZwYK2DF1p
SzlOfhgA512lHctJrUittCRhCXUrivjT+rbzLPE/VP8uSoi9N/rwYNUrh5B/Rh6LconmZFyVmVW+
c9FlUdf130AqmdoExB7oFkqvVV1ZQTq1Wkr9g+Uy1aSI6j/BpWvefZT6+eZ/hyvSwoGlo/571tNW
HR3E85roMSr+plg2fNJOLeGwTnTJ0A3a6DSkwgQETfdPJBbiuvihQotAYPfGo160JB+HKgzakJ3J
s95XQEKH55FXPvtTSJQ/ReMIXjjZwitMZZqg2DqxIjdaZkFwnmn3c8hQ1XXTRjRMf68gIuNo/Ys0
Pnoc915U5erfMv4O/P5B1jC2hSvnMtVfflhp7jjQFdjOcFkAS9tAlNAkafQBHuKPqdn2Htp+HJOh
2HYxnSSEshRGe/l1Ev5htL51ceP0R0Pni1H6rJpuWPZG2z8B3y3eUsDlx0aDil/d61CBmuL4/azj
XZNrj2cnQ2MjaUF6WT4ZMrydIHZNtHN8SeOvYpJQIlLkU+qI2N1wWBJOwq33/2r9VXBmvgsgjP6K
ts5je2Qo/bHkg1K/YhwQMFLPpspXpjaUsEWdlJyg3n195lAKG4i3vGe2UDX9U/JANimHW7aeTQI1
fWwobgkpZXRZt6A/WIk8soGddME0UltqdWFvMDDkEG7V2RbywSaJtMVuRLLBj8+uNK4ZZYmM6fcD
La8crBk237sTyA55Qg9NU89GjSpHcvUKjd0HmxkmKR6moCUHQ301yD8NMNLlec63ORrdOAekuvRB
CgYBZWz+YlZO4x2cPYivB85VpLn1+97U9wW0VVqUC0UpCBIYWMQpieX2Yp0n/esMrgoLAb/JStjX
z1VpOE3B6im6bgHfoKqGe3Sze4blxEsvy0ShD3gp7ULrWa7UPDqN3/5nQOCXYXaQifDc9E+9N4zo
L34mM/eH13BJ7Gpqzf9cVbXxEtqrELKMrdZdLEd0kjA0V4CaUHmoMOiOCQ7XbT8kGU5+YUElQW07
PzF0u3RE0mbLm7kty3SQ4XnVlZpW3ENY5ZzblxV3yKaBRsVwK4BOQsU92qxITV7OREkV4jtyH2Ya
+Kj0yKFNhLKJ0kHviqQ6XVq472lWfo/bc7o9OwyUyFRAeM4i9+y909PHL4pZnhvjMAaLaEydmNgq
5icMAsxCDz0SO47BHLwzkzvuVnsmVIU5iD7OGduVybpBhgeGwQjJkK1E1w4NAjeu9Yud7Ve3CMM+
ejrQSJKTDa37H1okPro6hXoA8c4pIaT1r4gp8OXpWTK87vKHNyKSpBfY16kNo0iiRMlSvO+FVdKS
s9yg1bieeQ8520fewODwUuVyB5ruKWhPg2RxnbryGyXJ7QcdBUxI02wlt90nKRMsEHETuOxMuKH6
x38++GwAFcvgP163qY2e7AUOkf2j/dIQO2n1X6fShR6ansN2mk2X4IY79eNIAVgXbuXHGHqB5tXR
AncvfkQTWdEw90tbYMuciTWQvlP2wSjaVu5wt0SiPRRNsKn9mGj1l+5mj7591y/v82/JDvqnK3lV
u0BGsypITtFJoEM4dwf++35TL7S9IsRg5RNKQqIriMD30I1CmCdRlR7UtTD994XqbVyqyy3iH7hh
Kp5R+g3u11/VEmCGov4oVRTWGE+vuFXz0RbByJZ9+rLGfabOKSnP+X4gBpiJq3nBKnyRtANkXIBY
oVR6AWVYBZxHB6Zp10bdts8xoaqrqgILKfsnnt6XBvuwToUHJAnxT9u5lBWTPg5hTj1BhpiMfE+n
Fr/EMMtQVTosPvhDqRyCFtgkgP/KayXThskZfvvQJWDrb4BgUTKaZzEy8yVLkVbfSJMY0GQavrYy
ejwtDwislEsGIIkPrg8RTJqOi9Sbx01dmOxguUt3oW+vlBwmsFJEh9gR0fjAjBviNlEj/UEQvLw3
SA0LwretSl8v5ck/iVch4r/yuYJC0JtUoVmc6Wo3PCSIpKkh+ATRkzZ7Tl6r6IQAuGnD2v/Incuq
sXVxLUoJeVwkOU1YxjYBS+HPBOAAEekZ3zaRsh+2k/4sh62xu3tnUpPmH8Q5lWCDFtph/NHIWR0I
DFj5Q/9GkfP+v9g3eBo6mMyISye9BKuLunIlTOG3sVd+9HVzMGw3D4GuufAo7Hz+FkvJH3v8QXhq
eW4+M2/sWj35M5zFkDUqXuJ5xUW3tHWuGVgO3AVWx2YX4NrRUAZFxbqKkYdOculGity4xOltZUi2
KzGVs3+2DotC/38Ov6+RAoNa0u3pwLZXshtqf4VC+LWn3GdTsb0MNG9iXgp4PCtp9P0SoyJaE5tM
/kgZ8p+FpP7ZKNt+jbCI9/pJaTIdaltiSmWU67V2jHIr9+KPLgh3jqQWiEhkJpO2R0JG6q7hwJBY
0muwKeIMl+6dmTOgotgtvLuZowxiSDhK3F3+6hHn4CASP8aSCzHIOfMDAN07gcKzD9Tmd8Z5ID1a
KOADEd9kHnD6vmAfXycSkaQU+mptXfKfc5ITC8K2c1u2TJMUABLFrjbLetnQG9lS5ZvnV4VgjQRA
INgzsHkvc8xbxH4BctuFWRgs4fguCMkSB6+Url4zYTwE2qwULmHHYlRZB1NjFv66gPYDfZbzez1j
6WRhaQuJzHN7XV+8lBsG5Ihsg2J0oHrNG+qwt/MctkwIN0Qt5wvK2WXTI6A1RzoBtN+yUPHCq6Gn
AwsXygLr7Ve/aEt5pYEwzbsl+j6nFtUJMMRKlLMbb+fsTFj9+Zywg0nm+KTXEa9r2yLM2HXlHMol
6DqELCk9gaezo/D2GGwTkMwGWF1lDRAoMPBXAOhE4ucaH/NRC/fr06DTR7wjgaj1SrMPBpPOrHsv
r0YKfv6I+Xgt6t4WqgZGBS1xGbsraEq5yU7oHwrLuf/JiEIvVUtawX7iLVALZm8/bI4aYKptkerv
oHws4uWypEHVwD5qWxw5lAONg3hmtn6xa6uofcWEyPO9C0pEVYBwYEMxyFp8Xt8WmHP1FBBAOuHG
14gwT48vkRWLI+hNrkKERfB/IYJqYfsUJn0kLrCtYmfFr48zB+dqloob/Qb3itjFIv2hAHaGiZQk
2LmrFrS5arYPOQaKpFmf8qeD2b5WxglsefMOvR18zBQsxzYNcbGHTD9SA2njJQdvj2ysZLL9Is5x
zvFp+xE9X/oXk2sY/26AvxEc/IkoyrGfPCw2wMmbDBgOLiuoto9iCZOUTFrXASY+53Cqo6gx0AM2
L2FND7nGI1EOCLdAxIxdGFNB439Pzgdn59b5mV91f5M/G3sQwR6RIqVqy89nLkRciEK9gSzbiPj3
LlrHYu8aR79dM58rrjx428tHDnTQxiXwqbZJNoAgAP5XKidKjK+6UKMKKoVerpalya58aiwcv4aR
GdSgjkCX/97TY9KBWDZPbJ2lQFz9fXeaccOIHfOEoqF2GVgJ1E4gqgDxQ3LrIMJIV3jtXL4cXehz
mD3wC5sPOhbXI7/d6jyzOPE2JrmZ4ZmaNSnP5fUhSbZsDVtJCIQxES/5AzaJs/XAGmwCV3AtOAOB
GbFHPRic8hK/Wmas4T0DX7heSyyzbf3IgfgKhzPbbqJDylIeYrs4aVrviVN+WuLWAQPC/aylupIs
PWLVvtnYRAUbt5fwZj/X1+WPFAsRfOouHvWyslg4Ic98bPFMVrmxIH6Lkx9cb3OiFXX9sq5TbF0R
hWDW8INQB81hwz90ZmjLxdLf0PBgOuddEdh6Cj/6KUxpukviqbSSGP+lHzDe09zw4qbMou7S/tMK
VZZH7jAdC5b/4ntcB5yP5UL9b25jOopo8A92gpgbW1L74E9LEdw7tScuynMVtF2Wn20Syc6L/7/O
JHyC7uZLEVKEOih9iLj5yGxsaE2OYhMRdOgWdX4/eFLk2d4OSyE/kdZRjL7MNeow3CElRZjpYPQz
xRyksBrGICfI1BZe3czSvzeoVOF7JFauBrVg93Suf72OiaRF+n4HE4OnO3txkNjeg/8Ut43qtRow
6aj6awOwgJ3OjXg+BXQeqlRDwXEPHO4Px1U15axqcXtAsSCCWJaSrJsiak6jwFwvor86mXx6+djF
3LMU4lxPg9S40M14liytaml4dfydd72Yu2wqOkH0qWD5Q8/tLMZBQxXN9Z6ErPPzAcChtiYVuJjM
ZpCbBWdDam4hvTE/tdQ1f/K3t7BOLtDANWPNdDvuHNkbO9U8HJpukCkajmJBpjkVvXI/uS2gCLoZ
NCDo4KeT2PMBI/NVrbWeU74zy1Xm9DeZSq0p8EStCrP9v1n9Dnl3LICYa5aCOvKJfGVUYrsfI1Rt
to5Lr4HyeskI5cB1LLd+vgjo/WKklLhSPIB8izm+9fdMZQ0Lxn4WVqZm5z0t7B1vcKKm9CQ9g0kd
43Xv1t05Ksy9mwq1jXfxfdjFvfWcFV5aa5INVOHzDQvSLMZpJHsN6SttuT0eWrpGPc50ySLzaZJF
alCRiPULAWrMR1SBmUld4PYv2azHOy5elvFMsHTiLceyhabSOvbw5hCeWqt9WUboACP7hCVgX2Di
o61s+lovase2qEWeO+Ls51+R9FBFIMnwrUsPlEw4uH/SrGyZN3PkBEgsrSq4Qi55htQVmuOJsF5B
yTtCk1cVHJCWEk13pBsZa+agJk0hDIm1tWThrOlzeGx6lE/b7TLreGmPOa/SjSeGsxf81HJNX1RK
eoY27CouZnGl1Dtu3HW0L8J4+odjYpmm93FIlUERfXM9OAF0YvNCwKH938aJZ3dc9wXMDux/RX3R
W78IgtbeoMf0v74PaUx5lLroynELSJhSrL8Dkx6WCRSyNeTSG3Yuc6uLvm6FQaEm4o4hNa8wQ3n8
oWpuarFvdlsLSS9CZG9eri1TSdsR6QVU88QaLhtllSF0p9fRkfLiRjuUI30egSWA1bN3Un57MAOf
hEtNZszOiWfTF1lCkPmY3ob5FirO1k6LOm+MBGFr6dSjnbLQqYHsfNhXPsukjx0BDxRTfnB1E3kY
ja/g6FwsvzXJVKVCz9goVNwFhb243iqzdUHTm4wPLo2amZso80MQ/S5wc++Xrftks7wfyIGKXQbh
8CFzjgkqo/z7CHQb1NYsOtCpZau58xPGbN3ptDBwFH98vy7WsEe4uhersyu3jpBnDIqizPNrOVQP
cEo5SwzWoX14tpAe63cOjHkYU6oFQWg7lDU3HT23JgRqReIeEdAyJ9Z1JZEDN4392rI3UmKI6+fO
LqgQZ0HVSHc11hZjpn61kFtCLbAyHCqK4BnDcZGrZEkkmfAn1n0VCuOc75Xnt8EwLAyreR5oUTtk
YY7ekvsu1d6MMdRP9KLT37sTJA7whhNsF1bLyLiZ5Y81P8fuk59q0vdZK9C3nsTZlmZUXvqFQggs
mndoUSY0jLqAt6h+1exUKu/B4CFDzyqAUOcKm/Uq3+Why6R+bwTecJ9rY8PqguThAthl0PhhPWJ8
0joSgWTb+5QyKWR5QUFfVQjnvIcS4WhlVA581cwG1iooAJkJ+H8tP9dJtMzBY3mYz1dBS4MQcP1Z
tRQe6KBdhxJLjC7mLObgZpUMM4Ecv7pxMHRbVlnLIJQZW04zqIZ6fYgF61scyjf6xDYB3sIL7NHq
L1evt0LVGka2RELvvd0ThIFw54rlhiHUanJ9GZSQqg40bprmQfJwMzOQ6fyb4At03wrXehOC/6w0
wWSeHv8w5V3StpWWNkSz1E0EPFin/mV/RSb1raXKQ0SsKHnnQ8QCYEptoLYTQtQT8XJnpDwYezTq
Wd1u2feIPGCuRZ7rRtJPxNtSDJxdkv5/ZQabvE0kA3hdH40s7zN/rey7BgQWhfo3LhkzvdW7OdFh
SYZ5/m+eGP77plzy+r28sstNQoH8KyMi8E1wNPvdT8jM1T+/YKLXthbpON0Jr4UbkOFnUuycuVaa
hvWNKp/ZPDu4ZvzhAS+YtuhRXBKcVpxo/0wjHoRlO0VJfvSfBwonCCGZ1f4gSJXwDpSafNs9Ait2
f21uAepKgKRDBjuc5ZOHaucvNMrynpRsj1dpKjxIwx+FZDAZbQD7FRsAC8HubXpnJ/E/nODNzvgN
fzLaV/bw8/rRTo42ET4wu+5KRdAbKA9gJCV8tjYbyA5yI5fF6uEzrcwNUsA0KaxdCQULxGqudzEI
ahnrBWKdEaRtaBZu55qXPe+qDc4FirHuubV7YoxMszacEAhCaYjD4y2oKH4GWi/WaS9h/+CsELHb
v97ltQsfbFrv+QPg1Sl6AfD3N/GzXIo8m4WpJAQEL40HXXESeTQkdlGkX4LnF3kzDFHERAIfTxqg
MNEaXyMBewu7qtg5nv/Ril5j/5jP1nY5VnzIkmDr50FPM2n/lZCMT3NwcHHeTpaHmsXFVC7g4EQW
b3XlEAReYn6De6kQr/r7oge2y2H2X2xrUFqtes43j82TDmWXwSVqXcTG8spB6CnzpzuHsJe7YHA3
hE81E55xfPBIpgHBqzmaXvA1AvrdwKXiwMlOjqALIsaOHQ0GMZwskO501PV1dlbKZHDCdMcPoJ90
KQAqMx4OsKW7zSXJypW0yZu5dSJeYhcCZh5d2vJNRW4Ax8TpUS2q94hXQ5QrTgsioAV2rrWTwxSH
H+GBnRGk8HOVeDVrTPn18cZU7/iR5+EyVB51rECMqsHR0KdnMLnZ/ZUCuHZuZKAsGqYen+eSa+Ng
0VkSmThdecE1az9P7PBf8egRVcT4eB1yshozbCIrw910aNeQHLHcmIyqqNFasVN9ryU4OeJrcY4W
MatG0z6xSwPiR9XPG8TKFreQYtFfIOVmqb94NQ943BHpoeN0YsvevAq99qtRh1HaagnNkm3Y8p9r
YwJ4vgshMF0/xzhYnmurEV0fgPicfEq3eGciaUMJP/pVt02etmyPCQtaA/cd5OL5+dJ+aHx+0YqR
0AvBqVz6qbvuq647dcf4weDzqh2qPeBPl1t+k9WL0O6+ejpv20X6/OsS7rD0pZRDD7upEePngiKZ
R2Pb/NOnVtgaPzpHqRUJbFc5UxFdiYa+g8Qpts+DUnhPzoturkQOA1u3j5m7z72NquX3nUSGXuPy
dn7w2aTcFzOCTNLRr/m4TBltRpyaDSRLE1hImYl3cDKcMoJnY7L+fiWm+dwo7gcHd7veECRcJV26
LE/ycWaP5pGeEOc25K8a8JCbn8bCC57i1PiUrtbLCYcuEtsCt++R2oauCkCOLEXZy3m8T6I7xZa4
LmLWDAEGYnUkxV117zu5ObTscI6GqPup6NVMdMpMJZ/IJruIMWpc8FCimYPiq5vnDUgESscMK+Kn
Pn1LRopHtWNwW8h5lUl8dz1f2/sb8KwefVZOOAYdLT2aCLsJ4KMo//WxD19O8VezPaCpuflUCEvx
CKWD+cco0RHqsC8667Lr52gXl6Iv0myroK5gZEIVjjYX0PHcdSqgecvkoPAjgoRRibbBMetnQSMT
ogF5NRuPeSuCthTThtxkypVoM6AIjRfwTh636VUrpiGTcKd697NJPudTvr6F2CgYI07IHaJpD8Ie
HGhNGfDh+3aVHSv6U9xHWO9gQFq4K5ChB6KTCs4KzkFahcS5ltrFapD6+W0ZJLWSaY3XtWTDb2A2
ge2PrOUQY1i90gA43Pliw7YIDwT39wOVQwqlSF95hUXStaj2I2SwUG99x0/Xc6dhCgIlbtOTR0R1
AEAkJ6vZK/Y39Ge+ZTvFkwA34B19sSjfd58SwJ/FH35mEVIDWuoPAFdy9y+VCgfdrLVtnWH6r0S4
56c1MDG0UOZwRghV7P5sFqxu6fQw65ecTWajEPujOea+c7metnqScAT1/BT0CAfTcVbisI/upQRV
saXFoXlsjui5b/lsvLgcM7BIN/RSzTUkBgJmWk8b31DgaSTx7LEChsbJMk+gAPqF6fLDmw5H7EPw
jRFJ3RjYM5lOJ9+Aq4NWGxwwQ8YQjuDw1YMdKBGpPysKnTpUzfLfKYhEo7K9mMN8ZRWxi0zC0FZz
fyKO5xUiKwBfSZYgrA49oBlYL3XwKXVzfAMiVFV3kKZffHZejUgvBg9MXzmPma1N29egGQXKlP6z
wwU7J1fZhe2iCI2SYjn589w7lQIFwbuKWs50S50uonK6NZ4Nfhumn6vR1z15ODmCNW3KlNBxTvJ+
KbbW96WBzV3umpFEX7WCXWcIiAWXDELuv0f5xWwEva6nCZ3EDdS8ZOj+8KWGgpl5jgr+Vu9hsyyC
27ro4Yr/+RRrj6UhSNsKnHwKmNeB5QES3En1nD7FzQtRESzU0a3gwTLpu/guQ4QPDSvd180A/Iw0
eUWBwKnCh45jwFy2sSU4XA817u1xXVluR6VEp0yBQDWFyqfrk68ZcRS79YBVkevPCX43QPgBePQp
QviwCG7fdkuDkOQVpAOE5e4ye6GbGNT0GJmhqZPkxpPGJj5TfhkB/SHbzkVS4wze0ZVjb1wQF9/e
0NIH5XUwyfHkj4pHy3yZ1U+aLYNtPR+u4X7bgQVWSP0DKWntE1XgjlSGOqhB2XxQ9PbULC2Ktb7P
7H8mPB5C1HJZMbteyW5kPmvi+QofSBzxjAlzveHscsegJzOKdrctCmJHiv+CivpPgAJponGblqS/
GT39w+cCK3WpbdS7PFj/yLFadPVXlzup6JHCbJBU6eHS11W8PzWAp8nGe5yvV822XN+fT82lSHfA
pyz8fZWwQSYDCceAjqiAjZkqYVMXWQBKYYvrXzMEf6NeXaD5ZpPOWKJ0pvyRh4ai7nYjFgPglASI
mXcsKwP9m0A+Vf247FbamV+Snk6FFW7dFMJebArInAsbAdlp3vPN2LXS1aUjyhYUZsC/W4LFzeP5
IfmgGX/VaX7O1dNZ3vs0nonDBb6T6VkxWiCxtvg2Ph65repWCfv66LXV3ieHGqd59cVOp1YzBPQE
UPnkJecFpGqsyUd6ZQoVKyULJwZd5Dn1T6jecXBGjcimHJtLqXJXi4v9ZUiP/cz/dlQbGEJMup9j
dkwUKIsIsEgm/jK8AXQCuANC5m5A9d6ANk+3AwyHavIDSCJcuphJ3KXB87/cXC07aOW4QPxTEyGl
Y7WhqTkC0W+YrzKJyPB89j36EZNd64SEZRmSxCHQyCmR1jXgFzXWo3F9Oar6zRfcYF1HS0nRrv49
JDAYaxyt39rwIdi578eRG43J3ogefWVq8gbme1Ot+INUPNmxu59vJQsTqxma/oBvd1ANXduyeal5
sAFhmGDUc8U/3LUH6wj4JzlcohEWvAzTdAeQgviUA7kjFbXpKwdprGN0XxF4W2pEIBMt+gQvLtVu
6jIpH9SFSsJFI43oCQdKoGysbVtZZAOZuun1441N32j/lu29N9UXt2ORig8Sl6DMZcpUdMsEf1/c
DRPuwRRJUPMqHsN70MuD1y480Ymvsm1WyzwqKBHjOSQ8CNAyu0+Or424mldY5aYF8CcVyIc6Je6c
aKc0a3K0IX4RzdQJ/ANErymVRtJwU+L80Mfi8ML0ArgxR38uKaYcPpzFxhcwFFFq3MTgz8fqZuno
RkbQ0BP7fpS/M3UA66JcQUUMblsl02P2iwlq9hoA5J7DDv9is09oRDR0sSONiuTydeBM74O0+/oU
N+7Brcy3DlKm4yQkMvAVNgiyfxDs7+GF0kdm5adOlaRM0VkN3dC1voc5/teti/foGOZfQeOKmVxB
ZAnmexqTt1l+V7YRIQl50Zq5SsyiJS+7ECi3liLH7VR21uWAQ4Jb0VYBKexXlmDvz0H5pWGu9dHS
vnbrB+0OielcWFB7/aSYYzSM8NT7sZ46Y8SG4hZzm0fGFS+Q4ARw4pf9nZiFxj0l/AD4PQnMoFWh
iBDuHH0tyeVPwxOg6XFmTNrsBrN7FWDhQPjHwdAHOWaNo8bmuyLX5s47my80/yPPR8bsfB8eJuVB
5ip0NNc8lUr/NWXLToiYJvFQuelKi0eiTXcMFPybxNrG0/vgLgMOOBhve+HL+7AlloiHruHe+thc
VCkUir/VWxOUUbKy7JDDrvk44bR3Q5JESr+NW/FPW4UUnhKyR3rJ0sb/BkZ18+wIXCv3vurPc4EA
chn3LLlDYzAczXMNbUqsJvcd8yMPwXi5qUxa/ifhi9aqcP9w1vK6CGreTRPJS/NGt6W9GVohWUrc
D/Hua2BOKs5gjvDVMafs1DKFsJ4hfLXc1LyXM097vq87y/KoY9T7DQi/Q2t3BXD15yUq/ChyOMHQ
5gEWRFm4v1nri4Aj3Ca5KExKWio7L71FE85T1SmfbW/vlH0NQIRvw8lTsW5yUWIlpHmjaCmI3YHv
UgZ1m/2yrfFjQzCBzi7Ya6CUb1P7CxglW0l2X+PV7e9TELB89D5y18/ziJmcyCiLzR9ImhiqTOXb
FFSLL9ZjvGByzh9n58Qjw/HF1Ge2zkL3xIQwAfDzyW2g/NBFvOdD3bnFWSjpHYbcjuNMMOylegJd
F7aFyd6P9/u7sjZFe4EHzmvB4MlJfOhlV2jBAy54KXrj1bWaaWB6f9xJInzg+bWsTxaY8hlvQMBB
fQ6jFwn5buNfvHHm0oqEg+m31fs7WbW9Fl2MwRBAo4+TW8W4/A+frwZKtSneyO2Y9DblSBCl4s15
7/z/YW7gBkCDYl3mZigwfvySdNy/QMlw8NPsxgg6SqKfpi1d24/xJnIlub1JeWUPGrjboZOX3pkf
+XH2sRdafBLXxC9ChThKBoNgP8QVrrb8Gu78u0+kjDSmSufKuKsK4gTr0nkXSUjnOZp6sBoE+P9M
MFLNXEk4A1UslUPawVeoFP9BRcKtPku5eda8qhNLHjrqGeNZmKed9qXpDLiSfZUnX9KQMRwcgjvw
VD/EwmlnEzFSYb5Rz2J4hseGU8bUlJ57SWGQ97u8P7z6oeM7KIvAl1uqDEeMZLix6f8BBrsj4XNn
MwTwrb4uOdi8oVmAenpgFj6lHDxf4abhWUF9R0tq5evHK2LoG8BuReDJdgyD/F1UhR7DdFBPibTg
Ypsf/fV5GihkYH+fxBn6sUouf8hpx7wxPBY00PqGt11fjwSjZ0AsXiVszdir1I3egw7VydEmojA+
l/gojglmmCNEMEeYuSMb4GzlNA8S0Gt7m1i8CuvJpp9wteNYOlEyi2hWW7lWMFTgNYu0l/8hIV6R
dYU/7IZ9c2mahNI95Yu06wb37OpINbYkyJTYoMlqxgJVlzhEaJa68xx2VCpbyFoNid8x8hptL/S0
FeSGEZFvh7FpXVc93kIdI9VRY2T4RPA44EwOKk+kN7pYzx9PD+bU3jznFPXStY7kl3wtsgX/7vy8
s0QZ4oCGmyjjXc+xKUnjMyeYscXjDdvPYgld+JUF7zVL5+Ldu/2PJqmiwOrGQxIKr3kzMIDX+paK
xx7UVHS7y7WLuvfIeku/fAgKwmxT3CeJs4ad5krRlGUsQSQzHth7ML4hYo/KwAeBzRzE1aG/mCBY
uIZs3UeLo0HcwyJS5ssNOeTqlRaSLi/Q79GsM7jp4S/RBO9rKFdibCfJcaqbO1hWT9fVA6paNAiE
u4ZoMrcpm9zf4JauOEQNeHylXZYJYRujTeFWpyH7fhV9Ndjcapt2GRROlfAMmtJZD8Mb+ugUxyIf
9OHcHFqeg8U7OtVhrwFX6huADPIB8R442GcWn4LlKVheZosR1T8Jfl9HozaiJDwiRpgGdtNJalvK
2QZAqc6+wcOXJnftbIR8Q7L6p+kmg5EPDHMcsW2ow/GxclLkk0mxOIIOsTmXObBmRHuZK8UsdI5q
FID/hA32ft823dmsLEl4++oQ4IBUmAI/XgJYA/cn8ztIl7j2rGDKE1qWZkRBmkAlNuz1FKnbP01b
q5+dS1sUazn6HqDgzHvJebREUh00OaICGXgV/XJatEGXPeBupytBoiZHKYTp8AjEF7vVh6mcmCHD
HYr34dtoU3ylGlutr5vsVunvyKMj6aNgvuf+w0cdkErCdEWbMzkTyFy0FpGPad/se9llmmqbBDWS
7q3s3fICQPBD467t6NgVkGLGgyo4x7rp6m4zyc3yPS42Oxr0u8nttA4szYRrcaCeM6IkD9YYyc7j
3RPXOCFjeFUsCumqOu3vodPqUVG3S+y6sufHPgbs2rHNAEgVNfeRLz8xJPfaVJJzJ1MjIGwIx2mG
gTjlAb+gj+w9qFV0hesDzcDolVue/naVl5POwLwWaV0w08TONoYj6xhKbt14T7vAiZJbQuZ4QkLR
b4vgUnJIZCIXRVcPLERhx5hxWk90GnpUVQd85vm7KmD+mfPn7YxyPjWbt5c9R7Z20XBEL7pMxT4N
oouhxDAgPbUwoxVNCn2EpWGyHtvLNtXZhIzzBba52yX7tSCxFCbCEItLWjLGpA0pTxgbfsDTJmGB
fXgrwOvv2r4MVLg7g0facDyVTcgYgU42g1Oc/jd42c7sepAnXEjAIVgcwg3RncDJAp+PofeRyz+u
Z0AuOuk0gmJxUnb3EzXx7RoRL/VXDR0n/vxbSCCQEvu7U+Gv1524PltpEamZ4WzAnW0xHeaiwByB
H329pisw0IH4GAONC6wKu3+HtoM5YAGJ4FGCOkBtbeHVKe6JEPwidXydWIUQy47Yb7gCoW6UuXWu
0fpVkD9KrbPZhWTkT+RbYaO3coaN23ENgBsvQY2hr3mTqO2WEMby3+655v3GWIQ8MTtWcstLtKpV
wpU+lx7VgeOjZNXEerCuPotZYM9Euo/DtkfeBlj5gKvCU9PQCAMCzSzCAJSqS5PK4JQB/04Bmsns
yfIuCM3QJhSo4//dNmRSyVeLkVpPziNiU274zG3/1nZyIzcjoaCioq3jdzZfHMMx9S309XW7mutW
w+6jcHjorODBFOhyVyy1ODaFiAhXXPT5edLAOb0VKhASGtkZCB437Fl1U04zeB6Ren2Yiep4avLd
xKeSXOxkTtSPmG9uXRiUqUdmi2uqpo7zKp6yAp39QrJmyGsWdDXOst+h9qoLM4APhyBuDlsXR+8/
5o89LDq/EQE2UQxq8g3PZynfctvX9clbO9khQuMOt0nVfF9c1E2HS58tDuWmOHW9+NKGyM526Y2T
ZoFkNv2QscvspTgCKTC2XoTb98hCG6c1ZYIzvAnkr7E8hAy72GTG+NLdihHGuUP63d3GY0LCuX8t
15nTgZtX/SbzxKg+cMVqB2rBJv+E+fy9Cpa5FLOEjrh+J7AllYv4QCNN5dVuZ7k2L134UAnUHGQs
1xCC6fA8L9beEKeQJoG9qSx8ONCUdSDykm0gCwKljn+i6PE/hZgNnAlt9SMXnmMGPSv7zDZtaLL6
XI5u8Ti/lHINYSL1dJXUrxwAcSWmREmUq5/HUDDYwSc2cVLv+v2eKVebDJbKRgrlEtElZa2Xe0dw
SGzintquUpIrLiUj8duCiA2Ks9husWevdGr/C3NNFhelD9fw+zKQK2CDJmnQbEoglbrql2C6JRfH
32fzlCbgSZjR1aUp0MeQabfqWIKLaXFVU+f4GHAbos0vvXSaxcToYj2ZPa7Mt5Sa/MKGn7OX+377
dc4RY+22ZsQXO39FQ5zDmYwyP1itR9aKj3bHu6uz++1s6MLZzoE8AOPvqLU3einFGenXQ7ttkBOl
zxXX9w3K/vq0EqhO+YZmS+IhR1ig6UmO0QuBhkghyCGRqQFOBmpZFU4UOzox3BcZkv0mgkQnTVBJ
crFdzaT5wnQG9Sv+2E6F4t+8db677uqhUSlnp/Rd5P6+Aq3uJHRv6KOFZEiMNwTSLp+EP1N1iHR9
Djk6rxuDkERWsgxacBFdY3mQToPxVRWTk2PkXNpY0f0lfT2R+RKOpYVknfROwktlk5jjcB+uxyYR
1u0le4ajd8fHs5QUzPFIUE2tmVrqb0yxFZ1nuesslH9c263DScumoO1BBAQXqcBGA/K4RpAaFheO
0hqQeAUMqAi2zvUnJJH6Ea3qgGkh24kbxj0d/vG2x6sBPF0/Qkn/SRAe3GUzPZM9M3sGyhQs1/C4
+D69+0VtmImJ3gam0Q3TKwYXq2OxEpjlkNd/Azrxj+R4VdLwKRO2IshG1wu69Ttkhf1YsJLEMkpu
MBwqmflx1duYinruWHdO1fP4r/9N13WEHuWVdgqIKjvv4AhNgseY68bPQTLD8GT60qTMdSJ6rPIY
cn0AvfKCMHVRC7lYR9wQrz/hOu2vu3oHtHj8FGmvesuunLOx4rCgpD08oGDqzCjFfZxMS4g7ruYr
XqEN+JZbMR+MjTyLTFF3VPZJ9eadNwt0IaiJTmMp9q+GypThKH/VkIt0ggJsqMDQ4v+lHa6qcKZR
vL1vLOMLS0wlqGHo6fkUqWMENpmpS0c9/Y5LAswBjQ3hA68gTwd9n/bsH3y43CGY0r0dt6rQUAyh
4fDYM/UVmwWVLdgkEtrn2ClhUq3WRyD6VA648oWlvQ1V+M1nnic2QbGrPMhmdjC+bDQUSRkwcPiS
x9IkfKUjyxHJNtqnNDnD5PN0Abm9cUELzgCCVCvkz/rmVpsiVBb7xHUr/s9duLKkb6sUAwDoOwCo
NoguTSjSnyLyGiBXsH5dCkhsNFLhFAEgeIYmdP0hMJ0wzuK9q12a4qFT8Z1MKYTATMvhVMQrBraq
8IOQlfi0yy8o4pOxpIvivJd5710XteWiJM7gyfgtj2eA+MSh4M5TzH2UFAgt3P9JB+2js9Ni1h2j
9EYAPTbUMs9+WPI7lUMesBP8Y6+GFaVPyu9/28vobWm8j1TgflZViU5c7/FqETQk9WETT6cXuCZB
0WpbJ4IYgnhBJohpd13lfkKnGG7j782QEYy32zRciGaTV/GqL6x9RKYIBbuyjpFNOuxTQrkCSOoT
/p+PJwJyeEVRE3QfKYESJriNiAXVLyhScEm61qXO1RgFQmyCWqjA3u/EwbhRAL5JaZzbKwUuF9Y6
J+x+M2mk9VDK3NhByJiR4S1cfuIqvEHSLagv1PZ93uwwZPo4m00OYnTsoi0SY7OOxrya8ErCofWT
sOFa424ZV6itNm7bFsystuZShw3JUjXmUOapmX0/BeEd4IkkVD1WYzr7cFoyyGEtCf2q7Pr1Q5oV
mK5VFUuJO+aOKMOKTtomSefV4mqSqogdvb6YqnvzQu/OuNzDPSEYbk7OUW7TRwh22IJVUbaLlrd5
o091gB3P17DmzLMXGwr9jkaUDEdLx82jU1zhLcGuDGS/26gNjMIj+XHEoQSHYMRHqMNnMXpyCSov
8W+jbWLpk5ZTeFFNWltG3mA06qIDJ6EoDhbjmDFNUnQJgv4ANKcvcqxbi0YaSwlWtMSFtYDAgjD+
liDSs9j7ZkC8eOIsy0LNswuJ9YsuPCsyUSgAzhNlOf78YluTh5p+3gShBLI1cvZWqdXiYmRRHTqe
gKv9ytQsIbsh118Gh8SlGKyb5fXJsM2n9/+8LF0cj9VmVJWZRmZOaseJsnCq10te9VUoTX7uydJQ
enwTw20eKLYOpOl4PzuzrjV69X6ci0IwpbpUnXIfbAg/YGiCoZyylDFcu4BD5FCRF3lxZ0WStQnc
P4phsJXHhJql/8tBa2hZ3nX7LxbFKtz+t9+KRlPSYzPxwQXcD0danKoxr2wSHHyOytlaxjdquke+
596RpspzzCJBLbvF3Njq+eIE1kXY5ZLuNeyunK4AwHa4jVQFZD903LmIs6zr8ZDS7MgSM8kVpDiH
A67sMQ+kbwkJmkDGV1Nk4cWBYaxYOpG5L+3ABG1LPUx3JMpTWwbk7LeAxH2Af+52oV3DTjk+SMj6
or+TUcBp+W/Y0wlxYYrKInbv5ri9mH5U6171Fl5XQvDC/KbKSwB0/66tPWTprLQZMB76NJieDghu
p6RQBAV9tLczcxPj1J/TAn2bWFDqpB/dEyfN9jAqAWaRyASpKG8W6srpP0LLxdV6jCVHB7F6e1J0
WzqjVCqTWb1rgHZEkIdM5+b7J8EVzvR1x2qiXRsvahDcO+GV51yrEDxuDoGPCIFqdN5w4HAm4dOB
99IO04r5mbeDOkYb1S1/UokVt1d+gx/kfYaWkzU162rutVBrLHGFPTp8jJ0nmftG7ZlA4sO9Hgj6
D59bLZGaGp7b1trjqX2LyA+UpG5Td+IS3AmyHU7PhY0uHe94EjgtdrRGel0drD5r0AB/8rfmoodI
UhVfv3W4N2aPpRINJkiDBC/GgBngu0x9WGY9tSLAt3sBxU8mm4nG4L3j7OHqgrhdaqH80SRburxG
+jEFgQ/VRP/bTtL4u6V8PWKYqOgc6+xz+Lq1BzY839QrjdSW4bOyEe0Q1aJ8KhTozbcKQ/f0jkxc
uGcaEaD2zpVPn1NK4Ch/dDILco+dfOX+88QTwoMoM2Be1CwmL83UiDKDdhLpAi9Y4XFJhGLs6bqm
ynQ5l6pWUkETxsRu4leU0ezHlZcdakSW1shsbUl1mB0ZcDqinFqu87U2cpmxOoArv2kF0VRIl5vn
+s4mVnQyHLcz5Sa5WVG/YBjJYGl016bDqC2UgVsrjB3WkbI9jDXQvJ/x2EWoxP7yJU63iHsEr9Je
w8/p9O4dlP6YpYa+30HVca7ie9jJ6Ozp90UPDkBHIulncV8b7ZRo+cBxEgwVvHNo2BnyY+oT2DNt
81CdLftCEev3b55hv2VtByL3dcFJSoJM9M5wC1qO0gqQ7lJYYlKsBDAohB7DS+B8UStauasI+crj
uqo4zTTyqWrEVW39FVIK0pw9w/t0/lv3jclQNFLjV0Fv/4sNmOX6vK2PII9xZBZUw1hrxSz1lynx
KlaVtbFKTThrwvfYC1L0z4dhBlzdVxKAAtGQHOchJazqrQ5M3f0mm5Wd7C4YSbQZtCBwqwtBOH45
9ySKMKa3bV9ud+ERSEV2bUQEcMIusANQ14IRFiPTCNImFjuQDnobh7hY2lKEwXHGINiGngZ89W79
kmtVKcSukCokdCefm6mZxgzSx6P5grpf8EDPfJ19YLSM3EkC35kspuqssmo9IAfZVl3fP5dXmIxJ
sny+Cb4ZPDvpOIR5dfeSYGWeGtJR/5xBIcPVuvWvXLRKsmWU4bcQwXhHSFiEvKfVi7lPBkaxOzZn
UHtpYWQdq309uYS0M3bHgdkJ0HyeisJwU8ZWC6L/qbPRkPyWGIQdlrbX5h5EUMp9FhvZKc57kvBj
drswj2Ds9MqRFGqc33z4PbHvffBq1mfb1aZyb01wcN/5mSbJ0c4DA4arF5AFp1VVG84MEpvN3iSW
evdYYmcpwgqJEKCgBekTIlARwdbdWwS9yXxl/jihViRgnle6v41KwR9qfOqlv7yLs7sNzt7e8aoJ
XyIvl7QhFiZrwsIRNvsAuVTIO38bC+bv8RwZdpR4gDqfDH8VaGirGcdKCqQjIefjlH5MIXDGBWZc
ijzAB2XKWfOrGhddRRNEz9qJPaIl7L2eGo1VIFX4OQ3meNnVZ08PTSj/d0FawtzZeuiEW0IbD9EG
KVpL6KOS3MKQ9VCJLBCzAx8AnXCeTyXBX9DUHATSYblHOgZv/V/zV2TdzQP/AwvsxtbP6jiM+Ooa
XtEeSVmWCUIIUHOVaclhCB6qXKUiMQRW60Xvc1LK4b1dmXrpl/eiIkRB9cXqtBCCxHo7LGxepvb7
vjd03NoVFcFVFHCIr8q0bZwJ5c1t0VW2nqShflO7D3aVQGL2Jq9GgZmUQdDCKManI8zbOmF8DUUI
7DCD9qtd4P1DBhI6tvddnePZx/t5oYyF+2GuZy/OvM47zyTBtFpruXMe3SW78ABujxiRaZfrisus
gi4wyKvdknkETI+m22vgJjNKQ1FIVqawvMSZi+l5TPe+cixwsWsAjh+wKraTkrqveJ7Fx93yVx5X
0sfPZ0kMEmEexELNLP2UJWaoEtJIvXX0JjceKLX2sQqDzUTg1FKY9l5EGmPicX/Xq22m/dSN8K4C
xUNt6kj5s4+ksuEgr2tv4NXgV1QWEl126Mkp318gycILyhPqfVY5Wk8uwRX0qt+QsVcUL2rdbrEN
24MPoy6zosbDRCzZyA+u8W+JXzL+PMisvlG8p1rmepYBKopxNJjlMKKwUHzg87ZexirMYoy/3BTf
n1Gw+th0e7vx0ZytYUxp+A8B5X4RYZYCkHBFo7pacAd8acZ7HgdTWTMMCicjJtRoqVnz88mR/TZs
c/6NUuhqYE4OQGIO4pxtd78YrLZ2Uxbm422sJy0fj9IJs773asZnLB+vgc28b3OFQI1SWL3yQAw9
hEFoiwBZIw/txnh96oHJFvNbwB62ntCk+NNCXnXWpjvVpgN9xy7G+Kyg5g/kK8EVgTiYjSaiXP7/
KwCrlLO9h+UWO7EdKYTbQgJ414TOLkqJ9+zEvE7miSc7VXeD7dUKjXcNeM63tfHRb0mG3+v9hLQv
vpmBs3cgrL54RMFZlCU+HxIpxcC15m6TX/yRw/EqkECeCDk7X/g9li3VmQw6KyT/kPg9UM1GjKy/
J23CCLDm93cOLbgXUUEeSXZdH8kRP/he0tboNwwo+jkiIOT8RPlHadJcHIymgzn5+Kgewa0f3lSf
M4YUE8PGBkBu+y/ioFT33XrXmdUAzj9cf0gew7N1vfOCrTL/MDYZTYMogRWKfLtSJWZiDyakPK+Z
4RawYjy/BTP8UaGcKRVzl7CIZuusH/Pa9PYtlDRFBJ5DmvBtlTwuel8dcEXrR7UYjPpTlHckbIFQ
KgGO/VEYnAUGidZcYEsMxkwqx1euGU3umbFHH7CdbkbjPwli6ebn+LZkukwWIbwrDZgbplsbUWCx
uxrOY7h6C6LzyRy2LlJJnaiIDn59nVoNRlvafAijV3VaWS16D3fdCwb3XbWC2PVVz2K9xUPWoy5h
LM/HrKLsA85m4i8syX8+TC/afAaPvM67drmnIGP7sHQLHulgJY2+xEIo5o9LG4THzf47aVGSFg8w
l5w49dSZeOyQE9CuXvKKluWFb+2/ydIc49g++MTcQn1aclkjYBEjb4D4FGRhU8lZtgagEZOejftb
95JZxoL9zlraMODOrrEYVitrhKUo9lZEj0wWZ9H0j6JZhNM7ko+PaX//tlUzKS5H0cCRWpmk3eKJ
/IGgUq7JA5Le/h3rKtkx3H94bqUcjNNKOzJRC78aTyRTS1tUwcFHd5vpq6EwRlpBKDi8uw4LhAM6
jWrbBCu4dmjric4VM8KVGseVDjbSyZDKHjUBkOC2ivTe93X4e/H9Jh0ohhlpayIxnOio0XQ0iN4L
erPOfGfH3s+IegLpoQ4p2tC6PgAGiu5PkrV+PeAKq4osxCzEsqUaRDEz8erSul1hDEC94WLaPvI1
6FP7Sd9pvvj87vJzrs4drGpXErHLn+5YgqRBc1a4rTStWkyD1o5+NNJnnhGu0xCVnODBKtFQj7M9
0rUfPReby/ad8VZ65dT231Yq9sw8rYrS/BwoFE6fWfGG5k3jlPik/AQHdTMGLL9rHBUndiEMI0EL
JnrtLo4AgQGSBWRD6q6lY2OTX0C0SZnNQv7iCaY1wBf2Ew+axQTP1ygvktT1l10ZeRwBfeqLC7YE
EUBpYqgoRaZcvVKr7IrtHoGNxeeSsLHw3Oo5tWFa1vExng8UIu16c4UEgfeHhtP//YoKtawGwJi0
beivYZ8nbwoj2TmE9yaNjLhbGy6FUvTok4LnHIllXd/oVWWkuR4923FhlMr2Ty5stmKlyvOrpbh/
M94q3Ix2RUT4R+2Jv6yfVEa+saUEYLpDl8U6qPxreh7FGFmSJ9SHgIllNs49TaUARFjh3hZMXS01
nT7q8owaiCHF1u92vSkGYMHtzD91QvB9BAe/9j2X9KTNRl7aMse+X+zmeMXrRXf+veEmatuS05Cu
Q4qarOb6vjs8yElgswA6t6ovWNXRIHTSRckrH7pLgu2cwULH/QtJrcin7dBfKYaR5jadq16KjVbF
wLBXZ7Q/5ULOBwaQWh2pswq0zbdJX2bRfs1pmYQ/kEvYLJqAHHdMSFu48PWXE0MYJm7J28Els42L
sO/073FEo2jHpHqRmaY9pRuFGdcpowiuPshD9VJeuFoOR303BpsAByNCdVh0hIIMEXxZO714zo6R
iDX/1ofPbreV/ZPp/u7h9g7eUzgq5YXX74PbC5g349oUDN4VU0DS84xuDW3nm3xu/cTYhbvrppOa
LcyJObZ0O3Ys7cHcDtfh8yl1sZBrQ7Qksh6dGRTbkQF6VJ1APkSlNz7V1iGcGH4lDYFFyqQcBU7q
srp4QpG0pytHQjLCTTtv9tVqthIRIeQWGCW6m92CPpWSzHgwJbfF4we9xfG8cm8E8FG+rID+fqhk
pVOnMnkapDVsJOHlBa3M2J2kV9yD4o+mYmYy2F6pKQr/GOLp49MJrwckqb7CRQ+Haph82wsEtOQl
blPdTB/fCZtWHYcDdrt7rQMfv6fxRofq9FGwEfJbRuQV3u4rcz/Q1uGdUMkNUNsoeioqM0D+mwhR
cgrgjMNACcz6gsSPYIRjOa6GskU4yA6xnAOmn6zrZX2kLson3AZhbj/LjbVpNOAfEG4nDNlc2AfE
ZaT5oK+1zZycf6L/xVJ/0xVQs/W07tmcnCFSdRTcGl5cbdOMgaP0b3yKkt8bcicI+pk0fQBC6fuc
gryButz9JZIo5awAbfsNSwzwKPqMEjWIC7qh6pMs9JOiuVhx3KRi9c+kXW8d0w9P/L21Tcj2Rw7r
9QfhFgQvoSWcvwpsrE9R88WrUlZ4IKW8kg7qmeOZlHaIX8//SowagYZUKoeb+IW515rGA/k4rMzy
XDCSDZ0X+tggJTGDXvKN7rFNtw6O+jXh6+G5nB8aS7NH/IbpSFZ6CVjfHsS7TXmrjqn6OOK7PWov
z/pK3zt+iJAWHOOGUZvFp7jIKQIAx9jf9RaYj8s28uS0dIfPR+fn2SRtjmgO8/gXt+vVMHkpkZ5A
pKsGpoxrUf1atQ+52yW5wy/+LbtvuPTUha6CBKAjqi6t+JYKgLggNuzWA4RVa32rr7VjjOdYTUKx
sJWpf/UhVqnIzAh+xgGt+H+YIlUxQxM0OPVedItW0a+tZJNAT2VQiwZ2qzaLdMxIUCMR0xWVgbXy
z27Bi4t59sC6619+vukQrCCpOZEyaFCi3xIftDls306z5oDIv7BUFFf9W9ovtina4/qo6+3il+QB
YEcssGU4hRk9mNvM/jlwyaourHOyXEEUH5JiAR2MYr2zILe3PDweuM5Fp4UV0iqO8q3H3VFeqGbW
ZdmgSAfWXQoBPI19tEXn59USRegAo8UCuAtVqDFVhkT/pW9NMVoWjkVfcZs0o8o8Q9FdQtGepFP9
mSPjBvtMoHZV8y8HZOv7xC7D5qOC7j1agHidYE0aN20VgzIA4JUKEEJGv8LzT0OoksguGfDYQY43
IuADrNlydTHiIntiB5CnjbvurlwYsFiHDsfP37sir85/iC9qcQUMI3JNs3U/BxBPW1oMDHgKB/Yp
jiLPmj5fbVd2JMvBDYqZ0jouRmxhV9G1Y/5kiz/VHiseWoh0JFaGGqX6pW5RUlzHXeTFvb7LCMxI
sGehmy+GGJATEyDmroZ8y49M5M37cjiybBKKXGmAuAiY/G2FIkPrLLjgRDTuFOZD7vsp/vNbR2a8
i1VcWjjcyE7HJQwsNz7uMgKk391uXwVKvGMaWmBUwTCWw+dt/bjrxpX09TiP2F5P1OMVtueA8V4s
X3RfsihfrHfSV6+ZDQilpD1+AzUzRq58RWAqW27F5Ri7e0fW3ej/ikgXZ4kqwtv5n4Enh2pg9rVM
XIYpmf9/u/0HmStoNp/pGgWzf7r5yb5Lnhc/56uaOJN4BlvW0WB2EFocscGMXlLrcmB1GocnP9/a
mhwxbLB8eeSS9BJzX7wUTITzvNwWCKrDfgvonIm+RUAo3XEKuG4f4b5NUdeW2Z8iAFnCi5vTjzZQ
0Zcgp6lQ8OPcUTKzyjosyn8apRILo2ZoprcuoTdGp9RgwaywoJ+GLxYbQPbDfCfUrchW1n+SfWTV
rquyBw3HrlhW3BS9Mas2BwwEX1ZFK6P9EaoxvF1A0nW6LEKRfdprWDAlVNsXx4lwRlv8oiJtsmkt
mWhRVGgU7P+5lssD0adcOEJbDOZIsx5bREpX/JzAyXn2jihOJh/nX9zXqKN9TaALCZCxGSglvKyw
fizPK4OWUPTHyjjTPpMbth89m2JfagF8vku7TH1otGEtY/mgdSPouopRxfhLUDUx6MHp/poeJYTt
uFtKBvtFU78zjIAknXSGDjSHy8AVpQlPGWGsm71AB7bu8SXoJ4V6yHIBaj56yYTr/tKQ3xMkoqFd
HCvVS+eaE9cI5mKymgZnmpiKhcyp3QpybU8IqcA0MmSa/L7B7hWjm40lbpMviqAAM05sPgoT5CpK
17D5ClIUhubaUtv7bBGjgDqDRID82zEKbBfDQ2gRiF/j02zPqNZ/Uyd8IsyfkVS0H7YY0ci44om9
QB5Kf9UxpR3ljgBm0RUw+c0f/kKX7Wqu65TSAmz/71CUyylsewoRGZNjaweoVqn2nKmjpcTkJFls
2ePbcsXDO3g2OY1Wmg266rkrvYpL5napGXJZCPYHopXsZNi2yAcpzwog24FQsdzneZgMO7b6wxP3
efUT63x8lmJtvwbs4V+6xBCeLWrPcRgaJOTkc97RyQ2lCKqJ5ouCV7z3DMhWGjiIYjD8wPApmj0B
V8VnNME+Ze4TPdIoLKzTLKenPki470VY+nCcQL5DehviEghXj4rXkWlgUBDbClh5ZOZESl1n+82S
cj9Qq+LOiUKMuEckwoiHWXx7JaVIpfFXSYZs973I6GU5ik07iJ4PdqQQMyS2D34fbYepMEF5/gHV
eVv1po3aBuPlItpDWzyJqhvhVE6ZCNEdRz2rTBRYwm5l35fzIzjyqM7ZKQQxz/Mj6UdnZayqH9gO
W+FieJ2PAiKYfqgu6OjvHgoxJtX88QXIPtbIZs37XZB3QfZ06vDhUIxcw3sX6+sIDORH5Fe4Iinl
CSgxuH9aYC4+T1oUpXzsoSAyNN/1RBRrNXiFni8KvPajYCa9SL7R7yEgcRznlAD4dwsLWSb2OJ6S
ABUN1ehFBrhVqezCag1ePZib0kc4/WM5OdJ2NXoPULYQN5/u4MrfAnSEEoNG6jNuFp1zqvMAl1f+
jmMdYeT5zDfClS4vwSCltyM6fDkENIyNqZzyQOKZP0JK6uNtFCzQLGoL9cDkrW1gaIfbck8YB9Hw
Jh2LDnLXMTgaJhNXukWSWdCRUTD5aD8AylLhHZ2cKn9Qb7g2BRHzRMYdpCQ2EqVrDb172ePJMlWp
Y5vUbxzsNSDC13Zlt+CNa0ZlnI5TAtkcCqRxxHWI+UJzF6I+f7kJU39M3qyOouezrwRO9wH265E4
sCuCr6bfEjV5iDmvBHqYWAzAihDzhTDZ4rtXJ7O95DDQexGeEpRX6k3d7Xf/zs6243VQegxhWTsW
fBd6roxSczqD9P6l4FupuVWTjBEiM+MCcOhThraepEr1yokzgDFqpWNlavp8aCtrIbH3AFn3KlsM
XLvqP1nGmxgIi3Z/NirsCrQzcDXBO+BS2fBBiT1WpaqLE/e6YXabgx+/gkdH57egZGb9gKy209K2
uvkn3xjFrfhoS9oGFYbgxwqSith67y6X/O+XDqDId3M8QDyK1DcJHnQcuYlktoRk3wth5MCQApKn
MFS4goPoYj2VG1X/8E39i/XUmlNWrPtmSDMU8lwrYQgq6UMSjuwpK642xBIxMqnOx1peABQsLf38
HEw1jGxND4Ov8OhS4fuNJv7Dn4s6ZcHtYtAzUK3ybIOIWAP4gC4Gjfbeo1eYzJFW/6gKL9lAn7I9
KL+H6LZAHiV0dgKwusTElqrK9/weR75fSxmeq1tAJvCGlTOf3AxnZqF4UBHOMzIsF3T+gMM996Lu
wjBTxVyMNOFkPmRu+DafAIykPycLqLTWL9Tfh9BJy76VP/4jVzch06cK4usEKgohrPGyl2eLueJw
lu0OipeTMb+mXkwMt09I+QxsQEi4x4lYmlzr6cJwdDCFzi0qApcJ3bU9ah0Y6pafj8aeMJP+SW7v
rfBQrg7SFYSXetVO4jgFs3tgdDmJDP14l1adGvKssZxlYRpmlfQY02MsGImWEjy8uMquilJ/tr+Y
dJRKbZY3vtxQ+CfU+H2hV6rXspXPWNpcCYzvvTv2WOxhQ6F4svEFCveB6g782tAVoeg+p1jCdetG
esQzmENte1HVml1fnrUxoX+RMc0ALkKFkEGd5b4z7xjvP0Xb0CIkD53FHlu3hqwucEEVfftDP4R9
BaH1tJmMv8X0GCF/RHadQVZEc+OtuhL685GngvfE3YT4KbTm83OVOkhIWvr/wF33pxi2QExxU41B
C/pQbrctfYmwR/FtBzGDm0cI2mesNUUZL4oSoN7VmUKZQ3CwnEe/k3TZmjKbK2L7RqMMTcLGk3s9
HfGtJZy0HL/B9Fgyso0xZE9F5HpdZHoB0pR7LR5czIEBd0BeNlaMT/UN/Vk+ws3O0Lh3RUO54EPo
dWo41MWTg31DvHflI1gm7HNvIxi3YvV84zMW2qD++z37aQWCK5pJRXskhYMvR5a78J1i6L49jFte
697ae6fwPBWmbphdPiOJTCPJTQ8Ip37BcQMPMscVSzu5ziitP74HmCvZXNxBoJ/1FhD3pzaq4354
Rm/+TtNONvy3p4nn2DigFIxs+Q0ezoNo8f7KQ44LejYeMlyFErptzz9VA5iDeYFSCFjOW1pGt/3t
qr6jPwMzlonYueKA7c7flcSrXIkrreLXjhxpaeSIcHYHp6SDR566n4hceHte1FvoMX3A0LpzInlo
h0nqQmzVMQbHZFbiH2w+n4uz4O6AVjwYIM10A4Sn/kyWHp5d8dWJ5vdPk634HS7daI5QcN5yzeX2
QszTr+oNAs9dw2LEh6SXwBXdBarfkqvtZ7Tvjd+TZFTxpNJP97SonEQJ6fOMq+pQfsqDnwhpw07k
l4kxQPReoQMAggU6gOen0dhSGR3U71KxpnJjEmkWRTuWhVaEeP3mCOe2FNl+ePMfZZX7OqncroF8
/9fxQUqPrdXjt6+G0BdEwR4nHqoFcWsRKikVzU01UEYOZek4rC/+TxGZRMGLKiWDB7LAhPoRxa3+
iYch6Dhv7bxifIK8Z9B4CBf/lOuDk/RPLpU0uai7QRmN+ivtkMna5DpVDZC+yng0QfgAGRby6HHU
TBw00qzD2O5noQEyDagwE5122iHDWFPpSqyLJjZ2zh/bc622spSCI0jlRezJ8SDlEIv4roE+G0Kz
0qvHw96W3Q2J8jO0qAO11On8B/9jygWyVC45fjNHRHH4S/NexHMsFYtkBUa7OU6ps4OIGqP3GsN6
DrIsl6YIdYe1582nvI5Iwnpyc5yYrOwkG/nx7z50wAydHiv5ERwt/J10jRQf5/uCeaNsPFGHSUqC
vYJxTvslPKLozVtTytjNZM7K/DxklV31TSteSFhi6fkcwCah0p0v8vNYtd8nxhglT/hrCLQ9eiXq
MpR2e1cYWAXjNw+1NztK/FP9r4xvf23iYV1eRthAMy6gMVL/0yAeiFJcwQz3J/RfRMnHhmz41O4Q
S5l/Ya8q0r9oeM4+CecZHczakpjL6YXhqh4oXrd5ThNE6Q/8mXqiMEgGio7hKKkNMMBPzPTWvsV4
jzv9/AYxgTXJFoXTJuavp/3AY/i0crsaH1PG7uwJ2FyKirmzhOOrxMbMv9O6ZxW4pecDfR1j0cMF
GBQdnEDi9/B7+8inz249PXE/w/iDJUjTq4ToIvd/R2A8vXQtCzIjWpL9zCnOKHtlEhqDG+Pi/TTQ
knN6rOwTUfkU8DnZybQWycY+uhdms3sL6qxqQGg4OFxa4wN6fE3ps2Y1adGkCEIy+kVFnros3dQX
PVfQUPqpMCnFujSFp2f2z1bwLH3CczCD4vJc5ydu3+Kr9SHPCtnt4uwIuDA41t8RqtBU5uyCUYYq
C9umOSq3pSrlt7/naY/lC//F5FntEnwcxgs6qtlXlzDDk/KYbhRX9kbCASPCSRfVMolstqOMjcxP
OHJG0lAUQ/Csk61DJNCwI4x0u3NHNPXDFS6OT6496i1kKJxQ0bCpg15W1P9tkzlcCR0O9lRAhoMn
72MfhDq2nR9VL4R3Kn+sHaXi3EBLQ5i4EnPr/V1VqsmefTSEPrvwGIBJ/SkVpmzlPF/9lgrR3xie
I92zemOBIaufqD/vcWgXxgKcGJlLw+NBE0hsqbJvKZJdyK/SU0RJ0HVHxiAnRkwT8HJ8JQctwAU1
N7aMSB9tH+s4OjCwWx87tjSsuMsnl4uJ0u3Qg4MpyCHLqvg7PUaqB3x4WhgR/Eu7UcUzwp3RdE6g
xv9J1MXILVJZHtdAeh9UWfgE1ZfKheV1vHv5+mTlNeUsIZ5qvSS7eeVAyH689WVxSXsMgMwocqHz
vP2+E2O1kd7Pk4f6Ok+SkHAFIMLBXRAF7UgWdWAli0obEgiyJx1ZmM7KOOBGxDjx3aMyDJKyardH
1UKUC5rJJn/xVfJSe1/vxjlmx9jPG9Ui8Sp8tKs8PiWEqxrW/hn/W+Zw3OVf9hA6iv2BRParNAuT
0M6WYQrPXcFUbZczAV3XbNnx0uBD9niV+6wcelVDVcGgeS1nOFnDCyf4h+pq5qPF8KiUjxsElQcB
p8BMp+BuQ8cmd2pb92Vkst7/5LYeSotz67YTrIn7o6Cb6ZGfUwbH0BjY5jD2Yh48Z2ggy7tHhrgE
tfKEZl0SGm7he0Btd/cjOSCfpxx4g71bqSrhj/s4fUGLkNsY0I1quxIeyzi9ITw5H3t84LLJ+JqP
xUbrCzzaIKccEsc9m+/dYnD7pmtpdr+UtuGgW8Z/AG+6LhEx5sOnr5uhf45zE3c5wSc8ihd2GJ93
3KCZuFH4RSam5+g4iHQ7XD/Jgv7J7DgiihCURPpvtlkv8wdDqnPMa6JW1DUE2kJ4+vy66s13IpNt
nC1XH9Ei0yfOTg7lOGf4SeZK1lAbczXWvehxkMcbYFO87FaP+UTUWuHl6EGfZmqntsf9l600MVal
pJ/tO67vCQdqxjW4CEcONV2yLSiFADt5zt7Fn2wc73GOIGk8dwxTZlaZmzpN655Z6kqzEG1KHV1X
2iz12hGumND59VXEDO/wlmIAvrSaKPEzXRhUXbLUBsA7nk1RXhlm3by1qtvZ0pAhyus1twpO3K6j
x/29OnQh916MoWmuLu9QwQJrS6Zn+TQlOF0By0Ife3H50h8dyPZKw7L2N5RDraNEY/iQYpiu1/kD
toTaRkmo76k8s/e/1fA6Q6DOgYohNyKuQzhuYLlZhnxosYRDWr1FX7/tHhylZH3GIIl9yJfWvopt
BWdRROfoqdKpuxy8AKemWkURB1PTkBzbcGpLIhJdIVelu6psZJNtDiELRG5qRVoNYQROMH4ffMP5
wYAFlIz0QDV/JXtgwBQzD63vWq5V3fPH10cAy3C5cveF8IN5i+QTqWtZBcwOuIctKHY9HGtfnndj
1hlFl8A5+NTQfxY4AqxfYmYfy5dbuiWPo9dvHu5C4j7OvMRo4Hxe2RHyXcOrs2sx44URAVK6iNw8
zLRvCo6ySOztxAH1wA/21iZtJl1M36nXltLSvkgyckIBg53nu0rxrGl4ouFuUPch3bUdwSXy1AyG
kcDI85HOqBmmXfIKnRrlNVqlqJFOqM0P5c00J4A9o/n8OVPLfgimQ9xWaGN8J7PpVbZfsdac/yyg
763E7D7SnDr9KzQT0L6f7QCESeznmiJOzG0trwU+BQeDZm0Ty8X1fImQ/iKrthCV9qA5WPIK/OQi
bO/MIP5UqVsdCIzver0eKXZ9agPeClqVlCNusfQk6I+2X6z0EcPdYyadDF5589e03BJ04ZT4uYcx
k9Uzfl4GlaCbklOAKXrQuXwKczn36L5DpIhYKl3JLw9jmvTwgm57k2ytmVFIvOZO3faG8zQUuVSH
CJl782KWS5cpSdq+gC4FFvWB5fAw3sAsATcEJKS9PVa8rzazkYWJMZ02RXt0ZnktNFJtM67B1f3j
rktlOSflRCdp37AQ+Rku4baYWoPosZyoJrodC9esMBNqHGVyifPKjVwlF9Khs4lGY9e+3ZTsWWgq
OBS1Ux2mebxXHNOd+is5iZ4fXi2rw9PNm808192sLtQBM1qz3XtD+QkiGrh3J4YMI/rD5+VC/9+s
wG2iy9Pn65tAlFXk0AIte29WEExn10QrRy5MdEcb6wvxx0jAFEcJCl7gzKRD3MBa0sYcmep8rzd3
vOtL8uWWtVED8lpv6ExT5hAwPxFHOxOWxJ9PKdL6WZuFsK7Ho9UnRYTD82uo/a9QrCgHtIH+GblY
dS9C4S6TuMeFTcR0Jl8mMX9vR1QFgydlPtuKAUDpB3NOpEFj5TLvsUaWFEoOAH/Pwp/0olM8k+KG
Tzg0XeuhRhwp7rMINuZU+vTxLMwltE/qbFI25eAVqGRTHWtQUOD0Vp7fBQ2ci2pvNPXailXSnM/Q
1+VqawipJfEsrQMKH+MjlpjGzK0k3I/+aR9TuOHk2tWBQJLVBSjL/V02H68SCq5FEGWfUxwYcUXX
Tt6ru1OlzKYppgUREvSbVg72WuepoOtFW+lx3yYw24d9XMNgQ22eej0Z7eTWN5ucwADGYjOXLPwU
9YyoUzZ78p7bsClxMwbfHP2T5V7SXyuRQ982cqfTyP/8RILWTbc6Qn6rKxjpWF/xHqCbieSSu6+M
zp29NlFFy0De8sZsSpUV8dvccx0X/nTOrTDbumOVxOz5cd7gYx/hkoSua+qw5mernkjWH0b5x8LC
RSGnv46g7qWPJPQ76GbJuzZmCAEr8Xmmk60jBWrRVaZ8g9N/OuRbznYuE8DSceqB1AbYgS2Me4Cz
dSPjTmam0yGzW3O6Pcd4iBH7RXAsKJ1VGNUA8WAC5mLOS/Ru9sO21aZWNg0s853uwyAJBagL+xJY
BMj1D3eZ2EvhJzDMOaRzBEfsFt12fZi1XnHUHHDQLvzyYbgplSik903oNFkFLgbIQkIZRYf4olHg
+apzrSKOewTLHNx7Vo7nOPkdhpyE1WrJ/9ZfRoTpJ4E9LspEVtAIdCWT98R8NnreSLku+ILTyZrr
u9yeMEGpstyGhviXd8Pt0dfXPQy5RZBVH/QM83nM4uRcPiNuOtWoicnomu4xlhZkVskwzNJUZFyR
904WrIP0LdbrHXNlH5k5a5TQ69BQRhvrlIVn2hkg7GVlVFvToXtJNbcnFCCNK/9aEiS1clAjlqWx
Uv9mUWDUV7fGYFuddVvBYd4GqVkl2eH0/QDBAA4c4TxMQrfuoqdTQicmlmtd0IFcpvDiGyjgjh59
L6LaoUI2/r5FXQGOWA6vZgS81KmS3LCc4AjlQHBoQ1jXATrlwBngDR9+dG/MDD7JzVsOX7gLxeU5
MMvW8/uosgthGXfXmh2QkDIRQ4JYOILELYu+k7WD3cfFSlFVDdNW/0YyvlHr9vRL1xDpqmUZ6SS4
rd785e7tDe9UrwhGoQgTbV9Wa4Gpi69crfNny0dmQkqmjsyg4CveE2tGJe/2GbJakEUik9METHb2
i225rEPv/PKErNNmdqwkVNib2SEQbRsrzDT0Jukl1EQ+fNFGA+GeQVagzV0mwB+bSqFvUHacy7gc
689VkrSDhhHw4u/Vc0bEHm4WvDdU1YQxP5YyBAObN9DkDUZvPqzzfvMuvTS/QcfBnmVZCZI7+iMv
rQwpOdEJPo51jI1WsexxFqfRPiPMSapZ7NZDqRyxarzFGF0cMLWMYQ3lPnsopJ+3GujV0jxhsDib
rr9V+YsF19OyAADCiyOeA0NfWgnxai9IkM+r573bLEe4sYmVD+hUTGEub97bE9Cly00XjEAnQImo
LdEO3Jkq9HU+AXf7xXQu7KhY7Iizp7Rbj6B0eyuYJSl514ApfdH0YcLw2xjJxUiIEFGyb90c/syr
yxwF7dTDlAc10XYATdQgT+9X2Hj89MH9P1DKoy07quRr86YOAq+rZOkNCNnizLkhDObHugGh+JTM
SqcGiICyHmJOF7CGGe4ByoCvleNH1KY6+GQAWmAlUHKBgvGLexyAOir8jJ3rEVp3n9n7ebtM/7NM
16at5+GlS6acyReyEOSo+v9gYFg3NK1H6eDK6bXbyQPDy7VCe8afwJYhMtu6tIOQf8tUzZYXIepp
2IfN/7uOsYgNFk5l/Tw2paXNqYhvH3LJhrgBBgSNyNwYlERFFRIjtRvTL521h8VZXrsjskeVMTKs
cJtFxlp5UIuDkorDm6mCum5u3G7xVxVWjlSyaylvZAp8FzyANmetx/GZDe+7myZG6zEJaehA6lrU
Fj0q1NqnMf8YtSp84ryVAwzU6z76bocfYhoaUG4pfN1ajlj3FYJ3SNKTkfs2x1b0Fb/lW5Ut18bo
dhDroAZWHrR3DUIhCeAxRtkeidohmDxyCn90ZIpmq4KEBo4stmSZNs9lo030SMWUFfZKlXU2tqrj
aSH0CQzv9EAdsM5cr04QWJxMwCaJubiw6InjbfllVWi4cZlZxm5lgSvbHe7dPeEFGrhBRPs1JwOY
xgI/nBc7aMCWfQQfsMnlh/XzWtdRl8eRtQjdpVk/nn8CpfuX4dwtw1ArOT+kr12vUBNcMcazzLFa
r2YLXa4ZOBPjn9pjelFhIJdFXoPckgufQv2DQ2Se4Gtuqtq6TzpSpY3NHS1cwnq9Ys+mQTkhBgeP
ohU87ea2nPcJqb3NY5C3LxjjVRk+yE1az/+EP7kSbFdf4UPF4WbFRG1Q1Qp2oFNoZxu4hbJ8TpGs
eC7mgxPLaTguXxvwLdsLoYMdK7RdWElO/wqCMAjzaRrePxmb/Kceb6FCrkwtqWIqKG3tXEhXrRhA
EoBzkwegZd7kiWqX9nANYGZjE2CZRZkJuB3aeZ5dVm6KyGKleXMr9Ht+9rjK6zgUdj6DFdWM1ZZU
Sx+l0Hs+4eOocSLa9X5TjWaQKnfwYya4dOyNANQX4lqYuNpYbYw6z8DcpIg9Aqkpcgk4xoyxeJx6
xSc731MjDkibrLm1kBkMOrQCW3ElpTrjFR7hiLqcfAg5eS9k7u8mKcu1nA2GjWcrHnicajyuWN9Z
QBTPPEdHU3nBqRAX+Z/HFu3uHVNy8E4Vyldp4qNdc9OiSXvdwDFon2G+43ZvfnW3ZLv64LfKAj2a
lB7/5CKSw9GecFC454j7A+uMqE2BzJGBePR6rSqRgciw9OPHbqeClHqEq73P9pjPBxB9MHh1vfWb
MrKmZQQg4pjhje0SjaV6jA9kH0sX7wx5ZQI8gL5z9i/aPprYEC52jND/S1SmcP8uqkAVuTzbv6wV
j1HBOVwTG/XOIUygF8l8XB+0hzvbG5GsjV0BBrjFGYcMWa2upY0mL9roEFnkj5IaAccNW9GmJkO2
FBiYAw+5/YXAEEoliA0r3s/Ze7rYehwqFvNXUlre9+rBYqJQ9DF6f72/3DQYCYn0OGu9iNWj9dwo
VCkL0W5eDNqdkFoNv2DRu/Wd19d81fymI4Mok2ZP5Mb4ZZvNdCInADGQHPCR1JdbVXh1ju87J7FF
rEY35YxmqBsm1y/vnB3Bs+lFtnKkCpzufYfQgWGQIQw3OnRHGiF9d+/C7lPfyjXa6xRAKfyTnLgj
iD80F13LRavbGDKiCwP84sQXOIH1nAYFFTC1R/FvqEIGfqMfsrBpedvfzLwav9J357oSI+tviLHz
mdy/YZ7+E8bzkEITHRzPYJPYX83zBY6o1oXyzBJURPpjJQq2/wreL8DG5r8SB98rp8oSbw94QfPG
tdUZYHh+zHMGALD/1dG9zPqd1GkCD4Aw2mGQWDg12kVyDZZE3UaBg+PiDClD4b+SApseOn7DPoLm
cdRvnCN9vCeTcFy5mO8ZuavE311mUrCqQjyPcSHw5ZZU517d6zLBQcvKIGYFNHVadIIpXaun7ySD
BQ0QMs9vzBMC7/PeLrtuv8rZdTpvwKCDr7gG6niqKfq4+txZeZQ/UyyF0ZRjKkn4IUgxeDb7XUxC
GwiJuWy3DIJfL6a1ygJzDOL897gGgGgBTOV5Gu3kkz91TIoeSrmy9LYOnu5ZA/fU4CSVx5yOX8v+
bQMtrPzIwng+IyuZ9tvO4DoMYh2iobCGNYRr1v02LXmRSMf8AOM9a3xVPjH0ULD0F13nBAJXTftG
TaoAKHU0N78ckz9nWvVvVC96kVC25Lfzo/ho0VdU8+PMTN3tlwmDtCvn64W1QPLSKL8BsLbWIJAd
gr2s8CHpbXgBeNIyujoO+aUBqJ7GCeWOBcHBX2WzsMplEuby0BrjN6RCQsyPKI2k8EVe39HpXqtf
qNen3YBTT9YkicgwdDIzwtjKeARN6T5bgZ6Ny96hg3r1Un6lt1iIdSoHLobuZMU+7UGW7flTzq3m
TJICKCKrdu8s8KkNGSSve9CGLSjjEpi/IdeZXS10puYh/rtRinTqtlstDsHhREYlSHTNSlFvI9Fl
jxO4SPgmjs2Dnohtju+ixJsIjoeZy2k+YbXNT+sr6qtHsToqPZlAQk6/908/HRFuJu2XSJ8n1tUD
5vUkVi4jjaW+qyh+p6qWD2idykn6iIB8L8a6Nw7AnIqmRE6aie2gRrNhWnBqPLkX+dspgBCpYhEC
UdSA/bG6320Yj7dvIpp4K9aSzOzAuxoGQIEg9egrUPKDqP9MtwCi2HRU1DW2dBnhlzgrBUCU7CZs
conXqEcseIh8auWwsRRe5SEmQLBBzze519EgxbdsmVB62dZZ4tcS9ss3UBulNh139qpTE7++2wOO
/eNaHfLowVfPGi2pz9V+Qa4cA+zrRpwKOBOqdav7eNxeh71LR+3XRrtp4f2ngKzNvU1BJRnE6/RO
SHnhSq11hNyzdxcGCpb+Lp8X8wHJP4dlGl1NJ1OCLDk4pdAGvUYbpUO8/6C/wtgyRsdDCw/ZQp5j
5BFIWYUkdKWYsboM73v7VoVwj4vJTc+W5B8ARG24tzLPnIKLNGEGnYDkqc3WolAOu77/9U54X7J3
YavPPNfwlYJETD7Tq7NfjA4gYWYiLUvVxE4XtwFSeLvIOpf/ECwXsgnVIFMp1hXDmzTiWbrmseIc
sydkC8a9VHtWbLIunyPX3Ild8IT/FfcdUSyQiVm2zKx+c+Fvz/gRjK0Fn8tFMTDCcXjsVAoiJutA
7iusc5qUl8Cb5bfvBciY+mT8hTnBRJh6bizRGEpfL4JoGJ2LVRzcQs3mzsFxovVmQX1w57YuHlz1
5elsALTYnEeFwq/gjKYiMT+6tV7MJOpm2YAOXvSCCdLJH69GZxd7yOQuTUmA5YmYZUhPJbH/GJR8
KBhRokIhsqNZTKdOVauzMHXEghZd6hHIX0Fyq5Z52P1SLD6ZUm8eeU2QCLiQ7uGtWSa9CjnbbCM9
9Ffdo8I5SZoKB+3uBcCGXiSBoK3FywatoSdoT6NwqU3SbpVorWiuMkTba6RNOxpbsQW3dORsNb8Z
x7+8jWhnNBpDzhEo82VEeMMR2FE5C3p1k/66jSPIKylLfgouQCiD5TRkMNiieDhvW1l5JDY2/h5y
WI1IofDHPkFuFUzXFoV2coPZus+s3MJPT06eyZgZX3hYUrrWR45EG/uewcXTMSPwDNJD+D/XsC7G
M3KASuai5NkD/iNocjbfN8hElBBVsmxwDncEsy82Xvho8DMsvOQCAFyU8zYVNJLD12fUTbf9LXI/
koGJKu5jpluAPrEcqiKMIe8Dp9CYYZ4GYhO0hhyDPJK2YBD086xUm2DdenQyVGsWM7BL0NZgp4Q8
p+U/k9/ATf3C8c6LzpIDYfe5/pNTeBJjAQMdFJVjPDhNsF04JnhjpGyBaDZhNIoASU7fh0h+aT3j
S5V+E8seJGSCMH0mhAJIU3MZz0nKTL8KH+j4IR3SJMt57C04impL5pEYerXGBsyT1+ao2UXyJwnu
DpCDtuJriuLPtciYGzHMwBgUL70qVZ2pi1iGzCyAHwrHhXEMp1zOy4RO9OAonEOXkDjhktU33QRi
QpnkgX2AUBM/uepGfdPmvaI6MTgiplpmuBDsykYGARbqSOC9+UaDuWFpbjgbZxEdkvfbNY7o8rW/
jAcOiQMgVf3Mm1dblR/iVH5E2hxQymEBBRqTXHgdKB+hmNfB42KiLI/OL/hyK1piZQy+r7DFBkRF
tQZ8QhMUmpt9Ev0FUvukh4+ZEeUdg1sgk1Aw6lbxcJvsCRAK8F61oGa1Pn++PrPY2RWb/JGz7nr4
UnvyqZ67dn/8HkuYw6Vs+ge0TzCWR1FrkLqrx2yVSWO/0acuiZpVaARxgkB/z+TWuPwlsad3ALN/
iDx/y/lN31FloG+iDm8iwame1oExuxfdOFdyiEJrDfsstAFq0YkpPmnKA1UWZI4Hq17iAXf/jrEt
ga/D+yUKnnrvVAFVxArrbNsi0NzYfn35/MSrnGg2s1AHo2/EMn/RzkiEf8tiNU6ATfo/rXCA1fzR
aHf46qvBxuyWO3y5fazRHDjNMmYmv4JAml6n86chrdw+E+lMGhVnBykKZwLVxuYeN+Xw7e5chJb7
cFJiW9Ue/8CR/NwEW+Gf2j9qZa1Tj7D61d6wzqk7Cb7di7ucECR6O4Kzau8zUYmZHlpJFJm4KCIO
VoLLs576iI9uJTp1w2DAlBA/05f6Kc1vR3/S49fVeviR/oAJm6HP5Stzu+Gv1dLnuID+R8WzgUxz
n/OHfunbkitEX2ZtWr1ABLSfpdE0Vh0UElwQZtl9fVzRzrel3fGwtv/HYgoaoovK6dDXaKUB5Z+n
i9MmL516H+dXSgMy6SWntxUq//g4ugfiJDhpskcanrAnkdqSWecmGfhS7pnNMmYNUmED5DW3KHJl
D6L/G6qQIiQBvUl6wCviYGi+0Fdvhn8qDzh9WlYIW6FOimBLyTRUcPE0Xm5KScxZYUgkF6LoX3gn
SDCk/35BhDkqMpvDVzUXrGtE0sKpsNX4dB8P7k2V8e9m7uv30XFP08n39K2tEpTxFc0oalmFhcDd
WrhVpklFEissCe2rMHn2HqTiK0DOkU5yj1slWyhPBU/M62/tRImGhOkTmk4cyyBrq9NTW3VnA1AV
qSIrYbLlNJhFKJapdIESSqxtfBWrttbgOPgnp9wY/tLhpoDY4Hoftb3T0Z77LMCF7T8P5aSzW/ja
VMGTzKc17kUqppEZO7oy62Id5bjGmqYeSvTPtqKNV2N/JEuBbPORdv2WjOde+xcn0JcTnzCLLYAC
UmhShym3a+UcO0YIWQZq4cbmI9QfP/dG8uytEaijqWRWVmmBttDFpFYdQHGD2kanBndZy956LTwa
0/f3GEBPvRqz1Ppz7msfWKmgad4K0s6NG8hqCqm98kMwnrX2DP7hyKhDC+P3Wm+0no1s2RcKLp3Z
mnuuM4i3kXR4W/ecI2tTDcBwHVEnJczXsHRmU2/F9XcxDvXFMb5rBZgBf1y6+f6wrtzysnPVhDg9
b66NuXAwXQdXJGli/zIgFaeW4L4jXb86nu5jVDmyEluwLpt9OHaD/GxdhhHqMO+AaCKxuLo0KXSG
xTyyB6G1sR8bLiyJXD7iSnJbr5hxHhqXSj15KL1XRIcBKj9Ho0ZSy0ufq7pyt1ZiA+ALEvJ92aK4
6E7DOKzjstX02kmRphksODEJVxOtLGhsU26B7tZYtylVD6g6tG+fee9GGZC41OkjQ8gfCpERKckn
alVxaBbbz9vGQhOqAHw7axl4kDT4eREG/1W4fFwgFdVe/FIRxwOn0mQA8Pbzq2/43HCThcqN1TQR
fZlGA6YrLfoMTm//lMfJRwdTxxIE0ChDzUQKWFyFMqF1h5rzWSLF21c8d7iLox87hZTgjA/Lm+Dx
sF6ODFcuxFtQ1qUQd+wSh64CsV82T6n8oVh1wOS07LjRGpuG6YIhiMcI1EiUSWq8h3QhAsQPwrQZ
R7J/IhC/96wGGMoKUiHeqyuPH1CWlw/Bs+sI2Xgb8s0qBZ5MTN3a9VTMBUhLi3paZvT51f9NpFAB
pr6xmLgDKyFs4PuSUduuhr0VkXeCwVKBy7sUFhJoVP+iTl+eqzYD6pYvmlOSKqKLWUjqeOsgRwNw
q5xZSC4WvBfhH6n8szrEmI9kD1xwt+1od/tg16v4stE3r0dqIA1asGNnyWl5bTQTtb0KkkNc1lMN
EASncoi807N5d5o2QQkK9f/Wb//ybd+7Kpp+jEYGsaRDdsfCVh+85sIGjQwRNfM8p4VbcTscFPAh
AhZUi3/mgZRfIPvDxcbQ2FZ8LcttVTcZacodlrNlNEXPc+FKVbxtmu5zosJxTiqpFJ3xrTsowZZS
OUfugIphR4CrQLeg5bVaTHjkjj03uDPxrNRiDdCfs7kzWNZj9WdFPCyxJNa2qbbGqEAjI/LN6XMB
mMSSGvsgZl/NwIyJkBtr2mjBDFeka9Li6UHDhOdL/iUHk4nWcrZ1OuYsBEGpuldu5AvtRUmcO5UK
nXVnrc9txMAdSp1EplETdFb+fnVSrTXt/qdV08qhbudYf8+0XWWhuq6QqQPnMHFFzphovQJ2+G5x
l4Erk7T2VnEEvebHklOz02OMDYW7UVJ5JXMlyWAeZX68ccQlccI+CMnaIHDCcrbuCUM9aVLTQIam
dGxt3l3gvWYSrZDBYgvwb5JhxwzJAJdmz0DWwE9PY3Gctwrb4IqrmNYhlrCN/RA23Cx17viD6dzm
0AXr+VRAPXLr0zyTRQP0kZKYc85G3WptUHI0tAtFxws+efyBbXqInh7x7l2+uvnbYjOhIj4vFXDx
YjevNXUvZulgjxD9UJfa+IoylLdyFtGtBiPW3ApPa0eDhMF35B2ga0yLCVMp/NhS6V8Cy5wh+9Vr
TLZUO1IOr8xlKMhm/+xmbJJZJTQ/b5C6s+rFGSMBsoy78CC+qPD3/2pL0Kfd/hxNHXJbhehdQsiz
1YsDVyA2j8fSh8jGSURmqP0Sq2MXVF876bxF2VID4UmXyqh9w8TKTHzucodItJ2o6swDc/plIE6W
Ns5y7tvPJa97fVVqttl2ImMnMe7HB0WJ5ZkDQ77HKTOE62sevAjJfDqWyVnW10w/jPnRf+1UqOI+
UbyKY/w/R/kc+lw6iCaVN03jEHHkjUemxT+eEwL7qVEjrzrRidsXW/D3F1XzLKg5Emf3gke8mO8v
MlQ3Wq1wFkANqe4KVTZuV0sT6EM6a+1SW1Sqc5ODwM6H3hTz+7GF4b6D05g/n9xlqnZ2Xosd6Cvi
VPC9rigvW2Ft47deN108bzZkwT3S1yr72QSDGdjIR11aFZXjHStzYH/BLP3sUWgEIsLQTNBfVGw0
F1F19L3BtFatBp81/X3zpjqgGC+UX7Z4Hor97lqFr+nJiyI6kIArK9eI1nXQEMfQgQ5TQIDlrI/O
q5KgYn9n4DCCI8Kz93UowvuLoFBFZKuJYgEMOfK5X+ynsadpGtMkMaV9vhPwcY769MLEkVK8e6yO
HsY1hgvPs1DFIoCnSOK0eqRwE8uI52h+tzYWeTdqztzYn3JOAPe/180kQrfnO9vIXtCKewJMuE8n
t2cp5UvuzKK+UGiCNJSKxMhD4u0DFY4lM7WQ+nmOn1Em2WVutboXy0DW3FenORqzEFZCgL+hyvTO
wfB8Q/KpxiFghNqS7yX8raKjSYgffpW1jB+4bPougz7PkzZx2f3pfMhT4x8cSG2gAt6ohUtV0/kG
i/meQmxDmwGt0i123v2EOUHbZNgdWcpV8ZkUPedyDZobQLVk7LsEU97hDTkpoJrI2yrcNr9/Loev
AN+pwvLs5dkxh+tKLM7P+gtwWZ3FvEvT3DVEDXWasTfeK0F0LKL0bx1mgi0UnU4FDf3bUQUEqVhU
WJPs2raKHZh4cQG51jq2GJKfqCDueMWgZhwEUshSFAv+J7FFIxZaa5FPRlON95B0lo9ATexH0eh4
SeCzNS2i4U9Y4L0CMEyVml7+c+mc6CSNHg8tB5eULptgtKl+qWXzoYAYYUpLRrKJUB9P7b7GYLrl
ihX8CsmDYiywrQ8SWm6ikQxt5w/EFG+O4MrA0HOmY6b7QQmvpzfP2QObEk0Kyqu1fy8Ysg29ciBu
4EnT0bUOCh5d85+Z+6GoQE1f3namlRJ8zbMLVsgd2PxvC8B9ftCJNl+up18U6lHyF/aMRy8qlAyd
AyBf6t5YjZmrSxuadEoGujjnqDO56mYPDEEMI0Rb/sbzuSNA8Mtx8tvtWroi/G/a1y1FZcn2/Mog
mRt+O+Y+VRCt6TmvnNyDB6A5AKGvYDH4VE2DfMjxXL6f+uVQAiBAgL39KF8rLCouu/wyZv7KC62D
TBWH+1zUk/O436atZyTbG8IgrSzxtdu23OXZhXYJYM/wLW97i3ned4fVkgruhgjVbprrcjQVY+Kt
uEmvxXnMqGXpqb15zvJtDfL6Kq5MeAkXcr8NIfkR6unTAVVqcTfqSQjKpTae4gSj1nBvKHLH2gmF
LapNF3mzF/a+wCHrG+FGdGfu6eTDnsUMn8Lbeyw2IAXquUSTZZeh36AxbzFb9Dau6szSJMGxiUOb
EV9+/++XoWlaARyGPx5LmkjPWouqhReJtjexmxoj0e/M3i0B9pndbqeXZ77yBWCoLENeq2pK75ws
wv4TjqbpXeBhbXEiZo41qTIhFcxxwQQU8XFcLJvpHsD9VmVVrFho2likep/UFKVRtTFwIpEsTLND
3BYw4mN7HatmP+4YVxNcpnI3RyzhE71ZRmIBGE+C3dNvfVPr5m+87ETlLbCVsMzHVW0FfbDFHZI4
LAkKk4c2Fy0KEks/8IvBkD9q2VYmiNbPoP00MiRqviuJTpcBl9St9E1jzBgXVvNwkupKQb/OavCf
lPk72tKTOrteI1fS5FckG57Ksinqol21e5ZrdaL3iiTy3EzpgsjrytlaiE2Z5BIuE2Wng46BXhlb
knFnuDwPLjvYrekR2jjTF7rH4pgVosJXiV8+RT4Z0Sz9fX/xpnKQHf/vLisIE8wo+NIFdPwOGYPQ
W7GIXmmJoFBm8sQSLWSneh//WuLPFZh5bDEOLjKprj4mxhdCX0q8PVYyC6mQjNkqvx8DM5xscAZc
f1guo8U5WGsUUK3NlimRqIKtZ9GzqexsCpMX2Zk/4kFMy3EATHoM6sERXEnCppFlqc2AC221aIRI
7QXB98g66oRt+mRQE0lAl95VIJ3xZK1oDQWdmZdn9n4CMVR+TsGT2ZsKwGD23nj4BqctLXaqVV8L
YnoHTecNDBVU1liVx/0zGc02RldL/vwh6BVtShPjWcz5wbe2/H4deJekIQLkvg2leWwuh5DhDaT9
rA0dCk7RtLhB5s+XHkekPZIsol2du3Ux4f9hxKB20YEpjmmNi9givEzkCkDnVdyOpbn9TrlObb6R
+2JoAq9GFB41WPIw3ZxDKR1QoTx98Z6RfvarHEDZ9tRkfPjvWlA62bdeay+mvVRIhcBljF8jZ3pU
o0glhQ4oZliRU6wiD3rJdrKp99qANnpgEJg+rhK80TV7SLz8e4aSRvSG4rM96OrJA96SFz/pXJTD
ZYPdRMvrkI9y7ACiMogmwY8uujsA6RFzgFRf9UE5iKCywOGJERhggfSTzs2+8c+Qfr1BCSv88LTA
TXv5LOBkw9pSmfu0NVhjhBiaBdtuIRnAYRELhR/V7njdxIFvMI8s54dzZvgYKkKZeGQxA02LtRWR
IH5UcbNADGdFGEPfjq9DB+q8gPkpOsttDbRFrNUrXwxcsZF1mDVkt8LDeTM6O1l5A/53e50Cvfxh
08P7gkQCR1gdMcdetkRCIM5GmFevrwdcFf+oUIg79kC/YX1y2B8xwm/O38dxVJVVYdWHhCMhIMDD
pkxv33aS9cfJUwY3lZfKF8T4HHuH5MrUNJSyfnQOZKzVNd77wWBy7gITOiYExOErzIDtKTMGTsMn
hksSmoArPxd3v7Z7XGLiX1MOLWx2+M6sOVLTA/hfqAMO7t3GibbOPOyPgJrMIUij2ARoIWYhiJ2i
ptMiu0su56zdpYgmdXhztJDf+mRNVK+/DO3XZeO+NgBiFQ8CtTdgzJe/afzsRvPgpNdtwCbEU9Hq
0m4JRDk6cCsomg18q8AqKmWp3Nx9hTzDXHwkSUtxBz+wWLEXnQjfa7/oaE56a3Cw+EyrokCKLmDE
NbF+wDXm+sf6UBWfIfZ3fzuuEhZ4083iNp2pE1AJQuPAu2XvUcU1dlmyscnv3H9yP65KaiHSUD9N
pCDe2bXE5UhRIC8q+x82nbvoNlLchC1YvRVhmWsDveNLwAZOIBjf4cSkuSzqM84h84VIAArH9OmU
r83aRUtoVujgKvVubW2ozlKnypzuUG0Gg9BnD3F7Y72cqgypvla3rMz0zt4kvYprqaDyqru3bwTg
M1i4Cs+gny01piXynZF0k9G1IoQp2oKROqpEfzo+kz4iI2XuuS5byoEEzLAA7fMx4E9Aw2Jnoh0f
hg2hkQORhugubT3wEbD5ZzGj7UmXZ7qSTeFX6fydEdLnd6u5KOJJW918eXDyq83Gt6Lxi8SQokNg
gUCIsoYHcZ0wPa+mqHeIqkxSo1kbvjJu9Zx7e3g7v4HhEVuAtSlJYoYhby3sdgHqlvmZHms5xGea
3oiSFybD7a+pvzIufnwFwxiAb231GtBE5AFPZph1c3L+V5EuDUXHjFwgsZy2HdoB5MzOqiEAb9KQ
VpRo23haRBpv1gbC/VPDSZEYHllifXl9sePer7u47w734i7qqoGjfhPAmfHatXLxvV3fGpmYrz0b
XgXL/jlqMN8+se9QRU2Yrqy27VtUwGIfnJjCnPBpjACBLcemr/pj38FRON4oed4iPangnbbGpWNf
7GIyXC+S+WSkv/A2u833URQPodOlBGHLQK81U6LSc11tQwQY+esURFHyzDNYgu+h8u1lTgBYq/uQ
O4XalOVbrgeTloHz98t7NB7T3hlL1Qevk+2uvdC6oiulA6EatKiKxz4hExxO09LqOwRF/YCNpUoV
Qb/G9pc8jfgN9/dPf3zIGr1awktUhDFk7s99nvFsAx8BefFp23kaDLV0abbbsWRT3ADFIJfSEGrt
ShNVW5xxUJlYvki/8TKHC3rhUTnqNEjd3R6qy+l4FYfECHj/pL61/PkF4FkygMcNVwCs5QAXMuVk
71LzOCo1kKjAub9cClf2zKJFbEBJWf7AWFcDT2jjyyS/Fjg9Ud2tvG4OCCcqcerZY7lX0E4SQ/CK
LkNK+HJxEepldkRjQwBpoEAm9INmw3VC+xK/MVtvk2i9xpuCoo53PP8kJ+Qu+1GoSJP+tFl+Rigs
lgqAhkciqGsWEWHSXHaN9Rto+OHSZe7MXfG6D5MaKG4lBusZoFALqGGKFdp/NKodTzRxa143MDLf
fu5FEOWt5DCczZ1eWoDhhnjODknrpmgtDtru7GMm76tK8jK4LRjyM1SIu+GjUt9pXrin7ZXUe9nd
mPstJnW3uIaSzMDM5Be20XF9mu4g0yJTbdn248D6xz8xuEMKxsBraty0s89gA2Hi9hAphuNQEVE3
ZyQeSsHra5F7ZgKTsQLGO+pJo76lXgX1KfqFbG/LNFHZZs2DEMbMgZCEL70nzL/bwtuRdbAF1Q+h
aV/DbFQ6y6YW2omfnu6yhY9xPnlmqRdRE8Q+bBJtokA6rMM3Ne7RKzrEByWiLLAb2rf4BinxnK4G
jafRe6/Ty9ddgIh9Iw6u+9hXTUmwgzeN4Hr3CRM+t5cFFdxvIbZKan3knw+yVCy/YEYHyQnv3kY3
uimmxQyuCPNSuBWI4TPBavvwgIUBkY/yPw11Y+3l8m8gzmNsHjAlapwYGoHDu/Qxr3DhGlpd4AN2
DNwPcv/9pPesIgZDrVIMCt7VAJqNFLppBU19gObf1kFLBIdhsdavqAj1T2AOyQ6eb6fqs2/3Zg/c
CV7qP8iNu54CK3fqKP9rFp6X83uau2ezNosg6hyQNJwxSjB61Bb8plIPr98HoCHMhWJKw4GoJW7f
XeFJ0765LyfG2E+YLlOLMKJ01tnKCuCf+aoO11YQR15WJN2yd52bDFnNUf45W0jLzdY6CmhTMnE5
QWiUOqA2rN0uA6O7JnONb5/we2DgnHlVyy+A6jFuaaCD9h+dsh66TWwnmzwwb9P+YPaXgLmul/+6
iqYfGv1DEKIikdt7SNNOg3PFLYxpCQhtdwfIT2dZ+zT1l8bClylno5RZtgb+QPSu2ibkSKpe+DkY
fSrshXe6AO7DWBrfxgItr7B3wG0Qjo00bVgruFd7ij9wc4NpfPjHsyoNSDLq1hwDlN1JKHoIHSJ1
bw0pd2Gex2LPXkGdHN/CqqRKmL1vlHXTeqGNO4W7jvkCWg+zIdGTlLJFOAxiUTMFsl+CfbL+6iOI
bB43CCpNgjpraIyoLPyvzeDiz9DiKyb0APYic2AagHYqsHNhEtb4HsHefEU/9TdDUwUx+F6RiZKr
52JqHORATWTGuklrXGz0+UBJO8zG+cgeTcTLo5D+WUEgUJfbve6n+PJtT0ROeVZL2mdNEwBZHYRn
+prW+DGpvL+rjHdb6x5wlDTOdyWRBESqp4sNqk+x1mcg3tLrQcFjn3sv+lMcAhnb/PCXzOWbTAOl
2fY4s6Wsrqi/CU5UFeH9c06eexcLdwzI5Zrrbc4yT9ysIJhUE/U25xpqn43FVkhbaXSXgRWy8Zal
FbLAI/HxbuxbdhFZ42pikfUlOna7MqN5uCYRtn7YEEal5Ow/s06AVs9g5dEhZwxhwRsq1FkdIoqr
icNJBgE/Y7ZJcsDN5PrFFfLvP5mqvllyLdczerF3LUfhQoHEJqqPqqjHsUxhn94Y5qEAfhq3SuIG
4RsUysWVpu7V52oFcM0qmLFLBJP5if7y614B4FRhDx2Yc2ZI9csStYXgqIj6j6HpLzD55AWiOuhJ
XsO60kUaIwk5wtGZfhVj1T/y9omesP/y3m7xhDPIDw3lXcljXQha63xZTKf+rw15inK7I8DkoK3v
hHY/VmFxdAoOjnO7+QMvdst/8WY9rrPdhfGrTWlkxhSVDXarlOehjiOGV9rHt5kZck3AfbyRKzWI
3fEXPF2fepzyQLiXa5Bt2oC5bJpo6i9tW5yMw1qKFOuR2FQeJVB47qlxhhkCxaw6fTcbX64yVmf1
1WUdYM7T0/orrp5qOctxEQ1SV5qf6yjDM3imp0kitem7/DvhTZrT6GTwqIshlg60CtD0appg9+qz
cEgl78HUa7vgYKzEq62gj8gwP0hDgWCtSYAiFfjmbv5cDwushvyLr2gJI9XUMCxKFgMofnULymhu
PzmyMxoh3H5MR8j/2Dq8SAOZFVKw/n4eMShzGXxvztYJ/cJGldYKyO742YKcAU5/mWHUS0NcDgMH
h+I/COPzy79uFO+KmHQfqvYGLWmlhbk4B5RDaWCPO80CgPwYC+6J4ba02Kij/6qkhVtANmphIlCb
wnt1Ifsv8/ifs18Xy/9cmNdJsV4LxkPjzdc/a1cz4gmABA+QjY1ZKkxXSxb39FrvWI+d9PUobaGD
g++n6Eq2Dci6UyjlEAgb0zN5STaSvqOQzGanDtdkfxVWiKoj5KQHhxC9bgbHlXj1lRx+kC5y9qlq
V812KHTxHPQC8rzwShS3P3qWYCB+hZE5U6dhs4OvHWrw755zXQoO9w5cdfNF45pob0XcJT6CaUh+
WZbPm0iWeWRx0wHnffzYmCyViWKDc5yhVTWmBMIN5yOYV1UtDXhx66xufY4h9/VuOSBHQDl2eRfc
vHrFL0qTq/vd9vqtkeau/QDjeV/rdpe8ocEMGl/q+GIrAoRqiKWm4ZGZ7kx2Zn1bNtJoNMPEV+Z7
Xg9I07aJDe+M+CqltXsAgPefmT8Jy9pJzuu3V46LUJDDpZsC20fKkljmzOEchzwQ4nnhTnCpCKug
wB3m2IPOCDrCupe5YwNOemYRouePmJWVfb2ezZtwry3EWZj0XKmBHXDClYCjR7kUQU/nQa2lqqDH
rGjBT3457EGu/+ZqLdIPoJlaKd0wqJj+vngZz1YsgoemZNccocU0I+QI8WqTyKrIeNArts2WDf2c
HvZkUmk8TOlSBADw1+dHAK9jXqmVoMrBowENXzhApNBTUpKe+8iI880rDIGE7s4YmdETgU9WGTyx
A7YsSNStA0YPSOx4kvegubjSEDtp1oqRvoLimwmzqWWWIoTbd3nlA1oeBu9ptDeXdis2rtWXM1uO
oTAa6JKgUYxIIKtfeuV928KpIhfLADqgGerXPUKMag70EDfGxFcuqRbl///NMV/5Phb9v9CbUbz5
TuKYLppGD2NPJkY3ZNPtkv3WJtq0ZxQU/DZ4HYR/6clQY9t9PmriyohCE4XKLm/wvcyfSKbVHvrN
aKw6McaQK5y0LVntUiPQRp+LqZWvHJkJWZNP0q69fFC6jUnLauoB6xWlBvcyLdN84ivfwTLCFvPp
zkUYARCi8/j/Qp0eilZXPsmXIvrBLrLtOtzy2VEcO/gSmE07e5OkPyo/HxtkCenQwf17XRtlq7aM
j86N3eDBwOiDJywt3MeRoW6QKBYAYPIGGG4KJJH4kOzxB+akf/1cMXHm+Fd/rUXZQhynvyN9+42n
6Jsx+CJg4qS9hHoUNws770t4BO6NFyeHYZp129oUjlovZuoqRM+ScGdRPtNiKiKAs2Dj2O11teoc
h5TQKToluplWBbobGjh0f6hLMt7DkIvTvOhcSJ7zDWUpru6dWncSfrNzuycTyn4vJQMQiVHw8kJn
EPDQ6EPTNqmW+7+haTXCmkcE1TkpPBBDwBwor/XtHtNZoNDoOOqQ4jHUR1xgqAyXCx5wOqthQHru
R4HxdnVN06xllc6tWGrcOIbY3CVcQTYbVYwclZa8MNoNu5yhSlETNsdqB1At3VYcfuCfJ7GvfmQd
vou0rr+mFST2qkV8zrw9J70WAl/qdjowUYOQZrNGR/8GeRmTX+iJZhw07K8Eb13MlEivHxCUO3+M
6UcE8yvkvczbTco5et3Gj5npV9B9ergmv8jwuHkg34fyeKMnpudhluZ9Fn/6SusF+wrg1iwzS82T
HGWCBQYr5zGF0cHPQqSq+ob7UAfVcBoYFxAPApbw1CKkVH4rFO9TIKOkLpNjpkxBODCkit6Nu1Rr
0M0zOhT6ti7mvzYj1iM9OsVFuABnydtUioQFs2T1STkAmiQk4/pVM5wS9LdQFJQXaYVnScjgmYZK
OUglAsrhGU1ks1uwNRkHre0qKt203vQGwaIiweaFFNHWLovUninxSslLyjD44zvnqbA50Esx9Ik+
WN0HxnUlpRpcdhyL7z/wP6F7rKGbepq92olnLRiqDUtEp51fUyIwcw9Rj7K8rNgZfChsc9htckG8
6tB5Ecykl/RMa/RJds4lqhoI81mEYFVSJsjvW8hT6ZJcUjcLh3xHUExADkle6LrgE4yFduQv7nx9
wb0YnQPrASziffTN2HnLdijsShhfg9LCFhV/u+ChHEH/nqal7pXpwQMaDGk/G5BzYAdH9xuYhwn+
sepihDZzZ6Sc9sR4/QtwerG9FWiF4+xyBUFper5V8Ns5XV3lWUb9TzUQLPw0Eh1dsV95fbUYoebC
E0fS99VJSFuA2pyXxnjn5JQrRDtxb16R5yeJKcdffA4U5lM9EASvrO6kvsg11E2L/ZLyijUe8rPm
9AkHl5MtGB1A81ZWjGjzE8pc42JKWz8IxxISfaYAF5VCxOD+rW14wsIJv/Ib3XF3iDuOM8RHZtI1
k6kmMGjaAaPswlBSU/Fqs6Prd9A4f8WDYx0cHgZjX4yfJeFxvtSag++sm9r9ZhV4bOks0wdgxma9
SMIGoUyoQSJnI914zNwuajn3e5k104e1OKsZ/oOk2SX0a/3gREB4dAZgGSsNWMZkLScWDYU/tsYu
mgTiT+Ll4J/TseMxi4vrPUst/pK8axRYab8OdSY2SZzFEW9EI3EL0WIEvLR+vqG1KD80UJKlRL0E
s5LK9kGa3Qyqd8+S3Jljte26d0wzVmIb82akF2BYAle0qNmfMMdzstEzI4mMS3GfYVojCVim3ncl
0zWBuMTnPajXTVxpRmAUhYI/SZSQ4wQ8vpYT/23x3yUMlGPtWRpWOEmy0nxg0S5uMnLnK5HFRW4D
cw+ibyrDesLhSxxrlgcKrlH6UP31+muTbrWMMpxNgBrovTdR+5R8o85eRrgs+GklMlQYVh7wrytf
HCwanMHmlg3H4GRRpZcmZMVgRqxG+VdqTkmGTk282OsSEKssoI0EaUdd8UuEEq95aqwHUq68xk5R
kLsg/TPv5m80E+9ubn+u55HetbCVaKNvmB/+ooPWsp9XlvqweS0AvGlRCLRX/Q3Jwi6t0opnfoKC
kPsn1e3OSpZIHuidkMp4fH6D7swpRusWxZPLrNWxx6w7HXVVAtSuaWCzF8QPUxDOYce3PwfuCeBR
WGwOdrHrgNgYmW+pvSsrM12EwqUNu2vua2OMI+ZSwHVi/oUJGwMJb98j22sF3u7xEZPxUKw9vr9U
vu6SWpmYCv8UI/uvXIezDhq3EKVu63Adur3HeJLXT1mKf1qAX5g38bPj8D4hBpARgNdgeGhwMybp
qMrqMeJ13NWOEGTzOtoAytBJowKhMvv1soehDHqivtkkcbvBnvKwOupUw1wi/3XrbO8bJDi+/dMU
MIy6toDwtoNf1oX1x24eYAxBxAO/75cmpwnmaOG01GCk/5+AWGPqapp9IGM737SMg6zRVkMktWWy
OSRWfKfowgYzYr2IF4++V/8VQ1bpHrlIRZkUEmiRLNtA0cWVYpCx7GJF7bhb4njT3ZAUp6ZVKLHI
BOW3bWNVeVYnCiNs9+0iKo2aZ36UWwou3K9AxJ/vJ6HIT1KabMjnSx01P4+rNxDHIhbmmZPtjhat
bnlV0vz/nudIMzRhcFJVX1UrEF3YgV6qs0lEuIyNOwi4kLuCxc21ZH0vZBkqhDnlhB5Lq7P2PYk6
Ls86cR/JPrYZFiAYK5maytnpr/098QwkO1OCdQ+HODlOHpw6CQPoe2bS9lj56lB7wQuDtJqYGVgH
rVY42ZKNY37tHPhaM0q9PG+QhhrFZye4KjwiVWzP9kY8wendj5GK1jzSXESbE/eO0mmqL3twx3rm
PiR0MFh/+aACVebjCZLfEM46aJB7JplIuSeIIInqF3uGPClWjMGKLkpHAnfESxLcCQec1sANejXW
1IvIpnTYwlfOzGQBjvEDWY+8by173jNsRFVbVxog5aVgtKpucXuI4yuJ0jTSVL6dZepPMOVsgZZf
Yd6l/VL0Ee6T5DSfyk4wDmX4BJO179Psg/Oa+xTeXaMrcS7f28oJ2z/Fqp8UdmufKkCPGtWgoK9T
1sbg7UW8m+WfkPZmg5uo7DZEnRvABQTB0hsMpcsvOOOO6SbkAHdcplmtTXijnPpf2ZJlNkzShABK
cZH720v7//ALt818uyJOG74EWnXLVxlvgC4tSBZE0v6lRyn94xjdX9Lh3wPJpjh2wiQ4LcDGJZml
zfW9BKUDoWYXyOWtRdM/2SVbG9noKl9oTU5EeLvOomJsdcAiG4rAlbg+sQL6w3GK34sk5o5ubeGK
YAWF9qINkFzLMKWfyvmni5mEX/3NTSgd7YakmMKjhOkbnnLhrDhErQaiSa9mAGHp0jh4Or8pUOmv
92kB4oko62PVxBGTT9E8RiC9SghxdYCv7PV9dK9luV8oMnhpiuDknsvixiI6XWwUjQesjKW2DinH
VJOTba6DuFcl0jzIkl5rFHHMBUThpKIxNzoAa+ItTizlZRuoxyb9SaZ3t3CH59xWmb+1y4P9i2XL
i9ltuQHhwTdX+VbC/yC6Cu0ta+MsTLsaW0TFq4A8tPaI+JugDEpcGt8EpnWuuV3kOdVHl03EbOTk
Y1Ae14NEKl50UNVKaKzWJGQVw64T5mmq35yRYSlrylg4z65GK8GTpyLFE7JdaRYYWVtR9kFLcee4
NvI0mxzatQfVgWGfH41XuoWf6lINkHeIqmptqEi2qwS4Uy84yQzjhuYqseaXVqz1ORr2V3sMXdZe
Xd+tFVb6m3NN6w8ql9xxPi25aDiHlbcKWS4FgLDwkXYU2FHu/+ufTkd3SNSDVspz2Kgb7i7b8EgB
APgMuUDnqR4/XK92bAJtOc4+LigX1+P3E6J+W6pkpDMn1hgv0Ag2/+HFpRZFxLN1Nz+7/QMeZl4y
4na8TSFYf/XjCp5bLci4r3TvD7ka+e2ngh2AOOTBxfo7wko/WF3zl8qpZCInR425O7Dlxyc8X7z2
sgscRv3TT3w2qBFO9CLMznMA9ru1jzO3dXmjIcX9wTAt21ZasZfDtbEQTtZjCAaom/eGJhtn/QVE
xiApxNMlgyOBhIhfpFKNJoN/6k65xTw3pP71Ka9Lel9YryiSSkpN9wk9wb0TpeD2JkM33fXoPhlh
wismUUSGSxIGe0wcTMCcg2B5gyqAz2GDN64KaLEGUTz5RggJe6pSvW5erRUWlpnNXvaVBiWODhQX
twhdBFFyFLwrDi0AZpbE56tgUqLxPAAIEQk4OP1anRHQDaQ/S2VKX22mZ4T2bxkY97NPMnqBjp7t
JJIKPrLAROKptXEikpRkALZ47cmUhTLdTrd5YVhjv/kN1eEgR8UUeiseEQnkZHL6KsEdT/iKaoWZ
Ry62Pngl0httguQvqSoygzDfTJwHr9f0lE+8dz/yMiLlxJqb267s8JnlkxCETu2zxxG+0O26lhbe
agVvfdJ1EJNK4JN7tlcE4/kMyHwur91913p5GLeTHc2m5JhVMN+AGuZNvpN9mp/pywawQWl8u8ma
tdwuNwYW4K+orDtA3R2VuyaHHEJO4KvHQHFZDZ3+k6FOyK/GEuWu77nC5+m38BENkVlcH6jQNOWB
s2jaKEaW2FocW7mQQ/ugMBCXEEV0wCBjDZw5aGCHH14LBQAzxvzfn7HKPljqnm9d7D2M4C2+0F/7
TZ4bovNseTojAH353iaq4tKSy3o5gIEJ+kZN/S+b8j3u2zRfC/DPQs6oL1RLs3q/V2c1YU9kiGaJ
GfR/Mev5a0I04AY6kWTXHY2r1AALfIHFefPg+VkK5MYEXwWzpPY//qUuI00lem7hSvR2w399EqKm
bCj9eaAswL+D6PuQYLYt3hEO/68gc/0cZ3bht7KRabw/ySr4gmEH//l4v9e0FlpSXYd3tXeNqRmZ
SIs5B80YSMh8ixXd98lk1Dyn83gL4+XUmdkV8+EyvC1aNsFcEttYX/F6rhIzHYMjnm+33nUhQf0x
/q/OVEbVIADFWz94iQbBy4BPDoVKWXq+VN2VJTfO1fhbw0LVtDa0Oz7j764fk8IBgZURFtaGYyc9
e6//kAJL+xdU/29zllg9u7XHXnen9lMRNjw6aR4nfcgjQAY8z9p2cEbHy9P9Abdyb/WyxzOKxoqq
/7Og4t7ejAdduW5xu4Hj5EDJXz4U/UpXivOncXj3c7MNs4up9+bYdhlKXJuOY2HNzxBQw8YJK2xo
kb9lY8fGVVgZqqz57oqHYljMCO4bAQD2a03trrMliqzg3z7E0CeZMoC7ACwi4To7GVvE+aJ9GmyM
luGvFH/bxIHgAyncqGtWD6vKopUdokTGsKzbNM8VYAlopiCE9W9EcYhzBJdooEDxcIPX+ysRCVCO
KSK7DrZ1mYoVf+lYIQQCwilGeiuFm6SPSGeYjnZY5Nw8Wdu/CuFlmsGaVTsfG6KT3bg0U4DEXDxD
Cg/eM9BXSrcAyWk1g/ajNqxNh5wEGVeUr8zC8ha7PC7A47v4AwzJ74ok/smVI6ExYRz4QW8npeyK
0fJsX9SKxLCgTJahtk3gY21Wr1HlxBslXFtFL19cByQiwkrJ7Aqz8nDNbwiK7wh5Hblsvf+hK26X
u+aq8ExIbyMCmhjZG9M7/3Tpc61JPtxF/ZvkeDBak1icBAAPYE8dbrUQVbUmlxTGMDCD0qc4SPKn
UqruCs+x3S4SKBv6L3napEYMDvN5RvHZag+lq6GeDfq04kDuQHPyl7zEQEoOh57uFvU+XPDLgEDG
tw1zaMJBK0EcAJ/sTOgW+WEQsG6Mkmu0uhFaGRtjMkVUW9hx2QndRA3n2ogXsOudsZmu1nHViPVv
2f/KFa9KEq79m5ifTOt9ag0KuQafbrrv4oXszS7G0L80bCMsJq1UXj+9tl4PML/a4+J5GDxyicV2
wwKFMkg/IYHPDTdkTwAxw77Kh3sVqOCbqC0PzT86kdOV+nPNEWuKJvhU2dcAlWXg6eWRft2uJ7MH
ig68jlwX61eSB2ioWyEhGH6v/dFYmMGhH87WmLFYNdJFbWoJ96vh+biaSgWmIC96AW6eRwlCPxxc
Fg39aVPdRoENVuiYVCdJEolE3QVbPK1N9fhvAj8n2bGT2osDGeTUi/Ghj8Mkis8wdmOwOmIPGG25
Kqx6Rt9GhrmGpCMcCp/uKFVWnSzADkoBFKuVkVmaoncIL4jjVIY/6/ou/CZhRn5U/097zy33+oCD
U+GIkkPRLvExl2bg0nxno/DRtctYX1RktWZGYv/L+XXor9smmNvp38kRfp1+77T9+6gRRYCMJqD2
dk/LAI2R+0sWUw9ihvd8lNdAevAJ2kKe3+lU3udlqpJuHgVDI9IK6KnnyFLHdzJTf6qf9IjdHYmO
5gwvI9IjztkO2TMoHvbFE01OjPv4vnNPMJNuwXCf2HYAiUypdwbCML8qEN1xOz3+2QdEStbc/8RI
bK16Yr+AqOiaIazQOWIO0yzLMmIZKkFkfB4m0LHQpJnpKetZfHU8GC+bD7j+zPepBQI7CYCWULio
4aGT5YkyWFVZal+dkcCmgwvmgpf7t+HCC/9LneZUJ+6ixEkALmN+qs2kNMbBatSihDL3inSLN0KI
xH5IZDVvpJKdOthtV+J5jzrNwTMrs3tHjfRKE34e3nN8/CST9KGc+GeG0oPHdyvsvVp98AQ4efp/
bQyzpZj00Nk1JEe5zXzLQA5qRUSxKUhMY1Usy+ZLYZRfTsXNmM6QTg4oUo9xzG4ro5LDHh1u+xep
+KEYswqhsGxQhqO69buU2ktJOioLxgtq6FpgmJ1hu+JkS/8oSw9GrEUoDPRHI3l4VOOjAcvk0x+1
bywvBthmn8/QebQDf1oat/LYzg7PfLWRPyRj85Nwpo5W0eiuGQNLHPHJgUkLQKfeMeuZ+Il+kvxK
jvwL9J94fLJeXKP0i3VqpSP56GRG1Ip+0baQSonwNxAhzHh4mSbXY8UhEv+sqWb0BSezqrNYUyaC
BnRIJq5VByO4YCd52PyzlMX85ZzSslN7683tn4ZL8wmkq13B8c8v+VetYz0YIc1Lg3BrGdgcrseP
VtY9mkY3wq+/p2tZN0xfoxHUzrFGtLbvW/8d1SlToW3+iURuYeAze7nLHGf7qVfNqKMGvHDg01/L
w/XWlRmtEWXQrHUjsmypdY05JQjrT+3KF9ljERHLairjjDydWiFq8yRRLyfcvHmnrazZytGL4Ywb
E81jmXMYN34Ofxz1snnoCLOpzdJYL8Rd4GVNZsjqTc8NRgtQwPIUy96nZ0utB9yZJdazAMAlsg1G
gkYUgn7ajdPiNMLdYlq8RFUGaRIC/3eyrDRIl55BHHHmq4rEGfstQdZv37iUDD5b3lhaKZj5n3rZ
TB2MMiMe6BARWBQeNpDtZDUiTCXakSOHpFvuG4iZXOYcziP93hlzfRNGG+UTCV1kXUY8ODKzAAZB
OLCYWu3zO5siKcqHn+E4bONUaMr5OpEAXnbAmnRkgjQ4G87jHmeG8IO9BMg5+s9IFTQDyRFBqnY0
4KLlEWqzG05Zb3v8AbrZ74bXuazxTcfmQAEcs50g8KdaVbt5LZUDJbiOAyM6XhG2GGfGyoEDQf/a
KYy85Uw/0ddnVK7TRK/4U9rQtqgEE145htwErAR1mUkNgZvcQogQidmzGoEidFjeA9PK+CCIWUrW
TngYQ77aZbfABkOb7VBinfmluNvWpBmKK1W3VXp82r5O+xAPC/mqvkv6oudzrtevLZghWsqWv3lM
VjRo7lr9KYbrTl29xq11DO6dA3BvVDHoVGek53DiL64PCJOaotbze8Hjkw08W4vhP3TLlUBaShn6
Oji8PF0I8/aGSeh7DNx+Y0DMEMWr9BoKM7iLsR3xp6zYW29vDzVbrvWqrj0HDA1Y7PVtMpqXaoPQ
4kESeQTt2uUr9lukyvizmAelnLWY0kwsKOI4facpLVkcHdpiOrnCNRlZO1IeZo05mD5jMsMmJTPf
7kC+njSGIK/gr57YPJq2+amroMg70F6z4w3xxEVJsrFMbkwbY7qyDocCYie1vJkRixnMIGl7LBMK
zYc+M79kA4CNjqJ+zIIAdjUYiQOP7Mq+eG5S3WKsqEaKvOs+cxhJ6dTeF7yB3jCBQQD+xoL2BVoD
OCJ+gOJ5cSAFAGIu5D3sFoiDXcRRubmXA/OBMeduVhUZsRtK3IffxNgNMdGjX7G9rq1NiEJ2tQbh
NljB7FoaYuuLBUvsh6CRU6gD+BIDtwCC410hFiVOvCoyGqVYsn2/XUpTTaDiqGnwQrIw9F5R5p9y
rx1YGBWR6YqQCXu1YdAVJQMW0jqnZBazypialeGNGLfh80YAgyzqQSsrT4KnfcXPyNimQgWr5lXF
hbKWK11vfqbB9cV25kZ11hTCojlWdfWUMRnZkkC6mqbFQOynLKp5o/BevuvcgVD/M/AHhQCGxIM9
k1ji8xHZLBTxh44jKHMiTYSk1oc/9J0ZpEs3MHR+I3bY82oGweG8zjJBg1zHbBXpNaKqisej8vP1
vcQIUt26FNVPK9kjQLne9+0EoyXidJtvX0aASxE2WRfPVuiAPZYL1vRYGcT3DpeUMbblJg1cjA9K
Ct+hlgUcCv4U+2kXPhta3bbGhNCD4u1eEhVvVOIfPrQvvBG/uAUK5zpwoSJbiowR3KMunu667pqF
7wWU841WLe8mLpkVIkhED5nuiFmgl1QyJVB4WWDIYORXGve+cN60BElfn2pnNQoV/ujjI0tAH80/
aR3h6u/CEDXi0RmUQonoADL8pi/Qz8oIFnR3wQ+ADZvniJWS3qigtbo6W//MijbKKfiBhoysfuVR
hfw/AG6mqUlKqSd8/wXyhegoGz7IdYF6C2umf05aE5x5W5jEG1+h5GhiI42G65DHjIxm92wqz3xd
mdRh4AtVBCPgUpCcAtsT+Vql1GjE1nb0RFNr79q72+dTvEmLr9k0mcqkqchmmOBEATker3TDS+kG
kB+1rAj+QAg6jaaICdBl/9Eg3aWI26UXBgearPXUPf0Th/ypLpwyOujLRH/LHYHfhvS24iZCyvhP
7FNf00LgsvxHJXnwxGE/N3uPsp7nGKXuGlI60GTF2PrPzZu2HmjbwefPUJRH6NrhXMp0wqI5TRhq
ymKsRp4Tn1dU4cyvOWBavyaEUdSUaui2YG/yKYm3ezmN2uHxF1EtCMrToNhi3a1+FFkf+jr0tTXm
dEX2EypPD4RBnCJ1Io0gk7+21gSAOyws/CPHrOceVs/fWQyh+X/rJZ9+P5OdHDntdezD2Xf+/F7V
rNKRxyHJ3oQeb10fGS23rYuZK0T1H2Hg+gROLp6vqm5zYSKRwnPEbeAb1iL6HDWC6nvWBbyiCudS
O9cCJOMt9K0QosXvvX2dcDFIZDXv1kR7K1VK2Qhpm5h7S7Yy7wZoJqRo4X1hkXzUEfV4jtOMLX4I
1kmGAyiSSt0mbV8p7ZikJZL0od1Bcr1Z3brodbYfx7pQrliUX6E6VuskBNohjclVRlP9VcU7sRRy
fNNfWRN3a48rOtufPdikBOYqZMj+YZjotfoc+6BeM0Do7AJFCvcsIQ4eP1zZ4YqALsLRgxh9sPhr
g2ooH9iT72cI+AkxQKxTd9CXrfahQS9tFGCZfVZpxKhLZDCpLsjnavAayS8LjlS5Pg8Kv0ATk5dy
/X+djeT2RXZ7yC2yDmtXIrI3amU9UaFYBczUy1aEdC0ssUth83C3HlYVXLvFW5nYZ9pDNjHg0HHZ
YPJNCZKXatq2OnuCDDhhSsryhdohg0C+15IbNng8bHrKpnnl4UEZsDHsrCJPAMgaKHQQx+pQivCy
Kk9MbLLoZQpO8Uhr4BNd7aGY0SZMthNdcLQW/COwiRpxRd1Ts6lbT07TPcB7ngBF99L97C+/ypss
XP7QsTSDYmLuLJkkAISzygVavSAWJyrUFuyt3qANS2Bio95pR7MT513BxRPi7kTQQRqhOmkvP6n9
N4OXivsWVdkrRt5yLrAdXfERaCcZpfIZkIKk7wqkW4U4AAoXM9QGIxTIxUY7sRO3hEEru03P3jGq
DUFSK2cGsnpJCkZglN42GSy5J/rPfjcALMNV0bTGHOUU3ciEdDLJiiEzf6X/LEAcjPSLU5wi+Nxd
KHohFMLikbt+yfVnqeVl011ahEnKlwnTvx4xtLaI0wXWxFqZJosIM48VZSzb27bxaqICjJHzBAOj
XdtwYtny/HdArEx044ctni1vFxdJVzwp4b28xBtX/rwF7mq9xVc+7S340vhwOdli1TpMsUJ4TpSI
ts5QzpHT0SUndbf5Uirq09f8qI1UNe4ryuTNjJl6CMJPW6LAgi5s6KTrfmY3AP6aZ1sOr9EzQ5YD
RFsUldffrOE8z+Eq1avBbjBosxEZSiFHIzaJlMUJgB8QWFbh+2H1Oh7OpKXb3b1u68WgodARh0Gs
TeO02o85zLfx/KWhEtWNO1lIG7zaQoegggj9mjDT9YsDlXkujuqgEGd1uKTF1SziXQQKg4MEWrAb
4JtU4A05Ei4QsH4pb+aIq14N5i2K+K+gM7dlDKOLit1900m3x9i5gkf63kGzLZZkc7KN+YRpIbZe
9tkQOytLXm5sY9I7Ibbl8OJgmg+F1R+W2LSSCgfl60B8/5OtnAO7jkLC9XFf+nZsBFkyXTEm9IrX
YLp/oBuSi7lhMlXB5jG98qdBGn0kI8wKqmvK/vlS8XxJU974o5Juwfe08jE9392qk8ZWSZ6ZEbut
LgQnE5l9HZEVetnArpLPs6hcuVCqiA7DI3VH3s9gPDwNJ/28oERTJ4LKFfllWyELXDh9MNb3k4CF
fn/GLU6U4U4jZFHgdbyjPi9AUYrJWY++vYi19BACA/E1ZGO+9xGenLiFHMbcF6M44UKz6xtk+k+e
Z2dKGJUYvnVzSVvoq8QUHma8HuTKnMZyCTN9no++AkW7OjBId5cuIiYXwJwTj85D9Ic78Tcy5wzO
g7OFjDF6UjxLix/XjCeP09p24WigYG1xHghpkI6UNr5IVWFBfCkXcFmNxpU9D8xEl8SgWXEj9h2F
mdjssZ1OcNXELlGaL/msDVf9HJxEVH0GXrn8CF5deVGqvgMmsHoQO3DqgCbMkpTzmQovYFay06/M
HZRF1iQTO4wE7B8JnS8R70ChWfMxZz+npSh1+ULfEKIejbIZLKTLHw+3kEW+REkdNAxe7OxUrSJW
SF4G6rg5V7IH6Zam/v0uOvtGb8Ay/s0GbMF4miI86U6lgdCANRpJyRHM8TLGchENk0sfXaBSfvnC
leDQL5Zk9H9Y+4evMC5yNnY7AKcDr6IlqXWafgvLCekVrc857t3pTWz0r2zRYMl+drCNY+eCJb2W
TUUaeUdUTUIhpFjhmA0QfN0CqAF0n+LPHVxu2q0kT67ZQZCpEByqOcC/cO75dnP2eXSdjDKYj0L7
C1H1rpgYvTkrozVD0vFwzYnzjPIT/fFQGluoXL+3m8Tns6v5d1cLjmW496ZcYWS3FDoNUPsKNTUJ
LatzTIaK9UaK+yzcnujUt8CXcX3TtNfLLjkujYFk6UMef3uM8FGkegTFQB6gS6B+3VUNxQo7MpWP
addy0hFiomei5lWMyp29wMOgU42UVPbbfnanNAUbkNJvx1Pn4mnSKdDE57o9j19KzedPidWbely5
4BMOQt3pbOW9i7hUXWsobDkJdO2BzDN9fMyPcfbcs9A35w5o7xkvttew544jouA46ghec2iDTW5v
rQdnvzQwE15apN70DjuE2qNZoCd5A7TnsRCKEWh+4yfDN7ZOzQr2jEISQQUYbUjalYn+fbMF0tJg
z2Ydn//pFQ2OiD8qxBovXJQ9PLxEv5wdd8mTNUHMwB/atosZKSElnm2VOKc0h5HraNteNgAQxuA8
24ZFU0dnoBloVEAGpNI9vfwuOcQAPWIEiHnoiPxJ20zN7YmmtbH9jz0AVvrLZ83RSkBFo0c0Ad89
hS5a61M4M9a2hq5dbxZZjsvCDyi7DnYh4GprXQa59NKq5pnAPW5g4wtWSXT9/rJMpHFgE/h99rDD
j+JGPiFocH1k3/D45+WyDNVzna5cynON5lA2o8pFnMxWLPwoE95mC0Lo24KWeRGJigII3SAVMgPu
TVefIfYFOzXD+cXs3NwBX9d0qmoGi/ZZ5uUvbkeSRmiripVjIxgQqmOG43lM1ctmAESXeEnJ/EJb
ylUai7CYUjqpzV3fRSvhktqInmstck05/uGPLkesL/gCAtMtV2ka+wPUY5rNL2e96t8VNGWYxYl+
l8aN3/OKdaw6dR0TBEhuyMoKiP6cP6IrnL1Fl3vvxvWo0y+BJjtQS0PAnbEqp5Gjn8OfNuou9B/8
4zJzn9vQsngPAxZTOjyfN8SxFQP5J7qoWfnb0BebJkP0P/HS1/kP923YINb9JnlcvP3u5mAaHeQf
oNvea7Dbgl5PDWr5nqiYqLSNsg8YMpXbMMhPc5Stg8Wp26dtp1C+Bmv7yQQ8Ag8oO3fOU0FMEJ4x
p78NEnZSvmseTuO3NpV4nO2LaVti6OdOUyIOlwawAcxIKUv0q5Sc9cmM6nYIbPl/c4S9oGLJLpRK
0ZLdRms9qvSV+OEnvQLZFLnXPOkF42o1jTVin6C2j6KDBUBpriAIdmY65tJsM+WePfiXhMd/YaWu
ASun47pXn/el2UScVI01cgEUsgXf+u37SCiv7Eyv2c/1vmqgwUXa5/YSVMTgXWode+aoLMyfYzuD
yhwARZMtyGIrwgDuYNqAfPWG196Ad3WAwmpfmAbcELEjtniZhuMJpjSG7QQ6m2nRIO8/taFMApuk
RGQYLw43gl6/9Gv5Oh+VD4JXxbAtDbXxqhStrCoO6ZGhrLozZNPiRUMGy+5BWHSPkovPZ7n/SczM
Jc2IbJnNy4cTxUDTHwpjBiDgsNEXhIcpDTvi6Uk1OW7x3/VWhfEKXgaI1FpbxH5aOZg4/xatRY5C
LkxteXT9Rpe0o//vKsNMwGcrY8PDhr2podq6+eAT+QxquaW5T+0okjAU3NuY9v6K7wxeP6/hNbGk
4ZQx949iV8+dHUd7/0k4+l5pzP766s+ePJtE30hn1SY8DDKUuFqIkB+UsJ9sPOktMBvbahie4zDh
tnpfxwICc7+Ylno7fjUg5WTC4uanHbYmT9MLQI2aIv8BF11NIpRXnIwW5EM0nNo3UbjSjdU4iPLX
/QCZMKWtq3BA9kpoY5T2e222oygMkc47n7Lr3hAoNjKL9XaYv5TlJKGDXSkPDEke4bMS1usPaVl3
Ept8PlxyZ68yJlRnEELnDcJlQ3W9dKDMJDciTOmB+q5S9s/cz8Vq28fAfnBcFS0uOAtgzjHls9VZ
xoQ+LYgVpCijwQDkrs7cgukWkjrRV3F0kzaHqnl6cjLnmDJc116dUOvUtGiX/X1psvjqSfPg8NY3
jryrEvDPYb3JcX91vJ9V/uvVrB9yiEDA0F9DAJOlHHn1XIIhvJ8cIxLHENjuCxFuuk7wxRX19eBo
xVCzf0z14tO6e1CX2X4O4opn7zr0YeTwAkX80gmOW4lzRfiiD4aJIdP6DIkMoQsAVNyC3yKSaSHt
H7apDuqIKry2yOqqcWp04A+rnbkDYGOnzNKR6kC6gyTDNQo+IUStVHlPbvrUC4ESRoOqu+UITv2B
OR8FARfaRQzUPPc0QU0dFqJufSRFn9pfnb/l1hJ/QdyTxq4Ag2t2dFfVS1PFtEXPQwMOgOoWvMTR
ermFrTf7fgzKzX9Ko9gkRAGQUecycBSov5q5vS9ucqu61JVij1nepWli2aNkmG/ImdVH8oHoxYdu
ZydVfTR/UI/4Xv0lB9jpoVF/XSSKjnoWQ3FzaqG607xZefOeZ0q3UMoMWuUIkSB855ULWQ+bFJ0J
vuXkGzP9fRPkRpaZrJrrd5CPPdkt+SWnISFA3UMG7UcXRvT02BkHZjMylzeFFW2Q2bQlrJpPwj5a
aCqDPZffolt7osmTUPnvDXFT9dR/iOTaJJ0jlxjWnQ2XtyjwnPbaZ+ihjz94lqF3ykPXl5rmFRG8
7INu4PcGmLBxI52JbXtS8VyVG+MnaMaVUYF7WMltOU48DN0g7TX86AZXyzcPhIaX4Glepq9CsbQS
/pTtVfHP0QGzHKTB4IRZOLDD03qNVfKWGHQAa5FMaxkNj1IPnZylU0kUiWDVsde1AVSHvUxjo7dt
N392nzy5JKuiQBEGENLJmf3tRFhHTomS2Ode66dDw0EpxQRknmS9MBEO1xorY2TxtdxGgHE2FnTp
96ESvBAHBMJgZYAzOQiwHWUc0fRAHxMTP/tzGebyopwYC3G7DpIOUcGOzy/YDq0raUSg44tZ03C/
VQjMUGSonRaYdPazCWKSwMx3ZWNxepjwMoEbDnEU5j7krSA5gOwtqfJJgnEdznYaYEcpg93VznDo
JvESZLDtguORYXrtIp4HUJDBBHTjLOVUcAkaV/wMLBV+Kx2L3gzXTm5YxA2P/iEwvqH/Ir4oBnEQ
XuRrNcXQzb659C5gfa6rrMaZxc456iHyNJ/rMoJodhSrDHT/2NX2dmWhSJNr7AiiSvSOa+AMtHJ+
EDAovIM4CG3kIGSPTafWWlCa6KRdJMwLX3LfI/yDg1YqcAzI6k+Gv98J6cYq1+l2sC4zOUra/W2g
OgcjOddMdvhUwOa9Gy0GUXpBOR1/4ZmdF7z0fjM8jFrQqRPZ8GreircvHOVktizigr9GI3vYHyub
vbZy3570KHKMR7MFQldPcXPYyzWNGIr8wEeGUJStlzS1I75ehXE1IFCPQP4gPkKlJ4NYJ5wGnu77
J5ozgU80eLnnRYR5LqtBdzUBaqAdUJgQQXA0JYvQ6LMPU8RDAwJJ/ZlWqcxKl3sHvYpN7RJITjfb
SJxKJRMFu/1D0skEczHAb4fx312ZpQccqgm+iDtZ3rHsCdC0Q/bMg4aAHOzJTgFW92MzJJbIFxyA
Su/+tb3ijRZ3EKnuDDynxveT4xDkaHRkGHj530DP06yHyYAiyj+fEP20aXCmuyDKN9+ejgSWnGJX
AGaBRbU+6vbrXFMnXiFYRbcHMTjzkIM02VmOasRUSeP+p1qiFWj8u0EDzFZmB7+CpcLXgZ6kPgI6
mqSNRY91+9tXO1Othd2vCKLj5BE/oXlQ29h58lF7A037P+mtVCdUQG2lFmNrsbo4ollEnReGci3D
SnIBCX9tYIRRQPxQpQCL3SdpF+ICOVhdAw8cBT0BjMUpLO4PsbZo8ZOE8BQE/tbCp4vPZrz3rurZ
6tszBgbtyH0KSKnRITj4F2y/R6S9McSzXXsdCItUsvXwal8d1L9Esv/hcdYHKoKRnG8aIjvndAAz
/gIL8CkFNApewrjkzZBoYs4AP23GXw7820jJe7HydbuMz3N2I1MpPLJsV1V5FUJ2EittJsNSQkbX
wuyc5KQVo4yuN7wvb6hZTaYVXltqHdWPH7EwWZlk6iLpPzqmYU2tSsP90j/L+028O6R0Br5r5FKG
Re0UAotop3TsKpdcMr8/FazOsFwpYNtIP0IvwPzPH1oaB/gLhLQSL7f6z1acd7OUfa/1R5Ekdre9
y5jK7c3LYE2CuBQNTDNflLxwxM80A77+AXPEETqMYgRgFbzBBtOHYPUr7GOaLqLAOGFMRMm7ibD7
suuvlDy9mL2hyBCtTHwK1HzNQr+auvvy7PLHLQSmA6c7XeY6ybMTdkurd6UiENX3+16Cbm04uIBs
/+YQKvqEJjoGvPBoB9TMXWzEdWwY0qgu0kWoSFhwk9p0FBwPhTJ6TkHtY0LfwDgG6QLdSOrbhMlc
e+hIgnigrPAgB0gvc5TqVZ3OKTTVbunyBHNLWvbujbxr/HYr+WU8D3WRK2UmDutl3KPuYw5glUXa
fw+SKRVE0ragN3weBLvu5DoE5MQ8GSJNzY2j+0iw8SnOVZWUZCK6gQQSIXsOGKL8cO2gDubQMZP1
11nV5c/tNt0yhXd+NBhU3m0upOrWHp6Qu75nlHyqUDAKabALa3QB4tNEL87mzfn4dQanNi91RHUl
uRtmkrObWQlPs6OJ5njiq6kNt4p2JGXHocB0Tru6DE7kI0/Dn5eqDUSeSHN35ySwGXXEkhlaxC9+
yfZ+/i+mLdfnkBpacjPX7sZR9WtMxBCiKSvRIc634CWK/2QEoS67Hr9MksGft9mje4t5jXzyDmXT
dKkkAiangZ4TrlVOqp+6NUo/qTb/Mit97G2iBr8L4XEZl51rJ7z4Qbqruch7mJdYIQregJiJCTRZ
cTlhdVTf74/Ex+Yb228dzgRhwqVnc+BPGt837h6sbjJVjl9l8ReqWp83CqT/Nnlr6EdXG22tu/cG
iZP5mld42PpI/QLfRNFiKMosS5dmtlwOMfx3ZZ/ojItXRjSttAncUXKi8jmxFe983U9biQgWg5dt
XLzJuHEl7ocgGcvwQvzEZu83LAdXGeNRzFtxmvRWZVSVOj+8owhyiPpVmMh4P1ZtLVaGNdmMIYei
pTAxpBkCZkXB6o/V0rpcpeL8ceG36cxsHCwyjJ+5IOyi8GJ1pNKK8bYAYtkklmmgKdp4duXRyAoE
zO2EqGbE2bJn553pDd4qOahDo3gApMd0V248WHVYw7xVOrEW23BkofxZwm1zMv38ruPkahPXNVj+
MW19khE48C0hQ4ado3bolGa3+MGN15Q55nAys2wmp9dKOYAYW5kJRtRR1kjLIK+JVWG7/8an+h19
lpiZXnRG9hwhXofpYiq5menpb1sq6A7IwTQT+0zbhSDbkfBv1bis/6JLNqxelCK+u7trhUvU3lNM
aK3Ov0ZtHUxhnRHZo5iYff2rmWRjFLTUiFCUqQ0YO4IhfwZlhTsjdEHsUsuhdZrdjpjYZaF0s3Gq
QDcZMX4CWGm6LXXGc7eMhVsLXx7GASii68RFaGLCPBL+mtYbYHTL0pN0KEjve1pV6/cUCXWA+TGT
6KEK4HWLDxmtkvGKGKtxas/5H3kpUSGf8iRal4KaCssfqKaq4oYBVBUtHtQrdPk8rmzM6yFl/M4B
2EyFzmtpIAm9TGeONI7k5kUUyj0n+wSQgEAQIvZTv5zBFpDqiuCewjW2lO8kKdN2vRmIkp+KsVAK
qcMcfQqS+2NcGstoNQmNSB/h6Ss+cFjjtqvuF6QFUEPzcBYoolTE8X3kysiQdvWLEBiKGaEVsM9J
jgBkWDCtFMhjHssv3i/KF4t+QN3QYR9FPUlssc2wz3Do0rJNXOem+Uj6UYMKLw09qYbyHTM1G795
dUG4hhSmi6xh/zdkw9wCYAkmOQ43K56qnReAl5NIH6Le8f+5tdKH1x6Njc5wuyE2Kjt+8A8hwI7J
urni3IH2HXUWdNAyDkDj8qOAJnzs4S90bry5bKKJzkpcTb736rHaXFu+mg/NCwQE3ZBAkEKjDlqp
4v+qFcb/br8sTE0P/uMGwiRMNcsugUwD7qFVhm1oFqO5/4dt5AcT5y3uIYhMC4DWPzqJQWyDa0pS
m7nZOizqr9IbsE9ULqvFk/kc9aU1mFEKHuSjZDAykbsQMP35RUz/OEqdz9d3A1Av64+9rYzLfVcA
ALj1iNYskRpr6Aa/nTa09EsuxjypCHkWgatPWK2hcuJqe7OwGkznD2OP4OtXYsjU+de4yBLLT0qf
fdn0WPROIXifdAL1hVC0/FwBit5+GBa61FMAhmX9ZdKNb1W9UBwudhxcioPPFww2X5/1z5IHZHQ5
nkeZ3Ia5eFPsSTzzcgpmQowo6VgyeHB+BJTkrr+lbH4FY9P9ksrOG5FQ7yRjxwnqcCuM6KyV2ukV
eRAmrOh5QvfSmzEOfKzg71ip6aIXplEns5/V5slI4VkqntflU8hb5F3psjVZQGh9QUlNTzz9mfCg
32edXeLHmUqDlj+3YGpHHaGq4QE9WSLPPZlv3hvRr0+m4rDJCffMguBtOyDwhsVFiSGwsEaro12n
1r8Nqed+Njb4Yk8xYhwaJ9TfTOlhL4rzF5ZaaPtZtAMhYikcvCH+5YoQDf5p/XWCvP5gFmK8a3W7
W/USlQZPgoYtPrlBiFSGhSbPdvm0p+HdrZi4LiZttNWP03sUIcVuYrBLXLxpa2BdNdRDq+l6RwPo
Rf+7i3Quzi+YolBoF4aPGl0j1RNFkqxbZnUlBr2rqvlFajFiW85Zxv62++8K2/BCbLRVndqEYyPc
pEi2PESkmjp7Y/M8HgOtPr3bzrTeJVp4tBl/d/PzFzwHT7UCbwZnBW7LlTW9642bdDy88Ls/YdT8
LLLWHv9fQE3VhheCEI7EZs8dDBzdKmrzTHrjb8BgyYfmbSAgMwypcgjWIKO8WGC416WEhmYhb0HB
WMRm5NTG9/wU9FTUnZJAo9W9tpMyER9wM/rcgS+ny4T0SFL0kXA65diuZ/4mO+xo6ErrxhlFG/te
2mbg97e9V8Yo46OE+IMQX4K4zqxDKAKUtTg9ZKjDsdzzcgDO/Mbryj/z7+z6tf75N7zJYG0Gh7AE
ygxpGzJooQRFpzkzx3byBGjoPARBUs7DlkCGor7U6ilXJI9jYSAAAiURkYpmBvL8OfWGiu+S6TgN
h86FBWm3pRcO/vqd1l3VN43TJp2OjjJZlSrlV8BDvrG/9fWMVjaFUkZY0gXn/U911mSK2ewe8Hzt
5/Xt32XjVyy1pa5+XbV5FC/lC31k6xTJHaLvnHaB4jm3A1RO7Qrj5xHtmmGzNUUb0tZZqmh/rEE3
iwxc7pEFSDml6OyrRClw97Iybp9VTexzh5FlSv1myWIaWeQ2zMMjhMoHIIP/e36LZFC43vVc94wC
3uVo2/bBxlim3gnPatZcANa4K16b73ftZn7WjAZhKGCcud84ajUN9LFkf6cdHY9pItxGzwKlbnYs
w3Ads27rR9SlwxT1aeIX6tqvKWRVidp8c8cRezLXvGrwbaagSPdeEZ0bXV1hoTQL5vKKSg7xf/M3
zLmK7ELBRWWIDxrdcSb5Acq7qJeUwbtCRKjf+OMOK0fYfFh5boo8UFjfAojtCb1snK4WpwoJfMTq
Q5OW8BDYpr5I8CaaRI0H1Sy3u1vxThuCDSs5/qx/kdxL8xE+ias3LDu7kGIk7bHM09d4YWAMsxA0
eXZOw5a6dKjnkCcOBTkX8LSXHP3rRJPwh0DIgrdw72SbhFri/P2N68J7X8czKMhtUv4lGWTK4Gf3
K8iYpU17UdXxfTheMmQAgGk8EEn/WCwklEUgLCEDpRReX05RYqp8RjASrN0XMAfGVgJ2UC05DjGV
+X7Q2uWowZNYpuZVET8fAmj+QLJnmAlEw9oMC46g49Hu4kClxHCDLoO2JL1mY9YAKR6+QHGgXcPx
24jMOOnkLe5ikcHVlm8ZcBBjeeRnglhdf6TJZxrONsPt9Lhl56pp88xCrM/b/1sXBedvsQIzeC81
25rNce4lQi0Dcr5687Z6IL5+qR2TBsfvv45d+QJV2Jen7FQL/NMrLXGqbykT1zeeaVBf4j/HRMe6
oDfR687EfJbj//aH1mkt3dN6b5NnIZ/pCKOAO9TI96Z5g042a+JVrpqivJYFvLk61jxFROgMZxqh
h0x8cmCtiNmgav4fPW0gdYFIeUbvfrOWmqHH0E7JRlv0ApnPCpTX5TTmEra/v5QEdnkG1+RkSBqd
IOy8h5lb4UEvg0HIWn3WIHIx+n1wKBuB95IjHnMMMTQhlTWCszIAbAswThwirBbSKokvvr+iMI91
cGa/eWUV4z1/NCujUV5zaANji1rDmrOPiYHsxvxEISBsdwb5etJ8GP+l4+GSPRdOAKWP+AvqtfW0
7qKPCtuGfq7HLe55Z+EJJsDQWg7EQH/3aKtDsVo1J34yHoU9Be85FT6VIAPejcVITC5dF6hqKk6O
H8j/WRg2UBAkVuiSXCsbAcyyNZxLtQcY5N+ieJQ7u4INir3jRsDNPkUlyariz1ZrV83lQscF+F01
YglcmviRM5Ggg+zs+k822gEIfhKSeoOLPJ8DgP59jjAYaFSOGrDyxrUdg+6/v/kt2h1dGBP45PMm
4Zou4j5xeUDC9WVLrEsVxsybqqIk04FbeG52KIzna+N+kesbUsrF2SKzPl69YK2cWiEVmjAQw9aM
dV+kJqb50Xs7kxLDsUNEdViKBoOgTaC1DBUYp7pYYN4BcbNhtaVBb4dRC1bzhNrwPWDZ27m4ntGH
ON8V3ZHGEUmP6nN7PxQm4jHeFxV/IerB026ANw57lZnAnLNl5+d9LsGYbzYjj8pniW9ocZSg2QYz
KhMlkvdd159IolBRF7/76yEXm16iJCEmTtuJFQJ/xd7b5TVLqFmFjrLPnsSE1ml7PB+wUVdjBj+d
Keq3q4bu4XAm8I2ABHfjOb4kuQ+pSn1kKQOwv6JRkcfi2gwhaQ3RaszQaeVUuVcSwN4wxAu/UB05
mVvP1cG/5yiaENIedXxLMt1R9dz9vtO5da0r5b0g5Qb5RsU79P/kDutGVDZLa1knz+Vf7Ygg5QVK
ND4WuHVhfsOzRE7gpurzznRCyB0zE/dlqzLncRSCT/rkZa7iHopbjGMOqxDY/VSdKV/SthAoZEk6
BJrh3enBuYj3hvdFM0XruEcfZdit5YzkTrzayDvXhlohlZjjhVRGtgrFHYFVdNvRWqsMl8McBcWa
4CWzDWIp6zJ9AER7n7COQoVYtiNURl8cpxNSabj84lkWwF8MwqQif5Qcmkt+qkM0bz5IceqMBtAM
QP4BZXnvakWXSZqAAh1XFowlm2jC356jqNyrJvFFbVbxQdvGcPUhl92R26RjtXA7NfEz36MW4LXc
SNJpw1lXy5BsES+As9iiy7rI4GnYocPlGXRknxNuBW09/oZwlql0kC3Z+7w0XQMUyAJOsj3dLScw
yU00h4zG9L0/dP3t3V4pRYiFKdI36P2W4OHB54nrw9Q7ONqeFqOwB4Y5CR86JaNRf4/ALWFLnkXV
AhTZUNEbQimRvwW+iD+cgBGw9or7bkEAHGmcv1+UP7CHukhc5RRB6TqVryyAj+HV07tJX9sCaKee
dvQxddFKzFMszWnbSmGTUS8LLLs+iGG51UkysSSOl+8osmDMd4wrABtdxQOajXFdx/lqgdaBdo9n
xmZ0hjNZEXmlVLVWNO9eRqhGCNknrtZc5f5jbNpK924AfKwzwfX/hfD4+6QBXe6/+swZc8Bs9K1x
l6dALHXdyy5oTu5oxc2OzKHDotvpI4FxbtBvXRXaSvcDmhyWrfWt5ZYfyz2CbWIuizgIJ+ao5XzY
UBPfcFKjpN8dVjMsaXBSg9J4ABtLx+4ltT9dE1AWnxMqIz/q9OVelLZbMJ+9iJcSPrQ7jwKfd5IR
WAkbJiA0LVbiD5aWOjs3vp2V3OOyxA8w/VeCDm418AIHMh2d1NYmvcroGshApjcN9EDLDQ0l+mXz
hKQJrrkgzkToiLqLRRnml38nfubmCwWnvxf3QFaYhpaZiLQtur2Iubd7h3Tjoxv+9FPLWy/5UvOp
YiZ6K5l/ojbKDg6N2I56Vqvle3DAx3i/idpnhElYFOy+R1176gU8D+nTlQIn8XTAWLFdazVOAvnH
Ht3FpWnh5LpV/tUZJAnYWwWVlmGsX/zXna18al8qdulPrZGT+ehktoUCxdkeX3DG/bqrPNyXiFO2
Q3PH/VVVgcmMcaYV9jN9CCOzRp+wy86wH3zw0DRdOPM2BjOLyMTrreIPttHd8KiW41HnTZBzZzpL
zjPE8+B2yHIBCD7YkDEAaaZ52reNpLVJ6yra5N9hHONW2JGStG0awQ6W/w3feeBaki+07dVjqTDP
BTceWCPRY/a7XHrWnX5LHs1Yyfz691G0eiF+yfymO2Fzj3W8YJ90v5euEA10c94WqJpNR/o8WUiX
w7Q0tYsXjHuzIRUkfPOj155v9fNEsg3K6IYmEP6pgC3POFTtNUWhQecj7jC76Z9dUKHFT0pITjGk
LUJ7EpCwJ2jyYwaq3w3RzQHcDAGQ5fsE3fFxKaq/j+s61T3bLKDodeRr+S573r+Or8dDGgeI+3Zz
0CAJKWX2p3iLLTSn59q/o+qK8pT45ThoBHl79Q54jAzhevpFICVC4peH4kPj5GLCCoUZE/33nChg
VEr3IaHOmXuEmEJgsv/OfT1mOcLfHOPx+BW23CNXUVzNhrme+MuhQpH3+d4so3EhCLu3BQ0FVAif
OqLIB03rpIZcmLshFHFh1IdfD20qdAlcgYK/ex3q3HDK1mHG4f9StRJMgYBcZvudJ/yGA/vnGaTo
atLIyweVBNDPMR737Evye9PYf5NuFQlHdoX8L/hY2H2J4LwbievzT+C2WjnO9/ziSZ9qHyVbeZ4+
H4C44jp6B5GR21XZfdU5KiGYPcyPQVnXyEp45N9rTXS1kzErfr7LAdXmd8WDmJFLpbm0UqqP8eSh
HnIxy/1KpnfRQybcHLMDw50WJySnhuuU5n3mq7EIFHg5cfjYbUQb2S511bHLZtgwkjY5Ds8fozmS
ReoH8pqvxAlb/amA7MVV2J5PrZGocpcj+Sw7krUKxO8Ij92YAFuTRqhdC+BPC0v/q6gFzdLG/Row
5ZIOCopSKr+IseXRvrNmjQE/HxP6jgmcJTxeO/LbPXFEG3SDJ19xiwdBE4UJu5I7fq+rH03izgvF
cwYa3RG/gW5WtG4kgzOS/RtgUHVSfxiE9NRNHIu+FwCS+v+Ka5z1Ms9ae3EhXfOUHP3EHDw1m4+2
WjgyPU1d7sdgbdYWAqelkfngU2vNDcSsOEp9+WvLVVVJeSfnHz98KT18iwXCgE9KXsHKL6QofIYo
mT4ajKH9ZcJq3bm339fyCOAhuKyZWIYsCULeJKq3nD0qyH333V8xq/H53QP6u01VzTwFIVZ6nQNo
jZstNv3ly1pck8QaAjLNPO3mzi/QW68kph32npQmkC/2TfCMZespJ9ppudwE4mQKYZx5VCd3Z3nY
Io2qtfYftLbxNNOrGDapI5ykqfUYVT40A8U9Uc1tqF/46MZtJ65gDTKmXIgI3XXuSRd+rGgxqmj4
EaoS/MTM2EXP8auaWpzZpgHaILiS+SjSv7y/xVK27SZZDi9KLcthDY+QpYFQlrM/rJ8iOXW3hMvm
Tw5zAs6Lvsjx6z4QZbE1j2+X8osQh+9SZWL9ciqkCWK/eNJHYUx6XZzqKJuj4wnSul4Dny3nOJKa
W/CY6TQ/xaapjKzzKq058/vYxhqecJHuURK1FiRe0wWPdNodD4fuCITGUfgr85rzUf22pFVBisqo
xpjmaYGdaa6GLI2AHFT4+7gRJdUsY//oFKpBHASu7YpDzy28NmlGY+dOzCSIBTkLe/W/D4y+Uml8
CY9H1p1FH9Z9d0iWVbnjqrO1l/36YyqU1dcjsdnUbTwGX8RS0SCyAonIb34i9t3pZLsBsKXmgihv
X0zTwhT1r015m13hssJDS5AipFKJwffAMWsRGWTgymua0bQ675ghrxRdg9kbWJSuYlYkK80grptX
2CoRl4arzuMCkz/QdnAJ9nFNGmDyS/TBhj9gZiNRV5CK9aqUQ/eCP+4TFeGfNIUy2cL4Ji7IwPdk
tiBZkaJVLhOWlW8LFXnqsE7r1TYSdRdeFHtFd7Lcxhd4O4u5D9x4sfVu/PH8NLd7Dc1cDkRW3W2R
x/MlhsDAiRWgpS1fLUyCr34FYOU8F0q83DTWB3FX++DQD4jMACNXuG79BryqYyumF8ICy5e3r0VS
PqBrcKEv4Bq+HSNdY+2MyUGbzHRPj9wup+5HYS6vFtXfv6N3wBvUydRSXCgUZlhFNTRievVzuJxM
AQbu12zZj/CEnF3xoO1o5V6sCesx7i/5aDLt7kCZCazhYL/tqIEvxju5VOli/2LxpHnl0+LsnKFX
Til1HwTeveFVxV0S036RvqkhdmgwbfiDK+ZaVoY/RpO/zweA5HR6QPP3caWF9baRnKq/qHkEucRp
Oc0FpJNj1TvWbGM90qsdzboYLrnnz0FP/Iva/zkrEaxZy9PMsxMbOPZHBbFL+4++ZdHHDofirqyk
rQCcsBsfNdzjmuhV0aRGGJ9g/JfnCtOMg7nUTwOkdlId1rfn2V8WhcOe0B493tKOR1q4VkfXie9K
5EE4PKqf8qyB169q8fARflZMx+rSwL3XI7NS6ieg13y7WKtxuNZxZOjhz2aXrJzXoE4d2DNsVxfw
fL23OrrdOes/2TVVsScYyTnBYBNBi578j3uEer/Dd0aE8l2b/9N4f71YciAShEcxqFCvhN8UXBoO
3fMw6JVjiEsG/Jpd85OnOrUFLFRye6WvflZ4EhzUTOmU6hfMDkVmfHORk/6N0lXKwNjSZqm2sAeQ
j1P2ZijDAzaZe/y7I1mMiyehBGm8Bo3TNSGVAzsrK0Pw2Qcff+pwbmf7CtLA1rm3KlXHh2i3mBpR
bdKlKflp/iR7K0NfLhv8g5SJE2sluKf2QeGfdduv8g3aGwVykfB3aLMqhIEapGCmGbs2gYhUQtwB
l9PDyxrJ4dJcqZ3Y4z5/DXkLW7uSN6rdss7mNG9U/4ACIHJ6NBj49bSZ40wjVH10/Wg5HI83otEd
HsFDWGcyxlm+e6BvTBczirn0RyRdLlODRZonn+Zx3E9DFpQADS40jUWddfnoveLB3/vUXZ5NyvED
xIWSkxLyLgfyJsaUzzuH8mooJc4J1aI6OAF8FrBJ20Vg7LCNCa4gSbVEamM06/feq/vdhbv7B8nI
py1/RG6kDqmt6hVBR7rSQwtCj/ceSZCGVMK+oDHn1sVQNNUYh6pwN8SeBMw6+aMthplVNpKR46o+
TPupUeKDb0oGEjP61bepLLsD3mcVd6L7Ycsq1Xy9pbF70AaKQ3nvh4A/azTAlt7ptrRJ8C0RmmPA
ETGVRfLDMQ7wYs+bzreZ7m5BG9MXfqYTX/RDc3//6ZmXmoQz1JvicaEG2bygR+x7mr+RKWrwR5wf
83a4XYyWHSxKKcOzROue08folaZxzcNbZc+EZFslLqK1wzwLBKK72JZc/1E55W+UeqOuc6SKCD1B
bzC+OAU1JubB/1Etz6VSgjHm1phCQdA87n/GMB+YV2ZDuVeMKFXcLlZLNzvQGMIiCBUnQvDNK+pp
H2PsSHIM2RfjniAfSI5gsbBjGzAAFQh4S1hRJ34X634GxDgsLTRl3V6GnA9TZA2iIJ9rJNn+ZK8z
mE25Xn2IxXxv8+jKB7cc7hGaLOvgHd+AYvdAmOhT/KCb5EN+bW5coT+8LMd+EmQAdxeqCBmKPT2C
m5O44ncfFwJvJ7fLV5yob3ZnbdyBo3B8VgY5WZ0zJt6OHhwZB9gmfPxy2d6HF7eq6maEFvWQ70Qg
dMZv0YH96c+WusjBoyVUg9pZP0d0tmKcG4gCvkRuGFzETbcOg4RVXlbwwsqr87/mffly5FyTXe5N
9Y1HqmFOZTi6xdc7FMy4xXT0nPksZ1KptSfVBo2W4Rc3S2iFSzaA3X/uQ96ybNRUVWxD8+aVsfLE
7SBtcWOEVmcX5BEetgVKFNPkgGbRlypLZuCgBProxzo6y0gqfIrmpIUzdpC0y76K68WR/nsMWoQU
5PqFkFwK8BidCD+DsavT7T+oVUhKMgHV49qbeI+JXrFXtFsSt1xj63r6fEmyBhxy8sLpTW5wH07/
Xpn3Z1a6BnGROFXHDMZQt83Ppu4KUYxc6IfD41pRpDuGSWX976Ob4pOLhNEDfsXO/fmu7K7/bwos
Qt3qEurf1am0VeBDGu7s3VPA5qVkHfpZ0e/dmvdoCmVQSTqrRJm3kpCgNi6rYkCPo6mT6r4CQ+Ka
cDlh+GFoQjUkdUnPcJdQ77cu+NQVW6Pkza99aHMT+/ctQipmCtZ6o+Rw0jF0NOXOD99x0fTZttB0
8OsSUoFTvazTPoQzzvZWDvWBYbcyJz2hYeXp774q6YVVh1ruk2sx5iH+Bc3RyoHlkk7WyiEagjns
bzfBx9WVhZjT+aRD6r1gmOcxi9ObCFVbu4opPCkOiEu/aywDXo/+zGqrNvAPyIiFBfTXCtEPppVx
439j39rXH2gE/JVXYE5zHuWNNAqd2LhbarTWFkLiFZfzk44Z74aClkd8AqxoU6rm14UliqJHm5ok
evCmVx8Gc+kgV7FtVbGLL52ziNFaYy/GYfMx62BlLzrjiChl+UCFRMvVd0kRnwtxBuFdH9ORPycG
ihMnaBuNDH96jqFwUqwR7I4h5D8nIp/fHPV+IkfarEdINCoc/Q9mmy1KJfYpdVuyXAatN3ag6GMI
x+mtSJwS2ZQhMn1O8EUoIxbSlTK1FujEW0wmDTwoFgEJB9gczg+rpYuVRwJxnrMvvN3F0RwnEA06
Ki3rP/d4nd1Ol2Qlf/XWS/d9oNniyfp0nvax+gdEJnu59ZGyrJlWYHfgcC+4HpYqjejY8a45aJ4d
+Ut1v8F5PLDlqPdq9azjeYVKjYvJW1s5xd2JTSkkGccS+9N6Jj+gEt+mZ7d0MXdstlnGSMBAw6Bf
cZfOWLHOnSTLaIx/aqh3uBzlcLdYP7wTrGTIUC6YVw05hapatARmTq+qTz91IZemf8OxGii7xRwU
Qe7eYsLs9kC7BydSk8sclnbZHhpFPK8jOMJQjbo24kPjdotmUpTfy0CJ7sPrbmHdaQMN62C12PW4
w4nv0LE6ZbSqIYF+OtJbrRforom8+oqORDgbd7fbNYtrANM8RlmKttwIFF1/lR1/C2ujSe+p+nn2
3ppInzq9PBbS8GupFtb7ua4eVwMJ8KZ1ugCG8OsQPh1r4OeXfJ83VP2vwYnihHVg2E17S9D6NXvT
bu4LrTtcKX/9TmYvlVX8IcQZmzOSWiP9pXDSo6tfBY+OU9djgR1TDPIuJ6AVbjvtfbTOhHQTkSIt
ROtRzCzTLpPdpAyrrAGdDHFat+Efptf2gWixX5XDkOubkBgK8CasumypHbpF2mnKpMo2Vc9qEVFx
I0yvoUcpdcXIq5FzFE3ElT9CtVRPUgGdYKiFhjH2LaGFQMLitkggxkqWPG5/fv3UpU0hm4abt5r3
8EHQ+m0Z4FbnQLDpRQokb2RofgyWfuFlNz5i6VMT/xJ7zNsYrCCVGeHiHS4xIr4c27OAe1mJTIUG
ikbmA1NTz+4C/B4iW0EQJpJ2OkXGljcn91WpDH/4A7f4PMgYV+z1/fbyidNtBeDKm4Dw+OoyJ4Fd
msxRR6Z1vt7wYXlWGR7Y+dsGCommD5M5kDfNqYCaUnUWLwD2aLqSS9ZarR1MsMcemXUN6A7C6UxZ
dwrDZYUMeAZ3RGSyzjCsfsT+l+Tbzw5BvzfwGIqMYGnxhtI3U8wq3eUk+rZIB2Lmf6y7OVg3xxdK
iEnH8W0pmdMBYOMgvxCIWqAU5LeeUnnrmtY+NwOJfWfD/uBit1nIghynqTrQDH6HnLeTCwEetyr9
vKnxvr9xgsVlaXrt3LTwKnbRPPs+RgyjixVVEdUPEdaAfXAf4F+WTwGTrU+OWhZF2+daoPDzfmfO
/1vMoyLZISd72k+5xIEJmTxQb8v2WdrqbR7sYWrMKatFGquyFkwgbygyXNDZewaV2LEnTvH6MRqK
wILj5wwL5NfX6SKv8kIzSp4flikkU/S0ixBmwhwT98Exi1UTAJk1F072MMYLDD0DMB6/0+XzN5++
qcBNmIPYqDesm4F8w0HdLR3b9x35Yz7It5WBrvGANxOHRHhBrvxdt5N6rRI48yppn+ICgFlqqYYw
RMl88vrzT2L5qDi/xd2phA3h9NtRk1xwSS7fAAbHpO8tccNBgdFLROwsYs04vxgU1EUfw1NN3w0b
MsHVTygL2oFH+OAh+p2N3gcjzYulE51nx7EMnGaK/RjwQrJvPTbXNJnhY6XSDAwyX+w2n2LrMuU1
+lkHlzApOq0NSfVas/sJ8NjqzhSbPo36Qmx6G4F0nqcJC4BBU+6fZdNczA5rRL8JXHjqN+T6/qdt
hTHU+Jkj3sXFOL6SK9wV5DamufziLGppRAQYg1xFsgB/N5gfCQBlRKToPovQaSMwwhCakd/it3BV
Vm+fAvGjIxFsP7dKd/JEjnSWQiCDXJ7rbG+i8V6hKCuR7/CE3byrWia6LajLxAgDb/LcdV8TaGyc
1heL05mZwwUDrd3B/6B5xMZKY71dD38vEyqw3N0bjJgSV+ByiPKLgGH5VUVZlpm4BSWfN6YyTbEt
3pBOFRMLaomhxLeQ9wYR6IY2wDAk2+PYKN75fZcB9C1IOiWLs9jIkrHtoQTiyMFqPCRoeFmEUpip
us9FqQxgpyPXJyrNGmiJ1FvhWU8Dj12MskVNBss0jkvas8eGNYirza/PZfROoNmO8cp397CML1BH
c+ZnSqJcy9NCWeObC5E7nTFb5prlwCTtEJmliZ/eqW+2RN4LVdVxXEMpYAHGtLrIU1cwch1Ud6uH
KsSNjbjj32Fjs9AdiCWE20E+OXIxfDsSfTG42Ps+k+s6oAvHpiuAiBn9EaViP+xuaOPgcF0XgJc1
pD0xf+yoY4zU0524VM00BlW0w3Tds4mHqeMS/qQ4wmPcEW9g+ObobXiU5Hk3OXxRDYcqSSklckej
jn3ie/NsdnO2sbEQE9Z2qATdyYydgIGsB5kSFKhm4hFrvtCu5B1ygCsD4qSOT3OhQGs/r6D2XZHG
3xE4R/qlL1vK9qZ2z9nfL65/xgWJVeDYJMjDXvMm6mgIF25Dy3eYMsV6zEnWOg/tDC4jERENjoji
fIAuBOJQ/YiyLT0U2cYtZTy10rbe+m61rWHmqS9c2TE/UxsVsfuMvgO6tOhvITzR5sRFUxUbXnds
BoIi+zQAgqXK62FizMw3+XNVB3m9slegBNwDOU5rcGnvjpsKrU9yjkDyfJdiVjFvLBuUU6KKJe9m
OjzqRYiShhyW/WozrFoHusQP3avQzTSJghWS4w5zGP0oBN87njLPfTPSNQzF5/ee6Udzs4XwkvSl
cFh639ZDZT758a0u+8QeJMOqChjpjjggrEwkgExDxhsiF9zVWIF8WYAd48K8bXuzjARAZaabgLuc
B88xM9CQoCEOzCMi8DuiHGHkijk0bfXyDh20Pzz6FF+sV4MfDCYGZH5DpxQ56DjMNYP/6G0wgXVs
Om2qU5lBR0wZxKBKqYREBNUMeHoQob+DC4iLmSS+kvuOz2+ZLyStuqzsa6ReLG2GQBTc3ATja6eR
mcao+XaVKH0pfNbP5pcoj6baP4m0NzdbpR1di+WY06XwfnYzqJNsUnwwYU0QZm7WW8dqN7DfVnMf
xctciuRK3a0uEHM3Uj8AEqO2PPKtRLMA97PifyBRtLy1cJXOEalqALWX19gw0jVaDJrLhMDrV3AS
RdphKT5w6iGvVlYtrW67KAxCJlL2va39bA9aAn/LHijkt8E3BeyYzXtwEtZWScLVamC3/AxhSYNL
nzQMhGp5zQIkWWTfmS/5zxxcwhOjc9dBxLAN+kCYJL7VASdQjUuNiCvz4dJxHHk/JSCICtahx3YN
YNEGK3Zcu+UjcaqICbFi2jTBalpQK2g5kk9vMqCgwc4jlTq5cvGQVLPs/2cf54yE/JnxauTxdzsd
l7od5lvQldEjOgdQ00oi9+xiqpeIlW/g+cySxXenBwNdI1eofdjyQR1W8+EVEkuvPPP4l6TmshLe
yExQBb2uBUz7/cZXfo6+7nSFgO+YhFi2SUU+W7KXg821BhZxcpXuRXel9jQ5L+ChRoZKAcDHxGYf
4mzSFTreM7IIwfQZCdzvV49gyseNP2yvJB4oikKuyTr8AFgaLus08zFkp06qMM/gN83+pCqeQsrH
Nea6Vx389iXSphtHNlraPvlX/O+UpylW2KOv4cwQeRA8xVscimzGyiy0Ac1wuaLWb2O98B6Ybn7N
XoIgrr7sU+vJybxS9eLRCf6W0DnCxWu/KRI8fJ8Q8eW36Vdazf+Ot02SjDSKfUe/P4Hu0lZA9pG/
mqUEz8ijpmW7kgJT1IiLt+qkMT1p8A0bhgh81LCwvCqsOwpUCCRCrpJMRCu1C5U9zyX7dgm4wN3C
m4zOx/WC/dRuFynPImjwJtc7mEI/kFebyw98vq5vTGOtcuZAe1uOU4q2RMCdShYo8WsC8yKoqQLd
swnQeBJduqfyWzd56MYRhegF7FXKkZpjzcqQkx/Yw0Bngfs5rvA0NnauNJtMjMHqwedTesXCMqgL
sttFD8KMYldutHYzLJ16jdqMP+xiUEF9UuFc1mtUG3F4dNXzLglu3E6wuUWT6p91X8YQkzdJSU3i
Jqvx0EOTfpXX0gDt4ggY89S+1nxJlLNnltcENqGGJHnpBdHomWtyQanUCI1VsPufwe7YgjxCnt9m
wCnshHtDU/8snEDiqilG88SDfzALtYVBDI4xzIfy4Mks3rbSf9h8pK+PSYOfNZxB0K0AdIhS9F43
aRYnemAueatCB3hNy86f0t6OWMNAya3xetTLujIbZXnXYaNjBiNko7mzLajkCms9rtC5NrCplrR6
CFZNT+4WuFjmtuLmq98Nz7Dg9g8kF+uxZ/XJBBTdnXg5XVY2s8hCcDBDiLuM3Pf7dmGHogpeDYaV
NQDCWEp8+xiZDGPHOCYQ0AEals8zWnhGMT4jEWFmh0YORATdrhBudTAPgkUztq+w3ETYqHv0oMo3
GaRc/7eWQxvL/YQMnfIDR1h/5OMWR6xepGaoaWAsA/FipvTd+lZnhOm+YjIZ7umhIY3PIAHfjJ6C
xo9tbxsSU+a72NlMU1Iicl38v4adkSrhtl3xtPMXLicPA9xBI3Grg37LISx/m9yegXEeLKkM2i1y
yYCTKoy4uAPPmKipoRh7q0Z6vfIfitYbiHwZlGoYWPw01XdMbqk7dNPKSLZwCq6BcCM+8m8AoV3j
wnfPeL6hq/22Tb7FWRYhKmFgaUk9bMpNP4arT2SXYkWH8xCIuQ3digJu6r3bOVoZ+1NN8yFm0jn2
SMkYvaTvmyGR12Tt7f2WoIH4Pacidze2+NV7sFZ5aMLzmAWeF6BQuUsE7zV0Z/noygcfcY6acO0O
lJU+MdALvev4AaBrRxkERMzLni5dV+IaRbl2WjQoOEt9j4zFVgNSb9+52IdrESu4gL41qFr7eY+5
AJhsyKcKeWoi6KUn0XKb23MTaEbTDG0Er5tlzCIZe0YzJGYXC+DXiwgOvscMV5QOllPROVrD5AVc
Vi0wgTLADnTbfzo49aOQMFFaG48tBXXBFI6FpMREytAJLuDoS7UnsFpmGwgz1g+OqDEjpo6+SJqB
T9yf5fF2W0qAHMRHGhdMrngVHJpAjc+Xwb7ZFh/xUxUrPD+vni0uLIPgYh0Ke7hDWhgW+62vtU/9
KS58c7YzsmIMHWKEWzK6si//fEIhBMpfaeVpXe9W7K34kA/Zjig2VAb/w25b9JRnoG1rf5iGy8O8
lzGUS1tNIhfgzddK9TDmHuhCL6tNfc3dWLkHxgs3O05SgPJAT7hNBG2OqnNIUUK25VVGKyNcNZdB
mLXtJFTMRzBoPOzwaY+BSlvIK5CYTSMfqNiM6sMOnWk+SA1ScZ3LhitI8O7h/M1Rg59rumN0g9p6
xJ7Y47z1xDVMEEsb5BByh2MRkWn86u3EvxDQgAjRRD7jvx0J1ZNes1pubtF7EkywDDOup1nZn+g2
JEUYIwE/yNn16Iu9FOk9bC4crWgFruQNCoxX9dHWCmAIAufqIZlyqmuAR6V2NCjEQttNzlQ1BSBt
Q1xd7e+DjnZ2ssNmHupdR6Nch11aFLNiQVRTsb0TNS65OELIW+9n7R+UDuOpZWH6OMPk/L9K2TGS
lCZI5OPZRhxJjVDq3ufWh5MeX5vdelYs6CzhGb3VL4nNGB/JiJ7AFgvZ4IR+U9d+sRns2baJjrRu
YgF/4eF3frriUHEw8ne4oJlWsgpY57JVrhDmKMPD3YtoroHrBpWihSgu96MiNFWwLza+0Uj8KwPH
ZJKVspm6R3QgiSdh8KRb6tMQQAestjPTxyaGVzUnqkbudMBFA86HvKgJfsXy5/KRfgH7D6Lz3Wbu
aJp2HSaVfJHxGa+VSk247fdJWsG4JhJD56XFnMG0BANPh0UJ2xjOG5pdTHVFXVH19rPB5lIG4Ihc
Udy7wNhnDIlms3Gm+D6Pw2rpYAfqEJ5u/trtQbTmtpUoE+naa2+Jcha8Ss/ZyLh6onvw6KniNP4b
HsIdFQ4QmuMnlP8FFF3UNyqXQjhpmIeSxhaGLtjbQhA2UPLgmZ4XKPA7hk/s9nkU/uvJo0u3n3uS
WSJhIF+cCmkBp6Gd0CgTtqBGiO7njgpOV35JJAOfBy+uRi+OTvM24vEDS47xVTewd9W7w+1Vt2nj
Ih+DKgopfgYeQ0MO1D7IKm71i2VU5VjvI3t7LjzGEccYp0XDlz/yo5bZnEKdve2MCDL1kLDFvZ2E
tcANKGHYOcSHe0t5Vw2PWYupivnWu7D1ozFHJPyQQZF+U7MEtzcLuwVhikM4FC+7bFdd/A+vrHiL
cxIyO6APUXT3X+4HhDC5SEXLDrl8C0DZsO0e+vaij1uLhaF/8xxNYTBnMMy/UzHWUOMf0GFQwk9q
JE3rugghFjQCr9KJJ7wegnvunAlIWnXr2/NP0Orb2q6OvZNXXWLoX/mbIOGiru5XwBuKjKoUf5Dh
nW65WrHvEpdh6WWmNIhWleo/2shjIBWUVRCHPjx2mz1KR0nMiHE5S4aLVMuC8rnO3Y4Hn7J8GcqB
G0hvkHGregf3Db2yYmO0y2/wmbTehvO1H2Gtz2ggbuntDX9K4oPBs1osB1+vAzg+Nasg5iClfi/h
fGpjxe6koSt3IPENQqUy3vGe+ElWW0UnTdr/yh84cZYZOTgfT9ObPUHWF90F/s0YFaYpf/1ydUXd
ThAW17eRHPRr6Id4ThLY2gXIgWc4x3I1rcu2E0uOM9hvpmqJwlkOYbx2+OtQktD5MEXpiqDm/YLJ
cqjOb9oBgAQXsNAiOq9YGD8cni7TBtZ9IgDpl2wChv9wwa2ppoB0xJO8XhjD3W1WQe197daazAWd
7mOagTW1c6CTv7kYA7FI+rmS1BD5pRdBu/dnGrmxskYnGiYwKsjq0TWp/C24Gkc8FoOufsX0FCNA
eGxLma4wTjuy5xRwdEJ8ro2IYt0sv6OUytOfbhoxsHAeB+HkNeohrSzm8WW3Tdqfz2I4iLjB17cR
K68ZZ8m7hrXdYvE5WGN9x0K1/kpA4LPB33sUbDqZkuq+4mEzhEHSMD3EVIZji9JFK6Un5zWuOMNp
gqkSfE9N2GihXbKtSQZw0km33yFpgxXTOJwCBVPjCfevYupL8UWuhXZUuF4JUjdIbLe1UnSNIlNp
HpjVVnnNkKkgi4c/1hpD+mAF8OCIu9++6s+ouiomMhGcPKHHESfuVe1KAvg2p5jeYLpqOWUjM3t8
X+ITiWrwqd5V+kKTgZeoLsOvc0oRt475sWWbO4nJDev6nHLLf5MpHGQUBPeRJ4aG+pgVKVYGMor+
YzIbsH89/3aN3sltDyZhkxnjAG43Hrek4jNb7yZADS7ZmGs9LHPUrGsyW5PomKc2mr6X+vQKYf5d
nVuTtbGjUaUjmgooNAMDFzodzqi+dNJ56vXQssBelJgN9nGznX802JtAKLdIgWxmQn+60xi5jNrj
+QIr5OX6KABhSHxtcth7zeNXVkZL6QwT++7cTXn4wqj+ttlx4O9mlEzTWfvaHZkC/E7sy3ZO8Vck
fbyg0uKIbzc8D8c3/0Exkn0YiwdI9kYbKkd628Yy8VYHFNoJ5/GgIqLweGpCcHBracoFp3uGbKXj
7ixS4nlRfac7V9WKjQt9UDz9HshK70m0eaVMtlJs0FNp1XN3lHg8WM1eQ0zmA5NfGOZL9//tg21W
soPwnVkaDHU7bBTsaB9y+O3fyM/eNujyCtxtYh4v3xqfqsWQedWbJIx+o7UyJINLeiezO/6IX3Jn
BfLrEre6sEEKTXx/uZGiSCc1yeSwAiEXR6EWqCKqPt59bHR8w9D+TaE3evbL4ntkC1DhFRaislPK
Ekf6H4YM+nasbr9oel+jrwY3WWr4NIaqxJ2gZQTOe6kXqtwBLYN/elLCerCs4762UH6H7piOu3bL
VIddI/EQloo7tv5PS24cOF+Y8cdgOOnMuhd66H119OA/SQfBqKDX7YwONgLllQvK04IhdVmrrUlz
Jlj1kyUqTH9Qh54tiUQz7a2aAQLzToVhHsPqhXxUELEfTg3CWUp1e7yDx2027WyO8YktpSZqjMcB
0nzvU+Hd0ocuW2nIqDyrTo1X8bm+3vc5N8fGrJHDNClIJOeSqfqHss+sBljnLH99YVoV7Z4WMMcx
wWpFxtbmkBcG5oTQAbRdqrHI+RoRSthRdYgXs+WeFPFqtiLRhCJiYectSl8OQhUkeZIHT28fvz/G
a30P7fLrK4NZqxXNATwe4a7KpOh+gK1iyXp/8gz3uAS9vaUAnVMtnWbb5PdK6X8xeTuYFD11FduS
hSDqNb/ArHLpJGYHinOzjyALf9+zKjmghUWIGLG4F692MXnUL/atZNz7PzWYzDs6vtTp6nk0ufHS
Ry4JGIMpo1c6Y1q3ey2cwc29c9UneBpxD6zPY196HK1LiFOHpOrwTclGpv5wJ9i92+0B2qPo4OTK
3JwzWl6MFpqXrAMOcVZh3+C46qs73LbSnBuRSyBmaL0few6vVRsWLuVByqWchxFW7sN2kVworMKq
+5KnPtRYfhhI+QEnIhX+9ekWdndZb8PhZwlWzJLEdesfToIMv/908Vsbg2pp2VLTeQboYlKzgMM1
7SKDPtXU9zDADtFPjbSzFjsOvBSdNsj8c1LOdovjiMl6Y2IKvYxWofLHJyE6DW1+IzqLuJDQG9yL
7kAElVO1BRavuCEV416Srg6NNjHDchmbDFsXPX71G9eKnX5bnbXbLeaJIrjAkJ2gV/jO4sCFu8+R
71k/OwcujYKJPXVcDxX3erQfaBe280Pnp2rDNWDyb87evL+/9t79qEQ7ymDbSYEes6zrvx2IWMPB
+txPgwKPTXbEeqY/UrX131eUhOmPTR+ECmVRDLZlR/G18LuAzWeTh5Lhzj2MKmMQNXdvtAxoVU9G
OX5mUEs46mZASD06mbY443xO+uwPpUAgUGXc2XP8FR2baOuDG6Y6MB4ayLHK16HKxx7GeljbzGlK
D3gzM1SYP9K2Eq0Gae1hAE/bL9qZSsLUqH1UfYcOUv7TJW4eGg+WmAjDHJo/JI3xLMrJ0W74w/b+
rHDtvvCNnYett0GqD931gZ+da0XCDKKZEQIzhTRAXHZGuHzqvYsMNhXOqay2DdwV7LWhKNB71O8V
vy4SOczoKXUEDozbppWGURBTg74CzYUqX9L+6FowY0d7BtpsJivlq/zQurDaLOXiqUZl+jlJXMPh
qMHNuB2aWtqD9aTTxIPDkZEELaLanWllVFkjrcncr9yvknTNj3YwcAHdO7ylu6hQuAf2NxyFC5mS
vwBoX7NjWZEDFICWqToSyqNCumAzk9OBJE3maP+XKi1RdLuk7h6wwKvOk8YixVPQLrlXpKbBEfkM
nj8hj//iUClCRbDFbrfb6dFiqZC4wFvANTT/6LbS4DXxXUI1zKaTu3sgcaIC7FB9CrBryo/8YPd+
msTA3Z7/fg7Qy5/XH7YMAI+cqvvoAYxTi6Nkfjpx5HKJDUR/e4akhDlgCcJNQmBfkgnyfd635XW/
89Na67GrFlZj1s5r05gPhWeKrh3YRjHR98IxK3v734uCwjHWBUnnx5e17J+xJWQcYuPDCoXp7tRs
MClduGFYR0youFLcqI/aeb/GmOy/OIpNr8rKq1j3gkdZgmHghGK/ny29iOWcAHSQO6Y3LfC+IQ1X
xMVwYWpZgl4Da+uqANm7SVd6KtPdUGLqOAmfo/E2SwqWpegyrIiZF6bwWgN2eDRswE3aetTwNJRO
4cd2HSbSaU1h1TYx2TmTyXF9RsHRUaYe/qt/HoaK5mnYO1zqCfm12TGrftFxjeLo668E3n6ESEJt
doD/leUQycegyg+Pht+1IoDXI+DXq3QUWdW7xY7JIPy9pVY3fDEJudrw+BXZ8+Hfj1omcu/89TVJ
f/eDDrzAWrRrD41TEn4FCGCTCFJj6x38aqPxDpUoHttaIxCdfb4p7jaosez8Sskx2jU/50A+9/cp
jryEo0AaYa1DizkQ7oJL5OSKoa9HFqs0NW2TRqQnY4P9BP9HwtVRks8J5nLIlnLAhiq2df0BI3G3
jqeSRIeep80HbgId5JhJt28SFWywO3svWlEAIxl0xU/RlxgL7tg4EAP7uO+N0U6LrB9JnOxJFEx5
CgFp2dd2I/0Nu2BZJ84Ra8W3+WDZd0DakaOns2FjVaRk1+O7anikZMBKXD5jKqQ8loWFPK7H01xN
lXOaqa3E/3ESqGi68a10rbRgc0Sehp5Pkw2wphqmH2MumHxUuv1PmeeizoXksVlTnddWSTM+tRzQ
E7PaHr9ZVr39FzS1e2y/Hq6UGcuXH2IujRqVCyU0IrD4g07dd7hi9C48FkZZT2479yxcv88yW1ej
Kh7gxF7rSqJdCd8pKBNBy38vDqBox9Z8/sh9doDSBMqyef5Mah5F02zrkCwfBsvKujFqIEryeXll
opsELeBVoMhnkVfvv/HkY5i8yMVCW6pL5D2d7tcR6245NUg6lQgjStP8uZQgKY3iht7hfkbF9mQa
+uKRuzoVPjK7ROaOrQWtgkjJ5DlUPGCqf7CGleycW5fcZaJJukiTBqMVWesWAYYhw2gSZ6JZy41+
gRqKxzjpvUe04gvTzH2zNqClYU69DePSX2Us5//ywSL+Gqe/l/aqgoctOmCjyfvOa1Icx15BA5g0
KDYcaQLb9UYOBfcE1SWeZtzegk4uW3bZMuw7HEp8dRengX/R1Qfx/xesORB3wvd+1niKO706rFPc
HafBtmre8X73s0udcgrRXJBHTX3QeFKjLKUxfy0YBFUskyuf94tXIrHX8iZk/VjoRQTjktu6HLG7
cfd63q4zaa8dT9+VkdP0zUJvMhvLIhznMcKJ0UaqueNjjRyNplkydZ1JRHr9AWlLwZUYYXvAhtqa
z7Orgw/WrHch/EkU3MWXlLjZizurjuo336ivlnnXcG6EG49NF1y2/Fh6d3GTBA1WW1QR9URN/XV6
D75GK9rxpTdNoIqSdvTEtUx1FB+xnQFunz7h0b0hYLZOICHSXezM4IqfNLSTo0wUlW7T3TBb1j6Y
aC1NFQ6y8Ey43n3gTmj94iQkBlOZhNM4PSn8yJgtURO5DlnZsxakYVaXy3iJ8AGxkxJxsvtql/H5
nYbvpFGFr1OW58UO4S9f0RcMw/R3HhKudW7GuNNXhiXcMCgmnFg5HJqDwTMJI03MTh51e/31TyQW
FuBSV9PXaBpLr/TQAOUomY986cc16hgJeb1FxBuiqwnyXw4U1ScC8ipN8rO3ihYboWUWYIAMAF51
e9Ivb29WNDy3Ba64wlgY2HoTTup4S+/17Lduzg2fXXFJgM9xPbn7fVr6EkZGiqkng1fjHXInGNAe
gPVrNj6hHib4Ly9Ef/0INJ7SByZvdett7zZ09VIPiREbwbjEL1OwEp+dQfbMlkEsiunEVaW3UgXt
49Hp6i79UKfUCcn/tTDTGXBjoQOTco1UQhXUVbAcimpveu2KFEMbNGQ29/nawXo16zv3WSopmoVI
h2FCNyfk6ArxW6cXrwPDPX3/GaR6GiCb/imLB6V4UcknH5NEPxu71Jgc9jRQWbkdWoCJgTNY29Nn
mL0gDzgjKaXPx41DegZPEAtLnPDyk+IPGoL0PCsyAvDmFFpA6CffbpfEwhHvbrZ2W8pRP3O9Ll6d
Obd/FatueLL4R3KJXh6Su++Uc2R19UTbkHmjcfBbIPgYG8yxLg8GDwnZqDedegpvG3ClYXMKc5PV
3wRdQNaFtStpukvZxZ8si2Hg17eD/F2HN/ou/kJJ8XUkjsHbS6VPYKOYytZ3sPT7zWhCMGuTMILT
sspNbYAVxwIbZCnRfjY2RmbPQJhuy5a0Y31IK6R1hk3bs2VKNa9eMMxy2sNTuv+IRRhxYIlvNxtk
4pCNqanhd/skqMLRF/f3H5MDzSwYu510vfsej8SdKqUoXlwWlZewlV62FDwhmbc0GFG+RfTxXPUN
+n2ObzIgnzpDs86DR/aeO8+VXSP/Vsw2qVRaAeukMOjtNX3kSqyp6g2jtLxD+JMnkR4K2jusju2J
NWM3/78pgkf8fS9ZXaOXEBSfVe8tl3vQ2nI4KzTTjnn7YnqrrfrhfBzWeXXorSFM+0nQ2jSPFJBn
2dWtFZ6XEHxgyo/bUCun/hszn9waGRJFrJM5zlnuYMymjN6pLimmuPE/HN9h9Tny8IuISRXtPf9K
ALJC+EO6xdQmXEmqZ57tthdJBHoTIH3EAC1xe7VDosIDaGsGLbp5nURhVQ9OOuUjBv+X58EGcuaH
L89GdSWaagYr/KuXrrU9mDV8lONGHB1vWSDiXComIMPwSTD2xSoi8Gq41E+71rHG38Yj/o9JsbEz
6GqHH+He7jkf3mgGE0XUHteYNqReRQF3y3iRtsHNifW29U2vnmQ2KAAUjgFChD6mP62IxW2Z1Xtm
/UrgdVSinGfHj1k8sfMhtWKcPQ5HNCqa2ITDUBa1GlSyKSvYqwnt7h+z31VJojkxWKpfTIPASPOk
1mGGKN4MtXcgIRSAoSPe5kPxE1/F4DmUKeuuw5ZOybZ9lI1DY9AreFjn8ecppg2NyHOu1cahUbwB
5pcYudFtZDzFxSEMYqhBfmbYDz1nXySCFSXGfBf6+ljKlJJG1q17zVHLZtZglW7ZcNPVlvYk55km
ghnYnrzjChwRi9WdDDMuuBq00VH8tPnxSOBkSBSc3Zrj/OJFJR55TBNMWVARbhL/fsi7Yf02/0NA
V6SUxRkO4BKGpA/crl8G3avZELdFy6GD+aoZ7nc9ZHn0ygIzrgZauLvV+UHmzGYT/VkgsXtrh9lM
S3DLc38P2xgiAfiNhFqRCZpgCkC4ebW+EM6JpB9EtJbLohKpD8Q4ENXEEKfEFaW3SU7fiP+w02+j
gBu4yJtyGFnQ8BslfeYIOWK3MrspUeLRTZfRO7ZnvsnY47IWSqCnmKbulmeiLMDQ2yW6WrndhMHy
MwZaGU0ATMILgHJvLuClJPHIF94IJ9EwOBu8ACa4rATREYFRqNPFS+fl79XSNa8HUiJ50lhNRqtH
II1tHzL/tBndz1hvhXTqMvhh+rxyo0FFYNVGGhtaXMCaTioN/YlHOnRN/dprk8BistB/U0JKc1jG
Gqqu9mLjX5gEBH0qTe6ckAyuKW7XbrBpiDFDtYkWDjSuJWBXYs70EYTWe9deGEcLqv1A9se9lCCH
dNtXccvStqsyAAc6I1pKv0Hd4IpEJ/q4sNZBtv2dNj1ajta+N9sVJ4dVrtHUVU5OcoKEhE0hEZZq
EHKqjV3P4NOfN+08MpozoIQ4c5gMVeWGxj2b/LYqQ60KuEau+j9KF+Yf7jR1BifTufbsYLgfjVmx
WD2cpgyZ4q/AxKnPbYMbTZlgtwERZ1zEjnYQQUc4iAM3q70ZJXvcDIvrAH3+bhuyj/NSVf6AxB4P
tNIpBhsGd6ofLo1E35QOKLOBWB1kjw0Lk668Q3Mmd8P52TEf7H8wgJ+APh6U9Se8f1/Vs4p+nNTS
t6bE99ViRMVKddU9AymImky5grMG8ztFbVurgLJcyfMam7hPKHKVPqi8O2hS2bnwDO4fGFVFWzqW
jGkM5f4Ucx7efA/uD8trdo2Z3iB1sDiCf76l3SX58Mu0CPQHUw+osBUA8e1gguZZtan6IRsv6hP+
QYMKmvJhm19x7PGjeFA90ZELHkz+M+c6MkNkqE3TaXlP4JtVp0SfuPmbBTK1oPy0Xcim9VO/xYt1
3fUyBiJeR7n8LSOhI3GblX6nQwZwwJD5jd/U/4cEy7qSTVllFGYCvyYejcgrrgm4cLfP2X0wjGqz
IxuWSG2LJQAz8TDKXFB0srpCh+4ySAY2Oci47mA3Rc6t+1UyAzVFf6JuPaZydHhj8bs96VvsKnY0
tRNeyT77QACf4PpR87mTtkhK0pzKB3DjKB2CcH47CRCQdISbABvSMppf3UABJuafx/WX8g2Bm9PV
5Gieitaxgw+pqY7x9ViXxTxEnIzYU3Y2F0hF/5CK+ywRr3w891B2ONgl0ww5ZMg6IYJjRLY4gpX+
S+SJ5YRE9tY/BPG8KTMf1wRTi3cblGnBYjE9dv7hFemR9+Db7rswLVd49gZkgsT2RQ6oBQ0YiKtD
cFky6YDSiAlWxfHUy08i4q3/9n6FMoc9p75lR4guMURsaBq2LQ5DapzF0I2v0hzWmuTH53PDOsoN
U+Lb8jinWHx8WwQ4Sj40/0sv9oZM/+0xVXs5JyF9NiBVRzNNBja+haI/5HYaDkxbrhy4hbtBpry1
7VdhkiOp14XR3UmOebGzEzZVf36qiUBrfxno3V0ZU1QC7V6/tWxE6UBxWA164sJUkJpGgr1bp40b
MygSLqXHqosbI8BKFk4d3q74MXhe4HoTD7MfJPKzuc4l73BRrLx0Dol+np8sr5w3PvWKYAvQzyGc
0T3pGQr9+tysFo23Rbk9G6SkaFeDVNpwiWunSTOU5zoWbPMyIqWELM0ajQlo1xuNrcyZHxiNqFHd
g6vNtpwppP1iXxqrdfzUjcKefCYHcwfYio1Gh3ITE6/gSv+AAdfxwHPFOkY1cEk8jdInTLjTtYMf
7gFMRuiznOcZ9iwf13oyukpkjUiKWAt8EtUnkc7iQGc8M/fhgWe2qIPGaGJkiPsywvLyWzjEZ7Q/
ovcWB4C2L/tu8WKcfkILU04HHu5pFbRjVV4npbHKuS+BRUhD0hjU+Lbe0mEViLLIcCGskJTFvV8P
l0I/IgXEbYemrLiZqJkPJP8izJPX3ncQchC77BywScLWOGUFINQZ6lwh/FIknmpOVOXYFTz6/D4m
Bw00mhDhHg5KodSORhYTAOJo4bci26Sg/mLAJuxIrV9MmnPZwojgZ6YBRRF5hTMWleWuMjkFRc+a
VyAoga3Ty2IZ8fRXeCGnyaUO4NE/wiSyRQlx3G/Fu9MHqmRBc6srrJdVpgWB79LIPTV/HQYX/CBB
InqiH5A6Ja0u7aj/fEND7/Vn2jdKr+5McpOzvUQ0r85gSOtmEM7/7knF4Wb3iqcm20fX2SOZHfwz
Ww270OhbA8shhILsAlTwea9uqMwEEHaWnO2xiE0Llbs8/s8PFIib5bLDPC+ldTknmJn/rmEXvVKf
f376/oCSD/U/rFyKQUvRb1i0nz+n86EaB0NkSq/S7hR0lnpdrGNHQ5ezY4Ws33Id3HhHLGJr8GVU
Ar/i6i+L5lYIfG8t9dx/03HGzf9OBeJBaWlreZUIWc7DdcdRLH3I51rBUCEO/jfVhuRdX7ev23+C
kLspNhxBaguxedqzp2umxFi9RmEAmxFPK0jr0vv93FGNzLkhIMoYNgzZtYrT8NcbDO4VpVhwn+cB
aunp4veXnxfHxMIeChkqychB9QKCEW62W26QMDimYEz4sM8rY0EOKxlztHIOxXk0frLBHw2LlRlt
Nsl5tZTT+ebLm7faKJnPkKcefy4vwKJE0Ry0NE+fTo8Bq6/v4cFYrmxhU5E5QnV3QZCRQnp1Uao6
3yUYOLMXK6XmXkaIDuOmB4fure2s77i5Nh2bZJj0EDo4ty3LCb1oDhxhnFZ/M3wzzDUgz3p0ed/k
7jMWPony6TymtXmclaPesZUX04sO8oNVfImt1z0TC5tuDxuclL2J9bkE1YX123UJhL3oe5OJ/XNf
xa0DeGnNTtbzubcyu/vlihFukvuXyznaWCc6vAa1ib2LMPPW42vgmCFR1EF3de/8b9omy2CIXzXa
L8wRp6eKM7fBNEqsigw88EQBhrNsqkc6Edu41rb0MEUMFbEvDWgFsphTxLK2V3/KAnS2dAACXizH
wH74njGFucisBP8z/I4JNTPcPYWW0FSvgnsfdz6c1QAuizW3JtOGSl6DJmj2wFO7F4Yo7XM4axcb
YA+oOW0JCknj9ZKLG2qAGoeCLXe6uqcZHUTxwqm6v0cHdLN6VYrHAMWn2gJt3uTYwr0Yj1K2NLSG
RmU7HIbhdgLdUrPJGWoIVtq0G6bJ9GXcVkFArbMqla8S/0gZzeA95XOJiwQIrStJbny7vLX8ngel
4NDJs9O5JA4ijDtROLtfWbvYHltaFP8r1FDnzXQL4U+1t9IQ2R7FSsI3lj8xXtcymSoWzOPCmv2R
hT3cGVLsCg71SL9ysRlI5CWW4iA8/tlZO/whOIQq2ZGR66adj1Y1E5nlxVjux2yRg5zBBW7OTG83
pLytN/wsy1iLkPnOFIuXK0KqPgRg1dH0TCbjmXAYuCbWprxKUiPit6B1RVRiVnYosCRjgjvCPzU2
BV77iYcjz9V9nSVXRaQ/4ujOi8JGunsjpPOpbaiTTTKHKy0+CHDlmTXpLeDy3VfY1s59gF7KNjuz
XAA7hhB5kZwQnAl8lhxduXDTDPNsp89z9peSFtHyQRzdvWKM/CzILXp92RmM9xVb0E2X88CcgEM1
n7btKQeAMFFdy4d293rXGC3FxYwTEtur9BJwZqd5PKnogzGR5uukSWhmk9zEzMPAe2/6CY6aqgj7
wlde+hwPvIWpiy9QVeoHw4IRq5r3H80rtQRagARxPdPSK6LyJTdLh/EclTLPc5Az3yPNDW8gt0q5
JnXrEEuw2QwxTJ0j2jF5qxeX1x5orAwlbFCvNfB92g49oSG1iczpzvX/C8pmIA1SlnhTaTejhQI4
etgedrtSIu9MFkdvOfsJ7l3iBQ2bXorm9kZIMf13bpS5CNuo5cOfO8BfPBXEVSOyBiCpj06zkIFU
qrDB9IEP0IE0DnkhG8CGMC7//XsCyClUdt76M5bLSpu+IEYJ/XEgcmjOgRSVZOeTq0WjGATn64ee
HxB/KUOrVRmbbRiWS2q0CfgNBgXGp40hjLgKo/W6JF/7wNrnLXfbz0ZfmoavGa0GKzjJ5x41SMrI
rw60b+t3xvSMRC+0IFrrAXpczJHxwS/kSdMvl+RnWxmtIdesMzV/eQ2lPkgs5m6eaxgB8CsW4bC5
s1CBbUT7emxJdPM1WrowdQJrGKgdY+pePsuQ6QgC8VWaKw3BgWyofD2JiEoaq7285I+/wcaN7i0p
zC666JhwgFE8boxf8GQ0zGLqaSE55+NirroerQffDEdbn6H3cjKvOBNzCz8fx7oAWG9PpfPy+saS
j9aGegvh0EdcPktFS9nwaBHyiuG/UzxpQrEvGEjT8d0UwtbyacnKJ10Eak35oT8dawpUig3PWiGw
zfswz052DMjs2Qdg7tVZ6eNct1DS6U2hHiLc5hpCdlgWWBWA0bX8xL+k3vUcTfgEdGP4WNdcKmCc
JW6FKTFNHzf18U+RdezvuLXChOCLt8v2OQnNDLLdb3Qj4ok7nSMbTDilXmdKMrACEhNqZ0nfJh17
GKiHh5Ym+lShxjpKMXf/otDBBA4aKKb1Six1n8LEzHB0ric1DcYdpg3ZqzEevknYYMDZp/TKrdKf
XpLAUF0yCg5xYriWaamveiuIBMSOYN5snxjg348OFTUO5wunNhRyTW6TVc2ql84gd+TwfzudOQUz
lfTQ501T5/BXBd2TWnpoReC1Xg3gZ6Pk9gea9Hd/NrP67vGG4/If4j+qnMlaOoravxtPabshFxCk
rBNzPfVGbMGDIvHUywabUQjjxMpfubR/Yb8zIuG7725g7pDTNSrZD0A52o3jEI4Wnur/RXGpcPBj
0Yv0Ledm6ZS58ty+BZ348rYJEFjSxYNV8JDC1XKdVPAMnryxpsoX6beQfhUu/wZq9rxPmIuEORrp
zMHVrDMGfrYcITm2e6Li1p9u4l8l2gDpnT7jWejK4sIbidJ+RaTbEQBTXzkeqQc6Cxz1stcoww02
txudut8JcNXiQz7+Jo++RMcKFuAMRZhkE0nHD70+SolhZu3pkOg/pD5BBxvzCJ0Q/7/CkSvGG4Iy
ai3loyJC+74oxmOLel3Ze8EynGvfqftYWeMTfx5A+Hxun3El+880ILwuyNmRp5zrty6mJLWOUcgf
rBv7A3E8ewFLrKCErWCytzz0IzImyEvRKikMkVIq6gq9+okwCpnODE4I0r/AmcNbwNfkXmtgkWZz
nQXP20bpZVYxBouU/OsdA5uupxHrk9EkbLogNPAFUx/wjWVLlRtzw58lAMcXthKLbGu0AHPiCmxI
9cvoNdWeIBP2Vo93g5+8iLZJjSMjgm5z+6NNtP9bHyYKDuomjBRf45cA1zySRzgNVzrTeNs3F3+0
w3ctbrp9YZ2s7Ve64fT+8IBaNPrlRtxPA2Jyt8zL85PHLMlqe6L0TKJZhKnD6nqJKO8Ux9Pi918E
wbQ11ni/bvI4y39MpVQoZXtWOjW7sCEhJE3tHDP+CgPZf6ryl1ZzdQkS90/aFbJMHfIPlbVrF8DO
peCzby2ZNNAdL0P/CihVNz+lpnWkKWrzQ83Xw/l9ViuzTTlaTYtFuWaSm1MG80gSe1m4IzynnNx7
w6Itqp/Q34pNIfYsR13GI6V4vd7LtouVFohaw3kaSPdMK9ReW0hwj/425cwRYMe7RrPi6z5JCSo5
oMPL3Lhkcw3ssM7sAGNUFio+AJJNdAMdJBrLwDN+bte18udBQI6JzoVXFBkBTtIANEZCDJ2HViaY
DyVjMrvcNiK4VxkD90I3cbXZGBHtKGJz6dWecthebabDHlA9YN+QI31pImrjOr8D6lg+jE9IVrax
Li1SLK1yy6Yv6ItiXhLzmNfNw45Pcv/md05yNbirdcvRbK85G8cQ9aJrjeDf3PLCdc7qLp3PtYT+
0MobzMixL9L3Fi1sbIGa7EfahFZYsR6W0+QW1hvR9VN5PGyzADBd48kiIAAtwR2NELjQXj5Ze5pv
+uJgc5t+cPdLqp1D/kOOoc7kxUdQJsVYe9zbz/ZyjZnUcab8EqWC3EotQCeCOWMVBMACGExI9UGw
XNY7QZC/SqSePydHEyxiTPMsDKekW+tATquab4BatgaPk/oLHmT7m4M6rRQfIeYNALdSmUmbyL4Q
9oPeenlVBRvDrEpxqqGgG/UbaNPHZAxu8my37Oo6JJwciqSHE/M7ITnRQwWOrZwIuautDZKX2LZP
B3g0n2TmILXXZhGHBqGH93N3wKybdvhh4/3fDQ82CyGxhB2rUtjki8ipsm9jL5h1z/hS0KXdkMUt
Y97dmvz3/iefyRz20DR3BlWPq8LpPaBuQUtNwhpbbRQHR4jwTG1jHz1waXGyU6WRzCesfixH1LfD
RDGFmFdutkndaQxSzJOcdaeYeh/jIhQtqIzsOm4mGPsbm//j/qvGNk7/2Bgf8bM3di28x7D91/IY
x8qIRgU3udDhOv8bycahmtGranfI+Cj2Pwy3XkP17pD2AKUZklb7FzsATavooU1tguk6pvtA9kzt
qRUMI6ZZ8noM+mbqgWJ05bTxIvytSXfEBiUnXpQsLaR+bbPuwvGSXm+m9peN/MZW9Zf3trqTCqe6
rqtki74E7e+lGnXWxuDG5hi4NFXTfZEPeB9YXrKEU/9dYS1CesyPtKME1Sz4OYMUxfo+hBB63GzT
51Q9HXmDIf/8SKmISXyo+Qt1S3Abb+9nJUA4MMWde7HJSpRjKNChFS4r1NNsSM+Bo6E++kPV4nrG
FrazuXyqcE1z8IjS+Ms8ExW4bpVl7lKiKuVroefCLlcfA/ZZrk9ke/aUiJGrKx8cnczad45CZWwq
/SzxHzMo40gqJ8BX6YPiSeknS3/ZEukJRV3+YvLcEnvYcXOSgA8kS5wx4f++KRx0amt/cdXooX8d
TtT5GXM8lse0sUmI5DSqnOHDMIQ/AoveGLAqORTO52YfYcVnJozqx6aKNQ7s+0qDVlIexxyTrO8I
n3sjoVppYhqfEWY1iWB+74aH7RTO5tYncXXaGkQBVvzmaqKr3QOwGJkrd+Tv6LR1fDSsbDOkk70Q
SEbSFFFiMW7Ml3+3yKCkg56KElD2cTFfZEyfcaaiLLHsFPbDVkzG/dzJC76ih17+uHP7+7HmG6un
Z5QkKIb0NeIP3AkQBM3Ab36uEQkIdRIW0Pv09rHKZR1ZxKxOQdhXFep4inJaOVKo1awSgMGAb2pZ
oxjGU2zv17BieuxUQn9pvbvEp0BCegq0sMU1uLLZH0a/3C+CzHe1UlEeuQ9HPm9ci9dVSK8QbwVm
DlcGPFGqFWGiXXvr9qjfP9V2nkhHXps0Swn0pDdTPyzY0kDb4qBFsxOxP1Cdzzt5Ix+iRnImUCWz
NQuOh+JoDQI+2nUZZ+9lVkK9oSth6F3eTuarfiol1vzWeCesjBMRuLJJaEC4xC3TwaX7lXbg6Jp5
rdNk00NILylO5PRPr4LhRrBY5v6okzkz0eVyE3XgpyASE8wQ2QQreNUvJSjte8W+h6xWLGbTOmfF
mlCn7F/9sbwHIkZr2I2DnyGQzFW/r6xK+ADeB+GQTX9maouOEvvj4H8Jq8Wc94WqVTEF8ap03JwR
VPTzStX2VMXCzfn+McfmX2Jl3Rpfz/05xHeJVLfJesh6emUTnSYYECsZ+54w5PTFXwm5RX2GE/Kr
kheUqZguelpM6u//jKhbltudn7/ceUkpojXLRbDpt8HHfIMGWHPDWhOtxezaBFw/pdG/wYyh2tAP
vFwHWZ6LTBHD0jhYe6LlhOi3SjbC0E4UxNfZ0ugWSZyIiBJv25++FCdY0dTsvAUTTN+cRW2gqgZ4
R7ng25/uAzdoI1Ia565JixdirWFwZXIfp2LubvABZQ7OZba5U8IZwWB/kd0ONrpvT3BL+wLnXPhZ
4FcgfeySnmh8pBH75L/Onkw4BmyJAbGC6NZjShdUmDPl5pZRRykxrS467tsjEGZ+GdNoigegKnSU
NhAC1aG2CH9Kaj5ggloAv0ENUhRKaAGTG8smDNk2qJTl9xH1fMn0Ng0Z1iC995IbZbBwrMMQy64b
/y0kuS6fydPx3PAxf3lZuHe1PgAbk685bzBpMyDOyLR3hvnuxsW2drzMMRZEfaXdo0fqx7cOYjXY
EKUwY4fjxJA2vkppcaLyTWKdozxy7eQ5G9eizUNvufeE6kmgDRMguA41E2VOSHmb/K/Mv1JRi/Iz
ELbpvpSQhjsjnmw7JgE7YyBMPxC4EVEbHiyjE2qDRwVXew0iSLM34nudsvNdGK7T36XFwGW3J9WD
ySfXquLQonkgFTN+OK45Rx0HzAWwsvV4IRCDhZCCHxceQ9APWfhB+fd9Ycm8tu+XgkfPh6YpaCK6
HO/lykSPpsPMHLHPlRctF19Wt9C+vlCH7/E4YBt9w42O5vAwksrMiggdwpiSqQGMQ21wEV8l7Irs
/G8hxusFIGpvi3SqaT86E3U9bc8pwSkBus958/Y2ubSfyVwfvQkgBr4SiaIN2d+yBRdkZhz0E0v3
tsxOvxSfioXHW+R5Ag3EvQMmRM+W23kmR39K8O3m2A+Hbm2/XpsWFDBkfpZYSz8w1M+fm1WxHdRT
ZvuDD69mmCXyzbpv22miKu72vQ8Oc//eI2xF2IVQATvKotRtq6mcDjl/s+t2A+W8pu14WLHaVeHg
1HskbFrux4NRLWSMpUVPYJELI7VLwbtwrYWF5wP/LaMWX8KpIXhtWFyrUxiMCwd4YCkM6s0+YQN0
PfluTaqqLDbCwJUklSY4Ywq0QSw9eb7qQ0GpaZ0IqPkrk7DmbiCWQvcaavr8dQimI+7fQsSJLCsD
vrg7G4HXjxSdd/y4F/8dtwiTSa3kTjjTDK8ZBSNZ2k3kNGOC+2yqh+ZnlNlHilmQPevA84V1pDi7
+QvfSozFqULWu1t1JFekIFoSnCwwpVkA1K96u86D3oSJm7m3H7F+GTnIIrlrFyyR3//fWP7ES209
4mmluwH7tRkzhUSB3/RIO0mz2ZVoDhhspI2l5FFK6F2ypkvv8rOpnh1WuAAscdrvO37lijUECfQB
hUmApl3XVs9GBFcX7kZJZNYGrEMfAcuMtAy2s+gwTeDx6loDAbxfMF2ktwg67jQIKJBggQPr9X6I
EV9RhdUy1iry4TEe4WTs3FMe/hZzAX1dk0i0BR/yGy9A/oYuPwzCF8NDxoqFCOr5BmwcljUiCWQa
funnP/naPwHjsQvGwoshz1OBxGzkEFiadnQ3eqjBtXngnuWOVNjkrUc8rJVi7EQqqIVvT0lluGEf
TXBTbxZ3T40I4C0QeiuRmbh6R3sK+EdzIDz0AF0meDJYjp1E+ytYAymmuDelGx5yFZwveho3Ene0
jBuZZ798/W6sSL74HHc3i2D0SBCDtwmmCjorXRbRJSWyH28l9LPNXLIpjSczad8RD48xubEI1c9T
z0JhaFPnwlzN4cHOOZUiICcJMsXAFKR4EUKf6LbkLsw6SEEPNy2bAPB5q+MfhEmJSsYG0RvEbgcz
EkOr1tifa3TLhB4DahG8YNTdk0yFrPyhN4pczDWuP6mnpDGIGfAssHhx7oIy4ZNAR6XN6Ty+JbwL
XL40hNZZBhmBOZ9GofMvgZ9jtCLbT6n6oXazM7ze+VV6YeN4sVCGS+eoI+8tPLhhf9ZPi/6WbFj9
6Q5KjRNLw10z9i46gb874y80PoB30RljuIvq2zjntJLT4ICBksU2qPcIzzKPHdpMeQQmNT72wh8K
S+kB9KKarKJGwOMxIswE2b5Tz9VPPXgoOmqEAvPOaSgKMrA7gMj+SF8mm5zUd0YcXZAtVgaIvpnG
Uo9bHFzaPP/2o+u60z+OZYr22rWXMjUvnrJO5Jpin9m7girXuhBWfU38B5vSKa/RTzWTwkoshK5y
HD80UF2sjCheRAGjcn+OI5UHvwFFh/amZXf/SdAXanuWz0sDBVapmBcQvrPADPCDdkmqaCNswEqE
vq1A8Vn3P4kvndPuGHp7lgJNnjRvh29hLBQryzz5I1b0PM/9x1chSbX63ROQHFNI3j+fYBIdi5yG
gT4KmUV8Q62nvZotKYuWxxbm7J7ESQxBVpAsP2cfTmnHg5oCNWHbH4qfOHL2sIIq7n4WDUBd0619
PLaq8hDOL8xJxF1LLVcx3oappD+ERmwetOivtBJFFDCahAiOyZ5i4KPq6W8PVoEbBNsRvgzYAmCt
V3793i6ym2lOTqnK6+/rVqH9ffYUoxBjarTzKc80k8pURcTdGwmL7n/sjQsYmW9YIKaWn/8DRReA
O3xCj8g/ttJez6WzLi5CHcJlIEEDd1DMFhqBmOkK+ql8y6z4q8+w5F9WqdRIg/daI8rzlGF259Oq
/u7N/4VADSn1u4eo5HRF+fQ0yVSWQlWwzyYiCEg1KdxSilTI4eFMjGUgvx52TC7oUygqLrHxXojc
fkyYZ/2Z/qMwj2VMg97dPUkwbxSLacm5AUtxzqVv4USaeUS2mHDuONvMSHaebA3ucUD8ojqpke+l
Uozgx8esfQX/CJYc7IWkP79TDDSm/ymWMjQxeD+wuq6MNXgsyUB9iYALgDo61xxlXy2RRm/keWqa
B39xlH3H3q526loWF3DLw1rLOQ9pmEkNI1YVhNXCGJc3tpg6hqBKiuzuX+NgBevS2L+sj23l08H+
qBkH/qczLAPmDJY+lXISPiCWIDlc/QHIrHJr6+awX1SgodTq4HaV4zlySiF2UxVWkm+CyQq/Uo1H
OOjafFNwWdNh17WveJurCK15qRjOZv80KFdhQTvr1/V6ixUDJZ4jQZqv/5S7QQLS0fCdduk5yhrP
f4ncpOeggRRIJOuN6kPwQABYtDvO34Q0eQsJlQUp6+lZxwx03rfqYbdDNjaPDFC2Z0Z8cU7qW93x
fu2WEucuZBKPRD6+Sm/V4ofrhMhLk4dFsu3cojl1GGc2tKiCqkE1BjeLlVCxXSA8rsHMXemhzZaN
lcIgas4TW/ewlO995+AS635pMZcCsqza3LsdMW5F2l8XeWoLVGAawCzN+o1Sl/vj4JXOC54t5V2C
uGKw4jPvFndsGYjmPF21fA2nG3pvcZls1Kgp2dzeNQAiBzPJyIsaKKmZYHn+c7J/OneHZdIkn8kj
z6qTkxMBRfYjFkdZKf2HhZ+Rc7OoxErKbLza9IsAtO23NSMROgP/z9Ss4t4GswccuTqOU5oWN9MU
UrwCWCm6qQbcBmzq0C3AD1k/uzsOX9GKJa0CbbGIezFxuVNURc2jidR3FbwIbGPaoH+oSxoK2gSR
/HeqdbSHse1l4UuBcHYUP1zNwlDLf/DFkH10EC8igXZstnOcUZTWCk0BoYzIzbgglhnBxL5+wbci
t0KoG6jduRMt8BMFIppllG0RkSnb35d6XnSVQ/1Ost8eFOCQTgLgYHWiiNt6cNda9n6yKIncWJlV
E9INEacA60jwgHFos9TDhEpXdPkPheUORfUYadjN93n2903JPM2TSTQoxw6y2ZhxFYMAJl1Oacmj
aNo4CZUkYd7NwL5PkLderCvJ9bExPnXR1fekrK4vZhewoRLwBj2+JCqwWXBK1oOa/6tenMi3EI1b
V48Y9BFu1WQmVOUtTsLxAbCmmWEHgUmaTtYOFfLq25FbwbUEyH4ghFueDUW4R/oQxcpJr0uSw1Eu
8LGkeOLBRJU8cfoCf2ECVBlaWFalm5dGzIFSmKW4mR6r5cwSAELUs2f37FSurIBa282YNGTSk+UA
K996TAzKi5JO41RkRxkHtzYzyEPBg5Q11TeRC/fowDmOaBaZPaJIxWkjeOBKlKBaTv11GUZWsBD9
Wrp2FA8zHjoHFPTfKwVKKwkO3PcAIMa4DyNx68TS6iwImwSSxBLtmlikCCNhMQ0mdE2U7ToaLsik
KNO4D9iP4nYh+QSThvIcdeaLcbwexDMzoVjx0szO//Ohwm3GbgEw2kl+bJQjSwXqvCztmDyZEgTm
XXAQhuNtH7j8dkViJxOvPgDqutVyL98qEbY0/omM0+u+j0aB5iXmIc9NKxUv6SNOF824088ULiVi
02vz+9gTgVhHYOg6HryYhlsMk8TmcnutNod0zdJdvsViunj9mGDEkt6GvyAk8ZvnnqaUeH0HJV1x
Xxtc5OqLzXs+xBbI9mlwuI0IXb9jMGDlPmfnPRT9owUqU4V3ciM7az0whKcKfscS1jB9hIMaYiFk
a+wdVvVh819SRwiaJAsOLEjcSllOYuAQ5bxvsD/hJ67+a8XJNcvnGD1eLJlqACuhJZXIU5oC9AL0
UROTGnh3yBPLyqdiNDZl/kKrOYwu9KViBqgIwmQlFboAgk22KNGr81EMKUlyN3aA+5f8k1Lnh7Gb
959D8DXEq+mZquPk+4xfoEBiC3VLs0KTUlcMcxsgYf4lg2STCR5i6YbJ11OBCrkciEUuCsY8Sbcn
Wk7lInBMZOmeypYwN0IKP181tS8Ow8Q+K3VAGfi8XLI/sFCYWa9U7FC0Rux/sw62D+SGn1tbIMHo
jqLTIi3BgdnUS5eygSBg1innBp4tsqS3tHrYcIyPgsH2V4ChMjH47pirsJloLKusLeO837/aY8fK
thkKdJHSJ8omcPrh1eXhTLq61oCLrWxDm89ayxXf1cJ2N80cWCg1U27ZPESqhod0XR+fZZDYxgBy
hk7OWrMag40T/rmVxtyMf6DwSTwbGBjCGznyeqzR3bcYM4iiDm/S0gkgJz7k2bpAQbdz6Sdt9uQs
fb6LHLuGQ4osCXrCnW4+B6SkmsSSlCT7zfb1FPyCoOXcMw9yULn1cSOmUaPdMu/1YMSgD0ADCre8
P+siMq6KzDMRwaVPaLEofVKZgUvHR4CG37pSutMCC0rTvYdp54RVHetEHAnxvtWJ742eCSB+pzWU
BizlXJRE5It2aaTOtjxeV0vpusZJaKWxVlTv5/h5qKBIHRoNa4a2uHpCbSIwNH66utx7oiOoIuPb
tepcnOjihG6KSAC1OUZYqjlvhEU4vBgnxeU2VvztqNNawfWq8Nn2RMbCa1vx0QjWo3EDHaohcRjf
7TlGxdg0jsg/66cbOaAAj2yg9m2jvAgNzE7UI3VPE1hk2+HO1HYNQFxVbRZjBAaCNbN5JbbMPYYz
oEsUWN54eZrjFtQnQfp0fZgLk9GZH42c1ytI9wldlA0VGwmyVZTVD7Ouseo5xZ7oGg9bXr7gsqwP
qx9AIDsKFBPSpSDypfB3Gm//asHi/bpvHOJX2rL3VbGjNtTt4TmZ2P76AWx8ggLJVB0oRrgWxU4O
eIC3xJkay29Nz3kWBGLWDSmwqiDVeoVFa78sgPlemhYYVNcThEoxL3fmng+SztY/pIkYFk7PJbzc
4WC3+9shlwF756B5s1B2HMzXtcdYKknq+yaSiuBpMBLgvqJCgPHXT4p+swlb2M5Kpig6YZixnxyv
G5F73ggGTcwZU1nfRh6ohcjk5MieFhUc53C3zXtcTUnvCgtC6LrkFpDAydBqLlopcmF0AEAl+d+i
FpjT57ifsQxxKEiFEVoDoQ5DMWq28aG9U9GtQh9CjMMPfXywA9o0FlWsqUzwRwpwPKcaHg/2OOua
GY2d4n8RBzCIg9dtrv2Hn0MsrMA554cA4Kdp+K2W19xN1uQw0mvUmH0gSIhEUMuQpkWISrwpqAlo
WVvU+iwbLUbKKv+jhzYYUgLptO78FjCTZIhrsFghBaEdnAs+WVOcEry0gz+hxbESsErPzomyC0IP
TjQ9vq3+0R7rh+RMfqe/la0o7YeP5shuztpjskD0yOdEgHBc4Lo1YCZbYm1ahxE2mRC0viXWkCbO
pLp1+Kyz/V3aoIfJee5yculy+T/2j6+DAUndTxmFdMCrPQZwrbDFQtzhz5o9oYdnHHbmEJQt30xV
C/urBZrj65r+Ddxmsttx78CrKCdMXF9wpEYN4BMDh4fwQpQdMVlKX2xQ2BAORfdcKgThnPaDrPjb
UpckkkOeBL5eyiYCB/es5UC2KeiQ3eHOWQpwvvDEGMgqPtZHIZ7CYlrAQip19rwgM4YDMdre4tGn
7Pb2YJNp1wl+n1+d/jtJHfpI7WItVzlEgdhx+FXwqMXDF9pKbQh+eczUnYzIGJrTq6cfzyKioySA
E9ZYCnUhDqz6Cdd66DwpqMIZwbBue0cn5IuP9x+hBUmw/4+kQw28R4MADpfOMXnqMBfYFpYY9UXO
1dNEiiZjwFyzkCR5Vq4gIt2K5xxEnrTdamhyB2oofIJJfr8YsNwoLpxuXFPUNHDQUgOFROz1Lr8G
Tj7y9cD2SqrOSbk1hSHnzq5/TdTe8s4nvxGxfb1cRu8w1403sMdDKHfLp1Inu1sE+zrD6NAO1pL6
pzCxUTx8G5Q53pqb14Er38rvGWaaxWh15MEsNWyUanuMIy5u2psNNKfCKETd4l/Gkz+emBzRDNWc
binC9KCa4OnY/w2S4Zmi9IdK6/lJqEQg0qlg6k8LrmWt7Z4tDwrRDzS3HAN4ni3gnOya6Zn3eULM
i+URBxkqCurXvg8iFO4r/JVy57drBJWWsLzvH8/UbxurYqWsYHAoCWhiC2zpz8jP0RYmBtlQw+r+
fuuo8asQCXaqBoM8bS1f0EkHQVbUqlo3fGMrTiCe6s9X51fKJvrhq/ypqdykDqxgTd/zyQKjt0O1
cXwzUGXeaozaP3AtXsC4gZJHJUqFTB1QzNqVe3kJN2sSrk95ibQUTyCu72NpfU5kGIBvcABWBJI8
itrZUV9ylctafBBnUH3eq6YGjD4D0yGVTZuxiL0MvJuVoB9++Paa0Dk2qhKTvrsGt743vbNfkCEW
itqMRqSptDUCg5aO//WaYJn3/v/s1g1Z5FwHdAnB1QUKxpMm5gTQXAA02NxxNogNIx552AeRgtXa
+k4w3TB3+/hto0TkOnPkVoSDbidskZMdlz8qPBQlciJWxjk3qqzzifIqBu0VNmxG8fiHRVrVeJaO
nXd6t/WL/hkX0AjWzh+0C5OHMkO4DcQGbu5+vs274YdkNEjWmpq57v8GApuLXYDQQ9bndAUuFVqU
nSgslBzPeOfp8IQnkQm95iVdr35txkDguMMXc5N4UE6H/MQe+gNsmiitCUqv7g2OltzHbUFlRtZg
A70CsF23HWYpmTzW7QBDc57z/2HIOZhO3xmEp/Y4LfQeKebuHq1Q3xlDJAdXKSSG0uoK7CpOXidu
7BZmCONyrNzHzc5pHI5elziQOUnZD+HTkCbLgtRotbgtzm6o4/NGREY+8NCbMh4ewryqxL7SEBdD
bw2kOIWOqF1p3p7yqKZOMdLnKASItdX2kXPdr1R67J/s25LFoNmDL9Mof3+MZOjUnLPOI2NHL5EO
O7o+OSC1UWbfvPICCO/YH6P+j2lphK0MgKJQM0qGiPfefMjyxXcOYW2XRl/iHiWAyh1Rfm+9E+lB
98QhXTnk7ZmOIRG0EMek4e2hYQegYrl+8y88plIDH/wFI6J1MolCfZjBqir2nrHhH5/Mz0LXYUrI
e9iD7ToIhaeZw3oeolScVFDo5u2GuIIte2gpVeXUdlF+Y5tAInX1aq6agzL9LOiP8+ZRIV70OnHZ
RJ+/Ib3ALUQEQzfPbA3XVGWuSLExaFsb0OCs0IRV4TaEl+g/85XBDjykxngaOl/9Sun9XhFQ0RWc
3bK7VTKoesr0jcMtZlQJ3/RqfdUIDikLn8I3nKoiT3b0OrrfFcs+ie7NP18XdOzT+XdTpS8nrsgo
rACbPXHYQxSCqjB9Psa1vmMF5g8mQzLfr7fhesGpMkfqP5ilN/UFFolwPW8bnSWU8vrGlQKeCt9X
Xb83yAyqxWe5aLXr6pUfGebnKvHf0pPeiLLSlBomupLRX6ZnxIWd3g8ql27+UpymSmMxmHte1Kej
pi+lv9jdTepZWMwK1zZXBR5vXcOvmXzoZXZlT7ab/xDr/maUmgDBWSWrTcuz2oCygLLIYWcdHmKl
g6TCNv1kHIHPUQLpifdMlfaKVqSFg1b/RTRLdnzv9IaAiTRoM8qwlpfGEMxwrCNRzpKYySPFiOTr
oQv3pJv8tdLM8L5IkZvgHpUoLsB18IBwgrUv6nii83Q+7na/iz9MZY7KkhH8KSdIJFrT2JS+jE9r
jRNfAvjrMtFskbM6DDfHB+fKFe1Wkjst336RS+jBGiBaNGTnGUKF8JC24LdvJaZJqGpWynG3Tle5
AlST44K28X3pnVzo5Rj/Ycwy4wBkw6p3WDRLbNfNy3Bae6NKpeIaCRQVpt5vSWhrAK+nEYendIxN
zjFODPKzNbkHscf0pDlymVJGK36lsrYySuqQbmBdIXFoR5qK0BMA9rjbnTbCywe5QHhCU6J0XV0s
nHQcBQ1gPKUZCOnZbge+kIsDaHeWogCWWItGN9h0DzXkUuOXThGiPQXHhMRQyZV4ytinvbiBZGFF
IakPrHDPrP6/f+ZWuFn6od/5bY5p91CnnWigHUVZ/zQ5tpOUG+2d/Uj8UQwhKqss84Ew91IXpsbn
w1WsN9ocGzt6THCD+fcrpu2HO1qhXFtpWCxx0/SQZoq9lP+7zfunGdIe/PKNtbEi7Vpr+gsb+jy+
xJDVdeQuxux+SC3fw2U8kQE1JVc3xLgRrBWBRDuj3Cqx/dN2spmCY8aPQZvZHbaMfTGPH4FLMpcG
ZVs1kp0piiw335EtFCLpievw5MUYFez+L/pQTv5xv9VuGGqeuUcmX0YSG9rEUBzD6T2PYMqqyNVq
6ayaHA30af5hkZWP6zjeeW7vsuh0xcGVATQFGZT4d9RfiFRXDztPGP4Ujy98TXWrL4Fxp1qLt7Be
E2Azp2z9lJnmjXrc+758QOM89Hy9UY/GMxqCxRGx2TysanzD71MSgng3mrEqPUbM//NM7SqiMMow
nu35o/HOOpw+CCicQzbxBl0TY/vFp8d9t66nrM3g+diMVk6e17YvH/PRE4fJcuhS25g04vOYRL5A
BGUkM6PZQFUXLfMjJcDwnqrAkZPWMD7Lx31miyYhAginx4XM3jsnzRMoZQLin534xuTKZvxX3C0U
WIXUEXOfvKT/BfCNLROSsrioOKTOPVAdbC8YEIQxCvRYRqwha4CQmunYTfWNryScKErF4P1xSB61
47EODDnveGDQMyFJ0fT0lCsIopMEF3od3PUCNjWe1cA70tMM+AWuQNN/1akPELPWMv7mxeToTGsh
Uu4+oz/eDS7OKL5U2368l6HbUmr2iz9wxUIyyCWUI54dRebOxFjH7uCkQViC7lW3rSqJ5tAfvpRG
876ZHLcU5Ecj3bFeD+wKvVrTnqxJ7E/JGyxlPKQUIUxQbgBQm5478UHYFBwKCx0KmJLwu7/DpSor
Octc1EG6vZ0hAyEKsp4DaGqkp0AnViiV2NqR5netwBWzdm4e/SBy/gqlGW+mRAmv4R3hFbrWwJTW
uho2sjZjmSVugro1oScM/nbInxNWbwJbYdG/Jm92Ur2d7/y5IDif00+U/9FPSLYNUz/Iq/EnnLOX
qpQyTGnTHMQ8E1rYRcplX5uSpbm9Q8Iq2I+QmKutnLyNkqdAL5Qi4l41+0Gnc7iuW45Oh4694P0U
ZzaJ0PWm650SWtxJpLOrtb18VN7Ho2dr/au8diBTWws9d3IQoHKYVGq8KYq3aRzdcC1rCaL+LQWj
5fmUQBz86sLMWO26JkpRr+0+UEzwt7rPRy/e6TzSUiL6i/9vivSgKISrKIgEdBykYtOGzLPcltnN
/yoRf9KovmwsOvLkIRS+srVOuCenz8xBnU3ua8znFtVENAuBbhgHpRtNlDb5Kw3FlG/t3YOENEgs
C2mfiHqPHNbfHfYOeS/FNLxPpa73P8HczwrCaj1Lk5rBJiqljO6v9L2n9KfQWfAHCdBF75suM8P+
noFEWvuzYcExKUTbGyD/YctHVELMO7omNEaoPz8oDNiP21v7XcLiZ0T4c0zaXvNmzfFnzwYy8H3v
wgDNAfsUtV6ICkt/h+0osbYe3Q0Ty0ntiirV3AbZHHyor6mxkLPK0y2ZdCCH4HKYnizF283oHjZ3
X/peYysAR6NfR28G9qyz6rdz85rG3u216ztPlcpIgRQJD3lgDqGm5RlxIQ0s/XqB5O0IMxjuc9ef
nCIkaSRVI1fTlDbEWcj2mYDkKVMgSCoZzU/s0I+DAovxn0j1PqZDhOZUXK/gB2wEAuOAiqJbwyyk
HLRvyopSIVSCSbDvBrGAT/WJCjCBBnk1uVE/flr43KPShUoBlofAkSDsE5S3tunfQmGTOXELpjJc
twqRAsKOMCd/uiPzqOKc6U4uqS8RE55iEo8CcTdP4HTPTdtXR0vrxoh3syYYj7ocBJHP8HHKrgvm
KeOxJfzmYFKJ6upVBD4DsZv1dYuNippylPWAB87xga06UEZojxmGLPlB7SfmRxp/9dK9qAKNwUXb
oknfXHlIN2YRaBTBSfqVjn5xPVDhKKEbM8uZ5ClnHSugbLdRIgR8xM6/DXtvZOR3+a0a23sZ5d3Z
srTxRJftDA42R+5UC21FFEJFKlHTpFqmT1iGSA3/2hiJ9tmlz9M7Y5MaBhcVm7cda5Tu654bTsZI
0IFE2BK3V9S9oLmHUeXWaPOnwiEfeNnVMLQhia4rJ5MnJnsmd8YI+C75CCSrCK3k/5oh2EYdQ8H2
n8ix010iHOmXZUTCOsgLfuoUiwpmTCnAmlLk2FHw62iKJKxk62wxBvq9jK3udJRttqHcVYBtgh9d
4kVMId2AWS5KOW6lqNfHAWp4fiTbk3tWbdtxciOxMrDQRMvx06DR5ZxsmELzTD+VAGKPp7gnG0UE
3XHiL3bBLQLDH1yyoUtkmoL1m3YN0KXUYWgl27GcrxpVxgwcmpW1BttA9Z8qGgQkjal0jV8Bs+Br
Cc2y0tbEKsLyvKp9a2rZ7DOj1CQi6g/ybR5SyYhib0M9FPzPHKU+YUr+hfWeV79lUUlzulp7+cIW
/ow5oZW3IRHWUql7n/xWG0O4NKDtmx+BkrAfNMj1I8v2f57stawsd7k9Oey7muyUMz5BMmxXg1BU
+0Wwdd3+/6nqSS0XR9jw4C7vDZPvgSARrgEqIg7mdLW5WIQi1HW1PAfkutTAyEv28baD/zS0s7cS
xZYJIF2z1fFCnibQ7VDyi2pD7vJnbKlCjOeKFxJ8/4R4hxdYR0bnqPWZgRjlG2FCfYHTG8r6f9Tx
mU+yLSwnBwHBrS7IF9RNrTtQYlxjsms8pDHLVLsJ55VtTgl57xu8MFaKgOKWvb7GWv8xBiFveb8l
t7ObvOAESpTLeHH9GlwxfAsM4VaEerThb95n0ObKGZ+4tdeJPXGMuhBHUkxgQiim5ctahH8tH2xW
ZbjNtVk6SdaOZcwmLJ7ByroM0pVCn4IeRfby6mKqrk5OsBvjwkrem4fg1h2MZ+dHEugIv9cPSqqO
9Z0c5DkseGz8fL5hvcn+/6wVVlkFGqYNjRWc5mdjqamsDH0uz5oOHzaiP+7MwxWNg4FmMa0V/Oon
g45yaZjdznmIY01c+Za1kTwciwIXhpEjJjrDdi/V7iu7YSExEC/F4H1YK9HF9Os2jqd4fSHWclH6
TNdJq35KBouukw7Hm/Jj9jz/FgFScOgArDxlRsuUS/nsvQni+Wy5/MI/u5VGRQxUOwmIvI7tSr4E
FiPg6FfXDaDzdlt4MdMc14hG8cy32ojR1u0E4ypan005WNMulATqFzoBi0PRo5foC8+AL6I2Un/S
r52Vv6vxe8iNduNbwBffPooGF5TAi9uh2zcdwtqElR4rae2PvsqEKQ7SZHmOWBJ/eoqoHFUuAB8A
ES7UH50h9JYvOVGZCQpn9M2ygJ/d2mepq2VJ09uvtwRmdD8R1QGGIQi3nr+aQfdjDfuhEasy8mGW
cMI2EaDTqaHrGzw4if78URs0CNhrwsjbn0AHMtUyNRU++9Q0OforaAl+Tkn5PXsm+/sQSkftW9Qk
kgGQXihyPDVqjk4GmEdKCILQBub1P1p6KMx6XNC8sl9hPbvatmWjNnXenABMbdLzT7DAWWkv4eLA
CLq9ELpHCNXjbuQSb/L5wFaa+QxW5fffCNdlbuYwmSi7XZhaYWzJoLWB39T59qQ0qxSG/8Wv4n1a
w6oIzn4oHSkEVpaHcDEthFz1F8/L9UGg4VhyXnj7shIQo8PUGmSfFnzsMziefkcogicoTFOaugXU
ekh0ssTfzQfqIQQiXyNY9oRiTMKquhz8l08FcaCiyGnn2zHUbsokb8Q6GchtWWXrPzJIc8/mpGnv
5aH3SAa06LecivJWLl62CiN74qXnK4V1zeEy8An1wgxWQFAAksR7+620SH2JF8zwAZKKtzJxMTai
POvDsoyQEZOCQibjH7RJGhrfMm01Hhmb3SjNw2uZbNf6FAJdlDdPZU/Yi61UacjX9NMV0AjlNBAX
pO756dqF7upXQIS1bOPLPtAbAsryA4FTaCur3F63UiI0zerpBoYXCmyKODp6xPYcP9tQvnrRoN2/
rK/tyFG1HmOkzt90oBlnrwpeJpgTcRo0JPqTww0Pwje1rfwr5RYDc6irfSFZrIB2knmhcd83JFO5
+iv4ILHVCRtqqxkf+/5/DhLiPFT+4qKm2YYmfFH9ZOPlRK/Z+87pggrSd6oZfC+qRRIgoe3lMiiM
IrTRCeHNJ9fZLDV/jK7f1MzlOrkYX+PY3kj0SrC0BUobi2valsZjeGeA6oUpbG6ZA0uQf7OC+txm
9kmhyrrPcIBaMDHHccTdcdcu15tWX2+fXc+RvHdVU5eWlMxCul9Wyo3SDaYTcFKDuO5GCDinVZpB
KDDU5b+QA2y3V0fmIxXZuJoEKC0Vk/KqFhj6zKc4ZFo/1CMaz1fw/evebELwaRXoz7cmDkPzdCer
AS/+9Ao1Es9JGRxjLg9nmbO3/z3G4Fg4gtgiV7LdbQpFYPiC3lFV0Xf+pb2h1ZXDO0QNtaYkNvk+
ZuLY4T1jKJg83EPPR5OoM+K7PfNSJdblO9a3q5DBeuWb8KSwVW4C4kS0fIBWthrEaWy1dsKn/A5B
chipAAMA4QNUH1X0elRUdoCMASKAl8A0c7VmqdsWoSnk3VDEEHjjMDV+Ixg67bkfQ6EWVgLmKt5s
EuSZrS7k16oQZjxsiinjqpMTDDnASdfWOcHBxZrOzf1P7lPQg5XHODwqrECxHZWWTaibcY1CWOgr
j0e/s4DFc2wsNFdczm3jDrD9Uq3eOtcLqoUuuhZVENR0GfbA0oVn4+trw1Ts2C93wUI0xf2mRUxM
lLz4kxoHWW2t7tq0msKpT1z1g7wjpvvdWnApSXS4rB7RYRtnFsT6xQZCwThXMQAXO/vFYIj+Z6gv
H7A0jNJeKdhBqadEU7Y6wkJtcd1c3RJh5EoRJr4IFSnFRhotidLvUODjpeq109BVc8ku+XlVd8rf
OGlCq2eSSsDbE8UJQx18422Rq0ELNqcqFJdn9DiQmC3YK+XDjoATDEfs6oM47OlVXDharRZHaOlh
A6xTAeDjNCdQ5ZxjKSiqvGUJ3yJUGeq2la9iE9Xmb16zV3YHHsOHYzTupCDkRnCXPQ4gd6o4KcbE
xaqbNUHEbAI9Q0jCpnwrPPrGcZOFoM8yCu++Boiu1QGy4R/DU6YGRX3Cp4KMNKQ/ODH17zZsL0mA
o9GrVJGjMtfMYDdtMUuv9gt/2fMRu8Cq4REPGgb+5MeZ1fhjD9sO6yqS/GvmZQjT2wk1daq6hnI+
3kZIV4P1SBsCj3S+JsYEFUnuw6oo353fUy5W8BJcKSE3Zs9qtiJL3ISZ8yRkbEktbzIuE96huErc
T83Ogou7Z/N1nfp/mzysiWGxOBIl3++GEj7cNtn7/E9KY1hDV5CPV82YqctK+8sRFE3/NrJgnEA7
YE9+A9UIlIG7rh4evljl5VdrPurprL/Gja54Pf64YDqHMpQIHlWmh86RYhCCh5IRnkoGUDiMDDzC
oZ4m3yh/0AGMRiK1VhBER8IjIqQd0hgVOvkVdrLWowZ0Ne9AWl7JMvc/yPtAXqw7jrt/ehIv/CdP
obuSTu3JmHVupCPPZoYKCTP6Ga1ZrrCMTmvzwt8GmHGaGI4HW6KtgT2rHa2YIVwPRTSJxpacdvH6
xFRMWyKdRDQM+pq1c+p611BXVn88d39LK1Ol9HBPWjeH1Kj4ARVlpjk7dMze/MY/JMC9OHvF8hlj
93Mh/05sGwFnJqL53g9UI+DO57nemjkATCIbMuZn4q6jCFgYwm9f8UTeim1271I3ONDsjmna9hFV
cFpH7V9Oa0tn+8/e5OXZbGFKf7gMhTHAVXgRE9aaKqpeadBzW/UlOg42HIWKK76RnrvAvVHF0Iss
yxkvfK3QUAKlf/2NuoohbDRXQ8cbDpJJXJu+qoZuYxCPIJg2iG0LDT3TVi1EizlGHw89oQPZ8ahp
W4FGezmjqunIxf2vVtupPaarsyncASBQnM7zKkiYiWF89y5xuNFIgw8H++QT4Vvz2/GypTtB1fmB
HFaYmbiMyfmkWrIcs/K5E1xl51CkTJQMB3TEdPTT3u8HkSC/DQCtIxlzlA+uPirKwH6YV9SajXvX
2y1+mQ9s950vcAwu/ftM+wTvkA6clkwh9jnhXU2iVM+KIACK9aVupRw4mMMOepfJjjMjCdjNEuE6
5asfHijdEQj5FUpauI/3eo6TKZF3EXXKYHQPpv1QizDKkTCRE9NUHqtGyGMV89HV13H2W9v1/pB4
3O9fQSyaPLGaNGCo1yKNm2Y78e9f5e3y+tKdCakcFGVh5wF87Jefxlk+xGPjOy7YIYC945dFQUAz
XQe5LpwZXZ+Co3hHy4qZDJ9OYiSblw1fCAUqsqmlvKyp0IqP7VrIo6ridvQYIJJGophOrUtklU13
zDHN2vKZU5XMlrrMHxuVN5v6/45DvLUA0mJ0J9b2E+TAHjil/8NyiTBhacAcuANhI4TMUI5xgsg3
ePGO7AjHf4uMkGqhQoppW1G+9obHD0PqOyCI5XcfelzpmMvohYwUY4DWx44HgwRVb1mi801HLX56
GiL9saJj8+3rAEqQO3l2q5CHDHwkCDR8i8oKeR/miHLJCaJk5rzSwp9RMzgvTS59ElAbKLxWcuO+
oEH3HkuoIk7SF1mS45CerY/sol7GDn/MOecZ5Z2HfAALfDSJx/r2jqvENYa4jSvA/eesQ9skDNM0
OKeNZzUA7NOuEcEK8XH5D729grP7dFRW5+hzDg45CUB2NfCuTyql8Ax2S6D19kq8vRPo4j3MafCf
G0sJTwjhHFCBn97rG9Zag3uyFpDIjrGbfYRnNaIUZuFzUnLu7S5RuQDAuzHLKdepRJznkmbD+uAr
OYHxASwIvL1ED1SjhwUVAEw97Qfd1HqtBrLUg9QaGZnM/RUw+jksM3WPNamSNUiCrmUVOQI+iNVs
RQbFpn8qcDEcXZdrJnAq3sT7S85w9sWO0YppAFxur4hggAVPliDsqJVy+cJIeI4yT1ZYuwXk1RVb
fhNFIvwJcIaAqFcOT9rItsvlYDG/HG3JvqqBC9/NT2R8fV0Lsa4bC13tVF+R8XjlmGxlp+hh5ToN
FJFwR3Ezo0IOyDTaE7xE/ZmcQI+Z+q+9pa+8RWK/HHUjkdC3RLWQzkVAldhl5YgaFFs5QZ5lta4o
g8LrirxhousjsQkkYx1sgDJTealBO/i+zAMJX35Qe6ZrZm1Jhkyif/ySjBSvZZQjbJDcJY5xp8hx
gFSa8KZ1m+3fQrbZNf12vuXi5I9QyeVtAmLuF+INTH5TaqPfDVELXWdI5bdXPo8kJmG9/GpWeAqh
fNXfFeYtbY+fEySwYgnLJDDJ1f/WfH4+Kz3pbvRrC3ikwaUEoFB2yV5X2Ii1jQLyyY7UtvvcLZ8d
eJaNHn5lWkmzoOOm6n40s5uyVnNaUUjrpDHEdwzAa9Y3NgIRSP8accT9RqYsUYE3QTeNHcUmM5YP
EoR86e/mrHArda7fTc8dogYmGUlo35qx7qrg8LAiiG2GNWOhw+ETwb2Ck4x4kEPgJZWtRyUQ/X60
p+K9tPbWZumLFTtJHx5uRvwhs4seMvSJQBTIOPEwx5JiEBcWVzHWmgf1xFhDCoZey4xhupwshynX
LBrvLwV4Bypl29BTZFuHjlpdOCJ2VU6PyhKA28qnGmQ5TRSDbkiGN20wUzpjCzePiKjMZhunfv0q
1/c8MpxTWKiChbVOcYFVDOSHXRKULz7kUV2jNWekLTJDbZIz5fHq3Y87vEqP4MbrKg34eehchpFW
SUb5VurbndAS0mefhVqYJQmhk5lIBxezJI2hHDDhKCOJr+fPJZOzx1dR4cKhxZEumndCCRhyF0DL
eh5aOunvaqvPVVAn18P17PCFoleNa0CX8GW7BqdIFJSRXD43Q7gZjNB0eqJXVoVjow0GsSs7kK11
LGEArHbrs+rnBJD+NvqTOzqIsp8Sdz7LY69iGvT26F3PedPsrG+HkLuSCnlDdtvhambdiXSDZv6Q
7TWknmQ7wjyy+XMS801JkSDxMFc8d2ZDcLr+vdmVLI+Y+L0oksB4Gqi4CrMhV5wKULbt5n7coc02
r2PH7hjA1GvJgbZr3PIH2Sks3NOYz5oQWhcLBKMqeYeKmJn07kX+DuMtNqiwlFPdDakZCvTmLBFd
dNNewKKjeRwd5NozfHz5ZlvZhavLHVM/kfGKlQfz/W9MpU6t2oITPqxY3pWMs/ILUcI8ZbkhmiXQ
sQA+pVJ8SndKJ0/EfXU/OsI3uHN+t/Wo2xMjmymctOhJkQcgG3emODgBMz51DqxCgXIBrbCTySQ1
fwUwgeIFFC7TiUwsw4htd90N4XVmuSCukLX9ceXzwHiLw3JxM9TlnUG8MIr0BHPYTAobw8otxgGz
0CKimh4Frt0Ambcz8EqDR2YliGc5MDCK7vhKxWMYXZChX4z+0yjXwcl7vQe/pxIvonYl7NnAk22a
PKILdGATNiO1FA6yY9lBWjKJzm1ZQtYe625B2HTeLdtl61xdsdxi13Yj4JLIKl3YmvWteL5tGvcm
P+YDWZjv6y6V5RnrbiKH3H7YeGnAU8Y0XyZZhKRjH8BtXuWY1CmmDFChlsLWPUgfmMNqE9oYckwe
HQpna6ZTkyHjN4zmIH3iQdWco6NrFCYwgKgrYiEuj2/iiB+t0J/7PsBQPIwvMWJKvA6EVn7WmqoC
0pq4JVyPSQR8QzGUCdNU/RSqYXuGXUPShXZvl/GYgz6wyV1T2XeWzWXzPIfJ+FXQAaTvw1j/rV89
IwtyZP/TgJtIxc33Mv+FFziWhwbLJgbTRKtdnx334Xq1mz7fdw/7UztSSyUnZTiJrlwfMgIzzKhh
riyc8VYs9Flua7KGyj0AiaHdESA3iv2vC94zcWQXzVwnsn32gaAuX4qMIqPJRTTLYRqxFE79kuXy
cmUeZzwMVTx9+t22CEK3/V/TOIt952VKs+7UrFu8ndOFnS8cTurc2gwYMVLrxUpRg8t8C33tcpug
rF/mP6dG51tg4bvmIALke/11qPO64oHhk9pXmOG/IVQn5WrUB1se6dmCqwdZUS/8XipCAeseytWH
FR1llYGnpPIgnn2nWnpdXAvshhhEcx6Zwp4y3U3zrbSAWmGzq4yoAHJ0EoFvwuEEJhJGHK2kVRQ2
1C++wFhd4Xq/wHOxEoeP9AAYOHGFe6V/hXE5VGixX4l9Q25fx+wdGlKRLSt8xS8VgITpkGjpKIQb
aw5vnM1SFdB1u5TvOo733ybXqrl9kyWG5Y9hv190xPmP7mUonVvxemwdFRB2klwPoTDBK48p8mjJ
Zrv5vQuVnkbshwgiU18mniY/fhOP3PsLVH39X8tBer5PGwB0SjamhJ4L+qp37OeiXOeRKPVinAXj
hAGtTMHuqCIKg2BKMN6TvJJS+/MDJQUsMmvCXAMvNH7U9XsOFMAszxUbMZIRRBumbABHb9XhkNQB
EPbOEa1q5TIrd0jfqnGkDbwRDRbGekHhIFxaqlnCDPip4uKtM9Q2X/fnpllQEBJHnEatdLygQRO9
VM8bLHBL2iYw7fPdTqsetdQeJnIzr3c6gEkM/djtoRB3/yXIBBhSNW/R7uIf4/6RLfQbzfXln9EP
wLdNBkRJgz+MFhEfES2ks2hnGhww3/0KiH//CKEERSxeU176Ow0RLKwRupSM9J5kyTTO1FAzV7lL
9n9kQO8/cieCiJopkNdIbLdsMZ8SHdWGhl23hEvg31sDJWLy5TpY0n9OofH4SOtPfuRueJWCo6Mo
BdRyrrImevk3llogTsXm59Qo/0jkCnOQMI/3pzkpDMlVqDnKEQnzsncculmvwHwmIjx/Vsx569ip
fp0YncdZyApQUwqgkYmH9Ev/PkO63EqT2GwhjRV5A7ApWn597+iq9GHuuXY4OnFJvrc0/BeEIpRH
H3sdAMW+bRXmHMNhFj/fkhH6oxLk6V51RBHf6IDUXfQjNGN/ldmGHVSV3BA0HkZlr6x2spdZqZKG
IWjFxl1kEE9iVRZIzW0sbGkG0lOA7qJy0PJNj/iYYr8tl/YFxEjoGtzxla9eOsgaSoMHdefpmYAF
S6r/4aHtd0As4iIklz830zksKYd7ts6ZuYXCSphH3IKKodaf7uHXtJVPnATsWyU3hu1sK0h0Vr8A
mH2iUO2RIUbnuA5xm4Iuvamzib5SSTsyDWpwqOvSHylbWdleyadO6S+dv9pEa+wG3IKJhuWUpYnA
zGFfrjrpb3ixK+RZlWPzL7XKGIMiMlp0oK/eL8JxdkzoKrFp51/UMgTEsMk+Ij4JAydX3nwKZc2b
8HkHxEiNmoOT8RkG6N43hUP0KgTAiMSxLcHwZsCdyj3pysj95QPproIeVBji8RyA+hhW8CA1Ac1n
efaAsX4qJenPYMAoL9rEgsusXh4NCHAEz70laUmfKLnmcOnOqSZGudKDnOD3QlKYGxl8aYKgpYSq
rKOaCBMe29xiKt7bOxsPTjcu262F3S90fmtwtFRZ6a3PYptn2g23Z+enWZojSU4fnp5v31vky7dn
LvMVSSVt/rkcCnFSHSHw/vDldzLJvCXjjMljC8t/g21B+DgYW3sTc48UkvNAQNtvSb4FSNHZOdRk
MtkFwV4gx5eZPpKwjs2+NvhIPUX8JqSrEfYquGQ+i70yBRfJsaa22ZiAqqre/FOH/HPxnyEVvrNB
Xa+XrP21TLzFyVmdljJtA7kX/fWOfGRxJ1yIVs+vHkPLe+6sKlCl765aHWu/hiN8S4DuJP/wtxbB
0o+dhTNdAsFin0PVcUIRHA30OqayV1TtTjxpRRB1yxlWMZFXjDU5orJKY2h2Q3NgWOe6rjjPreJ6
jpBCYlbgh9wnNK1feBSjQcjfYYJ41y2YJxYLJg0vo4RaYJTnHtbjQnl1Gs8YhooKbukh7JaysCvB
Hptp/ys7HuuDUZvr2f8TfytRzwA+bPXjeTgW5/nOhYA2F5i9gI1X9ecsqNGV+bUF8U4qmExWPN6g
xQHwVJm6nvcix4jMw4Nu4N3WQxl4VeeTsFV2OEXah2ge/ZnpHSzGW+dW8fCnEKA3l3+BfCMaf5S/
tQH7L2B0s9HkVaDdUIeIfKXNr693V/k8A5U8q9Q8UXAwx84Qb9P1xtzo/mMVcdRRUga+wkNutnYh
UfPwLeU8EWKVhKzUh6fX2E/XIA++EhuJvvKyFGv6PhBjo+1TyOOdAqeOIT/qd8XG+oHXSpmARDWY
ALgad7/lsLmSh/w8T5Hx1Ux1SJgtysu8wRKXMAPp1oVC701aVLSzdIq3MfFVQM685Lzvgy5UGcCn
7ZhWQOoKpwyqAQHtABX1gEV9RVUXrSCpP42FdbgnB4LONecydk1DTEj9GvA6ra33V6DVWiA+a7l4
zWSWf/v/x0bN9nDa6aq3rDL7w+49oc/Q8IU3zXQKKzbEGZBQWx3Hj2oJFzTSF0JLrLDgg9vO1Mke
cQw0ejJjRkOqarxID+QKwNeVG53dABCiESRYzrpZR8B4MyMKCVg2SARB15XEUTHFRGVlVk5jcrVI
Bivo0fyXoGPbzv9xjViX7FpQCcqzZNHqTwzVEuCDJtY4TQzjvGMcnGwromfyOfI7FDUJP9H23o3E
RJ/LUUAFvNe+Ub0zHJWiTWgWl1mOZBB9RuNmyuizvkrWwHA1uHUOziqb4UjUg+qPx6irUJ7zKHiu
TJE8c3ftnBL8bsukVbLCv3Qx48z5B/ZehwbA8w83hs+OSZtM+Cq3Ng9MYsJyDFSq8UL2vhJV8yGD
H3v5MfAGMBdMnBsQKnWeo7H9lPMS2Rm9OJaj5DgfSjYE3NjxTOBo8wr1zHUxrjzOp6tNwqgFwpoy
y7n1kksLS0+35ia/En6389u/POJCyd7LNQPJABREWZa0YgWwuhoMwxAcMYLhP9sVR2YhwRjxhXtk
LT7bsRCIhxW1LThbpcDGMxVWCUYgEROBwxAItdAGUyXww7NL5iLgvdxO0nSwwBAx93w3THZ11UZ9
QevKx2gLxipGB7AnOLAIO34HRsYshJiXqUFiTzHdGPbMbBkX1cLqFpVUV3X0bz0MyolfuG+4MuWq
amI2Gfhv6PRGHWXZgP+o7/gUHxlFAZFuhe1nrS8zQCqffWPzz9sZ63DpKfwJPsHkzaUKGIh6z2y8
S36qVrGypSEgjGzMsMzScRyCf5E+3LTY6nrOBWX/s7nlL0xuFHmWxQxzfJ2H2RHKuhJiV1MGLdNc
tlizPm8TKYUYN8vwD98mOgNWto62tgCRTcaemJ4incZntDbQjLblF0EbMPQuN8Kyjt9SIzzCbnoZ
l+hcp/+yweeLBU1iHPYD/Jy8CGDY/W+uursbTdf8n4UPUT7uO1zU7QIbKPS0Gm3vad6S9yQf7fkz
1+S/8NRls/WHqeQtTCCzylruOnN0TH2YrLcbnHRdiczJJcuMnzwkpzCCMIptLx9t2ugmdasph6aX
eV2W2eJlFLMawXBA2CfOXhiH8kaQ14X1f18GlEQlH3E9+Qop7VRdbeIX5OUEF9/yGL74kI547UIa
1dF+Ja8W2In+viLq6i6iZlqPrHeu6saBpHFlfl0GWM7d3q+8s5E/yjtX/UhEx8zsdP2SqUMyvcbk
t0DT9dkGLX4hgkr9AT5ZJTjr3Hqqsk8+Wtz0/to4ObaAYxcex86SCaFwavWsHtQIj6Nnhgic5maT
g0SRdj47B7VCTghobPaDhHyj2JsG+QjX4pcwH9v7NE4go8YFeS0Jc9YDPdalhDs6/dcx7tKSRN2p
RuTUr3BJt/brkvrViwPsnPKAmd2OMG3av3PXXUxhv1zXliuAlciL+H0kZOHN8Vi76VePaTJ+AtoG
/u5yzcGaIxhQK4O8zVp0hZ07mMfGjZbTP12mKK5lVm32PQ1m7S5AgeQqIzLLCLxrhcG3J7s9aWbQ
XDyZ36dR2IafiHhBYJgTesNBbIPtza1BTEHE9j9RR71v/8k0Op2tvKKQPlksim47CWJ3xRPv3bw8
srELvsMTctCocHmhw79+BnfI3zqRwTOTKRMiyKWjjHwMaIwVr6bxHOFI8KcTCMFXuX4W1+QcGiHb
7a+UzF+fxv+MuePWcz64/W1Qr9kZbP41gwUD8WuHVegN+TyoCT0CmUDU79mlXGO8Anf2LpjUOspJ
0Je86EBQGYlvN7AiC4heMXOfUKL9tZaPuTyWvdaGy7lfLKTFXl04O3sK7qSDn3zIsLXB4sjdzMw3
Lp6qHLIZcukKRSaGDZRx1tg5Y+OmROgpJG2Jp/28ZjfhvYrl1mt7uQXcbSLsolR4c0j5j66VnPkR
FujP5lHgnRDDeZMDB1cvhvv/rc9+wul0acTWeAC+woTu4eXwLfJFNwhunaGMQwT+mIbz8+yOxvf1
VzhjY3V1Ei3c0MCmZKbyQp6QK3JvXH5+In49Gnh76NWTALlYy+7QIJNi6dzgzWkUmEakKnOAnCMb
B4rlp7Uqzvqo386Ok4jlZ79ZC4c4IAKi+/WACEQyXNFcjVBKiwTaXT/8iyfOvSABRBnwpmBwPN+f
8EFi2NI8JCS2Y+O4GDb2BuKzdFLAc8mb1kVY8Yi74yudsbghtwWTipZ1P4oF1XVEZy0xvDSU1jT5
rFz4lcUFoI1+6gkPIt72gSuNHzBvvrL74n58HCnTV4czoxUmWk33yKvhx5XUYlqW1lbVuKb5PBVg
I16Kt4uvXVf/swucjaCaACAPz6ZTm6HBZ9N/ryDIULT+q2tqX02R86jw1smlZ4AjDELg5cJw8nOp
Do8i4bZSWwsT3J5XQ2swkD6uozqV3m160CSQh1oXC/BqkzM6fJKqs6ioNNO33pH1VYVqdgVhub92
XR/Yda7+riDVvppyMS1k0jmD0dIowrZk+/B5h6k4ATEfHBvHDcAqJ1AISeuaaMF+IgZq7UlH3A/R
hVKxMDn0uGlsJXPlLIEHLGk0iW9h7UQ0g3Sr3zi/RdcvAg9z1iPHlUq4hsansOJEQZjrnd0SoPyn
8Xz1LNy3Qs407SvTrVg6UZsPA2wGnAhvq7Bw9uWqPFTWyuqqA6XsYowIt7PV7ycPoFUAsn29zTbZ
gRlGbUhCkwS92Wpq4oby8UyTOfseX3zAB5Rprt8eq/R3KGH7T0XKQdBnFALRBqdEZoRc3GhVDbAs
oG5z5JlhHv6OIRJ1lI9knPkLo77SZQO4DEITKwiYBXmw1PcL/b/Z/NOWf7RPIs2FaRdn+jeOh7I5
lt3z7Ak1Ajz22ZGTzuAMMVNpNeTWWI1guto8NVc8TZZ8EKIHszUBxxAXiIyhr7nSjRtUilczFdDw
rZjhSVvgRiUibIuoCeSyNnXJmSN2BQCaV063IisXFtXQSm8ywfYqHGqCCyAK/fZW9+tce63nrVnW
KBWeShgV/7hpeA3T0m3nDtT+7cImVzKmse+i97riHN+D+mHEmHrauawkWFoTBNkFO4Jh2E+Mr636
durtYeG8X3zzqWanp6mQFmN+9AwRUCtZ16FPwyOCNVazxS0vWdZBY+NCBRmcaxlqFfYMGSglJTus
WW5s2hc2y2GMBRxnKJjFnPpl8ScagHBrN3E/RheTB4SI0dx2t9GW94lqKrRY6tyRaI1EBGJt1gU0
ZcPXeVYv/PCy1o1N1zzsXRhi+/Fpi0oLC/lLHVdy2Z8Iri97MvrEBHZhmezsNeXIjRtcGEou4l03
rBG5CKQ1ahNC0SJI070wdtorm6IWODCdxEd9MLRA5XFU94H0BPbl6obhc0vnSsMpfN7PiF7aesKV
3tRXvIffYBe9KjjsAjGrn3po45+EKvCRgKPa78EubnAQy5zHxGJbWYMkO36fwYEqb+g+OuAb+gQS
jUx+9mu39IQA/efFivOEy7AGEbFLA1+Y3wryQZSO+tBemetw40zpr1nhN8Kg52dZgk9q9OSws2GW
lSUx+JCaw9KayVqZuonO003QqLXKRb2NmIOGwVBu9b+PHknP0RUwgPjy+AVyNyOZ++6kykBYDYYY
Qr0QB14HokloPBWEzgECI8oMks/z0kGaPO6eMDzFGHtv0abMVh6OUepVPmCmF4uRay4aGojFjxwg
+nc8aK260ulq33TpOZnvamNPP5sf7FKEWH9Vi9iOEPRBm1RhXWxs9HRJtOBAWbG/9KTVIjzHrtFT
0vWUmwmdrGnvH3sS4hnjfExVudu9wjOmaN4QkiDGMwcP9ykXhcvvOBWb5GsD2XuGddcnwdPDBvUS
drCDh0PpAAF9HcS2iZVW2fCxCwy0wpjl3oiZ5XO5Oase/YslqHbd6lnWawJBy14/X4mkbqOVBWKA
AMxWWe4X3rz/nF0q/KuV2GPa5BuwyXOsYFH3jpd2gZ/Aufx+bQ86GFI4BSeFw0hMBqtLY18ZAMPV
jRxV6q3/0dxOAKwFle37iD8BPnwg2W10udFC2m7mPxMnLALMnHnYPqQX1KSh3Ao8PNlKSDn5ySHV
setpI/D5bIop+GHqA0FEw4/gkBUMgj8847H+DoBCGpHBcfuCd9Hq1JdDO3xCkRh1ECnBMnneZJ2b
Zo/3RLBggkNllE8pfZ5+mAi68hqe6pD2VuAQOiKKImv04WYUiw+UvBWXywJsTotgOwpYZq+DeqBw
RvcdYliY6mNCW9B3s5VyAAi/DG8xlgMF7UzwmzJx/ExXJxFA8k5bqqA2HXG5VcDoUUUEoSESE+yb
M31Eo6kfF46gj6a4lkCTqFjBd5WGtwOnumqX2OSO9URzZRW44Sx8x/aNxtZ2EECnLTwzWqb+/ge2
vBdFXCJN5dIp8OQ+ernU9zYa+UW0GKmFvGNzwTgeuUkjrqLf5pDzBqz61ZHP+MfEgrOmecYZNN5f
KHITipawI+WV5kYF8LZTBZ+HQOxbYgmsYFkSLXZHRNxLaxsUg9gimiqnswjxvze3ya4Xvj9uAfBY
NflL/i50eZa62FBgVxboX/Oh6OCqdIqPBdZqKN22fLxCorKq8HXaExyvdewbeef9RxktUtB87oIT
Ueyde14sPELIYzkUEk7/voTlHcAGGUZFFDDOcFSgc3YYrplgEJbrCbf+icFKCYV8RowVO9llBI1K
WZoCHc+IpDkuNBYOD361xWRlSTwkjbkXO22zG2yrNYosUSXfVHn+Hc9Ot4ITpzu+sMN9TkkTkPeA
MT7LQ8Y45QJUPNZK6WWiFCYxb9j+xUEdtZglfcQ0pxrehC1OSa6icnut/LwiLr0+yMiiNODXimgk
ve0nTGtpb4n8ks0TrgSPJ0uzQm+DvwmugKDBpiGiIJVpJwgPfW63gOB2mi0S6lcPW8Dg/3SE/ZqW
0HA0Di7wDYM+78FrqiR0IL/+v+JoGqvApS8wZvZdAjC9xG/taD86BvSFIJ9nNpdPKxLvPqPUFzsi
SFcVbzRxlMJ2IKeSztuiu5lxXp/M4c3oKlZEHz6iL6NiUadmbJl6q2i6D8Aj3VAat5Na554r34SM
N+Fkmm038HL7Rj/UZlcZp4J9FKE/LB17prLcGm53vNOiE7Z6p+QSp2xaguJgDRKMfMiCnlAY5PVS
YDjup0oddtBO3EdnoGoZnFMVNE53gMybAsEdgA8fHWIxP4hU6LIOdOKhHBmC+FhSJ2UwZu7KDnYX
b6YWK2rgktabA+bfG4K5BA9dlly2YYhJMl9RjZW+oDquJzu+4pBLbU1DfHi5/KclwEmXd3WadnHE
OkxJ0gSV4EoVsN5tgYPVyHm6OThQqCGaFZql95lW1AneXdCDRWJyZczYGOoYplzB1aF5fBIDXVTL
rPh5mmIVt7In3rnYY1mfmnh+zcpcttmpmLbtoX+3aYGv0zU1eD049Dl+nKPcpSW1yGY05dh0+qn4
3dlfMRDrOB0gSNLkmWn1AUkcM9n5aWFHFvxAUIPBLSV8uItLveHbzHQqubNOq92fgEbRiPJfIcmD
HASyZfiHbbl7u1+9qj3cQSdytBfkxKoJVg0ad1Pp+wgAHMIrmSsxslHKR0CX5LjChcMUiU4jybOk
DbAihZ/bcebT8+QgBblBJLWtyz9gK8Sn7M0l32IfYwrqxcdDqnMB/Y3ZVKaPFo8Bmfcvj+IcVP2B
8cDeT8iuSRvjqp0FJjMjazHx/6awnyV99uIqIqJPU+L1/bQHRSmyM6FJABosvZyUGbo5dB8wNkqQ
wGxP3T8S9cEU98tOayVVDsQ2Vp9ckXf1tTStbQw7zqbf//gDCDdwXBojBPGVpN62LuaFx2PnI4WA
gNzApR/Hv1/BLdb2dKAYo5yK9DOOcvspUI83MPlhMZEAwkYVtuiDd5I1DYPP8qGvATqVz+tz9sKJ
Hoi8M2zJDrlxMiCOZYYQaaC/P6cAI+OstuNvSk6hBlDrwf48+rzCXm0WGIWtVUI289ofAVsaDjZ1
o0++aDAfjh4RcEjWjBN051SLZ2lOfXAV6/r41rE5bDQNz7FaRbRSpoPc0iOyEjNgmIbZsDUzGeSO
L9cX+EHH4n/YlHvkSfKmZUYxr0gF/KpzKz5fjW7aGlyjyCt4NKDEAPTF/LqlzS4cidouxHd8O/X2
w9WLuzSaKBMU2CcAvYW2fETezQGNI87UmeN2fvXPJbMM1R0Ny5arpbdpnjim4v/ufPdEw1Z7eIB/
pkRcrYKAEeN5sJ3Jypo9dva4pKmQalq+GlHwl41fjVrWB03uIATcSyyV8/QHFZ8dUVUKUHnyukgh
vIpHL5SY2K9S8Z+FUjhVYzJ+a+Nng+EVKD++tEEYpssseI/EmIzrE3brCJ3GwKkMmhDjzCGkCPru
10d7AnwL+W6IV8HpVEaKq61lOLrPQ8oYf9W9JAU1wnIzB3C7MsoYc99GAFhnOvGCFXvNuNJ/Xied
fvvnWwCf0PLlg5YDHIgY8EVQmEWHP/0AOqDNYYAPY0UEwe+FTZr/W2FUMUMvI/0ibds15A1dGgwe
FOtD/SslV8MViEmBkM9WsNUm0nvVKDbZEqsjRXN4IikIOk/wNg9GVIx8TbX5zyFVVq156O+XoLsr
mu4zqA2IE9IdxRoh9EMRoCYjlHBRTvYXnlwMItIRCpXxbqFIS3QXlik27Ea5TE9coORaZfXvCHop
qEdi4ZD2EeWpRw9Sf43nREpdBcTbIgKP47Sju1TuRjBU8sxMlTfsndwbmw0AC3r3axM6vr3ZmYYT
Ai3In0kwSDcIVAHucs+J9+Na8/b0jsVVVdit8nUJITjmANerIVPl4ou+hBw0lniDzaYdcuJmcjrT
IxJGEwK6ahsGvtTaM8XReWXoLmTGEYxnnhzNcTDssxTHD/Lk3uYEYckZ2OxvAdSe9Nxn4O6xqgOg
6Laj/yIN/1AQU0V0jYd1OoIcGn5NWrWQzwNBjy708sase5AN14oKwsaX4YSxfrJX/IUXxwVPtYVD
A8Ax2Cw8ziKSGQolLGIJsyrupu9aUZRHAiCJfWlNi20qJvHuGMmueIgvIRp6c1p4oWM5nUolKv43
gL5oNQS4ZIG9CklP1f4Lrybb0U1wUzTOvC+9ZRA/ewNl9pWfFPbn11Lg8jgTEfmvo4R8RuuEAljE
f1ax9blBTvnLnhSUW9CQZBwTRyg4ilHucxRl2XYF5xNEUuvx8g5NGgSuEbUwu2ImN0YKHoY3Fqdh
q7rW8NWg7G+MMT8MyUx6ujlWnTPJ2B4cLtpgV+hrmlChBs0X5RRq4yAJmLbds1nGRtG+MI2kDytZ
Togz9iXZVRjeOnfowHfOc4Rtj1ITbEoOJftnd6U175JUHx4boHkJ6B6xlcpgpkUBikS8MBGXxKS1
4XLoOjw3BiTMUh4mmJA2xG6NIremAvJW9JucZ5dELp7nqVfqlesfrBZY+/7tw/53ikIMDN72G73V
QHp8dUcNs6txz09KIe+YBSNhTjKRfdB3j/IRqiu7k7Z5eQ0ZrpQTeUfowQ1SkVajFXzg0oeGcFUa
10xxLg1f8UfE+dTIEJ41wNy7r8vPG/LYI4fXnxtqqGmPRWJs/IfmHFxsNVsd3bAbiOhM3m0To6UH
9P2f6e736QC83neP+WyE++ewtP9t1TgiZjj0fUUk3YhkzXdW4qB3sShxz8yTWnLH0mBt93eN2tku
TKqm6dmyoOHEPTQqFw75yNX5U9sDgba+d0ykvi8q5Ac7XOWW/yQJiOo8HB1we72upwbQLlRHmWfo
idUvnoDdQPQlOh2y8H2VDL/js+Wst0ljQsqyl2aXvZtbHfTQsh668x00LgQcQ8pFHeivs5T3yvXj
cknn/DIkEz6+PyGBNI2HwWzHpT8F0sV+G1zfZpuU6IzFWDvAhZCNriG6DrN182Cl/xZAuARqPvWS
yf/rV3oms9UxRn7qcJ2M2eWOHczlll3DBkROfJBLPAGKLAuL3i6uunRM279dGN+e5rjovD7fsfJE
ciu3PBqExaeoUaxII1gtigFZnoEpNuDjyvqEUOqOINEnERJfpwWDZRKHm9cYiqCRybE3SSq/rcVq
tBRSWEroBXdZMeMpAh0hCg6Uac/lR89Eyse6xjTLoD1/eD3pdkit//OGYaYO3S8vSU4pO9zFnOjT
6NYLSBIvER3mb71d/vDS22wssdOztx10Dj/1YPYgzs/mOc3yx9HOYdr3aFJQsB05mqy4cU9zeoPI
5nlE96ANGCDIMIhuxQTofNhH4IFisp1a0DqGZxAIo+WUaX1Db+ZPrmC7UJqwHXuUzUbuLYyvflzS
+NZTU3HaqyerLYyECKtOLKQGJSJJ3yKR2rHjx3Q0NS5sqoGy57J2t/52nMWfBIzF+k+lf4rnmUfC
APclBXE1wsS0twRKoT3TXbkayB7625gzGPf0Cyn9275+AsiY5+4SgP3QM1gGC4bWpM6PGIWq/khq
4mQMqtchsyHFtXr0KSS80KrUekOVfEsLAZhslNYdZe1hMelUMgU+PMQYecjIfB1r2bG+Yg0Q/HI2
lIfQQUA/seUd1txWEZjXfD6cMSg74GMlZPmM+jmeQ1RBzf4gvFkP+am4fJXj6EySZClb7FNkQNz1
1GKjTNgrjoUJ6J2xrlHQCLUMH2Hwd4otn583TNOGCnvKr2Burru8+C5dGHBnCiI6SSIGZYyi3iFV
PrKs9bYS0RViS+YO6wHLpf7sukBgqLCBLj8flVxPzw6INElNFke8C7JeJ9stBGl+H9FUAl87Z4vO
hTZi1C06jUnVouhUrYRXHUWIWIow7gj3vd7YJdOQhoziNNOL89NhqnzKXDiUQ8EgVWhrxaxrS5cr
t/DhpHt7uz/p5puIA24FMghtjg7YOnX59ctenizZPWTZCRiH0SGSiI5TrwVKJGOlp5irt7XFJV6h
xOgYvszMpnogXIndCTMn27r7pL3mmide74B2Q3Z1M2/rQoFDraR+ZGMr0O23X9zChkTLHSBzW5CJ
Zx4xuloZ4Kq0C+YvtHnIEWtCq7Z8APCGWIb5jMdNucSVv5j7BDOurCCrac5eo2CyIU8LKpMqyxIE
AseKKwHcrm44zQI0FFEZHCuQ3YdHwzhLIQc+pSdl7gNtqy9LSPXHxkUqbIC0QcQGFoDnBIw1UL06
WoJ6nZeclag5dEjNhYgVYOzHgDl9IQvxdi7L6DsBRo/Cxgofumhd3M+FRL8dTjE5MsYQK9FJ+ZwO
QWBkRETX5ly6+hdcBiae1mYWuSfw7rEdoxpayjau8VVGqryM2CZtEb8xtQf/Mh9PmXknlCFcQnY+
vETmnlwrgHSlsyb5nACF5jJXFhZ+LIhOP6HScdbM0Lq4u7j+JV7GRu75G/wBWmiikNkX52uDxMX1
nt4WS6T+F//zRKNIi6ZZqAKgn6oGL208pIEPX1R86BWCumuKjRwflvUzCl8NUhmMR1JROOcV5Dg4
EyMDtCowWFvGlWJzQoK7IXolbo2uWdanaH8WkwLIgcPp/grLtuhFQWziRqwzqiQSg4Dl3NN06Q68
vqKV9lzHoSJe3KuezFIGqfvlZmVhnZdJZEFACG12TXN152Kcl8NTp00H/e1TuBC+oS1ttsI+X6CX
Aa8VeJfO5Nf2GVFCcVaxjfTNVFiw5jZakJu1dFXqM62YP+Ec9tvzdAi0+PQegkFYbffflaoDo6N4
MbNFdx18ZWJxZSNzceuZ5hK4411kwEEpPvdB8uuKJU9R/ynRtNrxQl2vSZV7J2beNMJ2LNH+Pyf3
FC8ijkZSRev820RNTVmefXf22eKjZdUnjxjVzamB+d0pJmlnXi98rPSA0hkt34pY8LHAsU5E4ZEk
a/0OL6Y8ePtf3em60vHot1V+UV77enxyEuiSXKISf7EbrZlSPMiZ3BrPzV81Vnydkdo6qRJ7DcXM
3F8iUPl6uT47Tj+HvQ0LhnRdgZg4dv5bt3kjL9JOQFeIrIIiNzSNiYKSnAy7nGU66BUnFQcfdn3/
e9vXX/84O9Kqrb4udlG4dZ0e8VbQvarjsMJC5YqPtXcSDTH/7l5FcjSlhDoxGjFRw5rffoU9d6bz
6qiOqXu4aeRWeq8iLkScIqoRE7vyqJii/GbhK4DippuhCH6yfLvOygcc7rhKZBeBVjIsCJdOdet3
Hk8Ph4TPSu+u1smVq5Z57bO52CourvUzYypLWFyYrsSy02zz0bAs0jeBoUnhxGywwk9x/+IUkRTJ
0cO4Ro43gAuRRKwbZHh84j3qsFA9g7yuvmz2QUzp28uR7c93v6PoET6VVXseS/Woo1ZKNFn0hTQv
k3iEGWLe7ig75p+mwLj2QdnxXTPOvgSb5Nnl0hpN4Nz35aX13GoxnXCoDIc2E1fz+RBmtk56fkbQ
QuOhAZy9P6lxe/yBU48EUGU/D29Lqyw4EhTJ4PFNRsBT07mAR8Y9snPJS3lAPABaSJsWcxQHt1sj
mC5mzkukOdUhQN0B3StMmXMvJRZ9WFZ7vS+gtr2gsLjtkz6XHNBv3anNwbGNBOpbHDI6atXSz9qV
9Xv3xZbw7RRv/edqn3sxveJejamEy55jkG5rC0EFip8uFMboJobP07u7sTp5SSexfng1M2DE5Nyh
CI8NO6PltXaopXjRxlcp7ZAda+tzpl8Ne9IyPvsi93LZBh5aIWArI6NdawIQ8NwwZS9rj4HzBQeM
U41+ZJviYYLWvTr4gswIyHT41U8oJEUuNNKJ73gFFZ7Ivc3xn17Qq41SYX+ghLCai2mzfcrnS+hH
GG+3pXJR9IapTgBCIQ/TropoO/k7avDuAsQsUTZi6aDAUFCFG8H8Tatmmkt/O4DOQYnBilE9RmhI
xf4GoW2bAJ8clig9wgvnX7WVblpIIVXvH/OifRrnscvl6uZWYfLNjJK73eAVlRwDQZGMqsKhC8BT
LzNLbN/vbnPO4cIjphWRsocunIQ0HtmEm3AFnd31jAw1bkdfnugiT0wr2eUr4RVDy8ter5OyMAKe
nT5Gx0SSgieN+1Ml+3x32jwa/hotP4tiG7k08C1olqEqKGs8eAk2vuhKLe3vodiswHZ/8nUCT8Rx
S493203O/5S9Z/uJFY3/wGSIk5xwsD2qVXD8P0eTkAiDaZ+mTo0jY+MA+o66tSPJ5bfJMV5EHbEG
vg3HX4G+Ex9QfrfGmwzJmJH5JclyPFlQZjuL8sSVv0nFGCxh7bEf2NnZs61NwXUxzR36X0vdvJvu
xYS2IXZm14rz7CwzUMnteBqxp6axMoZvbWtxD8g3UL1lF2H21vMUfEGv0DEM/p+FFxDT1kPxiu3n
YGvqbbr6rtlwWP4kY0Qge4iyL0PJycGca1j/YvB7mGKIBwp1g8f0gLvIGOSyHZGHD4G2ZIERqOPN
bLQW39YwKqZ/sokjJcaBq7Qtv/esMB8X/72xaTQxSbDzCZYJ55GxJQRuKMDzE3hF/lOpt0PfJkAa
Hg+In9ON/r4umOpywL50SPL7dXZ/OT8muqxSk3ztFlY5j6RKNpFDJtXu+tKw47n+dPQXN3Enr6AI
kBvYwQtcyZjISGjzHnx7c3AiqbZXmzW0U0mua1Lb+VyDWYoVHyvhOysuKdE1qiOD7iil1DBrdytp
7Jnb1RJLY08Bg3yiVrTs9uMd+7aVeiPDYyj4Bum8Kl+ddeSeGiU5vC3GLQBVQtac5NjhlMOlMMxW
7FVauTG23rm+RcDaGN6t+67mZZH+FqkSrYEizwECOD5P2qiuN3X0elpawaAs7yPnkCvXQg8qAk8T
vZUIDbAxAkbEymfl9t05SJiam7kWQ83zvMNJ80AyxsVWrwuzaU6WOt8nlIC+/NnVx+mFYyTdgvOe
wSnoUWrvnLftVovv649bGIIV3l51uBDqGWGuV+Hgy1L9g7hSxrKpz02kyokZcKBQ+KZ/ZISEkyPX
GN/xvaVPas2MV9PShMZGHRcjGEN9u4CguaqEnMoLU64rBOoRVdLnoz6G0t/J0NiFAtzuAG2VbGpb
6r2B81INs0yF9o5ZFb9Mb/v8m6FiHX1WiIMh7x314d8kryAFjB1rIoGqhZX2vm+i2Pr6ZV1jDpGv
L2DNzBKmp3USf/2N5sKVASfcoTY3KBgauP63s+z0FJyDKi97EMocceyQavYGGvHBN4OeqLVzNGsQ
XWWLPbBzW6k28PSpgs9sbupQ5ECPU5Vn+uRPAvHrwhO5R4xqOHaLoL5mUZZZRT028brvlxQ2dNv3
FE7jJapCZeg24tcPzHGdVdpLLzKsGZTN6WFNGsMUfhoVge+S1QoKs/NHRtLoSRki4ulinMgIXY0P
57lhKfKQDIK+bE1pvHz+T5LzQe4jhgVyp9icM2tj2yQXwefjrNmWiKFDNfx0M8iCIjbw367FQCgO
B5aFVG44e5wnUzQtsK/PWpNVedbN3kUvIkz6h7XdRgSDMZSEYstMW72UwkyES4LDNgSumAoiEofg
tZOL9V74zkQRzRzcYpZvrZY00aS/vb5WvwWwoYPp8x8Kjy+EpLHz7Md0R7v9ATfZvWJUF8ibKmjp
Q/YAUGwNkndLrfNlqOgfBeBn/1QcHpYmEPZr4RGT0sWIRcA/jHJMywzDwTU5Cpd5DV5Y7cFPDCAM
fHNFe4zSD4aVdXXIVCWt8WRb3TsDgigbjQzDmogHw1xeN0nFFP9qfqnEsFzkoAAbm++Wksddt6WP
vKkEsx5BqN8PlhlTjwy6J22Cw/ZboINyoFzhAuTlXPObw0HSdMYEvRGexEa9UZiHOEz8RvMwib+U
HzwrKpv+RnKPJURIXMLkJa2i+q5aYGCfeiBF6AvcOJLyrXcjbHrloYGPfZY7yAv96f/JFAnJJA2C
wOfL7GVqltUzAjIznjYvQCcqrjLYdaHT+80gPiKRvsmIleUNhfUeXd0WCQiiSfGvOWQo5C3txoYS
4g0OEUauXQ6TMiNCPf8ZjlgiAKKtWfD6Ndjhw3/nsChcK44uMmdn+kpeO3lid39IJY2aeC+u1fJL
UPGuYs3us9v0fEj2iLiNVY3F/zhdg5EdcI+r+7q+xyiUDXtwiJQYy44oNLxp05h7c4xsBch+Nu+O
AiAqs3uk4vRn1KO8cWdF3173vHXE0x3QJcOTkdt3aoAOYzYxoeUQ0FWvIem3J2FdwuY0WC2TVhdy
Bj9NYr4aik7BU+NgFgZrLBcBi0mxMYCHPQ3wDSYLjiMUjh87kleai2Q0IQ7qDSFH9TiZUnEV0W2l
nLnLy9xc1h+EQqRxynvwUmV+mtngI2zknr1j6njbb6kcLkd0x1dG16xkrl4L2kCOez8MvFK+ClOX
qCIIwEvoF7F+FQ4PD1d/ZPf5PUOIJmFZ/v2ohcgMisTk0C1SLafM1CQ6lBTiaSz32kfuO2vWVTm/
FGA0/oNIBcXT87QG13XGkxSfoUdnMtGsoYgItOeW6yFjFec7Ebc92ECp0kChXDtsZZBhfoKfmGO7
cg7ogzUp34Um4r0bhfNzqBPVpqpkNNcJG99KXEtSVv4G3WnddmzItkglrjdfbfs+vxV1V5VRvsU0
iPBXepAkm9B1XEnLKQYVRd8EfDPBhOav0HW6XJtPbilYMbnDfg35WYqlNeYsUeesb5SuLWCOQEZ+
41XqSG84Kf3JDijhrXrwYe+UeiELYbSPLwQVgAHSBamKz86ziUras7L0Qtl4meCFbWX240Eh6CQA
52YdQtQib1MoZkIKL4cq1pNvZcDGkuwvj+VtlWiRjCycoGr0oVIWIilniiY2W1BIP30L0yt3K6O0
mbUCPeKBviG70ercDQyIGzZeKMJ4Ue+iZEgwrz5i3MU7gmsvZxdze7pmbIZ5drvyYdWBtS6/eN4z
EQebEp13i3lRwLfsih4dpZLM/igwyqA0mO1MoEAFfJ0yz2cnZffJPxdKqhmuFdvSJ73HnS6q1VcQ
m0s6IkTCrmzrS92aN+8NISYLhBW9uaU8fanF+shoBX2vS/2sBFd2UabBPgE2WvhVy+la9dueiP+n
7j1mVBzOam92ig8v0smJVYKIIhj4aWvDFAtjtmUMFR5fe9xjuE8rWIgfRbwlK5LA6TI/rZr9cjgy
oeGMERTF0HD9G45emUJ7HyLDIQIHOKDgbpHny8UTLsKTNm2J/6EejxbdMeD25hrN3EUTjm3vmH8y
5T2II3quLyy0rK6VpfV4LbxXbQmjsqkju4fv95ZyG+hIhwh+ypZlTRPfHRL8z8K/25GaeXX39OtX
VSHMpAffh3sNrF7+t/iEGL3x/qudm1VFYHyhPSOLGM08jfdDGtWng76Gc9ZHadBntrIXzHVm4AJC
dxWVz5dwT8xjDphMlTYNQ/+WcwJFPdk2ANJ48LGTN4G0zAbIECveGatJlLwASoGPoC06FCC0GsjH
AEQxi0rYvCxtI5uzGa1kYxyA55EdCfnFfd13Bm+tInsQjIgXbHhSTs50QuWvQwt7gV6gZ9+POSKx
VJc38n8JZkGhXoxWE2iT9OzSmJtWV9lOZ2QKach5Vtt06vIcql5Cnpjpy1KnttwQcWXTxnPjfrcL
7V36c2JFYpcTqm2MQ3A4IPUlzoc33JMs87zsIgM8Zfatjy9IrgmVyXDMomJ0ad2stBuWAANu7wEu
59poHh+NiWNAjMBHV1+bvGrz1RE9qyZGSxakjDvm7A2yTl9BuGH3Z3onOnZyLLQ96Cg1ycj/K+Jr
n35ijA14rQWyGLaLkjLHxxSyxnSyoIcfcbReqOUFYGO6u6kMytNxJhSA/dITXgDC728X/bzaOQdc
2fVVt9xoRxrIar/sBavGpj4YpaI0/5e5zPLgGTXDO13lRq80lm3cPenlRpCdun8xoLZQ0rtUoYD2
tP8OWev2gVQWwY/+GRcnl+tALL94X5hHIszmuARS/ftC5ugEmmGUGV+hsHQ0BiWK2QrIhb+YJ03M
ZZvb7lq8VVDMfg9FzxfihWb5ZKLJm4luxVDjI/p1xj7Rpz1UvoKDHuIGh4Ro8Z8L8Gk1eXVrJWXJ
GnE1y3qUL7g66Kt/2DN6xrQOXTWglC5NLLqBUgfML/CcQDTCnfNNUKEf5vGRbLnSa5cEKWwWzOCp
W01xyJacVkxu7eZ/czHZvnCLiI/XQDmVF5CeXenQb78Ny6IohIDBUxTZhNJ0Zff8MtTPfwU3jiGb
XSxZRJvnvfRxVF0lpnijIdNiYuU1yEzOtr75+3nrIzWvzKoyx2pTDv+EK9j70LYQXKYcDe22rT/1
GAWjwkdtxDk++5sr7vIZSHOMWhK9s5AgaJykZJAE07F8Beks8wbLUsoY8c5op1zj/3MDQDWxzOdS
KTqCNs1ara6wY9pjnhPXsFjeq7OT7zKd9R/0ljHTxuT6aB0YMkb0mu5bYHymXljl+As6B5jiVPXK
cAvST2/qb7E2lZ1tHrgcg/WvJV4UBpCf3c1ufU+iybqwMZvEVZgPUH/JfjZnOF2Tt0FoLCPEn6Cm
JNlHditGPahx1abPRM+ufEo3V8CAjXvGkQzXidl9ZOfqaXka0sDD3QvuL/7/rczM9IzGE9R0boFa
7O7hbc5FRlS2G5dxQSel9psLLfeZs9WwepW+AbgPw/ITqcDzeVr8077l7aCm8USF1XspEfwJlSB9
hmlCL6jkdJ7mR7ClaCnKeTvNsm5ivzn+tngkFUGisJ1E2YTODms/bN8LXUIGC9h1thzmkbo8HGd0
v3q7TGOBBLmqCnb1zv2KC1ECDFIawQWqp26vKgratMYId1j8gZOk0aKJMaVWgkj59ZyqnTqs5WCn
mw6jIxLUJAtf/QV96BrYaJZ78BKU1jaaq6VZ7zkWKrPGrVtECsPrG4Nl2lQgwFcnxFjOaaMrqIcr
vBRotlgS0oV9fMYLXwIAs/XFMkRTW+fZ42tU4ucq6BwKKVc7R9TmuOcInivYEV+l0BRPj+ThXdJE
xQYa+qkO/pjavZDj8McoHVPQOgBdr+8Bvlsn55J96xFgk6kOMNC4lBFKdtdLk56CiLVxuiOUH6Kc
VHowdPNPS3MAjMmP6Rnqeo63NhTZRRpAQ5Du/fUvJQWCFfp5orBWbZzQB0b4ReVDyhxpd+P4Ahlj
BkiPCsfJ/p723dw4MdZqLQRsLMiaCHEh7xoO+6614bgQRBgPvEDUdIOz0YCO+g1RoTnVXS/yt/Go
i9PYr47ReQ7V81Tm5licTLvfz6sSW2duMue9OHRoeDFShCOd8LUckSzuVC7A3OtsKaQ0NwlNpUVi
lO1e65HzlqvOfnTAJTgoBtBc1/XRcFmEkWib3wzUYrt6h07sgztidjuZ+XLI7irt0eHuO+KUNvWb
PFedetADd9LuZmjBTRRHl4vgFz6rwJhRDSh/+yEIR5xpdM/8pGpkJqZ8mmOjFE6zhQmITghgPQdA
Msgd2PchXl6gd6xj25kYV4fbnG0p/5SoaZho/AdiPaqyoCPx77ym8WwLZur7IEyJ82gBy3RlZ2eC
R+PJqyESd0MUs+caX300CDC38ZWw20/aDaA1y4SBmsUzd+5tT6x05hyTfUFCGBppagZZaL9Xtw/P
3VMIZAv8jadPOVJLtAj3R9zhxpGmXIGdHVXlIJfa8A3tLt/V7k5Rv5Lx3iFU2kpt+b2kPFugOx0V
hIYWNSL8HaIkitKTIC+oRpp6pliJWK39EhUS2ujbHcgCDUq4bNUcsH7AR56+UwNlbugUA30lmBgL
uyirusunWuIVKUQ9eDQSN5Gh+f/9DWD3FZ7lkezL+b0/n4LhwYtF0eQ4Ruf6kQiP3RNwIe8rjOKH
Lb/t2MyltL+0XR9jVSBwzyMyWhvdD9KJKzPnJ1CtRodD3PhKK7ONhjSTYZMvAMvhUZ/pvxd4VRW+
ut0WbKNVTFMls9NJipBjPNLEm7uTDqJtQkzQJszhwUVSn+7XBezM9QFgtvMKt3MGKo/02LyN+UiD
aqtH+mMAqkuktXlaNUGZCf+ViwsB6ySqSYMmPHuhfAQKq3GNuPUN7+/7GoGxzil5MWNHIk0quQ32
HGvq3En5u6SptrDcWiQUQtLcG38jNnITA+5WoERRMs8lJvapYUcjTAGErl1qY+4YlQKKM7/9XLB6
TrAwxvKRffKgRGEUATIGiuv1Dn6NBifmmdPZLy5oK77TZUhd2lKMXkquwdZUUcTX101Qy4SmRe8X
hubFML2N7aXe53bfh8TfrThc5U8Q+GIjxLtc+qiD6pmIk/SEwaGIGo/hcfU2IC1qvSErs79bBw8g
t9zJEAC4+ZVqRuzG3IetYjElnk8yWu48nHbtgFHFzDVrk0u8j4PRz1Kjvk/PaVbjv+hM1yML7BcL
jqU5J4mghMi2wdmKWYgcwkUnIb6/YoOc3SSqqKcXCngBgvQOvk2MpbvDfmI96zSfkdsWY2AP6jWY
Az+eEy7oTpXcE2awuM8d9j1a7U2hX6izMuJv+rLe78ZQHQXIcMEMYX92YuNhOqKDoDnBkhr/7y05
QrBDlu8ihfOtYHspxYqOu9DeUKO6k2YOXJYA9zt+6qBNO/wNpxBzXJyumtU/oGsG4dPjIrQY9A3m
81HP/UADn10P/fBdMmsfretjHffEIUy6kjzyajEGh4IjdiRLRvn56TzfoVaR9h6937h4tBMjAHIh
lpqosDJXH32ij4y937tQVtfEP1d9Ibp3RmYjBhY3gXSeoZiyTogWy+nF05QmK9Ufy3MzZvdVT/hR
575Rhdhb1XBPgmgWve+WrJEC57HSlW6rOVxk1zVilrQnS1LKr9fOSC/a4fFAVL3xoh6lELdl/8uk
J2W7RQYDoi2BZI5BylRHwUFoFI6gqj1lYU8vPkiBLsfV39VwXvEwDj1MLN6KZ2hbABgReGxQWqSx
ePIqUf3qPCDbxASXldVFcR+rvEP6UDC+ncVoQUHRDEUHQ045NCYs/rQOPJimKFG2LWhxdd1OFMzK
XIM2kZdc3jKC9YBM/2HM/7g74U1hV0MjmZpm+tB2ko7tJywvuo0UKyHjVQLo6Un4MLEe4yKqDGdm
EM+5mF/n0OpMLhhLDWz/Ds4tYYCa2mHCFOz3Oj835DIOpjxUCZNc57QXOoMXfVrqtBhIrgEo3Hi7
7m5Y580nqVkXWqxZImWUhkrDp1xMiToy6x4l+hHybJ4FYc2ku+GWj2YwxlI9u1P2H3m8ve2SO9eM
ltv5LrAFX0+daoeRag35QMxu+6Rz5ywFzn22hPjGeZs2BtbNqai1qm1pERvCOLCaAjHxJeRiRpZE
z13v2TzIkciwsME2dGicibgbsgQ7PSjIgTYxCraFcteODIMlg870BT4fKXf47javE0sGMa38zfoP
voq5paYlSt7PtrvDfkn57bOJRbry+68TrLVDZup0UuJyPLRzgTjphutSskHOpKNqoNochgd4EdoV
Dmab6HOfvOdyV7PP79MuIX4gkR+qAqQG+bFPXlGV+kTnbrIbT6jo90AUHKB8XCaMTVBpTt56aMaI
/IEJqwfRtb3h3Ks7mUD4JrN90yPU5rER+0LwCiV0RfUy7QAxEYH03pgFlzVjDV4zUMOk5NrvNHcm
FEgqfbK5M1n/Y3Tbt5cMG37lSgplsN1jGSdHSwD/E0BDpcTdTypN9P8z4dKjY/Sajye+9P1bmpcK
d2oELGEsZWwFduPSks2yY2FnfTMnv0SMJedftgNWF2CxHd/1CdOtbIkeZBzdPkoOqB/A19MVF74q
mPF/9yI9vsr4M4+1m9nluNkFPH+rwqar9j8hMPLajZEy3PKwmTaQwTpBd7QuGn1OGNCMqJxWmFbu
QJbLrCJ6N/1PSJF9DnGOA/s1guLDuO5hBjIaN2bVGLne9ZORnozlqNYpIgm/VZKt3VPIGBIXCjmw
JfvG5oZ9owTs4y/j/AM7uNhHoCyacHFtGtfpv7jgvi++U4v5BStCWeBBkvt4Nn3rPKNsZb7odrkb
yt/s8FqiE52pgPUedyaNoHR28RI2duSxdGZJIG5VsaYjTpWrveOlBHoR6MVwpcDrqULEYghbTjNO
Cr++hkkMtbojCa4FRy0xi15v/BEzQN7JOnGstcgcuIvCrWwFbpLFIk+JkXbDbwRi4oXsYPRz2lNC
hYlfZ/czskRGmVGOlcOfcGx9WIi3OxMJHfkHzPmE3JdEyJ7Ub78fGREqCO4RpQFJO3emuJl2XEOx
6XS/d57wqWqj5aFLXpFQXXUG5AkCoDWNULpOkKvmKfFL8Pe7zr2Zn6H2v0mNk2XthJa23VG2hZ1h
VDDZMha8LnaZwW/zIfzziNJysUrhkepoizV2GOIn6pFktdLF6GRvjH4ti/Q2yGpLiuQFrUvGbyhg
m7jBU43iQzWvi/ni0EH5y7wEObsEjmi5kN6uUcEj8thjjqcgxBo0jlaIuNAjwjOHic8wTVeHEI+r
v1gp2MCDaw1TpbtyPR1OtFC9pu1eAH0blk5dBF6m6qYWi4jUrGcoszTgqjwSfbsTacLdXnH9GzoJ
mCurZ7BXngMEm6Tv09nelLHMiaaceTk5yV5ygnSimFOQzRDTY1JkyXgGWNr0mzxjqN0qJZkMPkVQ
hmPQRbW203vo+Ig/8euhsGQ32Ik13pySDd/ArZ1XVZKMBJ/+ReTdrLqXNao33az6FdduAg1OhXg9
PmTczYWMDGXi9gAPDxkXALbOKOmkQNaIZtzur5Zdc+R8rYqVkTKm5O5j1tv1S9yPMnpl7QxaMEmg
FDwtsxN2x+0GXOoxS0Hy33mveUhbrZpSq06JBwiN4H/etFMU0dNa8uoro4/Mg6SVWv96OBlc60d/
RrNtc5W02eooI92/rKMny0IWq+m+3EIvKwJNBoQ4X4MgvtAvHggfwyHG9/E6QFXHiTGUkw9puY6o
tS6VOHIjTlpEF+8PoAKRe796LUmpZngxYG4wM/KItsuR4H8zLoTuIh13tMRu899V6OKAEaUV2Dye
JPvxypq1lEUCS1V9bADF5hid4N0FngiyxVuEJBOG5F4ghjK/JXDGry2l9zFH6ybq1LgPS+bupZO6
a8Z369x3DHepk+Smsd/jBGjuxNk18TtBm35wIqVLWoueOeIUW2+wbaHHPcCvfD9hvm5z1zQJovMF
iK/MSiR2dA3UTgJnlWXpJ4pWhw1LZUSWaZRoPBJOI/Ek7qQH0IRa+BpyG0N1UZkOnr+0LxcxyKmt
sIUCItla2v7Df7sOYHgfob/THMusSl8qk9aI/TqJhTaNS/CUFptKCql3yIdAurk2kIWUh5wNZZ4s
du4QgHkXIlMspLUbBi1Z2vG03tNuOHx/ocoSBZSYAtBAdDh9fknDq0VfdqBZs7gEQn+iOKDmM6fs
K5LnmhT81L6Vsfg40PJExM3AI36epUWlVKk7gDPpHKogGBLZ6IbtzeaMBJK+kAQznK16wJ9Oe4xu
PS0s815Z/44AlQWvcl5yaqi90jDsMnK9c+hDoWJTP9xWkxbxgMS6MdhS/niDU7zEe7hpBrh1y/el
Im/RmGbqJpN0MzYMtGtzoDaPdY0QrEhLc3690VRwA1Rs13el+WpB+mBRxNRl4+Wc3Sen2+ckgmJC
EDHxoX2YXu+r8OJFIqjwv9L7uBDa06G3F4v/C0whVXA8RrJ4f8tsJgUB/PiFcFHE2Djk3GWBWK0o
OeXSxabyCDz1YstRCnhShlR8tmljel0rcYwz/e8/nFz2lGQm4hg4ua8wai22mMbGTbBISDaXvsU/
NiD9UNk22UTecA1vTLYf/b5Q+l5OxzA9rLn3pn+FPy/kGV8Md9j22A/UCGm0WPKBWMYuKM/gbLc1
q196QzWNa46zifmxp+tg19OY2u2dQ1a9rgYL5ST8PXlbEfgOuCvF1/uplrHPxZle4Sbf9lsvWHZM
ZgzFoqT4QnubRUsjdG+Im4zGdw4MIB6hwARFxKxfRb4YYi9SVL/9rT+Ta0tOTYwsdXf7yzMDgFVa
j27Bl88zGBAvBq0HRszvekaGlEkBiBfPnJkiTFIyBbMSK/U6lKN+c1i+SUW7EmTELeU1WITyB+pu
66zYbjsGjaiwW8OjOrqjp4f/G0Fe7lkuZbJ/IBcfGxeuPZvRCs/oRoaTL57f/exVR5MHvzC7Mi7s
7Hzxw3AtSANLcSbMPWlQWqu2lwntrJM2CAQ7UbBNHs+WRK+RhNYSY2Z+SEYLfvfkp4oMC1im/ju+
R5yeN7qChfKGA6smuBL7nTk71+tMt01JrBdwYjeXAzEGpEIYk1eNwso5gaqg/O3+ejSRT4n6gJ9d
y90rlf9w63IRbzrzQ5uzg3SgL4lfNfYRTZCvC3gzjtemp11LI2ELgM7xaPeWUctTM/Kx+nckSLgt
y9EzrJAU7GPr5h87DAmIt6MwsTzoOBYyxQV7X1I0c3ty4l8tJTjEmvLQ3JuY2K0jkMiM0gP2kyDs
yZXoZGtDf4+akYJk2rzQgxEd74E2MtknrgpGNI2kDLlKoxNUtt+/JAeIprTzewvnXGVC0c0JC9kS
Z2Gli/ZZPZOfBL9vmwmlAL3eX8vfAx2dFSMrqAF59uH3vujIn1ZnMLMlerttFzzxh/hEPloOEI/R
aMpNRHAMJ3c/18Ds2WvVuC2ejqVR6oQvkgeXxJbbdRDlTrJK03jKOkDE29S9BOmfwxRuTGacrGwD
elKwu9wbFSae4qloAaM3+CwHCbdlJawAFyzO1PfTkf7JC2UyqwR6SM+dDP1pu8gz7Ez8AQyajnXU
rbaiONv/0fss0vckiD//XOXyE52/QFcW3Wr6fsuNBvypBYQYU3vvjvUeACaMMbiI7v/srtxakjbI
iWU6+EA1Qkndo9Q84D1HCdt9EWblxih5eVCy2DTmLvc9NX/DtUkzMq78gd92xT4BxKIR9e+5CBm9
UTt7dPIiwj/Y1zjfaBhmivAZ5OJsMSBIo/JbYEJLqgEqAKLKVGVvzc9fQ2txN97Tl5xQAW7mQG/Q
Wjvu6ZkuTBQSxEagIQ1IpNh3vcoLaZ9bjOf8XPmH4qE4mJFCwhL2pSWtF53dyBjyy6p7YSKTUpZg
OWMdYE8cUnUkFyEVnruGrYb80qBQNkGwPssrMd77QAzeA06ccD1bgDnSgGYw1X5krvUW5uDzaB+5
O39bp1fbpWpwbWYi1msWOqL3/ICM1YS8PbpCH3TfuHLSXSXt2x3/sG3fRpKVqPOSOwKPofyVjUks
ieDU9aqYLcnTjZWkqMGHVAjKWV1rehxL7WRvpGyi8p6iPXlfNUF7vOGn3lNQ+lhIoOyeKrzfXbaA
BrmJx6BbxNvKl6m6BfKUIe8dF5QkgjE4HxmUgUU+gB0l/fmkkpvnTzusfkJ4zb/Mud9Bw3oAeB7u
4WkhWaqOI2ZJS3X9jthOKvmpLmQJfG83REPu13lB3JhJJfogeLcBhbjLKxuyYf+v+54HkBJMh+EW
U+CH9Kp1njJequyz4bfazeRl+DfiJsUSIiYxTPEEiMbMQ54ujMReHwOZwgqj03rFMC+zn2x9CQky
3RNzuVnfGdgQHcBC85hSMC20AHXvQ/3lpacW2bjl7AKeaGqv0kOWu4QNMaEUfe03/Gk5jAdJ8PVf
P1I3WkR3t/S+vQFk2FAcIYOceqfUmAM1sSD2lqD2tCveJD48IZQPqK2huWhQ68KJ9yzp8L3fdVFo
4+6DdLibHe+EoKrkz9M45g2SpmwUeukLrp++AQP1EvAqtn2nzg6gFTRnGtdMDSDqsqgwI5hznBaQ
LByoG9cobbemDEaVc/FvAzTz/Xz00S3i14/w2Mxdf8KqFUn6ZIUammp3WXuz5IimypdxmlIY0GOA
zZ/N80nP7pyveyhJ+LYc/C8EstWIHns4/ae6ypcOw6gwbbfYp+0pk329RO4TVhLsdKaMZQdvalQk
be6siQ+wAtL3yAdeypI4AxJWI2juU252QUgk5iWaMCgAQkgcyYW6iRPrUtE/MWZd6jhT7xqU7S9B
Pmd4wwOupl+8l2wjxk25KPE3WS6SZp3PN8n85wCqj/98+yNIOW4+uso0109l9zLU60MmB4myIw1C
SUS29dqvNoaf2OKqwBN843wP3vrQxAwRGa9GvRON7lXvcM/T+8BD1AgnRLxbFiW8HOOEwPse1ak4
Ms/GFFvevCc7NkAMLO1FwVImsSSHlVirY6v/33iaqmzsPLszcIHDphuuwTiOi4mRlcoRmuPjtrdP
go/32qeFGSeH5k363CK+YDQbQL52ZTcnw2gBXl80lwtkkZF2gwKAuo8uwjLQ3DArz5r47rGwf2xi
NMmg4bcTx/L1efPIhiR75yod5pWGiYPkUBdpVkXhEw2NXazZTRiVcPpN/jR/SMEewDOtPnP9uxVE
dugzt/BOmR24p9WxE6ID0qZ5tXbht8RWYuGNVsuqLHIi+Y9Ghb+PF1k/3BOt1vC/rem+gpKT07YU
cCEjO0WVhq1Z4i2/iVg9MPbKCzHnhyVHo0pnqBEBSOnO/+N9AVkU0HanwyG6wPpO2MKWYE3Jc3cg
pIywRV3+UPFx91XrdxcRIDSNeL83CnCGEYXanPEWbc1QXAbzvRdyKEai0gfypR8vDSrDvBqJzP+B
NW7EkE1+ZaET/dTzZWWJc7tGjd+jFaD8Pc4z/Je5EPxTvA0jG/Kbh2XBKPNEAtWg3nhMYsnWWGWK
aSetMGa+SZCMEPaMUz/uR/aVarbRDHV5tswwe5Bq0q9fbchkSLxQ2mYWCHxOmvVHF5/YC0+nidem
xpXTnEUZBqmBISpQ2Xj+3AbZih6jibXZQ4ad942l/ECPVR0uBZIydmBjWvMKzRd1M1mJbN1U9e4e
2TDSnHrD9bexnfUQJqU703kr4De2ThF6FQ3NqJsAhD8OaazePbRNHsHd8G9vmpwvYLqQJZ/peUv6
PdiCAX5iMb/wKTffT2PVLnLB/awnSXeBJnFX9qm4x35lo2V8+Zd0mdkxKCcNYrxixqPpwIGeGhpC
Ej8PkOkYCKoN0pqhC7cs3PAnpDfOEIqQd+UO+Y2mZrWwTU8pOMsv0Hygibdz71SDpWqigKddAJ96
gEZqbGjhr1PTbyr4d0O7zpGa5sDUt0q4hbBG1I6rxGD7Sit3MzwXqUGqbAK71uY5HzeP+jvQg9dm
8vA8LwfbcWC2Jvy80w+FiQT4veCDyOTwHU7WNaxbUkVS3ghVYJgOfNZCvQabXO7YRA1B7HgEssVn
8/4Fy4HYtUtn+P9mYlhMMdMs5jmfIE5WD41yyNy3OpOvpx1nPLxCWQxW9A2si93XzX391SgKoITf
6yph9znYxqetX90ambiHoabkTu1one3h8Y7+j+EPWzYttmep5Qsjxo/zsqf9yqaWHlpXvmXAfRGA
hmmQlsxxzcNw1mPWA3GKSgNc04Ytzakxi+eGlxyn3gVcgJDzafdcCLpwsx3MTeV6XshZSh/eA3zh
cslu1+7WfzxQNTw6seLquL6Gye3tINl9AOMWgmkqRVtK9J26yOYVqacRSexq0b667OmS9E32Ydud
v/R4bdMpm+otZTI0uo+ZiCZx9IUHiUK+BPq59e9rCzwjkVlFAOkTy/4LCfRIl+CuWWwvQkjWcKJS
7LN2aH0hq1lbhK/slFsIwoledB2ukTj8mmIzkmFzphBPPfwckcqsyNum82bVBu42NhWPfK0nvO+e
X18x+UOqnka5wwpV5fJ6PzOzP2WXwxywVDLz6kBFcTLMe8bv9VHUEsXo6HjTGQUBpMeFsWkhOc+A
59TGYQ/zoo7qMJM9AdO42ImBRAlSAKncqhtmCcCJt84Sex5LdnP5tWqTtSoQFjkZu3hMT9azLDTb
xQTcdDQtKUU1Xd12kCLKM2kNRCPOAakKfNVc/TeXxhfPca9jYuk31vI7WH4m2kJvdFQ71iciYA+/
Cnj458AgyemvlfvZcqiL9hTZTOMih5YxffVB/HcMd5qBlpOSYwb9ipGaQBp6SwJUuc7CGG7Di2IJ
xzL2YllOdbc4ldIRjlAwxpsi/f+zJip4VxOkRHl1zMl/sXPMP+xDYKVJrlhuC8kojqZupD8ofvS5
RU0XM9d0qLobvyEX+nmQGSRXEZMTKbEcAsFGeUoYOY1IbU41a8iVL4623sBtLTJiaaiCUZCHba86
EWoiS2qeJdrCmGs93v4CwcYml4COLif7KRHhGmfwesFCXK0PQvPu7W1x1rJoeEC8eplKj9ClDFUb
Ofot5QeF+OcZUgBj1bxAfYPC4JWcmoyM/zYiSaq2z6b1rEPtbOqROhb5f5TOOYPSQYrR+dQWE5Id
ZEw5kyyrx3KTTBP0n6GsCGZyMcBmshim92BBEHOS8yU/zQIGh+NF+/nUsILjfeF5ju53gzxPz7Ha
cmcJe4VtKB89f1d4WJkZW916UB6SHU11GzvCTHjBgyUDzDOfhAShkN2dndem0QbJ8RWiLb6FDt66
LkiEI9nbxs3YXve5eLUYCvgHG6yGVoN57jOKD5tbl01mxSDBnbFwqvS7DisctPa5lYkR2xGWmwl/
2vSmY/AYcJLNb024hoM4mi4q905pxXmg0tBn2HvCkzXFfp66dCdR48spoz2+FEBtdhzugyly0D3v
bEx3VntsoPE2cjMy8T/caOSltgEOwgQypT7mfpWMuRzxV9JjnAGsBT/eBT3U2MGsSEIWor+mN20m
Y12yGHPvyQ+zskLQZHzZeH4fWYh9i1PJ+NbtwIuGd4Yk6/Jjkw/+J1FTDFTQfr33Sd1d39IFFwUL
0rGwVTDxgYZxcy5xQU/yDh+c3g2FlbJN3JrxjBt4qAMh1pyEKEP9/Hi02CWaKucEj8ifJzVyEMtu
dZ4TXCYwdCtfrupR0S/QkzvG9Nv8PEQ53nLIiMJaUZ1cumXQ8a7lB5A0Vg/5h+bSKnikJVCVZCT4
AoXf1Ambs6lQPHz4/rgrWLEDnakvwFO+7zzyGZb+thEHiLEoBNW7l4KKBnZZuopc5jEBCuUsKmQg
5NxFaMaPJawk2BYZadlVo3JmIpRrkTrHjVHd1Hgy2ghz5dhZg4uoy2r0SZIoELgg1Nnm8n1GKg0s
ZQmJ/gAbtd9dTj6/VgMb9KmRH9D8EY2SMT6ZSzeV0+FiFT9jGBBcGRFJ1hVWXahL8ip9t6jVLQnP
Ja1i0VJxfY1um3HuBlcuscFLUwqKge7bLioG43NBqG9JbPkGKahaho5g3sAcn0g0kkGyFfU3S9St
i735ycahXoJKxbI20N5vaYdoZqMpkotye3IFfbIzWYbWc5b12oqtWqt4JCv+0ITbnUKemL+olDip
INZJPRVxsojDmxDHRY8kYvEKptFSda1v3RUtJv3bprIzbS59nij7gTsMUS5vpPJg/YAWzkZ32lCg
ipOicCuWtA1WAWN4Sz8O2v4ni6PS9TJSh3GOlTzCq13MDFG1gb/mpYdXQfixp4/MYKbPmBTGURjI
Qx1KcsPJYyoeaV4IZn1kI86p+tVCIG0dlB49VGXQ1S2OETjzs2QcPEM9eCM84Dq3sdYFVgDITTQH
xZfMVehUn0dCGSXsOtcT/6HF697mNf/BezjHpcPROzVcQOldafkGeSawY+aW73xtyIVHRnhBon3A
JerSWXhBDjM5cAr06lGsvm6p+VI3ROCraK3ui/18WKrnQqtAVGlhKsKyZGGtAh7TRsS7xjXqO9My
HXgDoDuKzwqZu5/eoPY+/2tatN9fe+T6GaKkOl5cj70rayuewo50wtiueZ1rDqX94BQXCHpSVINt
S15jI/67dDHjn8cLdLM0IQg0ne4k167e5kmvWm7PqkMdlTGFSLOEi9O3BUCSSBGfjUXN/S0o0Ffv
tQ5lQvVhK+gFKMHZiScthgwNyhmTRHSmzuExEBAHGyiRUwChbl+wCeDe+slX00ydK0r3rt9dA8iL
At64oVOOhWUSmWQeSk5NYpbw5XjAzx8YOXopsX26VJARYDbLNHS0jHsHxyKNR1ZpcScqjvturz78
a7noHtbEQssLnMFx5t0KG6+b078XY+Ie7cKCm4b82UpaAEud83BUnWtxKi2vJDwMWfp95TBiCjTQ
I5VArdJ+wks4VHx0/UXfpFzhCN1kjJw2l7Mv65gkIJk0//2E5ClXDbYZN6bTnltWaIaBDeapS610
Ow7NG29TNjlumTyzxHfRFqThlZcn62En+eM2kMZ+F7Tb6ff66fyF92dCWRDLIlAsB+vdA+vWlZwD
yNoCO135OZxV+YxSnYKItAlE3rk+sH1T55MaT8WL2kibAgNd+E8PBbeQdS/wwvEogt/a1U5svvlw
nKGAOqyFxGBisKvrpk/peSvJCyg/JdL9+KMqvN6h2Z2RxheAU5UHrJjGt5KWGGA+NpbL6DmWhCk0
qDj16fLy9NRfNBRbVL4wfAL1gfdVJp1y0yePPAdj/A+p16dBiniWNPqEr224EZvqsuTzHOfF/w8n
RCSR1QlUQqoZLcMYeSbTqze3S1X3uW7tDkStVW96UCNjcafi5VUpcG/94tvZpcjojpmM5rBufz9x
BCsAbn++Xi9LlwbbVixDpj1NWOrk6yK9nUFv8WPN2bIge1A7FckmtC+vqKCuVOxVNbuc/3xjTy/j
ZvP+c789FyUYxFDavZETHVd3lKXr4aWsfK9bQBKnFJ03brDlNwwR/KhQTXa5AEHlXEbCgiGpzKN0
WqwWGCuXXsqNAGKrYXLXQq1+aWw6muHzrGczpX1pN3zskRltAhXwth6+zD2JplYrxTNPcu0ykeTO
MXjHSrBZ4uZu8VTb30hYObL0IRB4qlszUgOdF1Yhs5jUnRkVGtKRiHuD53HSA4UcCq5jYlXQjI1r
AQZfxfcAQ3cIiBOG/46KTjH6u3bklsLm1XkJYDcehFnwCPxt9q7iNm37/eQxav+RewOGIpe016hk
1bPpHF0DKgmSOS7ncdXZto3kOQizx/lS0G4aLAjwNtfQ/naXs1DdHX0aRSXwpYZ+g6RTvXz8LVXW
3fIudAOY9+vRmE+kj69PaEhiCNrHPGsiSesKw7+rpzl9Rc92m1KhWbt1QdwEEULcnZwlYMKASGIF
dz7c6lBx5p+4lqyPQ3VLJg2ULeY8pabxh4JQ6UZsSry6UHSLKOtGHOVYaqkfKnRSodOOm6eG0KyU
e3czHN1zo+sB54YjGWv550QaqQ5U8M8MbLl18vAywqWbh+9yIz2mLfotWgMihmHFYddy/XVKer66
Mgnor4W7SYANQxsBaKXlgqc7B7uxncs1kexD+2hVkUpBIMUXPO5yV9OWkYerLxR/IAAIZ/zzx2Al
21n3zrXFhvEbMqDFBHNrVjVYxnb1IHnPcrLTwlzh1f0/1LXRfAKv0cC3iQw/GTTUViwzSjRjPZwA
mk4D+SXFVECt0P8H+oCoFlXxXbpf6E8oVK2oNEswni+oej9fzRXtJ7bxm54KFG3EZQxikQrZXg0h
T0uIxHeZn3ZGgQH6cjeNLZdGVkreie3MGBdvBqNoZAS9E+TkO2Zbvhvwf00xXSyQ/26V2m5O7JjQ
nGo12egSws6iW5qvHuCO6amAobZrqwHy+Bc1LLYxZkHwjfALN+dqZ1eWbMq8lMXtgrUrPfbDnYoq
TZLMGoajxBX+DUreqvGezgFlBJUkk8FL9olCreMKFMuOreYidp47GiOETy1fgQVqbv1fIrLxO8hp
xoqK+VqDa9DZSZp9015KKu7mTA7exm6W2/LgoASeivh23pTfOZwsAgceD0zmVDsDHcd/fJUl8sme
TlH+y3pmnz72D7BMSLxW2ZLvocLZcgg+w/t2tEQgp+FS37D+KmljNvbkRzo6YZcNK30ns8iQfeXL
Gg7LxQ7lYcZADG4a4/hQUFlhKkrjeT65oIj8lOLqsAWXwQ+msxVkyFdNfeLC/z/CtFlOtnXVx5TI
kKT4LXAU3/uUoqtRuCgvYpYF/SIuBN2e6P8xBkjSuJa2Jq+6zUA9YZmL8/21L0xB9SMDc2UnRisL
6L5tqsNnNslnckBVIDnpx+qaNxugA6f0oyKvLxK5rJkkABmTi2MxJhsu2QnQkSsz7g5bTRKjga4t
euT1KnDnhHiWr7mK8/gIiZmW4sGDPi2OtuVf3FPpc13CuDFv3KJ8/GQ82RoKDz+fzkLjVwrU7gMK
mAp4lS/qx0ROUgFWokTPQVQSG+7ENpDacoBRjSJVDr/Y7/+67UGcbpQbFG2CNfeSFimmrcM3Lh2v
UDXehNTBedQBjbHxnxCTOEhKYFJN7Yr6Nh67OA5tqNOKGi6h4Balgg8oaJBN6GoBvR1vrh0Qs09+
Fd2TS3xqOR8qZkwSPZwAsJ95Cbceq1HD+CRJyf28aZ3xiNHQ6FnW8YWXxmyEDBwqHY1movAibxzm
4PI+va0WcPd6WB2Tu1DD6A04rMjrnCCVL5GR0q5p5iOz6ZakvgwF5fU5BZoueLnq387INqqv8iwh
yIZ+dT4DEv5XZjJ8Y+nZ2rw3Hto71kfvWV9dyg85mv19M3ruWYWgcCtapGEnqS/Nhu4QeuLdCKVn
vz4oTFm2ogpYpLNiyCbVlD/9OIw+at16teE3RrXodHdn7lEaMTny6xtcUie6mGdwl/SL7Dt4dUoZ
fHYisY75IwWGsE6s4IQ/2F0QA/TmZZT4MpQKKSpIgK925tg1aYso7wrvbOj9svgvpeOKKF5sobtJ
Dt0mioyPQNv6Y4cppYnJZZW4KqSGnRRjaFzsBEVu4LKZ+EqoCmBLFmsyYd/W7vfmhpdCnSmDl7T2
b3Nh577HUZl9I19o3nowFaDMFS20N4HHLO9H3QgvOiGs4cfdpoOK4WRBlvUL2NS2AWDaSZ4VJl06
xagGfLd/CHN/gKGFN1Tyo0lDNPKQZ+30n0/0w7Iq9HMBW9NNpK6WQVK5iJ2U28dIfOBN5OtU+ISU
MFZk2vR75Dw32BprgE3kz6BZMib4c77HsIEa2b+VD/nOIAY/nvvNrmjCOkJhIfgPVHwdPyf+4ldX
9auoBUHSr561DGG0HgecIdsOfuRwAD1nIZhMEI6ZngTRFozbOyAEBkQg0egRVmrmBVwcSVFkAJZ2
YSPoYCpBzbsjiT3Wk5LcDKAe4/uxGeA86xSnp9wCfAAZGsF9AMVhlUhfTaYpt5IZGth3FQurP9n9
eNZA8WPjI+WyOEeysdyBjwVE/fhq5yLiZS8My8LjFUpTwvG5a6uGS/pd6LzfKED0ulUIgVe9ZnJr
La1tHJc/7SPVwPLQI7vULl+l/NUlV6DfVqDJNIHlYytbpNNxFi32o7lBOrSqOGcRF7goAzOEB4px
7bzLxy0//ylBkexWH4dhRMTWLe7vviMgdsTd4HALfplEXeLFFWxL1jllArcTEYjUvN39fG1bwEDy
1ZKtSHd30arxqjPUrNcU5II6QmKM5ZeJg2oY59LVtkQEUgR/HySVehqJEKuxvlqyt7aLTJrnk0L6
f8E9y/sIHZAYVlzbWpUFv6cVdFVFmraejbdRiR6oP/jHu2GJVZlnshvB8Y0t8vhd8oe2LRLRqRsh
G1BY6dxiOsr1RyvV+JIC6vK17P9fFQ+J+Us0p5WmXJuj0uieIUL2jJK2oqi+22rqXrbyW8yG0tSS
WOr+nEDsec1b7Gcvm8etJAoEk0xaJNuK/XA2nn9vnYARnlFEm//TezLpPHObNRGSum6cGEyfYfcH
m2EIo7VzNz0F0nxYRdLwAlu0vehEQzA1ssjPHN5jHKxAN7yYzcJ2a1d09bG0czArXyrwVv+D38hN
GRgLVJ9onMNMOp5lltmo9lgnHWeTnb0ce/SobgAfXwGSHiVWUQJQZFJ7gqedZTzel7iBjDr2+PKD
0oqTUcKrZKmT4EuWZQC9pAtsF1vhRgWiH+4MMK/VoYuQLy8BNolHU9d/6KSYoE6Aai2eusajjz42
mGoxLDs8aa3sChYknE11m1CrYcQpFtcXGhNRqsCwwUVbzTJJuP7NDWvo19x90CdCJIRqo6b1+Y06
tPqfcAvz71y0kgr7dgIXXQZC450a3XcgKPE07mGMT2FTbza03O9/4EgqN4sH1fVK13mC4umVqyZU
Odu4t9TTa7XbxMSp27yGXyi4/3iyzFnS2ho3JjzyV0qWTDZJVt99JY+xPNIgeWlmmXvbOYciQLaU
TWJwKyQr3Dc5XWnX16DlcJmF0oAMa2Y7ZikU9BG+rvb6LMvSIHg+r2hVZYGtxoCXABxbb34pSGt5
nzEngrDQcCuly7B80aAnDKFEb1xald6JbfhPg4iV3Fa4CRmCIRiqfbZY1pMBw/PJ4E5Lv2p4FOnu
5z9WZHvblnNbomflc8HFkmm53z04c9wElwUS9QU5TTTvOz4zWisVeW+/m7iSK69W3lgFdaHZXly+
TB7sqraJVzuEKLwOnA1u2UQpqAZ/OfzD10pelcf02xG3khMifyPhTkE20TIIQ1DQC00SOXIwbmH6
7mBzSuckwC/roaUpAHmDVWLBsveLsIlfpV/zgLwDfTv/+N1kwCb9fxrrawElZDU2vbNuUyxJtum5
TcX32LKmoe4Nxaji1PCjzOKeylh2YJstHk3BtKQ6SZJ1Yn+aWxyxcLz3uzC5KHVlIioii90X61p3
vQxAxEiSng5NsTPGgjVrtQoB+TLduq2oTLXv2cMBZumcSlQ2b3b21VXb4f5AuWzd/ewEFfWkFXYs
JYwaRPmHEmLgC4V3xcIxGeMdW8/QCWpDwEHbhO+bsx8BrTXEuWP+iNKKerEa+E7KIAYlIqM9CQ5T
vDi3slVKWLGVMKlcWTD5PlRfiQ1xcISdmopi0Fk8zuSpRgT5+RMX4bahgrEXocRqzfS2laEiMH2K
EVJVLIjBZ5YCrRSz+JfJgMLpJEnZGkzVz3gLK6OmFUouuoj+LWNvybV1DN1DyzPEW4S1p0JH4AMO
Bb/H1ySzL3C2L5RhXkG4RabmcIHtMv1g1Jo+EZf4B6RJDOoDRPldyVf7neXXNLMirYuBrEKtiE+F
gTdc1ze7fnQaIBAEHfgOqaNKNcggp2N2oOtao822MinkZSvwDFynGXdU4I2yqr5EeDUnOcrwLQAD
NuXkajX2Dx78yNRD+JIb/DWHc5aohqUktXS2sUXpKLQQTK9cCA4ZijIug5DjuLfZclx41dH5K3mk
VIz0L7qF4mr+UcF8skbBp/VBKu9A9vBAO1hn6r1E75FPG4EZkoeR7pdNpJ6+W39H2/jOeWOf6n7n
b3QIUvrbB9JwzBryd42OcRrE4MjfVfiYCcSbygz0iRXtrLNZ79eb3xjuiNbxvMBHgS1742RAVngk
HupEj/7y6qDfF96uXAodZ7wA7IehFiwuHnY7HE7vU7FGQixSqmKcLU0MfqE6HkDCD3b47iNM59Q0
SFXJ5HhCcJr1XuBihqV2Ess/7XE5GfMLLRRNKajnBCdxqW136pTJlHBje5l4gTTpoHVWjA1beFod
vbwi4541ELZ0iKrAqRX/4b9W5cq89YIwoNrB8aBycnQ07z3hYTmfaPbPWtuEK21wLOdt6u3ttqno
a46KXBkzISMH0x1rEK4/shvl6F2fuScyXoOVW33okxgCjlBDNaNDSSdi3nNELh7BWfzrAfn4JRSi
mR/+psrzopacm6vQB3+/p3e12E1WNqHN2MlK8xFTlQS80tJL+dKXSW7FQfHNY6nQeFyJiusVzgu7
ttQh/Dz+gT91QxKmlADS2xspJp0R1FblmJAAv/Kp4KNvy/ZnPW0n28/h1MmS0dRKaHwim6YqjWud
ioride47YCu0YOjUMOKI4selyru7YhmJBNyhP9pvioR98MLcfYSv5vYVQJh8GQjd4doq1H4NDqpZ
aMLYQS0PlpxG13MNR73Hz3n4qbUtCl/WIQQuZhPtTMJdic0clxoRgXmNS+p7XknlznPcJ93H6Qq2
sOS9Lz2EPdrS6viD+b7v13xdlIfl3bxhSruipsBGxfP6FEy2Lbupg2fEPj5jTmti5Zb3v1uFixSY
Dn4SrfDkiwXCVhJoOlSFoIPsJRA8H1HeeoZE6TU46irD1qeFvWamNpsBlz5nygg9yY5aqiWtKdC+
+jjEeU8PO0eIoAUFn9Ka7/7N2qrDc+wPhRmsI6DQDtp1NLQPywPQQM/ifwxOAopaA4qpyhKWR+g3
+TQBsftmw3xvF22ljKihqyuMkW4XhpiYVHWekAchH9LOsMpNqzjI8oosPTkd/5rsLlY3/1ZfzxTF
3wTWrY1idwoxTrea7MGaTypiPExwLkaWxLEVMRge6a+9SzhRH6uv7dL8VvoNW1mN82AGHhjrc9JC
GuEFCHkYzwYWEuOqHwfraXvrte8VGAZehduMVZpo8CbMNnMHmFKB08/ezfvULLzEkYS1f/usps5N
wj30FB4kfEMMki8Rgh6F3OFmADUjLVi9twMBigfK7gjKCt/h3hvuWfO/3vx586hqdTlKCi1qp5xN
izdiVSolaMFQuAFUGvbKdBmixaNXdRQX+KtfszcZjL57/1D0j90W2zQoB+z8aNNiYIJm25DrcxZN
T5fyTUiDNAWjbQ7onQbLQ3gclG+GYH7oxcUeCZs2t1cw7sy9cLmxGoBt44T0+bSAaubMUcE2hfrZ
ZbO3T8kp7lR5tqiWUtkpyq6zXBHZ5eMSStGudVjjjbrNOr+GvGgYAWLzmfRZJ55v0iONj9IZI9eK
wu20GhoAJhdB1ILMjg6mctC1bkU/2dzEgekon0Fxa8TeerZlC26Z9U3CivwiB0yXH+CS/oaaWoG+
dA1HshPJg/jzAG77coPa6NCK+zdUPFVytIikW/1vX02CEJ7t+3mEZgEHBgAg977kkyMscXlgkd4y
0Rct/npj5Vw5kOqUIFBxtlss244aNou9D+eoEs6jLlZxZGdeSkIVrNyMkTqy9d4ZDKZZc29vZVz+
Z1ilD/bOD17qjiBaqkGonEViMcrTmRJZuzQKvH7nVaBsF4vMYAnpwN+u2bBd/w0Fh8U0+MaO6MKp
u8VTdIWiCd77dfrY86N4REcSA8/1QxkzEKawD3HMIqaAnG0KNcjFO2cnCFxAqPt87hHkV2JB5Bp8
TseTMwuvsDFWx5Wu2CokZGjP/ZA49hdIxOTZDStp1MXj7m2vGl10hXYif/+wEW/V3lrEnnl0NIc6
75557bnaNjouhPSlLAaKPDdfr6FO5TCMN2syeeInSYClAwqOmGp9MUnLwrk7FBVewXFS52KFpbga
sU5wKvEoraWnTBrEgpHVMbmAjqcYIVM7OWbWM3WfXeQvm7u2CC+sJNNOKs70090Tki/1QSWwb8AG
ABLpdA6SvSUuPWyxD/DIjcfOxNTVv299PNcWDHKQYQLamF1Pjw+YoR/f4wTLRezgEJ0AM+LC6lAe
TvTODyH+550GWt+3gtejt40zN3iv8TTmy2oAYjmidTxO4kriNHZs3aM5V1ow51jKAy2PmeYZ1gXk
6WMDydSs2P21+MpNPPY41Jyw0T2rsNB5ruVVBNvWSCf6D1qcqbSguvV6Tenog8L4RCnLnV5D5AZJ
jXhAH8xu2eza4bX6eAYsFxrq9OvAZoHEL2pv5K+FeK1xPmoA5xtrdQhhD55Jwk6je/hGCjdebt/c
/S/+bdb04tdBMH+O3sx0JRNNLfLQIyfHiJRHPtMHbYONwLG3gvGn8rUpJh7xFM0o3bllTm41NT6v
zn2L7/LlQaLU0pcM6lJzl8VtovLwskbBdEajtb5eMtimJv6HVY2tD6VoZEjBJxCWM31CPr39lKiU
PgV/dykq+aiL++eUHPOOnQzN4jAqZlfEOL4LpQVxg00ci8U5UM81phaLFA+w2iCbDRryfTxlHhL5
E6RZQ0e6kIq7YH7Ugo67TDv931542xan6D/iy9pZkTwzpHqA5irOpFrgxkoEpqxhWwQhXyZWSnVg
sZ5hnZC39LXf4zUJOogJeCQM37uMtwv0hRoQ7S4mwt5R6AokOG+VY8XV2OMXSr5amrcCrkz0H/Pb
ZKBF9IdMl60xFwHqtUNbH0fIIc1yHoF7MPX3800XOJ15KOuOXDswHcNpPIeci32IYJuk2vFE+McS
06fc7aWeDiXtL4dtSbcqBqcrs+oxvzI6IzupJfFipMTK+1hFymaU59rGzVXme6V9yvIDjGxdDrML
7nneAKsa+PYRgz1XP0kO6s8O58y7pZS9VMe0vy1FJuzkFULRGeq1zX4aS14YVUZoUhCL4GFljM3K
zW2vUiP/q2zjL7lXT3cy52L7FLzgNbPCpCRgGJ3SOP0MqvDwo0tOhjpiOFdcaqyD5GGEoC0Di9AA
g8DDVN42Y47HZIVcKs84ieErbB38mXv+T9Cl2i/L0ncoKZvIByyxNEMCkBLKbhB7up/gCrosarjF
5L6MJ5iPnXEAaHqwatXhKQ7Oucqc4duZQDXC2++lM3YDXd+6awF0PsvFv5AGXjVm+JINSNWl6aRs
tzkJVIuY8pRG3uzXbCiJ5nYQBPrpKsssq4TutS/Qz9/hIYJ8BJUKM6+sLMynejzLcZl0miwhMYCA
3u+WljIEoskWo9sDZUrZcHQyirWjbMA6T5jGID0DY/5zLFuk+QhdH2aFCGgoAryDqGOwYEkEbtOX
rjKyq9/0X1QTRa70Wd7DJ6FZjSwOBEZyhwcb6XgglSYRkjvCCxgh7v4PR4xM4GFRAD2PGNBEzAet
4REK94e1u26uAAc5HCMioDyojFKsAqXfPu1MiRG04bWykocmCqnwXRj2s/jM/3GHDIb0ba+eQj5g
zxSgHGzJY6nUx16cG98y799zIqfIo5NFsd1Xo8I1wjaETrCxkZHrgVeo2bXMC7qcxc1flra7XAA7
EJwFl40k/KKjoDuDOX19EN2ZC5ram6odz1L3yHnoRmdSN7DHNVwceE4rB8ZQHFECRNGaRuwdEp+Y
KvTNfcal0/CuuZz6Cc7eakOhRO3wchrRO9uR8lTwBXJrS3wAzip1qzDGp4wiqg5+57xozq3X6F9O
Qn612HYhjMnpMjMy9ds8IR19677KdPm+b5Y7DvuxacLLV04RRgNfjh2sDGTilQEb72xisrpjC077
Sa1ewcf3i1/BmGKqzmj2mvPdCNtycqC5rFmNYDJDtAw7hQrvvgTINeJo0b/nTs4dTr1TP+m2N9BV
8hS9Eo/tEwPoxDUFaPPMEPrhFCM4KoCF/6jxwX3gbXsXmW9sH2zENXXBmRwq8FZMPK9m8QrOXiGi
lEZwGyEhxplEWe59MvmZrWiR82C3iNWhjogixFlA++bQ3xY9eLoLNVjyYn5ptalFmdwaD2wRuN7k
DPWZhLyKaPdtWBjV5B9cpKkFQpHYRkN+i5+i0DgQwEL4D4yXioUGV46pJoMR3f45BDLCKQA99/p9
Uftfa0BJEQvkbagqUx7wDXS8CYX4hVQlVUj4yeyh/qkJQq1fhJanRrYYpyvlyyhPr+4FS9S6aSV8
7ECdXnlunWNkVxY+dxVEQr/QdfvvyAsbMMdXmcrZ4VytYldHCS2PZbbBvxHac3YWdWQR4md2KUyx
efsnBu1DuWUWT4DWxpM8oOA7gHD3P1WLnU/BjkJb7JGbxqvTHZV+Ik0udAnfXTbYlD8eNbtWOaaQ
uG7lyOf8ruw2VioXtCiVrCBG/0EB6SJQOJh/Yt0oABDb/tEAaZiBN/ommMAT0KE1XUHF1scEk7e3
NiPfF3uCanjKdIvXuHFdTntRXM63NPVh2HJDMu3CtJrSX3zWA0v+LibQHQssQ0enXoETmaNXcIGp
Z2IDUGSsQuQvA5rEPa86GYMj+KzGj9wPIw8uuP+XRKCv7kL0xbai/fUAHk7aEHMcHY8esoO1kWcy
KnzBImEgM/eDUQmEi/PY0ItfGgYwkCGJRybEYJZuOSJz2hezFA092yHbGghff7JBdso7qF7BaENL
R+jXKJjPhTmVnflR6+Drs62PRHvn1ZdBseb5Qdut1iMbW/mW8+ppnJBn4PZ68zvW0Sdy2hUITexs
KTPT1zHUUuDy+awQtBpmkPuOLue+icwFELKcKjAAEw8pkk+D6PmomOLn8zfO1PUDXhp8Y6EsPuQC
9orTD1c9uYErrAytM9Ze02WnDyeoWiSWrGb7VbV4WZDC2iPVyKUlLn6CWOc+VBcSpxfVOcsGyhP7
DX2UBVxZAFDzBXTgWT8dPaeJ2XHDTnwdW1v0qz4PqiAaOHUpRPvUOe7STY3V95lNj5mYOS1ICXsf
Y7cpkRAWi4HJjqDJGi3NuIMZSoA+j5L2b3qslS96lInBknQpSeas0LggeMzl7OpLhYL6DgJUwCiX
9RGGYbo1hvWARcL9TO0FYGBvmPexVuunDMGj5mOjlq++XNSz+iAXZ7qiVoXiRf/fDUBbNaPfVtFP
rZOeE74ntvKfvjmblRQagyfVGn53Rv72K6NdD2KYO5HtKKjFMRt2EMAd7TIyHyvGn8zhQycHV8/u
MyG6FibiM3wvjVVVj3GcOO5VYd3ttZ1xhDCSkCLL00mh3zOCqBDeaIhKSDulmo5d/rEGLcGhiPPw
B/Xtpe1o8xAGTX4U+gr5G3B//fDmmOEnh8vZ5xJS7R3DcP8h9DAnqj3XnX46hAOKmheM8CNiCiFa
6RQFznuIGO3cX3MsThJvGGmxuFZk149QUB0Z5VMJvzsE4HbhJSOxSvnsQuDSLxbGhtNJD2OEK/IN
Z1Kwp1oRm/2divx3PNf5T2ZDxE+vtKR6YNJBbTtLoZ8TpBKNnQ71xRHUG3zlHOkv6kQgBhy3V3Wj
JOEyOTEzmDKcLn4I3jn6ZZXA+h50OXlLEgoLK/ct07W/DXaP8HzoMMAzaupKPdseignIhyL9cm9Z
XntTAIFzDCnNMH8tpcUJkWdLcrvRayVuGQxOyx6RGFNZ0t+mfSQNATBCl5dBxr/AAUoNuXx7pzRH
GhnwP+3l+yrTtJWCe3niUTagzKCI5gE0SkGLhKhgf3v1OANnN4VRpmTnVQCnG1XU9M431Va/KHwl
Ccg7lC2tcYNrUX41HQatvUeiV5bCw+feC6Wp211OYfI8yLo26lOQFabP2Sj4Wxbfrta6EYPZAI7l
VRYESuxfVPXycfU2kWg2NGwK7Zwkt+MGqfvgf6dMB807lUTo2arR/K6ivLd/IoePzgX635BFB3mL
HcYzcRnuKhoR9vHYqJpho+si3jna1t2pm8O4HAKEtWerBTEmEQgzBGOvdkrFPGoqEtOK4Q3qVajm
yq6QsuuGE3zo23z/LP7Lwq5fGWbf2LxCdg1qQSq9K9DH72j2vBe+2XAUsQq6e06x1in/iV5o4VJC
0ENQG5tVadckcVDG573uvmmAy6x1pFMKMYGxhLZxveR0Vz7BsVXObmHGLKKdimMhpoNH562HszSy
KF6GgsuaQcK4/n6rFnxJIThtiUcAU2PjewEOB5lxrsj4ClwCbnPVsvp/nzwdXpqE1nsXpuyv7jDi
1BJgVmKwZzDLziCa6EJYkI4axnd8NuXxrqjRfoYNEL1vhe7QnYlhdCE8jzdu/sH80ySRQsEJMY/X
c+MUIV1V9gjRKWhjTGaVU6nBXGlNkToNwzh+dn5AvTz4c6XHfSl8q76rDMAZbXmW0HVhd8Xbfq+p
mXWMbIYPbfNin0e9S+nLP1LmSdakuDcH2SDCxZ8Kt9Z8dk9EvGv0lNSPZKGrgq7cN5tT234tQypb
6a6RNSdZuiU5sQLkfhJ4ZR/YpF+cZq88mKcvvwGvjtp+1TQKCbmcNpdc8T8FT/Joxfa8M/VqjptU
G0Lzz95OIHtoeo3lbCMtPWl5OQfL/EFBVaJByTW+6ApDSVzNuSrHLLZGuvcRbp6ZtK4ETZx4FmKW
Kw67o6Tl0/e3816oJ9uZWBOjPyjdqYydobWRGw8vg4Spy7YlC1xwWxMJvQQQU6E4R6tebxOkAoNM
8Qr7MMD8mZadUUwmwgFB2CwqdHJj0BI3lLcmUr3lEkSN9EBxFn9JR6omkETTjmnk/Ybnd4++De1y
ow8N6FVHybz1SImlhUcJx753sDU86gN+6qlvWnFyaJ56yzwqW/6Hsn7IChQxPoKsvvTwOyLex2ku
xd764+qPI8hisiZ1P5AE/Kq3qYVgx42Jgk2b4qkqVZVoWpHdpAJV3/etUNZM3L6NQO+wFHmsCLbw
Iv1VVw8lLrHs6++JY08eutvTq/4BlWTJCgKlOIr88PEQmR5FccaYo2ZlxpEkSbCORPI2fUFhvxAM
Ebke+yPNvjdYxz2rUBawD0GdOFggYJdM8QJQcZG7SI8Zl+P0exyhDI6bCTBeAT9DsfQBt4O/kpE4
Gg+rSdskSYf1I7xVj1w1x9KH7K/pSXL7KIcYUy6ZfGBRrJDxjcfRdCButv5x5/dFpIyv6fLrYFD4
Rl14eacZA+MyWlDR+wEo7wcpNTeeeEDHu67Dv6AxcI2UcuWbdpwdoZauJZhmCS14SnwMkFlfQXeE
rAY4kNh5nz2ohmJRa3tHDXNbh2YLtoG8x7gnIvwUh84q5GDcEHhAFTmEBlXjfXiE/aDPbWjQ0HEq
wbLmtZIGhDZ9EPFD92vIyxQbWZneHmC8I3fboVqJyQEcQ545ognF78Zzu8K3fFkfO/W5f5s0WSDi
SzlPBGdQZZu98Ls1NCjddzljiFGmiuHkeaV45/iJdK3JPAKMoRPU3WskFU6b/NoEnAWYvP1FgMX6
0ddFd2uswe77gtOoH7NKcKPzhb+L+2WwWtxmCeGurS17OxB/GMPBYKqjcOYutkFMUiRuFpjGdzRJ
nJ2tyvgJJkZ5+kBmynbJa/fKZcDtoI6bu4S/X6Bxfhn8DkXB01gNVARLqpM93ytaGeigBOvXyBq1
zAU51KMlPOYXtNRfIqDbPn5VXsn0EN5hRnBJpkr1yIRQ3CwfX2yS3Q6IEFAn84wjK9zsmTTG8gx5
9HBF9iW1Pe1ireW3vQ5ipF0nleUhXFvL5GbliHaWxwBCuA8zAS3ZiL+XsF2vKlJU/lsWxX7jgWX+
aKu4ypeKiNp1IGTnzX2TDSNa8OvwLhXYrJqkgaXtjJL0bj6FQVyD6GO9+y36puE+m5os/Vv8XhOC
G77fjJEKnTNBx4SjHAWT9wzdZ6gHmXPHFnwBsI2jTt6X1Z34fC+h3HnLBcU6vLxRVjLH8WKFzcSt
M64ymaVRtocMcBti8z+wb/mykHVq0txnyrd+aFssCz2BNHqpZ3xfQONohRvi79JNmDpHU98Qe7A2
BVL1f7/BrDwdaleXxTKKYOr+rS6pPw5fI9I+E1Qq+UuF1WisSsFQbTX3SHDtLtPtXLsU3gKD2uxb
BHCFAqbgfUt0/PipyfO0tzKpYDiUj+8RPpfkAQici8DgjfE7LgU93Rd/LyPUyHDd+jovmBwga23M
AFBn1o2hwei9ap9xXWkXbrW/IUklq90SS64Ybo2O5qruVpe54vmnFt0gk/G/i+ckrQiXlw1k+rhI
6jMCXnlgSRldrRPBLm8VxJHD+EBDzq7YoHrgFWbAC463es3TTtDZrvh/wHIUV/0ZSOecVZzwfgkw
0yq3XPxf0V7HovrJPWsNtXTq2jshizZfjmQ5rJnoYNtEnwLC3MrGpY3JSIXDw7hw9r3HwNhBIYP2
M2SOiH2lMUy64UzPsLXiBcpQCjZ3Ffty+1ECbmzd9pQ+nAgX2SteBiQ/6BHtzx8G1YGAR4mHZRK2
EzupBM2HxYjVBrQqHIG8hpphDxybDqtS78md4HNA8NyjjercO/hLbYfa/A77wHnda4ektkDYVK8n
X5BHpITYiDtbWOcFWrOYEADW+pmghFyT0REVGzE2B7ieiCtBdnwTOJNmn8P4mQuYhm//pul6Rky1
gy6B5+pUGAIUvbCVdhmoMF6tLXOI6NpT6m5BX2p3lw5WMKelijsU3QjiP+cbF0fczAvh9QqxLnMt
jnV9sb6xccWNWi8J2TyY/Aj/h6l5/FmICch1x2mfHHeS9CweN5mN6N5VJyyF/+BF4lfWA4Y1YA9O
+QsuVT4kRpKE6vUtvAIGtjCokJl/WCuhpamkdXUYW2ZwEtpzsOJuRXZkNjuYRRD7GTqPZB4pPf12
f3RB+4sHzv+y7CGiX18ij2qSvAqW3X58UpO+AQp/scezphUJnVOU+c7bjvGirAiNid1WEt00HNov
RtQ1Ggpr7kwq1le/LhjCwYfGIJZWO4scT092itF86e2lgAoTCjmQIOdpBjB4dq3D85tk/XIGhF+3
ahgVwAh2QHcM29wBMmATwVRdiB8qBplKmSHmrE2Q6ILx/+YLMKvQ3iS+9MPG5B6dKOajcPrtujnX
coOJm2ASfbeSsM/ePrQKLXxg+R+bsxWkn1Frcv40LJ3Yvif91j7RgRcxJB6XrAskHZZrnB/gJrGW
gx1u58gCsbiVzzPt5rmqX0MY4jQ0U7WPUPHevQw0pdPykVeO2Om/xgqouTWYcnxTJcF97XO4JQTs
JPlzCi3Ae3YqMXh0W0QwqbPcqqnhxWow5bjnCMpaO4i+yCTAmbF/mfSgGhqLFKyrFb2VRBFL5p7d
cAqWN0qowBrfybM6voqqrzAXCRaZ+ov+txhIExdmUXY+E/S3pMbw7VaT+0joKHo6F62xsaPc0H5v
MNbXwxhXw7dIw5YeQFcgf8MUEKVFL8vw0xYx5RncCi+4lGPmq/AtamVbsHPqAfZZ7/6JlWW7mlnh
HPxc1WZuHez5CYlfcgfxqi5cH1Vh0eANrupcDfEJUtd7UcmTZBVa2si2W61zIXQWin+uEub+LJqA
hCvJogW8EE6xt104xPzqvJtbFcgoyTBSkIKZ7k9F8oPDfKiQ2xJaVSrgxpYNn1ZIX51Ohh2Rwg/Y
cKvCFKBz1kcYompqpe/oHzrE3/YdAbOQubon6/A7rYj8j339Jm8AWex8NRAl7vxtnVi5Gf14wN1m
90yGWenMLj/j1m3P3wC3dnfMuaPeeXseQNvYcAHMp6p08OHcIUth0KoiMuBSv334MgTRJjabY1l/
M6Ce5dWCu4BjcE1QAD+D6APnMPq10iZiyZ0Tccwp17A1rLg0t8IhL1Tlt6f44Dqfwrsu7fUqBlgn
MYRuwzfrILN2ES/gX0LYrsfsbRrmkNnesr2GIn/SwgvLbCdauZ8UasjIqZpDq1TA5VE8qw4L5Cxx
aDwFmkfOKWbuQzF02loZtQAxQTS93Hn2moGIxoQh0nJ3FVQBg+ZC8mI+c9TsX3yzITSXfpwrAgjD
MAEwUjuYsLloKjrzCie63TXM4GlLFFxERtSFybZwERGjSaRyhjY2u9ZaGjSKwyMOThxd4ymBbAVr
rZlCN97ibqUVA1YtMBflzFOYU1tH8iISDybRPIu/MZ5KUF0cz2Ke3G5JdE3MBKdGECVAk15G4UGo
OiG6viJee9MPm/CLbOkneNNkUX/tMjbbKgixF9XlgzVpGesAGbas5oVEkDeoKC2qF9l5mhZFBfU1
7vprG5KOvm1Kgg5bukV3bZfXfU0ZbBO8ip9LPa+/APsRGEo26DqQlAy5Za+Bhpelw5Ylh5TGGOjB
wUap+VNSWSsoaaBtVJ/OWyHsEMNQ0YeYM1GPzR7X29P6dxEnAUEv9oIc9dlWZ7H14uarxP3MSsPI
qQpm9Qoq7svNhOXV1/pGpf6gECIMbjyQHRiuf9H2ztRv1gUQQs/TAtyY4YSgulh3cc/5bKcckFJp
WzuZMEj4AcGbXdoREf2xCRhxF7pr5s6BOCoMkKrLFGmzHflRPVlSLflBDp+dHIyXy0d6wx+tvYxm
irw2iWZm6JUgPej05SLXnCjy73nGMfAqPOYttqPxGkpXz7S9CzQsnkPKNv4CJ/8LkJTPFi256a7D
X451MSY67tgFC/2cPv3WMnpPF547Af2oxmJxeNtfZ1oOg6peiItZZMLppQMRVzCpJ7KvI9bZJxXk
EsSX2XZsdfogst5apfgMaMwhBo+Elma5g8dGD5KblrfEPjHHQib2vpQv9+Qo5+QRj+sMWLm+eLNf
hu6ugWQE90fmbCEwEbja/6IdJFo7vuVNzlDDtolHkFeWysOyDbYYPJHZcGvEorxEIk910KR8MLRE
49Yf5LVcOYdMUo1hwg3miRo1qlL4bjqRYt40sz4TlzaGqOtQl5atpuPYeubCqC5k3oF72//JqKFV
aBJTtLQuNq3i2qHOxf5/7sLb/a9cEHyT7EPX+rSSdi+cmhO/41JQtj1JkZxpXmQlI13+JKTP3vO8
3YBZAJvG1WnLGLe7CY/6UjCcGxbbALD3VcuNyVcGCEg5EPuNt2+lqsDlV7zhJ54OELiSKcM4GT6z
YCG4UraSlUA6/rTrUVBdb7uZJhHrvwGx2p8JqKwxzXe+eVWIfBY5f3Rz1T4zaxa5jSnqQ+TIxLY5
NQ8u0SFvzGfzBoVDWwOmOQrhlb1Qenlgs0dKRo/sivI/VHAR6Y1b+c2IUScreh+eCWR1DS8A1PYM
3PcT/wIa9GV6j81pDEwFWODNstLXZZWVBUqWBCVqAR+TuXr2SFd96daTPSa0ZKWX6jnzw1mfqsIC
vT1N6Vqf3tvigSuU1nLtd5L9SpiEywlwuJBwSi6m+lyHMU6xqqPfKY36VxrJeDqwI4jHxIVgWtOA
njsV+IQxun18nc3NunVdnt721fSoTMwtixsJszuVyPNgQCS5khRAJq5AcuD3R/mmR89o8QpSkJZX
atG8pmDU2YHMNPkpPTPROhSMSzgLbg+qibd0PzrzRDlUwg2x3Sa+P1KI+CIoJcstMvKWdwU2zZy9
T6tAo7zCc5yobOeHq6D0Moliu+zQ1JS1cEceo1KX/2sFIBYj02HF+NPC/1FSvQu8RVRDsWQA0/LS
QgSNxjDFDo+zS0BgbhrWtrSwtaa2D/Z8mZeSCTaE8ZQuELLxnVxKAO+cZuedKgY7uE31a3/UGzSQ
ORF9NHQWm4sMd2z5v08QDVtg05O4wD2JkRvDheAPkweIkiHF0Hb+egRQccHYnp6KRHIKF9syE36s
Z5fIq33OXIzBntLj/ZTSxcNhCkB1sEovgeuN5Krg+lR34hpWZSSl4MvNT1rqPmMbG4CHb713IBLl
dwL8MbWE4K/5qM6943dUwTOz48EzSgrH/0XUbP/URFsNrjcGhJLrZKKy5Ku7dtWv5w5IcrfkpLjX
4wWDZuGjYTfui1K4oDQ6IYdeFV4k+jFcBBcAtHYn+8BQs+U6E9WhFpeTnniH/lfMJv020E2YkLcr
5lzZHZ2ZBlHvjYwmxUf2gakPI2ZaxG/DD/ThPxDow4B8qM44VsraUJ/VO1c/CJOBUcnB1mFPfdXz
kA+z7JaBrtua5csx0mHwQt0kQzBJRR67mck72uCkVTVfsfQxIraCWLgN4dG/Eny3999KNEfvVZs8
yhfwevSx8V4P0cW6wA6HjLwdrTITB3rWtIYjASle0JYXeFr/A1TenGq0pO9NORvtipgeN7a6xZZd
tPehm7KOiBNhB0/VQqWjt7FObKjEwF1AYH8GPZTPrOBEZXwdDIOOKRhKH7b+xMjh1J9JZl6N5LgL
ChQXZNCDVbmjgj0yKhnkq8qSazmAaLRa7wH3iS6HZkZhlVko28owCe/0QiEWDQaUOwEJrK+z+hkY
w67ECuoJ74alU61bAvRugln+9/0VPRw31hQFRYoCLi7ftZfgWFiY2wo612bZ7S++L9TY2FQDJoPJ
6rjK4kBEVbchvp1JSl4tFybqR9nHw/piWrXNjdl6ojfzjvQ4pJ31ljZkw96lK8OhqCnPOUrjTbIX
6LhyY4ju7yekc7MXF0jIX8SFYklJFgBVaooX4XDEkB962BUIkKYpaY/743WgboOjaQc3Q3LjMk21
v9RGA3Sf9HSqgTy79bKwredsP9kND99cGiFyAByVQygg2sSuKySfXVybMD4rwjP2HKJqIdGn7Z15
ZLR4UnsGbQnDmkZaIA3+nG5Z7xHSjEVOv0YmHAxY0FzqRNNZfE7g4rYFOVYvkghQfI87d9HwYW7h
9BotJEQd004COEbZ5kyIv1MQJbg+WlWCZS/nRgAAPs5uGt5UUZl8UcD5hFgwEp6hctGufWyOfgQE
jMojD9Jgj77Hl1rjwbqVCM2aXYwAM8Giang5l6R1/v4VwJn2on3v09S0edB5bszeOTXsKfJnCB77
pMXpEt9Ibk2HFXqzCzZiNGHVUYsjSLrujvVvqjTMQ4GNGjOWwuW5VYLHreLqelK69mUE7TP+ZIby
+aFWDC1ptNULiJyUmtxDRyhs+Iue9OSj1ygGldCCAYwJ/TfVALa3eT0zUV9QormddiKL0f/alVtq
WQsPJYYl3tocfDkpyrHSbIboZoPdirQrESmH1Lg3suhyIGMz/V33wT2mn+JUVDTp8oT+aCY63J7n
M0qqthtO3J2XqcILtubf/g6ezXXiM3m9oD9iAsKi3vzuwo6vQXonnHdxNim2OGgFW5m/snjufE2U
wd8yLQFLNhRaNjPbTVV6cnmU0DmPZnEdl7kAb1wrV3xT3NVgHCPk2kj9s2olcwRqtwb5xr84ykP3
emLTdgtMLYPu4HtOfQ1THEULI1McyFMV01aN3DYy1jztIq2gs0M/E9sop/hVMNH9goDCOX5FosSc
wpYMxe3lQnx0zZsMms3+GpwvOV5jtE1yKNSOq2jbLY8+NELXR3g6jQot1bLycLSMpzj/uf+lX0Hf
i6mlznq3AcouyJkmF/U+14eoyXgc8PAkqs547Q4bXXTrOJyD69AWkvEHG2eLQzB9lVBKk0c0EiX0
U/gYEKHCxozPgOLJ3bajasGxQ2ho9mhy88B0IwJEt6A6twNmNhM/hacQmLCsz1CwbXci7kpLiFlt
8eU5E344dY+hVd7Ng0nPvAPIiJ3okryBupwic72zVjX6z49nxL1RVhHR7b9u5E8A0i9OF2gfkxOG
AvMq0A3mLnPbfjuY6lXlKNd+vFMubRrS/d5zV2BQAC30hP38muFujCsYdL8MmUUcsb0Ofd3DwDqj
sFRKALA6WidQiy8bNsE9yaV3lMMa4ZlD+excSssbN7djnk/xYo4Ni7/EBLrEdiPPBuEkzL1f9BTk
HRxpwglW4l9iVPLrdi3S85S9rmdeX+wODY6vVWdtUwELsuUk7ZlQpuK2CkunAwiav9p6gYW4QHU6
S2+hA0j5YVzBKSYfo40CgjHUjj9OwxgxvQWL+fy6sxqkwne9chqm+sDo9WJxDPGyay+5NCAAjMcD
kxDZ2CQwxeiM284b2rTu14vMAoafgWjCdajHnQTwjVUV9ZRUTB2nT9E5Pe9aC4RvP1elfL0wk3At
eYw5nLGhZRKXdIYB9MM+EqhSOM2hq0fGpCjKU4N3IyfmBZRFnF+cDURD2qe+SJRfh8nM9xKO24n8
x8XH9AbG/4+sS7Jo1aF1TwL5VMI+8oUfOsTsr4w0o91ypjsDLR6Bsxw1NSk/13Sw4eCo5oDqQAtR
CxScWC+/wNfyA8mtRazE64ft1fbs/Ss4VV4J+l4tcVPMVODwCWC/T48lCAxXMdkXpo51vr4/DoWb
LgumrbRe8B/8m5xPTP9Ky5qtIOjQ7xWPW6uuqfISbHsx1dpQknCEAppJkA4c/IC91kEhVdIHAfwc
7+KAP8zyc55EAmd/LwCNwpf/4YPpVhz9pPFnLoBFWMZWc+bsu+XkWH7+9JVDyEUS+Q1Bw0tPXd8l
7Qps2zIBMNUWgJ87Q+NjtfdL66jBI05l4P47w6bONvY6tbxFD6PS53VwDk5GfhYSeeY5Pq4yMtSH
u0l1EUdVYVypdSazG+l/4pCIhOAbuyYHZDgUUSpKB/IjOdC2vzeHu+KN5sFXJItxN2mVMGzITgbW
LEYPcphRQ+F7e2wupuitoeHa4FDhXAQvcs5SP+Cexw+v9mVAn5NYc83yTdd+gS5B2lCYvSjmV+UB
cwsLREQwWRGz/GfataK1c083bN9jBHzPhtV1268/3kb91i7lPpH7RF0ZiDDDzvuFD0ahhlFWD2xQ
LvmgGdmE9qr1Fvs1NetErKJAziIamNoEPK54gZVKdK3iulhOGGeFTAstFJ8cAUyPZHEe0wboRTDv
8XKxv8O1ZaSOlojK60RADf387ZmFonGyLYUU4KSh/MtbskNX5zsxMGp8FPLtgow6j/rceflHT8VN
zd6skEBIkU73Z7ayBH1gG8jUiiiufqhfP77iWQt4WmIrr5JRHbKny5BHJMdtk6V349JjbUGdDj2E
TieZTVHH3Osz2wU9sfGyWJr5sgidqkA7PV93KOhG6bLUHm3A2HzIvJkfjs9y5OIP+U79QMxYOyVM
aY9aEj37H52i4X/CTIgOPsguxuHmF1r+u6o877OlF+7Q089QlZDwvg15dyZuQKe/6m6yKIdJ3aZw
XaK1TQNIVM1vKMjCo/2ejDVBOeLGuqt/CqOi6sAKE/+ZaPHvN6VPEa2Q+emdGDYzwVtYQrNhFli2
9jglw9VXei73chRGEwhH/LTUKc3S5N+/0hNfeKqTGp6uurE/awGrtvS5jh7XZTyQmoeMIgwEYxnT
TzMa2He08igUaFSrlH9h1MElbH5CPmvHEcE09+rVATR7ueNYdxq/pk7U9Rwet6SsVC8qiAKT5Di2
7Zd8qofV/HGnLU+PTdOEWBcqnaoZ/Bh62pxHJVMBd4kEfyUZf8U1i2XJx7ND+HaDJ8qtjiJ2D+j8
zlACSHNa6GjUL4d4qpanj+mPOsXK+RZTTF1+sFFA4RCrrFck7hVgq77Q2+42qZ05VqNkQPT3SAQF
7GpW7XzqBiRXQSRsgnuHOIjD3tEBVSbonMRs7VA4iIFES72yK97YaC0pHsB3GiP2dqMlU/4llsx0
7hXeCOBQUQg3zHxsrU3h2dsXUw82CmgAgtI+e+jGiBQvncq3M/F8a8mGN0obif4qFc+DR1SuSr0b
UH7auykCe1od/GxWwDXP5rrNXq2MMIVoCShjCh8M9xOGFuE+UUm+qtimv+YtOW2txGxg/bE6uxAK
ChubF4V6EdMsmp2f23oLhpsjz+ls+n2T6Lp0AstDlFKHVNmLQSViKWWyz3MnpFlLRohM22Z7wYn2
Nk+uQDDPGo12spDBJhGXgoRyEbYMxqC/x+BSsEvx9bvbZt0GJX3TXM7MgjPsGovP+O9BSQNtCcU6
htXy8rln1k6G/aqUfT6YD4oCxf+FCWTV2jckufuwSIyZJ/fx34gBWNIjWWsOUr6ZKUhqyStr1l2m
sswG8wuuXGTUcLzNzP9ParTlRT9OhpnG7YfkUMBeek6V71vSJV1pXC5i8FQjPGbwjfaVVWSyB8Z0
0W86i3mVkINurXHdX3bVIUCFVln3zVfTmaN6DG310Xno6yCKbfSGpPaf2L9XldJVY3QCiYiiI3/m
JvMTT0yLh0NCHrMws0oTiWLMbzz5f7Z2MhFWIlMTO36a8IbgKFvTqoaqPpi+hjRUlF/gaK3W6w0L
zrAlf5sR3pKYFnYEZuzu3dErqmsVIoeC5WE0wGjt4MnbFpTYL6ADetdbWoT5KmWIaCFYpxqbJfz4
4EwOV1/lC/rtckWHg65lUNvvnVyf5F26W1mlbabra54SMTEWi6ByklQCZ0mLbd2ijffwFuaWa0td
cQiyKnEh81/N+45JlFhdikQ3GF2whaqzL2PdBhWesqioJJ+5UUXadTFzgrHn3JBq8TGMvlE1T1eG
9DYU1u25BSThWk8U83kEZC5Fcy32Sg7f0H/0ywtZonpgoChQjt/XWrSCRWYy3yO7WJEWfuY+WcO4
RnNy1io96LBzXoR9uo2pnYVqtO1w2Afap007yEE3hMcBnC+HIw5CWjxaZLcfnWxYclXAv5YS2DxY
6Nd3eB7xZrPv8JqkGb8gmMIvOmOb12bd6ary+WAQnDq13K/ymryCydsAK78sG09V50T6qUqIylca
R2rGPzULTsd/CSrSQJQNw2izcq091ZHgpPNKXoo18Db9tRb3gbiGfltDc2/pf5K4VbUfAmHkSx6Y
FMqrjyyZVJXaLd+gl8MmrLdYrRPpqECa/1y5h7VN1ehFnDFJwje/OuvCK4ZPLeyJJrSDz6EWE1Op
4zLXFwJgQWyds1vvw6d5B37cm+dyzQkmaCNVk9Bu1MbqQAi+KVwJFNGjfOcNb9piZTh4bEVcCDL+
IcpWNwQXBL1g7WOyXUMAbkJMRiVxAZQBO4TC/1eUQ+lkk7/Qv8WJmdkgQ9nuFQd31j4m38FFn2wZ
AlqFzm4AXnNWecAkNJSOPLDex+0M25HGyhv7MepsfS70qGzhZB2mfxLIasBmc5ulquUceHERCBdI
kvrjvAMJDDNTGfYklbIxgpK+/9xTq7luIUxgPo7TyN7si5mJnJQY7HuYTJkcLSNd0xHnECXXc24O
JR1KmB1Kj03ozxTndrNaEkyURdKW+R7Y44p90RXrE4OFcXt9md8S0BrfnktLDjsTDkWAUDgGh6Lk
NUZYiVQqq6mahX+X24ry3I/SGgoMzU+IfPBpLxcMSjmHYY/tHbpmP74CTRmMopKdbNmYObnJenKI
075ST2GpPyrXyN3QiSUyF8PxPuhCj5Cy4k3J8n71273wedBR00JA1F35PkVnlTh8ETHRgjZpQHQl
C1ij2xXpi5FLfVZGMmqEWT8izND1h2BKA4gvXSada97aPeBMPH2CbJiIVkRuZIACOmysi/KuIiU/
VWBM/tqvPD06wXDrUTCU+P9WztpfOIWMFI4r+Cprflrt67V4azsO7nXKf3Q8EzOx6Vk9C1rbEA9f
CoInEYDckrwdSARCZhlEEWnBkTvYn0f/YJi/UB+Wepi8VeKkJJINzPQIciNOKoC7dkAuEtWsA5Ct
Hslxr6xatspqFwlUibLrYinzAUJD9Xrb65FWOkHIiDlKSLO2MbhXmyXqwWEF8pnuZCU+6yOvQT3G
JYhPl/jwAlRQ3eV6IUk0uyEhr8NQfH2H3u7sl19yIlpk4q7qc943eQGqE0QQPIrPttIRqp9VJy8Q
sGU5ee0LMlKOr966c6UXfRom3TxmeSIWo8h4Nfbn3b81/I/XWsir1WGatkqlT4s3H9vKjNhawVB6
EB4mr2unkL2591sANrIlFY6cLRrHFij18iNatNhz4xtvzXF7M/3NM6QuFWouzQEJE1iQmBvsKoym
XhqHL0rjUnFCGqCfYoe73f3kLOmEuDwg3yPBXDXjx653RElE+FFQXFBqdo73whBDzgsFJKrdomXX
6oSPoDY4PmCjhkpUOrK4JWOCvqNUBix/6/+VivBF22sFwSl74bte6LBKABEC1KpeIpbCUt7FQX0s
/zGJLbgL1t8fjwnXKkXNaDddeRt4CQGh25Y/Z1SxwKhvaoXaMWC2HAtcWmUpAcIsTvK8xn1ZhKO5
5/d7onNdudHsvflIJuLj7Ccr36Ps7kCBPsi7scOOgQWEoBqq+OPhaUbWV0mILOrkvMlRmC9asVcl
VCevnNfXYhwPKxyXmbeMH9GjstgYL4zie8JPOKe5lqCo8s/DI3kPOMPaLStl33p1UTMyRmQMr8GR
qCsv8CfsagxRRKtp3sUjVCuYOU6nt4d2+IbD6jpcqy4hyk94RcekbFR/Mk7csqwHsMOPW11geVUj
fXdQEGy5AaFaraxvTFB/VnmT/+AhlqWRVULwe69qB7jRrgnh4QvqMTob/vZFQhQG7UJdgi5SevgZ
TrfAels2IkYa1BLKe9Vvd/6pA0XmYzzWDgPHv61SfrGGnIQu953NJN5h7a20jhMIahrxp6qs5Qu9
SdGABtzmZ41oxkw6UqvT9eUaLivlhkj0wHYkVQRwgv2ZfrQqX8oQ0CFWVfFX2p7p5+l0g/6hjpUZ
G/DYzvr5NMaP5Sq+DHtUApr4AKDexuZYLHdQK5Zb9iVFstWkUQ4su/dQzIY+TB9liW8ZJAASTI44
631PENbjfuj5Y1Wo0tLjlrbOHWucL1w3DhInJdy2cVk+UVDyXtSafrOzMYxGuAu7oHmKzB3hYdID
G9jD9YZsknLy71ujTqCUmZQS1LqJrdBWn4La0P+mhuaqhgwoTYhQ7bkI50gmqRbh+FAhGnZkzv3u
FV0VzAEtQmUyOq6tQAy3O3YjHRmKmgoXiwkdJri7bIfW3eq/f5MQhvAtv8uN3u9InxnNyG2t5GK8
foQhvPYWu9jFpY5bxZBo2plWihqrz6ygch7VygqJWFTUz2GFcbussXTcDx5SWUIgnVOKcfiqBS5N
tx/H+lGJxV4wCryrrLmPL6a+WjTjR+8ifQPNQdfTxj5Rh/aNLG0+t6opUqZiXUmOze8epDKKyku0
aePbYV5AUwOgYMoswknv/cQ7p6T8+gApWjt7FPQT8poiXteSL9u8KUqzo51ax7roYSIQzUB7iywB
8s4waqiosmApVPKr7422NN2b2is8QBiy9ToSX6sZLAXbR2tnDnT0XHQnO5PNdvCF+nsUsXy1r1Ap
UnyOFw2h1tXWiVEbkJZ9t5MxZ68avN3XBY5+H5cvipd4W67O9+u/2cd8det1g23igU+yQ7npkli6
kULHIT9cPJ6hW3Knf+nQwO5dDr7sAOk94re0A82Lx7ZZ1FeR6nNDvodNI4cFoqiOFh1QnA1PS80I
2bnSnOMAis8W2yndMIV3JvYDz1xw6u4FBO2jvGv3HLeUK73TqgvLAw1RDUn9N7KN7x0OGsGDXI62
Wd0SR8FJYvyZsBrmyAYV4ujqV0/h+q29cFWoHk+YD6mUt0bhFaoZJesGGir/J/NvZKfEFKoSztBi
YoWlkBwPMGUXP3zZrErFDywF7TES21GSC4qvbMBwuh1Mwj9/ek2PmZ8ggcBfka5Nm27qTrS12Jfa
8TMWVXqDCFvuZeyzK7T8xjktxG+xB/GJ/ZlyjRCt0Qd3ODbE50KX2cPuuwyxLtazJFzlC+WrB4ph
yQWsFWcgWqvlPofT5QVdd0UCTN/Rp2id5T8xlx+1gPVAJmGLxV8A4mJM3hoA51rxiheoVKGTgxJS
Vxb6iSDC4AeINCvbAJB1hyzedsviF3Gtsnh+uSVijMl9QbHwRmFokICDoR8RuSm1Kk5dWp5IgwJy
AKqUBvkjDaBVd/KyOolCdX13zIkO+WI4G1FClhqOowY0u4fx9IjeSw5M5jOwGyPc4/bbd21J6DLc
675dgj5JDRguo2xpF6VTsv8tDKdbnQPrihKYX1uKo7KfOYV5vIvsAobgtoN1R/PcTSVTX/PQgE12
A+frXek24ITPg3Eo7VcaMpUheM5AXh1P/oSeOrcoWvAw/C/3F3J/hPFg/gQIiP9S9h289EAAM1bn
r4nJCoTedtLHhc7UI8YqV/m26fsdvkSAOPI82nEitei53kXSTr9/yc2ao0iCIdcMAouXLsPLo88k
Dh03KWR3JXrh6Uj2eua7FoVvHjqn+LpT9EtZeHOhV+J2xgkIQ1Gdjq2kXIDQ6K8jcf1dlOoaFKp0
oZCp900iNhKf2+FZQCodoIPMpjMiAIAwlMP5uzGU3VjEHJTyE6p5qwNPSBAPfnGRtkeSeAtSrzQl
JsGEAS6ZhMT2AdokyThiMxfRR1sqd+iYA9ovXWp8cMIBshtv3BiD5ZzXmUQlK4Ji0jwLishQL2vw
HqRS6UoVAX9xA1A2LYh6BM7pBytiku7rW+uNRwFQW9YTgsAZvmqe/bIPZowMzM/B9dZ/KCf2ACgK
FRe+Rr8ypaTTVfV4ieatkS8bMicBUdViQfUwXsVwIJn5zy7yBAehGQDPqL3c3JuKAjlkdqWJIGh4
ih4F2Fz1Wv082MexYKys2XjdVRp9gYM4De2/36A+v6CUvPGc4wKNv+zHC5Wo6OoIcqndEOY0UqLL
wCKuibL40KjKZvklB9Za2YcJxu2X4NkmbRsRlgm5T0I3wSZb0vjpsshiW/RLU3BDL8ff42W1cBkI
GEe2PF5x20veH7slmxQVZA7bhJQiv39+gi2E+fkkql/h5nbnqnDY8Tx5uKZQ7wLO7djiAMMMNjbu
TNpfLgRHTTcCsAIxfKMGG1erC0Q4NUu4RAmHYdWNYp1yS65yRZUARuDPZi3P6Qz3HyQ0Y09g8Byl
ibaXmgqYQPXNDdQY3ftR9E4RckExKqcHn53buEJNcqnL571Ni3Pql9qi/GksFHMghbVP0Zp+troq
ct5qwkkdfJo6ge658/2/EaPmh6SRJg8BG5ss7XZs9JrAFWczAePn8gPH4AUSCokpVLfHyFRAL0g4
g6pCWtSgUeaAyXAHScmml3kmIG4aXETeJ1fNlUETw7+iaaVtOAgboGW0K51lVDzK4FcSVImZ5idS
tXgOdMfVQNQwTX5Sl+DEfPVv9VhWY8kgn5lS2w3Cf+6OUclygiEXuhezDYRXPU5vTbQE/Q7x8Rzw
PyO8E+vYUUX556/rBM5Zg/VRQXLRDA9J5roImNgonOAV6XiYpu6Og2rFs9u79Fn/wWANIV1a53Wd
s9NRWSS8ZThEUOPooG1mZUbgMQtsl9kqQOu6iPrkVMEtN3CgeeWDTlEPlY0LCMTIhQmFMHFylEiI
BkjP7F3HLjjRnG6nzO2cgQYzGw3la/PPx/b8ANiritE8Eckn+F5RaQGwkNWuwrn2yy5ZQDjIy0qT
v1lobvfLqutIhF4t0OXVLCiAmjjA1HUo1Xghtpdo5hnSRpXjN1R4n6v3dcRmgtZmrFnetUDRYaeZ
1blfd1jVjtcnU6syOfR6zVWF554Xj3c8pxMJ66yDkyOPWp4JCIcGf8r9Kh/wT5ONJTLviIXFIlev
DR3k9mLj/g25+RXZn4ATmIWAb+gsYVaKEWf6yjMdQ9ULtNZa9OyezZjZB12aStHbUzzllqxvCBf/
k/Gj/9KqglLewXU7Ifw0oz4sMFw5d6Cq8TG5tTztx6nhauyO1tTvwDbRsbX2xvtv/3kH/v9ik8yy
0uqQuy2ubXgPFB16U6fRc9XMjE6FOINPOiDRORGSPBTkLHCe3MAbCu+SNfye/hQkCOGrV+0OCAJx
fdhi/TYb8q2kI8LlhuxGCih6QDD9tMNfqi0q1oaZOo5ZWX9Am0U/HxyMDCcBJo50JtvdnN+elCGy
L+G6+w4B9/w7kaUg2cnhBS+AFjNlWNPF03NJ0v72d8KWTA/0YH3dWwbn4dAm2dYI77fIg9+xHaUR
4N8VYBHH6FAyoUoEFvJQKRTX/1b1KqS6khMOM7Rg8Yv3FIcXWdKGamocDbFJsKesoUWtt28Ewqtw
4J4tCfnEGJZYOlo/NADWDI3qTsLnxQmSSZFw7SAn90kt2Z6DEz77SEHXsm//n7Avv3dmR9Gae3Kv
Ek3DbODJMVsVKz19bhi4VJogNC8BXh4BKJuwT419OpWAyrg33sEYCWZk9om46JyTxfT59leXtm1H
moBuvWXc9fyCD2l4OlryjdptPJVdK56MnkVjN65tJXqe68eBK670HWgk/M0UfYDkd1nPnS0jM0W1
0CAbmQ0Pstd1LoyQcJS5zaHACbDO7lA+c3TkoIdDLz/PTrh3MQNT6ZRi3XpWiR4jCp0gUNP/OYci
owOYIBAkWIqGu6mz5tumTYjgK9tGvY7WPdClxPm6bqWrCh1kgvQrM6oFhAe+H9+8Ywa5GQCn8C3G
G6HMLW5glbSmxKZEnqhoUoPplTynphpD3L+tDxFF38oZyfsw/p4eXdgNGf1gp530Hve6bo/qkXu7
1NljLrc+LH0jT5u71lpfy/0BvPWjTbLVwjQrb8VEx1aLk20L6Re5uBRJq+/YJmU3j7ETQAsdrodo
kx4/j2m+z3+KYVyJP5TNuyOY1HgDjaAUo2mDQDh4Aa1mbIx2kWke/Tpv2FAVtUeBAtBTv3ZqtsR3
zDiLyP29RgEZNq7vz3RSNdbMPrYb0E+n8QJxrJOOWBLIP3v82fhlEvJx7B8fz1unWAXKyOxtKTAS
/ZEmW2IGRfRfKnu4+NLi4YOWHPovQG4xy0Pe+KGZUCodfF+8BlhUVOLdBC9LAhK3En+PIfxbeusj
yM47SLRufBM+lNNb+6LkoKkgZGGsLFdTbV7d6lbmyym1hR6yPqtCceBALQa+dJTALlX4mg1S7i6J
iRtB5CCoG0jeleBL2MqyrHlIbHZmRTtcDmKnBbKZ0Cqh11GB0WkB6BmfmFp3s0Dy9UnL29UzjtG0
V9qoLKdUxVIfaDppaZY/UmCRCZgg7K3Blwvm+g6bASRf9xz8m1lgrYYw0gvEliU4wRNFu14Kj3Mo
2NZkUFvl8ovuxZ6P/I1/TDQFI/tGs6XK2puvWrgQbQ8ZNOtoXw9Ow74F4mbbs1Q+cP418WW0FeXL
rRKjyzsvFjUCPWfDZ8yb2KXLJIFWZXb8qpjmPw4TtCehmfjGom1TWej/QXpfzMVWD2+f03DaJHmV
WFhnc9gmkq37BF7XrPJY1SuZB/DN/Ru2/8y6+pnd6twbZOhWK6QHckxc9u6cmq4XNo9Zc0hJYFje
sU+j54SaFnIRjGPJNzhpHxB/k8s3YX7t4Byl6sLubqxD7CDlGqkmQ96YP/LcBWBvOgpEG27iK8yN
260QcV3AWlCJnLOeNXRdjE0LQU4jiuOxjhK3Oflq/Xm0wL+WP4jf/FDUq9mJGdnVrqNiyeM64IcD
CGQmSQbJCfvf1FP9cmvt4RXZposvKZETkVAGtEywdSYb8NiXR1uhjv8Ha9EHMK+0yHH2fNjjhqLy
NPJ6B9fSxWJCqyb3IsJy9XES5lbDxR0cTA6EY3m6H9ruTJZiGz2Og++OleXJbZ6iPn6Ktj/pioYH
uD+jdd7ekUzffQVooFCcAxdlpjNe5kQp6Z10rxaGbDDP0tNRPY2ahHrP4LXpJdpuTSKPAonfkwxW
2czHQ20HTBgF/6xCQ2LGhBoanYUj70nfL9aN75bYX7zJgWnY9yYl7k5YK9mVzxWIyTj5ehwRSRMf
q6EtLQboyDg7Civo0F6pvldN7r/Ye41QHJQOjGaFJpmAWHERcHgrweP+kOQDU4JRdZELheRJdIf/
WuUWft34KMOih8rsVMKoWCnIhpXS+GdoQVl2LsUxYDlaCKadCneXuzTVO+QKZuEH6+qWBnYnHUah
9opI7K7BYSiR2Jn7T7KMIJWkMWkBpLFdMkPC6WVFIjZ5SsnRhGfRBP5z113ZWj/Uv7FMFwx52V4Y
dKtHTDJcjhRkvaE/kSios8JBAIJ5uQfCvzCbRANGpEhk/SzkZ2wZb7SxdamVj2JumI24MtZovW0n
J/h+4xaJeKJzXC86lSw88kfmhRHsg2PQA/kqF1i12w4hs1pLBXu/9CvTY6V9Z7z/+r3143M93++q
zJiZUEZRpogTlYMLlf0zA5dXFkSEYGOxX29dNpSwYlG7xKaDcsPJWeAXjirFewLLb1mx5bB7bkN2
lcSthkU8tkzUlwNfpZ5Kp4nREl5rDCAlo1+XoaksT0vT4Wgo/WeMQMUX/xbodZWcJr+u0vj/uuUm
b0QODdVSZ+ELpW/TvVtzuXaL2iS3a7iw6evst8EDwfD2g4/TVxEj8ATPW85pZLbRK24vSPo0rZ/k
/gXzbVjzzMBw6sYI38HVQeqmqdbohorXPTHXm/5xqe9OqfkSpgzv/ez24pqqmYFfFu3azD6TpHNu
LUj6XVQWU0C2vANH/I7GKgDv98aHZQtaa87R2a6O9+YswLqMkpVHHM5UIUUJs4HQzLc06pvR84cL
u16QYkz/d1+V3crAMWluLt+r1BWzUPVFIS+shEaqVTPw7OPWsf7XF8XjeEUYZs58y7KiaCMkDOKt
qF6bLPH5FEVoirmO9UhK1vMFRVMLnFWDmbf/uNSMXZjm/oVmVfy+kX9A2Nq6s7u0MUAiqCINJ0Hv
3N7Dt17RL8+3P2GELyegs/AVun+qyVc2M8pWvW7Wayc+prmoJ/jqNUg3dLJ7jSr6JpRTTOPMWhAD
cOzA7tjk569PBQ3ooJP05mDnZxjne4QwPyVOCa57yDD45ylXqfeH8Bns7h/NRGdN+pWJ9NqiaUo6
La/l59PfFel4P5gFcH36nyYNbO4yZw88/sY2oDZ1icgITbH/0/OqbdJy2vaDTM8g1Hsh3qwmoFzI
PFduIKeI9jDRw6YTknp9t0I1FkJvLaUomNecnaCFBMbWTWk+wByGn3uNpHl+mK8qADOkZvkDJfPY
j0Mwit3vUfTxzUxFTVAfs+0QrUXZbCitwDH5r6POiPukBOQUttpx0zYMQnaxm4Svt6AOKRr5AnZk
8caseGuFDzpNQ/wL3eUo34Kr49Cd2ZP4qVHPYQ6Ib6B6MlXJxRkM05Ky1F6P3ZksetnzBpIl2uoZ
m+Y7KV7/6Yc394bAXH4AG1xP0uKDxduB+DmrzVg7UB412qld5HIzdJ08FQwSfcPN/UfZxrvqzapI
DbdnusZn/Ym3ivXw2JcgOQ69O3/RI7pmRQWGpUaHKlo9ahFfk2K8nTG9OqQiHyfyLTH4L8aJfaP7
dsm2NKVBbEN2IXzXpCgPXuAxAf7NVSw+wNGtz2wn9S+mNJSFTiUk9zXyXK/RUP3vpslrYo9v3iGc
yDTkhgY3NvYks7ZRC9egWJGwkKqthTZiiPt0rsqd670/EiHx18vIZAy7p0TYGN67Zykr2hPTrDnB
0cn2UvgP06kpJveyKCapNinqk/f/+o6NH59oDk569OUcl/vIFNSnFh8vybgW/SF3p40Kv0AQG0Yz
Qg8ylPcYNExB4ag4MR0onWoC3IMzObSF91y7v4X5UZveYsUC5cQajxwIwrBPGHCeWIstBp4bui4v
DUqV2mighYFZyJr35gVW7dTblPQZ4hDU8tPdC6dMp8HXTigSsUmuF+BILW7rv5Hig4geyyFueOR2
xzV+ZyY+bn6+rWeyV7WrHY2V1+MezlGe0PqW3Vh2Hp+7bSDomIM+A6js4CsJuPBIENCOIPTs7XRh
H+BR8PPMj3T3929HCdnvp3cU4QUTz0uwZS17HAta6CqRjS0hIh+3+c/W47sQ1fDFWHNhPNkzEO3L
gVsSX/EOhMF0GA9K2W1q+QlgoRFscocB1P+OjDDmi7FzsBU9H/KiyodW9dOHDhx8hSaY/U+XYN8m
vfcPZeYXoN/nQNQLAEObx9S7GVhQ7ce6fnU4uVf7i4uRGAgCn7IotCD7jgTIbSM310g360rz/K2q
jrkl7yyvE9A58MCjbIii9IR4/LmHLe9SyHP5A9ef0RhAJe/yqDVZMAYavS5QUAe0CwlzMJmYcyRh
QyCEgHLMPb/ImWeP0EAXcVTZQOcowdvJziMB0DEGtD5nTDu44B11vVzbi06ymXXbFIRCewwIVtV6
dgDORSvWCTwgiy1GrEaFZfYx+VP14He+e/65xFdI7Janz7R0+IZhLSJDDm/yTREePIrh54oD65mF
Z6EAQzPwcqERnO/AeP+b3GU2B2nKRH/naAnD2r7vODY1lyrJuQNxgNnhRZVSQOnrnY6kc9wUoH2E
1R6BdEy0ZnN1fN63UaY4RIRoCJBtLKOQfJqO4ScVLKuQDiX+AaNz4CHJK6Cl4jefTB1RlgBBax4L
gInFTnec2eEwVRhd0AFR7bO1ZliXoyvBQS048hEHpDIQMq0tp0tPX8coFpjiIxQPkNT5O7/DlOOz
LtaEss6iUIKg+QLAl26f4kOWR34Yq+0AqD+dziuPNRkrDoX5a0TdQtfrtx9rnRX6DOTGFij6CjWW
+72bHUqyzWdt/yYzO1bOs/7J6roLUPflfk1FuFw4cT16sbLhvQL7hDOftLn2azeIB7eV77qbmY7T
aMkjwBC7I74TTFxkpR/dmTjk5JBqw6ysulMXyDcMnNvu89uK2UD4h3Pef6IT7w7idZMmodlRfQsn
wL0AF1YVX8mTJkp4PY8fY8NA26ThXSjzwD7ADn0Aq6c5dx2tvtrBH1ocIt4yXKMElLBhGk8YjbG8
UDHyZjSjN4xZLA1ETARfSXJEMkvKajFm3e4V//aeA2Dv2AUuAclp7/wndqQ1QXiw+mxiGEydL6uU
gX8cGNy72edNYw0FQoZFXnUcHH4ouWZNaXYwilmllIs4xhVkvMH/VGZ250aCcvk0yv4dCG7l0M9p
4GPGW0j4fLYVxETOInUEVrW+Ouhhpb5lJiq4xrPHsLeeJ7rC65Zkq9lTmiCkI6GOgChjwsNPiPaS
i1vKkiiQWCoWhj0Junn6g0qjQelCEEPvS0OeuwuYXR+QxvPSrWmbv54YKZnbncE/ypzkQ/z65gcI
3aIYZPW3UGsxhEm7959otIV6GTsqJaQ8Y0LvXLSZn1erMtNMS4NeyxzzXn0r2REVTkXPg5LGzM1L
R3LnaFjKqK4ZLuPNjL0zZRMoRC97x1/MPDKN2h2wvAukj92U+/NEZwy3E8Hz72wCHhdezHD9NzQw
kQF25o25UHktTtflk0TE5CDj0Y4PAAMH7kDFPgDjUscWiXd/uU1sGK5acecsfl1HjSWT28XX3Rs2
/obqSHOPfeT9CBMU66Xvl1L4r87J8XTOAXwCdB01KwWcA9XZaQF5jj5VqBAG6CCr+jqHjEUakg7Z
MM4zCpjFBPgVSDGZDM6adaPUxnbyltGHW5+dhMtDGw5XWeIjpaWREGcVQtig2b3IGW7uO5HsRoDe
Vz5CRIh06bjXVdGmS8t/oaShXmgbhSImpRC+0FR/+NjxU9o1o64kO4XNeWjI/d9Li1feI83/j32X
c0GgFGu3YIx4YhS356vxh7iVe+Hf2FfswAmAckFRa8b43cOQ7JTrPWy3bZVq+9ZLBQOcBnUgkE/D
m56XZkA4eynFox4Zn+kUEezZmEhdlA6EquNZ8apDKk/D93kdZuaBl3eD8Za5nJYh78dPT+077ZM+
4GCb698ITjH+NWrSDlnxxczkkRimrnlXzT7rKTaH8q9flAQCTq2T055NBQDIk6E818ySZYmHWGhQ
oHwvhdzTJjpFsHgNPHV/7ISIdN6tuzJHmMXjfA80TpUp0QyPrhU76510RlBgSA7O1l7yDEOlwQPf
7vyom1mjt6ZoH+/2w8b6FqflwzkF77DRUtgkvElC0N+7YI5kKuPNBRAtwDRA3G6OGTKDWc0cUzMP
azJsejVy7KtW0R8itISICBaQpqb8+DG6b60fdTp26X3HCRM0+IOxL4vlnQwKp4/0FQYrB2DWIdKm
uyvtIc7SFESS5CpzQb1+GK6Ixe0siANzUIqpjx9/QXhOv3HVQ833/8yVkoSvZYgibpdQEeMkRDTS
GPmW0dLfDaxWwFyJZNOSlsI4PmvJMoJHeAYSHwdYTVWsSlFVqsonoJLG833bn6vSzZ1B3pRsSyiW
c/1YnDhdk0HQmfWv/wERbaii+hfmwtnrSA2aprPsC0D2ztLo77UANMyzSoub3KKFR+tdsIZQ/Ghf
Pk8HuoESYcEyAPaOES0V8BGh/KHBw+DRAon4XnHbEW8kHNFLgzoFGth0FuY/7d7STB5FBL8BtFFH
Ghvc0yV69TC+dkJLXUYDko+pPQ5eJ0UJPCMK/xiG2/r+cgr4BU2Vr8DjhPAmu5iEnTPVM3XS4PDs
/IjFYaX0xPefppqhGNDBG2csQDNpeDILwUcmdCqk/j7ibrpvsMAsByuObpjMujHzPumB6WnD+vOX
i/LidGBcH7eCfCyPzqQxi53vArC0LrXXHEAsrVCufTnq2S0p9dOvpArtITkCFkhOsRdt63/56pq+
jB467X6DHQ4SdRCFRiI9lSGT2KMGbmiMx0OZDvJhWyABmsk6tPrtkLUP8gtPhMDqfWx3dVpRyPy9
ts8oQdP8I94KcSQ8T0mXjKt0ekeJF27/ZXH8x/+2d90Gnwx8WB+Wpd/PgwccUk+HU3luBJuclgnM
GDqYyMqtgmKHMnpLdHowd961nWH1uGHZzZKFl37W0IMoZ7uZJkeH5i2KtZYxG39KEEqwop5JdG8I
nGa55ohT3LXbXAbgdyJCskNtkSrwyWWIzo3c72Uz+QwZ2pBy93FoWuWDgHz3gu0A7SPkG1lk+vRK
+1QDRPZKm6wc9lJ8g30PcV5rQUQAsbOkbnAPnMz1ifRKZjs/jxJ3ixWBXN+ZeijyqgfV8GPxrejY
3tk1XWvBtMR7zAWS/mWVxCALGfa88Q9EkovKZe15V0TaI2P0/r5ofe2ED1i/oGdo+LSlnjtYsdz5
KTmHKVp+Wxo2f9TmAcX/kF0rbakRjf84Udwkc3TvzBnNIvNYhvdOO7Wn6Eo3OHiVBFaRPv/ruqA0
lN4LMzyr+IqtPF/njKWr2/LQYktGl4hT//B/HhWYo68TuDiRp0dDizEubvVnvYdYokvmMXo+NnTl
e0zW5uMErAMNWP2e3gnEHTULOdzDR/optvrALqVPDTC5cha9R6G5U2GjYB4MjTR8PSerW0/Ov8Dm
gZNbx9ihxKUDwQKlVSqszVtpISS55ueNroFthj5NUA5z8skoaxoTqunejENLxtW5NCUFPLsERsL1
huUavnl0EtBcpKUawbMn7GgPZguLLue6LSHS1a8CMmDILAt+FTo1cPu+81NLTnDBzl+D1cEy/T0p
uhdpTk7virdNP92pWeboZ+v9xvrUpJD+hlNUQFAr0zaLQKrnpfQ6XmVmnswch4irnKoFDEKYhHy4
CECD+i3b7DLrWdyIo87lPLrTT8zQCvNpP1RVFNMo/RhYM7gfdpqB14geprqsfl0WgWvxp/tA3wms
21b60HQgpdqSg1dsWzx8HhRz2rDuy6Y/NLOti1HRKovTCZz3DhssV88x+G5WzbA0operZgPvJMFW
QMe7jbrR/az+o3CMAdQOOuTyFFzx4WmXCeNJMmElWBa0n1lKnq/oV36EbSVkp8wUHH813xvCjvVF
Eqdq9MjJtBi9ikeQ0BILob1lUes2J3zFk+y0Rs/C8zhIxcJktmG+/lRtVbZr0NBrotN1SVZCCSNc
HExCRZ8dVJkO1hWRR9Vf7uU2feCHu/a+jn/BQ3vvhALSWkd2FVg9a9tvtDEwU+1HgJay2Q9x4x3G
BfEhHG5H+SCJTzwLqD/nuKBpSfLAPCdBIp8BfnZ/6Uby/8fNFpIv8dWQTILF+aHcyuThV4E4CFCt
z17BtHcMAllMwJo8iH+xc5sQmfPCVyt+umLbZ0jptDL6pFnvB0Ryct3LYvVEY0OqbENWgSYFIk3L
YjbG8qcpc2RV9W02XLAx1sH6VdTnywLJScIEIO0b0qrDLI4psCf5p1lh4RsZSpoX6CPhrMPGspTm
A+iUHDFxLV8Bp1u2fK1yM4sa5uUY9CR4HI0OkPtpV/BsNaIOWVRUP6WW9VxNSVV02qbWDhXAI2Tq
h9saAk5zBp1sfT9ZM4LCobqDKLTHl92YWxN4m/ZFL4pL1dTIAHqt33sGp5yO0QNaZlHpgnCGhA1L
tfFCPo6L0CVVSs2nbYLjgtSHZEh+aNzaBivK8kv7BImKTXVNEVOnQwlp7JcqE2+HqC82trUoOMD+
NJsjrF8prorVFITo2h451Z/1XDOzKm16x0PNO3zowQpvTT9a6I+ODqnDluC1HIChQao1ZwxkqTlX
RFcQIcU1+wEd+arrpnqxKZtn8+W2tfOCk0DhQcM3tjjuOmvs/gbaKQJGud2FQmlDv4XEDX7IHJAr
X6vZ45EgDhoOl0c8SP1h/+i3hGSDj0yPLLFHkyJp1NFyboKZ+evx4i/w+9v4qbN1ggtLmuhkmdKO
p0O/B7IrmzpOXgPI2+veVWQ6l6WoCF49GzLP1HbmxRKLXRPIwuQ64MxGwTB7CKhC9Gt6X1r3cZTh
HtuAGIbIio++ST5T2AZTEMnRdALAS2rXpS/gQRfIXMlfSxIA49Fvzqf6DPukhZjRJ7tm6zeiusXq
3FewnaucGv6OBfHOFVicYAZmOj/r9U7l6JJRM+/oFEsKvuG6dPP1UAefOqHBXimFae/++Vvq/4yU
26lFUaXHsq00aowM1117cEuaqu0K8dWsa5fxD0Xk9sqdY0BUeYOEk6zb3dKg17k0omzNbOtzpfMx
Q16TOvP5OAxJXWPvFveZhk3b5+vC0NmsTDeiNpkr1AlLZyWhPBEsFg4jrh8tB9VWsrYyGpic6B2W
+4xLwNiNHhg9hIoTKAmbpe0O/6f2Oz8SxMyBf9qQ3uEIp118WwcGRZkV6LB5KMQe9U7/RCdnCBFB
HzWS3qPM+vl/3+ZcZMFVklZHRUbtUMvnr1nE1ZDaPrSvM2G92t2ff4qHw3cAtOBiwmDZ7uwJCShn
E50NntURVUhAIbgV63ghPheE/osUrilhYr2+YNNTnrkL7WWR6xzYwXEUTDaCRoPzHX+eV5nJKb44
/D8Oy6caeHT7K8CLqevXsKlYQYKlFJJXaFXWTZFMEdfnYZMnMMjniiGoriWvPEANu/huwsUxhX39
0nNFgjqIMahrdQL34ZiZx5bdkLfYkIGURFuu2E5Dl054rTEzz1GvvvucUyfbU9ML6VWDBe8Hf7Wy
qUyLojewWZrCRa7zN+YNSX8rmdXHCOKnXqxqbYdNruJsJmFwscVZABx2vLhDQTk46ap9/EGZ+R7l
8/zuAMuZaCw8XTv1AJfsKg/qwDwzmHkeeSt/viubbkUv3sAyiazPDBuDE2pDOB8HQSF6/yxeOiKd
9jwsnMxg/N3z+EYmR5Nu3iXWsDEoxCwc4JgdmHJE16SuQGgNWIueTu8q0vO8bzZuHTmV9+iXZ1Uv
xnCcBEUB6S40ELlppmpqoEgHk18UKAcLLao8MQsKRYWR0+LDK5uHtMxqr7h0rH9EFafywOFUoHZ9
4aOM27wAyym2NZEEJP5jFqdy6G2X68/iMBoH7JmMaJsmtZ4VON3o1GW073nMGNwHRNyTqfukmiTr
jGTVqzq6utfn3aOvq5tk+nJMwQK3mQzsRai5tVb37Kj5l96WFmqoFgwcVkXewYQGArv9HWevBFJ9
rBIeo5h3uwR9r/WgEGSw3yZu1FVN+3YQKiksLHyPSmOyu/WKzAlTGzFl8Bd02A9Q+bFkymjLbUPR
C4yQIVKnwKthtxNHQ0nSI1Un1ReeoB2qO+rc6fpJO8N1uKlmofThs1jtRtgaZvS5KoNtZftK/2q/
VMMmZ9WLAuhgau/s9zmwP0e7T/WFy1WIJ4ASnTc7gHy+7SfMxVKGllv/FsPCqNPaG191LviLQikX
60jeN5Scgr9efnhCDCWSfhjhqGzdVe5HLbnxkcxi4GCJwCBJYDtYsvqYRl5ZonwX9qAHGu3HtPMX
W2quPbWjSuWE9ptVIiF9a9q+Yndf+vOT1EW7BPScmCuz0CyXROnOgim9ZYcF0dxHfMr60UI8RhaP
2xlvBEdFgsJ8qsdsW/u/uVVerI//kT9WzkpiXyqqNpkUX3gu2oF94njvSq/mIBX14fmhBCkHu6MZ
ROTNKSA/Myrfl1DLlcWNUCKkexfrP0V4moywhzONkkLmQ3nN20c3BCGekh50z0jDXxnAUp9sJ0X9
vhNpOTH6TvHZ4E+LXA6pZUWUgRSvOX2VbXSoawTEL+1nOGiOc8k1l9yY/h8AbkdiNSjkgmAHL6Mc
H4X507PcBqxLb/BRuV71iWhg19aIdH1lxHmHoIlEBkQ5+AJu56PL62EDYuzo/yZQgXNNLZFTIs6g
uDPOHaNy95m5ifbKavnOg3kEnuQoAouRdm338nBhKbZr0i6jj5TFBH7atB7wHfXnAMcups4syk2H
pO/JCRW4VA9N8q1KkwKU9xlplkOBWoOw/CPNYVITyl3MzdIq5KqHjCx5Bx9oGS2Aof2KST82bCq8
+CbumUx4ShXGq7vbBEC9Vd0czMm6z6ntXL1WWPuNA6Wb7KCGyXtZJaPX6BTfzPnel0+AtnRXe3xT
tg4Xcud5GzwcYSzuIr5hmAMG+NK40uxkCwLCVzd1X9lw0reqyjdsuHnIRiAf8GMTWOCwXlbTJy4x
FXrwzFJSPxlS1hquk2RX1KZt8emBN4+CMrBUbCNp0s1JxniUhwPN51Pwq8YqLYAmsDrGvWXwXvbd
r7ZCeRo3AYUGUua+mpoEIRxjfXNiHQY7tRpgYVpbDlL7gyd47zYzkYwqQouF7qfyOg72SzmfKxVi
bvjF8Aep3NbW/2qXd5wUOU2QdiDhmhFtsylcMwIHh1jxYGHDMsTV5KGjNycbZ43KigC65ecQ/Ylz
tIdZ+MYZ1rgl9K+3WodyecEvHLFqgXLtDIY2HTG+dvM6adoCsWgYA6+YLIzbwgEKepSla4m3jsiL
SvgA/Um1cBkOzU98/O/HCZRd0R904nzky404OsaDOKBd7hXHJb21nJen9tzxKoCilhWAR5pOcwCJ
xmDuYkn33Wnfr8lGz+LLeSB/9JudXbGgRlUevRoCsqJGM/ymYQjeQjgeemknD9semwxOkSmM5NZs
E4MD6Ch33c3iPxKESa9yFB9eYju6L/Bc80jNhr6hchnLG464eY/yL5Sd2eDZGKCQ6JJJ45XGeDR+
IryAOulyRW2ivr2wVaDaBfmOkbcpyQ2AIA9XRdV1mda1vRcpAbS/FvBPykU5tBmZJ96t5xUsosWd
zI78Y5O5aGKpR0+D6QMtdFnfoN6tkDh63v3Gu9ud+ESorTE+7SWyNKcqgocw//rGgHLW2QLX7SQO
js9PicoehKxtP+qbj6VxKUsFDtn1qfQ8SdX5xQJvclLRSJQxNdH1KWb6WD+OJfO96RYHsZa1ED85
7ijgin7ih0L6ECXqLHmPgzz+EUMt9PgW0X+9wR6dnstJtnHYF10wYCRkM3SKH1Af615CT9zZewpp
Sj1PIB5LFBQ898ufNjbeLjyTi9ujJlSV28r7nnikMy3r0b0zBsZTiR0VwupfoxioDx/mQSzRNfbp
OdM1jRrBw32tPnJ9tEQXObzUWMs9+c4TLJDagzHboMdPCqLKMsBeaujmCt0pqWWH+VMmqzbCrX/F
E1voW8fTeHlYqU7BtcBJXoI97RHEXkmhE3MJygoEU3IM8irfjBnkHzqjY+LyKgLa/flS0Ze6BaLm
MQUzqHkVu98WsZU/J88UbHZiWQ3OAIGSiekOi9k4gynKZ0t8mJy/l1akJZ/lo7+gr96Y7Pdtp7t2
9L8zl8eDo0lPxzCaZroh16b2D8R+Xry8KRkbgCbCPnkRMcuSOI0cxb79lBWqj3gB/Ns8qXc36yNR
KZ58AIjxAIIR9wXogTsY0jYtKLMs13XEVkyOOXocJANVH3QBWTseVfWjbvHA4XJA0uHwbV6k/UVs
vSM22NuyInAv6nQ5lG2kUBuDIJcO+ENPMLkGZ/2t/dJeSloHyonVf8dATIkIKJNP65riwdzI6VgZ
EvrU0tqcVoC69GZlkP1nAVKCn+oApd0X8xKVsTm99mMrmbGweJmEnKgnEITgoZ/j31V9ATsxiI3N
hQTPQdhuMv3/f+XSWtkGNBaByiSBQ8Q+w2xNTUlFGGgXMd7InMWP2WK99pBtg0p2wNE/l//epIZm
W8DzT6kkN+QraGhRP84Nch8q+6ThdF5pNmAUnksh976l+2FyvVEewT1jMYS/5dVlo6ZeXQ5JfQZ2
19IrF6No+7NiZ8J/LolTph3j4/g3oJnyTMuSECFSOgRnukvjr3xk6/dKjO2oaNYT7IrzomlITq9q
aOT19eMFnzBHyzEWJ/EpcSAh3EhgleAtQBhjnbljwXQMMO3k71FEr2FUFjZgdMDk8JSrf+qNSfA1
g90oQUAQ5z7pxv6GQurZ4C1/TlCP7EY6c/wTniI1d2jEGIp1H8zDLdW6iQhBNpxQn59HYBCaJ3j1
Oe9QI0UGJKOxNPlNxi83koUt0sXgKHME3wAn/Ge3t5FDTXCvcZvgacPbJ7pqsuJ17maLoEZMBV8Z
oDRtuDo0S9ZRxbp9NOTE+/JAM/waAD1OVxL3b68y9mj5yAaPUgyf4ZiqhUlFt6gIqJIxuzLoDnnX
W8hAsyxwnRb5U4XMjX6DW8hQqhWGmK1ArusChV4T1v6nCdiPfCFwz95/V6v06kh434gwt3WW5ues
vi8rlCB9XwgrjtwkV5Y66Qg/lE5C3VimkqPmYN1hs5SZ+oRbAd7obdOdVIFG9W0wphZWvkljtq/o
PrD2C4RyMisj0WWWDBfoCUGta7ri58pA1w/dVZ3y55uCOUyXnjDnnB5qkA9vRxkOjtUjggOB0CkL
eys52v2Bt7St1Bsit1ZSAW9eJIRXxDvEjYgySau7Q/UnQQYDGnDhg4/Majf5AvHMhCuD4O8by04/
scR18gi94hggCMPZbb+QXtm1PKjEbm/P9mbBKuxXkKTbnATFXjYcs8v6GzZFm0/NiLuUCT2jb1XQ
qPRDJe7J6RO8z/LKBPLxN3ixntcfpKoeoG2oh0dbZsjmkM0ZkRdYAPnelRofFU2Lhjq+rMIMWoHw
YtP9wbqNoh0vsDYnNga973neqDY2VT0nowLAeCicSvbA/Tu5U5qxRVS0wJDWbONWcZeFtSfTovrC
Q5J3YdINpJMM66zV2MGbhHPJ2m+0WxWTTN9Y1Qkj8h0K4zgUlvv0KB1E6QHB5KkCkdn6Eold7HVG
/3IdE1bHwoGMLCWaxzh5olqs2U8jYEjMKUmOHN2YfXRDBZh2iQuv/lkWpdBke/kRv2M3JWjnk5ai
Wv/arY2IHcYRUVlIbw3UIx26QqDe4T1/zX3hjlHf9PCdXNbF0PTmrB9nTM4DqfJ0B/BAQ7XuG5Pz
BR8SrP4suFEJGRztHC1jzC6SzjUwhNCl5fia4tO7WdMvgXvsWLQSyQeJX9AmbIrZImylqwJLj9vD
pXEuegjElUmBr93m0nX2NlKXIcR7LQABFpydXzEsSGI9Wc+RllDbT40/zHnDApQAJe/euIdYy0tp
7yArX/Fl7+YpD3XYptvmVNfd+HlT+zppPSmKcGeByq+H0k25oukbkR0la/v6PKF5ZdkxvTkSOCbR
x//ZpluHwqe9kSDtoZ5o7kddODXpPB63vgGfsjZfYGk6ygJd4zxfui2diuiErZungWPoNi5cQNip
fEjf3YZT5bO5XnXwXIG0e9dVw9zywGI7NskExClK4Hfsi6EjW3rf+ToJMDlKgQJnCH8g4IFw6DIL
cz3YAZkP2OEkaI4C6hYVM6kHcFe5bd6mLiD85n2q+w/y+hyGVGEejdBljjFr/mFuwdhbTPPu61qV
2/JdzazCzgOjHWFX3wK2zq7dFHAQT/wLzfoutlfLDMvqKRPJ6kEdkfjVTqIlTgd+NCJ9BYZTtXUa
+T+s976OEJje2rXJ7eP1KWEEl3tt0wnPXTI0bhOU7ZZdyWpDaLqLVMB3IBSxoljIoyIqIdWb77zv
x5G9cUIim0aOUMM/R/HX+gAS2ggqAkMjnJ16IpKPUUrTY7AR7GG9Y3vZNFjslbLVdVeGhcBYl/LV
IvDIguix/IovjH6cAMPYQdcewuTyWF+hth8UkmUZ3KW9SXVtCq+BkWyw9rmBbqHYqnbbtQC7WJLi
dJXgycLXq8Q+93SA37K8El6SmhJTFgIZ8ia/bUu74DT54Xr98oKHCTvu8UE1oyR2oZs+OGAiv0YG
XsJRUR9DBrYJho4efayj9AeFExyk4GFWO2YYaEVVjUFX1HwyKb5mGzQw09h1EOw1b6bBmZI5824q
72Excr2m7GyLEosQitBQbyOT+EozPEZWkFb5JB5UTJpmv+CFIeryp4nErGRyvCLW88g5b/q4lA94
00/MIuN4pGXW8d+qU2F1qRz7UBTuGYfIm7X+o3YhsAHOWK3THvEVC/HjuMyq/winVDMHkJru3Cwe
d8g97OKfppvMUUtcNSsAHlShpcYa9CnhIBHfH+J6fl29vSPkXfqpDl6fQkXheDf2E/J3wrjBhmIm
RDLP+zTJg9YRzhiNQGTb7nQtalp4qel8C9buWij8OpqJa8JJp6393QQdjig6CLMW2P24gZ2km5ci
suD9qZ2vOzkN8JEEUNMIbh66aEXm2DRdqdKv8ecgeAKbdYk1s2pR2c0XWOZMrE+lg5piffCEeW3a
hS/7Z+ul8HdUxXanVdupcEVMvpmMwNVKR64nv2NFA3uwavcYwDM3iclYlA+YWPQtdjjADSXNWHoX
zwEDLdoRMc3OdLiBnra0+LnEvSyQvgq5cPvRyjqiyGCzXQN1FmyAHZrkI8DRm8cQQ26PKkq6/NSD
F2WOQ6WpEzoota+/Z6QHOoIyddIouQ5hNTJtgJ1D1S/rFj2F1IBN4ONfdMy0t2VsT0ekbQxFAOXK
C+Q0wAAFF0dWli6IWqbZ3Ytg7z1Xjcdx5MUBrtrARPl4+LxbtoGxvTMvw4oLRSpkwLoSsGIQzVh8
V/FKrGmTqfYLur4CL4keDxarkid8q+87EzwxzkyBtaDExihjcF0PeBKmoiKP2plo5NQ778+sKVh7
Q9kPd/ZLfOPjZW/aodp5hKOTcOG3TPFjczj7oDpEIW/wcEEgp28eAniYFXSi6ABODlnvHe1Te3Vy
FFxi11+DljdMHi+aekv1vDumb3jPizn52HbOsVHFvSKk9DE6slrB5UIw6exuXq3nA//zRvZ9axDS
D+70demP8t0ydwuuj3k10j4KKDHPTNUcsj8V/zR1CXPR4R12SYLJPoQQCeHmsUzyDZRRbgQdw35G
l1GWMJmjm/duy/NSuaVAU1Y4QB9zjiaDDFqo7dOTqs2zYeILQg/Y2g3Jv3ngrwoevsBIAHdsPzYZ
PEWpKeK+23DNm7bgKg7xZxXWfeCjScy7bL8L6+AHRPhbI7HCofTRSvUCyd9ILDHWtYYR1cEw9sqE
4D/KHXw/eXDK63dXcL5gvrQ7CH2hPCjoTv9wjif3B5PnJbSrabaRcxXyd/E/IBejQlkW333K81dg
hp2cqeF+hRnKlz7jE5/GyyaUOls9fSJ2OmnzyKEBc1y1QcCr18onHCBEzJsTVFClUdvQCdB4sSBc
gpm0XxuKBCxtAzctsYlzsQDehU+nSeV9eGB64LwHk2rMVeOUUOISMdF8G3N/ae+OQV0S/Bbkqlq2
Lc4YFs68wI/9hMMI3BGpBFDqZp3K+8w4VMl5t/V8dTUmZolKIe//tcsug65L1Devp1l9Ur5+ij1W
WA17/HwzU2u2uWKGIgtvmWtH9Dprz3qkLjt3bAuveErmO9fVXtyHWz5lQYOglq+0wBvxFHKj7hHA
ZkFZbtpbnBDOeg8t5tXplM8eviHMSAD2kuZvhR+MsC1tFdpWGUbKpLuql2KvtszolvX7hpfWNwR0
xQMRiuz0h3EQlSn3id1Sdy4AbGF7ENbhzwOE9ERvC7jVWtpxE2OyH3Bd0UFhwqRwzIg8LblIOBXT
VtNbyPCyGDkNonvskkxVxHvcYgfBAK5nfQGXlHuj0Nkb73GN1/zaGtPjYvDoNH33HG2WBIFa+zaH
lSQ/v07VVEhNiysG9M4Ect6T+eocWpkTIjoLxVyzhcogwa3CLHla98BfeUUVnf0p9najHtynAZDj
GY9bScW+YzuU3YPDvBH9ZrJrAIijbhC45sKo9V1gsZj7wm5ACeXqTY2y4dBOPw8fStJMlOHTm6qC
4FuPOg4nRY5Cd6MBbp22faN1MQRRpj+jt23MgclX/6mooy/Kmj6PpoRXAAWV0wN5VHHM7f+YLXqQ
6yZmVEXot9wjlA0SF2Pap1ae1AmapQMxtQTMEHH0vTtPFdLPbzLFV0QBC4YR/x/S2+TPsq82fFu3
ZhIA+wgJLPnMVvhkoRk4pjEIt0xry1IJkZ6GmdS5nw8IRmOj9KadYVu1T2nRKl4X4ExdBkDNVSar
UvSmjV7PZH2g2fiy1N0ZkHBl68GBzRDMj6l0tX9PVswXgjvLC0keDJ+LfLjq4YnCQhGRJ/dMdfYM
68jYKsYKqa1GY6mRflFLsxtO1c4afFddDitX5f/eTmTxYzjnbrMtx0ocIpLnI/rvZwqJJHFrmDkI
SFVYanpmlcem7JGq81o7cCkkcW/NPtR02fuVxsY+HNUaipqx8qWhRKXe/DLBvsyk3VvLJPFXOsLy
g42Tn/iGIOr3pHczg+d35TyRtziDhclWHdBEY2jSJVIMVbiYH7MchhAyj6l9cFmuPfp9+yAj3AnS
AwdlQqsZyUaVABJLgmIi8dr16wlah55VYD4ARf56tF4gvdj64/y0NAzVTo3KDB3BVaRocR5B2cV3
bIflAxTjVNH/46uhXpHTCuhCRmQWtXsGZM1nof8R7gRlHmXNZ+n6kaQ8w+JuYtfgB5w2JyjDvabg
4bGXmL1ApP2LuiPpk1OTuHArxEo86zLf0Pq67LMI7exNBXhP8cCg4KgzyQTw9vYeo2oCWe3jSrV0
XM50/pLjD/hnd7fwCAnZ34o+L7NZv562p0TitnimXreLMdY8kZBLaXTgJa3BhBF6s2xR4wFL36au
K1ff0MF6ZBzHvq8o7sZH4HIl811lVE946dga4cqA2YgyaUYUw3N3eYTAFu6DwY1HyYld4V1dxZFt
koCTyCWzeI6rOe4KTJRh2sypWXN4bMgDNtuk5I2vU5MuKFACKFEp/nfOkT79g09ofTiFKFGuFXN5
NfvBsCLgTlMIencxfBagNEdnvYJ2DMdR7RAcAaYKwWq56D/MyN+X5KcR8zZrWHWq3IWqxv3Q3h7+
jf+RFappOxBt4cQG5EaUVe8CPs5vXhd4YnNqcQK8vO8V0hzHI0CKIS7j19kVlEk9UEgFOM19PTp5
tSV7WDAPagDCTpPUFrTcWXTyfUHn3Fi0JFmGbo7auyeYXoQCZdF+zgvBGKRKPNSs2llCpoHgQ2g6
kUR+bzx4FmS8D931OTDL9hCrGtB0oYvlgvU9/E+ByQRw2axOYF+PsrShORTqPv1ImIfR/S+b28NZ
fFAslAV+G8c3cFxAub0fTMwV6BufTAjQdIzVmwNuvTqR/3UoJq9YUApTJjp+tiSmyCEE0eHArG7o
t2UIJeiGBGslX1Tj+sgWhRi5qRnkxqrf6mNAG2mopflPmjRUmYsJvJNnRRzQBvVabcpYz03my0wG
0i8MLj2lwUzfEYlJhrGJ9Nq+MbOUt91sR6wi33OprKmfranv8KUIeRJf2q7aj1Z7lP3Jhdr6H+xm
qeIE0oo+9wza2HQ0jIJEVnARh1g48TSC42bEadfOZqysEC6SI7Hnnj1CLuOYP2fzA0dpHMi4W8Jk
HVz/h41L4LqkMJ73uyoyv6xMMAI4hlff6msdJuF16+3WpkhYSjyYQ+6agQfIIXgNzp/LiguSDUWP
u7ueKO4ZMugPaUD1s92K5yGVE6zz5Ep2LV7MuH3Wn6OErlAE4F97OgeqMCWGqNnpG4mNAlCBRZFR
/gqP642kC+SZJQIqhK3DowXBqDLHSn1yOlU+FaVnRib8N7mVFvCAGJvLDNpdFwVNOoq7yxPLUbUi
Fm8FMajcAXo83ffkb3BvOk2S/LKa0Kl6vApVINQWui1tWfewjYZCdpEidw0aUp3zz4p6ycQu8Asq
ATsw1IN8sekzxhj1VUr3YKUBJgwcxO0xFBLn8AFGjKf5ZsKXFRxXMS3WGScEANroQ0AFf2GCzpYY
TMjydCVc8TFaZ+D7H2xj8GQ2FZRsCXTCzw9uMd6Ol2s/UgH38+ve6l9FwGraLunPim19HIDzWg3r
o567unzepKfYWOR4D7j1qOlDVvxd4heE4Jk/tMqYC/Bj0n+MZFs6+Fc12ijRKV5NzAfdYrddg40T
mEpllOy/LYYaxQA0hobZ59ij8NF8ccpXVRMr7Dwj1xhNVv4X0aCtBZbKl6RvdzovXriuVYmRBoUM
oe6/8j9Wy5xvEzvpmOx255eLtzqfwAZEOi9yZ9uPqY23E5HQIX3rD0HpQ7Ne3m7kYtZE3p1pxID4
YiofUsbSV0y7QV5vNCz2AQKiPUZJZAHY9aGH2oZor5XSrc5KQe7M1I/75Gv9+bovy3gTYLM8qQhF
yVplQOs4U4laPhDEYqpKg/aoE9KHEEqf9evxJ8V3wQXT3B2M68oWWFXGqNelS0sBl4fURDKa2pO/
WrbJShNcVvr41GCRbT8HjzskVD2K0kEAIbSD32PYYbXo9XNIe7JNz7VQ+d3QD14CmIKRpMMWECt4
T1hTBMN+tHQaaODrEI1rMDgQ6hZgA0WikA9waxnhFBsVuE5fwgBDD7KGEafssJAz6hXetE6cBIw7
Wc8+yXeluEHA1v/CApfNooN0Z5oJjhsxS4vZEcG1lmGROg+kYtTjUIibyeDmhcMkhd4GEEGpBgqt
6Cs3pzdIIFXpSqXSwuj07qtKtIPNOoGfjaTdrT940Rv7k47aBCQDNQrUlBA+9ikFwEoah2mnGVFk
O1KiSo09uQhGC2v/XviXEqO7GBXgNBKN9bI4p8nWP60BxEaLac41ki0kXH3jazCSo7hm9oCIVBE2
aPhEK9332W5EHK82aCzuiMqF0ei4CpIG4At7pjXU1wjRy1dAlb3WVyD2xtqKZ8GVQe3+zmmN9WH5
ag+xChdlB5yjxaOfXJDy+r8l/dOXtaBAhfyrrbX1hkey+hotbkhk6ZVnJWAe4LrJthtsy1B3WH0X
RU1PPjudE4KAH5gChH0je2Ss6viKM+pAsKipZ03fz/ck3Y8WfHH4VHoARPWldVILnrAyLqbJSoOC
Q8FFkSVmbH6ZakGqBZCOcsq1y5uTASuh436G6MdFDGBtlaFBQZqKuh3VAbVSYF8bHSIIfKNeIsl+
HkmLxYIqqfYNuU5wDwd28L0ya40gBk0J7L+IYRpkU7rntlxGtjuLxLtSyilvrEh82pq1zXdhTaP+
rEwbhN6RqBSAohex6S7zVjfwmBOHbTQwtA4jeAM0gUgEkNLKI6mdFA8Uwg1NTzbI6o/cxGIlrwrF
QISOY03bylGoiqGtD5ZjCEjYTmk+5mxu9NJskmA+BEYx0nCILWDx+TUEJXsf4XHKPVb56/1tHpiY
k0vlv9zKEVY3BG3AJnWOKGuGxv1n14mAGSp5BDanKnFcZfnvhFhD55iqAmbQ2a/RC0D2iADHI+3a
HH5fFlz4TxiVdmbAAf1HVUT/UQdnCOPNt0v9piUMSjOPW9vvYHLbJIVNLP3wWj0fyLybq4Q046ZB
8lFYyEastxNnTymdeW6aVLswOy7NCBBuMYLTEM+H+JAsuEAlIjNDQmE0Ttr8/knHGNz+PhRueZ79
1QtuMs8wrHMY/9y7ajcFo7TWK/hMM6u+sBZU9UNPNrF3vdAN/k8vEhHIC6J8UDO0qE+HfxLhBUkK
YqICyQ/EGvx53ai5Zyn2Qz843nCf+9nQ9Kh1H6Dh5nUz3VfjLxx/+eIDuwn+AhP595wNXmv84plm
vlzYJCwQpIZIS2RCV884T8dIVKxuS2UM5RD2bbroxwH8p7vwLaghyEPuR2Lj+XluQ0Liwvr8QxJZ
ZmUa5bphRbvsbHbeSwlgKAg+Nrnd/IkQGufactUwFue+tdC5U2aIyqLr0mDtuHVeNjvi2O+TwyCL
9yyHOicuf701Fdm512OJWN/qRi6fBrkF8YWl4FolbRB/a9Ub1XN3gtQX+6iAhcLCdxzMIrP6J7DS
gra/0IogbQrB6uG1ZtWpVs6ioTlWjlTUmiiPGrBdUE6S8M22vvxB+IdU/KhcHDcgO1MDUhv6PYpV
FbdaljIdtWIOjHMC/nPa+Vqbqwoyz3wxpE37pLYrBsFyNgB7AVWuUUr3VQhzVQwbQuKf+cWCo9go
/4LTPrUjN5HrrEXQVaGRzC2SDg+o1W1kYIThRrjxboG6OmbVHKFEj7iAl9t9dwYr97leWuk0VMxg
eI0GqhEbNIG3LhNo4UbeFl6PuIWyNpf4KSO/LkvegFN6+lO3DjksHkcJJl861K1NSp3vs9g850ZL
Yl2SjCtEp6FeNlss50xjXEztIpTUttF34XGwmYSvKhJ4R9GCZfeJ9oT2LpxFXPPTKQSz4ZOGHnwV
K8Gt/z61XFkXx7Bji90aSb1hCDkzttYdShzrs5ebpz6d+QQcto2/IbDNRK73NQau/E3tTufFwpbz
wnHIP28/hMCXVDbWnB68N7Ubfaw02MPtiCXcqWxzMUrVUXzIy6rvG1Fp8S2U06fRG/mYtmDlbo9N
J6Tj4gA/rheJxw+P+Y+1f6weNpNn7L9DSvJ/MwT65t7XOfeYA3A+1RgpTnZt13Ms8OCWCuNaSDto
wWEgOcdJLSjbHQ5PT+b7giJcI9yMVyunEX1HTphoveodkikhnyO9pie9h+5dCSf8TRvn+cPM2lua
yHZe2E4k/BDMDJNSQLuUgOlZRmFFRbfdLDqsd/+lqjsTCjPeUPBeC+OSzRJiMvriMURkQPvL2wOs
vwGUd0GxXO/WXLHvn2F4GEWvnSjIXVyJaKnUSIK1khdW7jhce47Q3bkMJCpiGGeEkihY8GdyNVUP
+zG7wBqLWZjXxIyR+3WWaKFfs+99ca1iTqrTaXlCTuIqRbR2ne7KXpLdjsN8Y2pPKvZ8GZQMxBMy
CgT+er53xZqK+YuDgQxa8ADIJ+UgPE1/oQT88ViuUd7c2xN9A+RqaPO75Q5YWPjboy849QCk5dHP
r+dLbvWFogEt5PGluiw+fR6lG8waZCrHEC2gRHqprnqKwQIfHuJEfU8ZYfYpOSM0g3SInrjbDG2n
IduQods9/+8wBsWWsQe33yb8KF4xtiSsy0X4QHquy+BUEW5SutSJ/nO3nYpiI63O8jc5WMt2od0W
/yIXL8WSF+nbnmvWbT9+HZb9rrUvUQUPbxU4nKnqlbHkNM8NdatIymO1LVch1extpyYTP/rPLTkb
3pzg6507zVKHh0froRLawQVkx5U+ZbHCIP68Ma6MnNeAq6l2Oge9DwzPIvCLL2LT+MdCq7hWjF9d
A3JzE+dk7+HNvEGP+BnE2+1BboZ6Ou1rvcfZAsUfXaujv4KYPSjlWzEEJYfIi7FdJEwoAl/bzBz0
V2P8HrMQBSyTXJX8i3ep5spfromPN6Gad/TJZGBJjqdUcxmcT1EMDp5bTZsULQijAgVKWUxM5BDk
VsS9PagSOoPz2T9oJu2cppP4hlWtOHh5PRlgx9rCjjZ8Hs218xJ/uXRdrdzvq9ruhQlO03ew+8sl
dIwpdoqWFsnq/BMY1TFtgA+8BzqS5rTTKH0+yJGpSniZZbxSCdQoz0A9fJ2C6AJV8Qq43ZvtpofN
Lifef0rkIhajJUmzv7Cb//trDrpy4gINeyKclRnR4ZpwHd9xSeJFYG1vRt5b6aBAtNUJha4eYI0M
by+JikN9U3WPF+LPT8uHbR61ZUsI7KX8NcAYfoq24To4oLH6yrlZvGrwDE/D3TNtJLWj70bFh7kb
th6UZOfLXqAGTMhEJLHviBIib/5oFmQk9TiP9wsMqibbJmKA9Y6d4Nvpgd7qgDfdO2tMsiTbPlGU
1ZGh31fHsML6THsOIUwpladAhy9tvSXQoKYqo53UyNf7UF9EtGzd9bpYHvBmEBZlxtFhKo6svbPD
k9G54+EzrJGdUSfkcVEnPPz5KibUkdDeiHKLXVRdNb6THmHNUn+lUVajPckbuRZgh6dqaF6o4hm8
CeVGp8OapR0Q+79VeBbVaA06zMZy+khur8g0ayBDVKkq+AL9mtKXWpy5UiHrFOQ5X6a/PAScer1K
lr6rvwpH3NCh8DA0ujHnCEAJcvQFC15I1Z6dVu+LjgAjr9smk8GZr8gxFNFe+xvadS6P3fW4KGDA
Ig3gInCbLl6gkAQFWH1nG1l/V9l7RYpOvp6zR/vnNLJcgbd2djMusfy/cjUjAqlN0fqDZjN4dvIJ
OgusyIMzeSnoCq/V5Oc+rtEkvCgH5AGlfSH7mFAZjgxw4otRQW4DE5UxDrlLveUrGn8w5Coeg1dI
gnPfVxNADeMYlAROXylQ3TLCN+FBkhfCGbxETFCYg0fWRvFwdkKdTNQqs3ezojOQs5Pwu4S8QYZ9
tozrytPdnpojtvVBLFgs5oiwMU/w/uPrp3IZj/4EGea5sPcp7oEAJogfD8xK6/bXIGSW17CUOzXm
bEeVpyyGwEsGvjEsPygfshnpoJQtuugPqenY0/gxShkJT1pQQNLfngSYFKQxMWmOk+vzcfHEmkcz
sTdYbagldjZj3oyYpEoRSUEAbQWBV9x2f8MTlopz++tv2uvMqKqR7nfhlhreLvcKK55kkK7COqn5
K+imL1waK+Yaty23xW0j6ucoiWu1j61dKr20WQry76IWWkXR8ZGjrwzGpa1TqaMtY3/yrbY0R8VX
p4HQAGMbOJC4oPl2oFjL8jf0gBE6GFI3y4YjrP5e7Igjn63BYy1ikHFQUcY9Rn88T/t0efzvBWtc
CdNGpVe/YeTNO5accxhwGkph6GeF4J/Vsy85vUir3h44MAjfoKFJl219Lp/+/yhQsa3vQiJ1OVP9
DQwJP6mzh3NXRd9G/gjC+D/CAx775d5nbOwIziAB44Urdv+BbjrLpfkUsLfCy8zBxaZ4JiY6STSc
dVRpJW5wFeMvx9jfJ36fKAXXQqCPPmVqGxv4bbEMhmwJTcXt7ayrYoKg/zN45C9PmHWyObHQcnQv
RM3cp3mH1XJipp5lXrV2OasowdqRhZ/mqlrMMsvHSKdj+vNvhLEBVkwiRhAV6QuSbKnWsRrJQQuH
UxXsy6Rj1Wj6U8QKK6HBXUcmAaWVCCQnTcXK8b8svS1cRwXNpoEhNvOzLuMddKIRDsmDYA2ANCmY
fljeiEu/xRPxtYFJHo/sVdOtCzm1c5jiie6gO1P/WjVoCsfa1993XyFBZcnCuugdDcNwK5kID+uY
JCp3ub6vDPbL49fxTt1ioj6plRLs66mS3dkO5zY565JKQOwrTIB+KmiE5CIoYOJtAU7IqojCvS3e
IvS28AYMVob5LBfjWtiY/6gyAfh8JykODrD5k00I8M2PBf88VHEvuMMfUSHgnL1UH4zQRLUFZfvL
fcudGPoSMCDP7sswwzc+z9dgsYv86P5kkqcHCndYPmSoHE3VfsjH0nvHi2cqyjk4HQQ+qTloXPz2
fB4b91HyuYxAvDkoPAKACkylQ6vSCU9M+DlGkItfVI3o5gCSHjgepN70O01RIcRgVV6MtUd0GVz2
FYV2lz+tYgHf9UtwdDEyQoqVFfQw1lJVtjNqY+SMF/GTLFfgQySdicBDkRTnyFxaimV3OqEnbPmG
bUOVren3T0l4iJPIiqLdXXdJLkuP8Pl0dVCPBZKmzKdGtXdUeJxNO4vWrqL1RWj7Y5G+iRKiodqt
2EEP1tXPZ5wJm4L3BTOhIwm+545Xf0xERTYYVZjDMyPU7jVHbsIcMIu62bW79/pORcXQuOdaj4bu
7RRdJzJJKDOukOarWYOj/eIyB6A1WdDD9YBt93cJIN2jsYo/tcFl2l0WkGIlhwR1FBvvsLwgKOt1
L+fyESbRPawnsU9DtkoKKBl1+Hb0Gshmvnw+AgtIYpmY+v56Hmmxl8q78OoCaqBxoAORQADWJpw0
l2C3ZZ+G/cBBAuAg7Rk57VZbyaJwfpI+bwNn2YXsrvDdZ12GxRpHh9CFwNrbuSizK2In/Nd9n09l
Su9xiViF8YR9DtA9kqbEddYhfJT1n3zL5NKJekpRSRrE4Nw61DEm4RXOlqk3lyYzJ7zsJVQ/a9HQ
J3wJ/mbIVRCAYQ/IkmXaUGynMO/a6KljhJ7jT5e8EoQtRFBw7JFc67aVHsgszkhjWfOmstQg1JxD
uHY5xHRYOteVKvtvUnjqt4biSZaX5FCnSqEb4ZOI6/x4zbXrUH1u9/fhRJU+lQbEy+TgPj4CoL2z
woTEf3Pe5bieJ2+KOjEMprNaAYpDbtKjYd+mx97VMHuANwjwYuvfQFLOezihxyL3LDoy7Vpr610M
3yR/cw9aFqcAVjkcSOD6BxSsIz08/Ok2X7+4eMPKUbJDJtSYGrd3L0WCiP68yLThcUM6Xpk8z0IQ
fGkmH7QVdifssLbgKv+TKMI2M62W7LfIGjNcZdORJkLK0wDSOeGO1U0vJzxyCToXsqZ2gmkyKm6y
dXja6aHJC/AjQmpmKB/8G05rO5ZRfwrI7uBPyxZETqZ9IBR0EPiFt9qutcEJoeG020SKohiKHOKQ
ctPkD2NLUsvPhNTmRhI9+y4VjBqYKd+9w51fQvN+bLKOl0da2sQSpAVtb2ygbjvKIR1FVasLlHi5
Whgw5GYGdYnOJpKClQLqjZlXDEn12j1sNK2v0mgx4qP1uBBMRm24Odz1zNdK7rqMAqkSLo78bi2l
ApiZfv7UHdM1Eh9Nn+WDqjudE/KsM5YhGIx1RJH1KIs89mID5iZcrRXh4VOXbztdwcwAuP+5t29r
WYY6FO8ObJiDXgHluDsXxcEB/uqlb6SFSl8mOZT4B9KpiwIlJiPbcSnCMQRErcPSkyy9nE3yTX/0
eM0CS1MRnap7ZPiJtbQw0YTgl8A0nh4qSuxX7l4wG11Gaa8v8812kos2ymbrIahVjrMhZV5butiO
isOzU+iRJMos48muZYMTjL+VLf9HjxXcyzOtSloXPkSQCH/tE42PKKoaq18CZslcFFqZ+VByUMSh
jwX60ALt8JpGKfWl12Y1kKTVRcegGk+Fbh5txiGUexkBpULm6YJIJ/yh6MzMK172O/YMIwtZGnvW
ymAfoByJ4sNHNdgl/w9k00lYjqN66cVcdvGluyXeAFo2cg9I+drHW6VLA6V/y+EIXiANLgRyIUZU
HzfoUJJqdhk3dmVaf7ITPU+avbjnjmhgYFxTYrjxoHxJJknoltC9si9Eke0xnQ5YxxHUZ+cltPQB
W8ogjCfWMZhyGvRrzgsFauMhSqmnfOjAzTopAyBYZ9h8SVojkZYd/tM6/FtMMs5ajKi7UUiNRsMf
F968FACDwteW+KNQGXueQxuP2P4F6aoPasKiHXcjo2cs21ZlenTkMMPCKyvEdAcERxPs9ttscHt0
DixTlUhoXG8lbcP4iuxWbvoiIUgRBXeKGv/itCGY/CFhJlJ6LyXy6nrhGNIqq9xYOkEITfRUdHgp
Jw1YeiiNwfqHuF2lId9F4i5UtOchryEU8gM26cJ+r9UKTU1Ua+/W43CxnqpU0jKv+oR5bKZa4+Jq
WnK/tITMs9IwKNZ/26r9v0PaaEEAJvWeiiMNA5YyUdJO2z4CSKPqBr3ThheBLYf94OOuWqTL9D0a
A8GspCDphcJr51S+dPo1xYh0NRYAd+o+MffMahzbQzvNmtMNxbjEWLHd1qo8qfUdaDbPz9msr+3V
eu4mZPuPnJfPWDoDASMe+Cpq7oRLeQJz3UDKe2cnMQF7Hiix3hz9dplf968iXXsjU/ua6x+YCOO7
mh1/igCJPvOQfqsokPOaRM/3BxlD+g9A4nW9QR+bKhELBg2H0tPYdHQq6UhB2e3pRXub+ObgBC5E
Eojf4hgXbMBfBT7NOA2s4NS3zBztJmxw8aGBa1pDnDt0uoEooZpJ8vgNb9fim6amqOeH2nzO40m4
JZPi4f+ecHRNb/D0wN94/PUhpFesRgWHZ/xwh3jMfak8CzYc4FpfMSUv7tzNIKC2VtE5SjYVWOcX
wDzKvaOZ2AZ5TG89DaYdvNTWhs7t6C6395pphPfCSowbncixlINYD4FGetyDNsqc3vH7dLEcgeww
X49qXGssBeBUlwU4WHaqVg+zyKQzfRUHLbM9lLW0JW2Jmyrh4SD1XyZyQO0gGfUOmLrjv9rvugpz
UUl/U+14HNzuDtUXubyqSz3NuUGsJKK+XMl50d3MkBtXPyijgh5h3GBVQJXeehcUzNFPpeVVeYnZ
5WwEmNddUam/HJHJ/flazoCbFczwHEjrEv2NYklch42J3jkLFde54Ac5IJMRmDE/k+THFXNS2F++
OtBRxdtI0+I/bsgZdLskAMkdrVoRu33ZaQ3hbepB8GS/ssqz08iLQ+mHq5b676bbghhMI5DaOyxv
cuMb315Gchn7jorxCfB/2xReKdcRYlj7EgMF6RSOGlnwhX4HQh3A4bI0/t8KfVqHCDdoEtaegKYf
sx+PypOaGH0/CXwtxFyjdRfGd9Eb+7U+VD15d9a5M7iIlQ30J7nq329NW67uZEhShTTgDGTG0yGj
4pJ8xecvZI/J8H4re5B+K06FM3o8FpPxx1gAYvRDibaU2HaQd/Vo3HOwnYNFf13yzhM58iuL4YaE
ogYXKaNBeWQ1HZ8yt8pVBNfGgB1TkXFKXPDwJoqEX0BpyhvaMXjahlXoyJDJUm+pV5Xl8Wlx4NzI
9/+WbOIlS1EKzY1B3uxwkoJSJgOmoYZGlD4HGcVz8Jb0oUBCZb9tkzg50gH5cdxGqg/MIcqhTtUe
S1urDCWpBVdm2s+ayRKCFSoYRDeS/E96Ri29rViIFe5CIATceeWQXws1vmeUqNLLf0ChRutm9GDi
5g0F1OSSIriLLulGn5t/qpeTm7JLrj6AtSPGj1nZIzLQEGX5939Tym6UASqfvJ/Ide/vEX7MxWnb
7sEAyNIePlmdik7eUIB4ef3XfqAku0V+nlje0vz/GcMD+FRKgAXCYTUj4+iXDQ4k6cHYCBuZBfhd
7wSEtaa/vFR0jk4xlWprIBK7+w1JHHL+yg+HGyFKtg6ayIa/9jaNaIH7wQeiW3U8t37XqBy6+yZY
dwTUaZgVP1i8r+Tn8JWLnOm37AGDTvWFKVRfXTl+TXDhtmLHUo0LcIwiDbonuCEY8YVCNJZ557qU
Dqcsn48AUaqzJpzux/LJlVH67Ogj/eSTGPqVv96kRdFTyjCQfcT49N9nn9XtLfkSbHNZb4Mi1Ub6
Ac93DC7pYMAnQ3AsNUYsEzyQPEfYoebCZM6t8stE0mH4NsSRKfNj+FqSTaDDz+r4+3Xd7DyrTlQQ
Kzat5htaXzLo5wxOcpKAeJBNOPCMiu92bf9aqB+ZgX2m8qVJ+CLad58PMxbkL4A97DIDmWjsmt+j
PsYnpp8671f0mBXVZMPzSY3NgQE+4R4C5SBO8m09CrnzZ0lsEkahHg0tnftgnE7Q/JiGwwxburbg
G/1oarqy+n08t2/l3ojS3M7+EaUgnFI75+pJhS5YDXnBzU981mVMwycL8RuGR7dJ8BmBMtOyWiMd
yQ9fefA2+KwYXSTFUGwAaBFx8f5wlfqCMGW5saerCrdkDJ+95MiaQbG9Ng1AlHI+EbGBSyx1iIcy
81AaBCXjDhiCEF2l94suplKVRKxopSnwrQBiutgpmufGYyjAtTcPVD+0kPnUOz6ORYAJjhW638xM
z3ixFj8SPJjw6+D3g2xMto+7vLIietFRnRJS4R2vsh3CJa/pADe0DRph6DHaqylFuuD0VvX7YhDA
2guABns9WSLql9szznP7Avwto0RElzfUau/cAL55+qH3VPtq8IRcNBLXzC9IKF3xl8Qgmu7Z/H/P
b8Lqz1uhDL0eW1pNU+9ONY4/AwqILDM7AasPxBHKTIT603GEWe3/ztM/L4VLFeUlnCe7VQAGT4bf
ikV1DPhHcUfSSfNXI9BOwHm4uwaXnVZTl2164HcZ7jaQBq1DdQUtiBg4bE3Wiaq6a1ZJEX/l4Qw1
p6NZK/XRcSsU3x9Vffi72hiX9DpPsKrJE1W4zMYszWvE6jRpU4gMFWMl/LeZK6Sx5Eu6u+WtP4F7
6qvAtjzfDxKe3JWP305yZRUAJV+ygrAp9F5UVF2EhXE53VSLQfmGH+APiySr8MatMLK1QoFYIchI
YZuMe2fJVGXEYcodx6HJAMYdzz/sXx9wMhFwQz7O82fh79y84+09L+PlMX72P7Ms+J8c/caLZmgB
aAfOYto9d91qtkNtPh250astABJLn3VmHJ4G2+psTALNWFgmT18/5h2tjFln0cBQOZ7Jc/R1LH3k
AWTday76NdbRpSzBfjyUNfdK8iqAXvNQ9/RHOHC2Qg8bzY9rM8oET39aTKnGOk2aTvgCAQkR0J2k
cpOswZQbYCI/xz9jRFUrEmCqFKDm83DnKXa9+p/0eizIMLhHVf+kyT+HaBHUa9N69XA9UIbkmEH0
pLnefp7nW3iieCnfk0AxIHoaD2zvIZc+Qmeiwan+vOjmibXLFxPQbMmqGGGTi9Hx7jvAhgz96++R
g2vfsrBuF35MS+k3QsZyCmNtA8ja2ZwC6sXkTPQaSSd21ghY5VB7c4FvAtVQI1tid9WxRyfnTLkf
THF4M0gWRpD0lLdunjclbj7BausxF9Vsef2flUcqslAAEgAPDwRbZLRdVJ9mBHVhIPZm2d81UqrE
lfsg63TZoEUJ9riYbendU0gXE6OSTyLpeo2iBUIYHTcr/kGvZJp1Xofdz5t2eK/t4sjw0UXxwccf
A0GPYAjQ+ZCifdRBQdgQBe97hWsKr2A2zifl6LeFZ+muZONbeenpW6m4s/7rY3JaRuGj0GSkXia2
6bfZ+yZUM+LILD0d0XFTr8q6R6r9cHapHcgkv5vsyqysKjSCn/yLcCIIHZ0lGQEpt1q2Gx+1hivL
JDswmaOzwR42XmK/C5C1d1R/DSJGT1z7aftatGJutfyxZEJbNu54NaUD4uArTJKtB9EJcIIBUVPo
ytcS4aqB8DstctWcPzfZobWLovv008WirfZu9pH/JVbrGPkk9/BkcEveUXyvhBYArNXCWydwcbaT
Upr3/n0BAb1QQzzFh+ssQFt27PRnaFnE2Zl9nJPpIT/fdYRrBFFU2omkcrxRdeKSR4yTQrNXzXcz
GXIsflm35Ht04e7jm8Ji7qWuU9yrBr2YRdBej5wqFuibXebD4a2A2aAo868KO0XjkIiZH6o/nwit
zdVCtQ22Db6QVA+JyZ5YZMjheOiqtZUj1K5w4hFh2lSNto6Q6z6dlXe7SQizSjZ4Tp1Io/bXmR6j
vW9gyjaAx3nLkFap436mHFLT8dBrm25l+BCeNXJTMXleJvNo1/XU3z3atTz05CwX8YfqqU9JPw8F
t28gnwyJmES8eWpj8cOShDXEsAJkBQbe58zWa8TOcDRZujzSTXJASar9vMTmMKdLcm/xZc9GekvG
yESzlx5bFSrdnD1+PCpIUcpb30P0S0kFB/p7JWFdjRp01MKCXeb7+RYP3ERsNZDMia9DDeIH/705
9jLEtI3BGxQKfZMXXsiBZZ4QUw2YIEM3J6Xety4qHXIXoLe7w39hFR3Sv/UTr2dcz2/Z7gslBb5l
jZD5Z5J1AtfHTavwhMTvu4fwre16GS0mWk7ezHF76x2Kfr04eyh6M7JZ3l8+w6Eoelqjn6XL4/l4
nZMVA0mD42V61Qk1aqHcLRFmao9fkylvgQlEDsC4GsrwJ2jbPQ+2UjC2eecsXf+MLjdqw7cn7UDd
qmHsQ49FyXX4UMuFb8OEnB9dLknhEldUzwTUiq4cZrXZZI1ZFPT7wyVf/y8tviqNYwxY6hJsu3Mc
SwmHvZMw2lV0+f/u3e7/FdA11vONilAaavrL3H6p+VPm9tirW8yVFWooil9Rw/zYVhI10yJ9V2qj
UobgFwgQDD6hzCYfGeVw2uqB0zd3EKcn6SjOlzXctSEdG/cQC3drUaT1SZdn+ar0iFHNTKRL7L0J
8KLD5Nt+HF1defWPd6etA7WvsN8MMILUssmEZSUPJW7fru4qBrQ1/mSwo292imb1wGh4bQ6270Ug
zgBTgMVYT1urUYJIttouTVU5opEiJ8p//dc7JIbop4pdkGNntLmzXhcsnNy4qE9RQtaCeEq5riLM
3SA2tTzC0GVCQBmSJhATwfIfuSFgFLz8Cp9ukLhZBcDssBDqat3x+/Yh25/yjCvF0U0oajyMG/RG
ekyPLiEFZHHRiCRkyP2iCCwt+EemMAjODDHy2WNWe83WLUe3tEC+JNIE5vQQLInbXXcwhSRfdM6m
7gi2GzK/tdFAMBvUlXfWS9cikFnvkfs2N1usMOgP/c2DVOKlpmHbLQfOQCb8fN16NTvya+1W9rU7
W8cytHZtBavFfEqAp051ly9sIXcHOwOdltbP/LpjOMOnpsmwVTDiqXLVw+4HrOFadVYUR1ogb/gO
kCm+tdyid0rG+Uzo1LHzj+58zJR/D63oMX7jAYosSdJVt0/8NsUJxJZokknQV9P9pZoyUJgjXoXs
rwGwZB/HGN3hQ/2U8CGcUUGo3vZXtvblRs3q+N7fr4PvPqzApaRGED6KJ0XKVem1GZ2lNZynFhhw
1hufnJYH2xDzr4tQYYlxpOZCCYohmltq9Wp3fYKoJLKBqhLDt018oTvnicP+kUXdtM1EC1Ob7VAO
nbxKibqqUtsNdzjwVBuug1YeRoZwskxhumQqx0KhUA/iLUAq6UnrNBlEV2csSJ3Czux6jho1X1Zv
vdO7TbEHLiUZmjMEn3D42jXmU5UHcHiVXO7NBfFoTtNvj56tklkvrnCgP4hOjSK935FbUbLDdzBg
emXWF0Z9b69J5/tNgfb6IGwZFscXyUGj7W4Rg611lveQE1vepkGHO1bm3z4JS7y0cxOpRhEY2Wn9
qTO9P5yib9EqUI7LsdYpBsDlzdmKDGwwKuN6wOmK3ZRukIOsouQfSSPvG/mib/LD7MUGBkKU8bFY
123h1jhTsUvN6DMJAhzn7HXxV5rOO7+QPKZEkyw1BEEcj5LUSg8weRV1CfqOTRDq/fkMT82KIHux
pzNaZJcRcVUe1/xuYqzmCPUY9iOgyFE8nCdng3sH94Xi0UTWlFzIKWITcYZeIr3amX1dQZtlCRyy
NiUwtqV1iBu2UGxUJACcQFaca0UvMjg/dh3RTmnrOUULlfh0tEXSfrVHh9QBEtSQ5MHlPqdfhWe7
nCuTTDtvoYHulE1QwbbVAiUAW0V94pFfOz/P9wozZ1vDwINZXx90QINGpXCYcPk9PnJgFc3mNtVR
lp7QS4jLanfBsndywd5s+LAaXq1oI7xhlBQd2cf/7W7IImOGc6QNQduB9dZkBPArrBLsDiznHZ8C
YvgVoWZEL8mS+vD5x8H/VMtDIOrVPTfsNruYmQ7yObi/t1MtzGH/kqLxrYRFRZgoA8Xh5H6/7eJ8
qoBDcQvJkrSd5apsGkE2u+gM72fDdn1/GxWlb1WpzAN7k43Wju4837uMOp7OeX8EyZdr7mqI6hfz
5Ofd8KMxlMsvjWa7rPP/4jgzBrefBGGSYwxaXQ9eP6xcPLn6/rV0mGu8GlDHmfUzviLPtixJex/3
56bGqQyqv2EZZCNJsRt6ve81i73Rt/1Wv0napy5Yvg6B/DSwWYrsp6/uR5hit2ryn0mhxQdlPekw
N561mvyGFj1bPSJwIb82bkjj67jAq1SRLKHPgTZky6y4v0tRvgM60lv3rQrOmGQyK6ms2ytSMakh
3d0fX1QkE2SqLjJLoQqJt2QjmgadTLdbcXr7NT2OcJI0GAcREjAawkl7E4xR4+VJdSlgTdfGPlGb
7D/mXqgFNzeYEWmXjSq0q1XkxqmLr4DW/RUg0yIVk+3omdcvmWE7sqJGkRhc1U3Ca6LIGekV3rLB
YAEKJwZjbdml+OPLgvtNZds+LUaIamhjs9l8GnUsQsISe40kr23jZ7z/ORR2ZgoKNQbINS2Y6B25
fQVME5Lnu/xZWHgAU0uhZdKjPCW31K2B3bBhcD7Z55HnHkHuzp7QNcme534HO6nBs/TdOJVBjuwB
+Cagf9azV3wij3bvsWQtw5D2JxQsdIJ6vupdzuxlFf7SsklHPCiQzIdx2Lm5jgg/Hsjzvh2ldT8H
K9dLIuIfDOpRjfDSpzQTmWPjl1yBNZn6Uyjayjj88FVUHeEwTaQKIJVug1w2rGmmHcrdToeU3cZh
3uCRIRi+xpL0xxoZapzXPWwRRj/nGfc2yGce1wTLUux6T0xVWRJo8BpFIy7wnTSBQ0knb6A6W4NN
4y+3stXjEBRVdD5jQTUymDhrHtALs/CqavugRPushJ4wcHlEkC5xSg0RJXQG9iTQlALjWbN8MgNo
b75FKVoXeg4uPDmoWIP2apfnigOrY2R+kgyExh8ZWV2GOM4qxfVnOkoxaA1LE9iExrhwzUByAU4z
CipY4KiBZzEVx5K5vQdKmRAN+qO6EvvEwD5d5LCkRKGf4KLWR2i6Mx7A1ACQBIIQ66oHrjSSTyy2
rCD26oepjcGPV1ie+/l6JX+MATFt0fE6XGCn+m4Vll6JE/jicw4k0iFOVnKgxT5lrvm5BPLn+PqO
nssrJkBO13mlzYc3zL+alAK3SrhCiASMCHt5eEr0fYYA3SuE2LqJAcYGm4gSMVkELeEwCCwkL1UC
1QnEhiLGB33WUTRC0UC7kV0zn33e68IFSoajW3phXKuAErg/mNGEoJfI12QGwaXKu2sIwmZoBq6+
g6ZN6S/azegdmKQShjc4e5tWKixo81kbXCSqqQu3Jbq8WqQiw+CDrlcizrHzv3WXIxDUD0Ngx8LD
L/D5v7x4LuzLPxR40aqLNBBU0WKZ3/8kblx+IKsH1el8Hz5X1yd3qcN9pHzeGc4iswHcftUdFhNt
pd+4y51GO/T7nvOgs8T6Di7Wp9VPp+brcRj81x/fHlasH6LnF1LQxY0gdOOtem059cQBZ/AOeo5W
RudfFMcoPt89Hq7V5+HAZpW+DpPin4Aqab9Ynf5IwX32U5SkpYH3GRd2JG99fqzoAJJg20Yn9vPT
BWWXbspgDSe+1mzSNyB92ahNGvWrHLvcKzSW3YajnF8PgCqGQjvYzdWODV4mxxy1ECUfYELv/xDx
uLldv8kVog3LUcjb0fVnbntBxlxAOLd3bxa26kTaYBdiZHKO2RoODAmK3MvbIxARcW5xwF3roEHO
QlM6O3JWo/E9H5cFOmAxA2OWUy4Juu8hoSf/Vf7QVsBXEiQULovVkAfH2gYpW8ou1VRFWtiocpTh
2uo9vaZpPfsUTnoFWL2zpdzGeAwjCELKfaGQcB1ltvqMTRtCPJ00c/b6WPo8h0SYnGWHbnC+JSpn
9dsduW5Mn8MXl2nNMDbYtmGwgrG4vaitEzS66j5xhoPjrc40ndPSqOlr1snQ+maYwo6VhI2CWSen
C42hhrtUN8qcPAOAh7ZcKtaUP0JLUrEb/pDXp6XWk21M1ig1K5qHI9zqXmev5MFeL9YVswPuGfbK
c+f/LNx5bknQDaDmsvSiDNffo8FZ6CI//s4q5ey081jJMJDzPmNxetukbzdC+qWK53jQ+pRX3R6l
LsfUxJaUZjmwcaiFgNhH3gYFJTKMVK2YN8V5N8Ix44REPJDxjbKQjp0+To0y3AKQsfO93Dhe6664
wR6M/iS/82/vY5Q2aUzbogdQni5jDMW4LJuRPmjmlVvyc17L6N2CEYmk2aO3WEh6Q309+4/yxpfR
cs3aExtvxY9435asemtWY+ZdRu7Jywm8DlXasvBOtKEtAs2rx57nzaqpbxN2wVzZLWfqv+g6B0uL
dLDzSk5A6G83epdCUCnv2bjC3iG1u65gJ5Ti+8YKUPqHXJyggSeEtPIq808cU0erkq/RUeri0fJn
jBe9rzIbhSVSXcCxULtgK+E5K6GM5LvJMqt8rRWu6Iwm73EcA8NT7D6OTwulRumF7DgfYhIBSDQu
DUWsTkQjboGK5tPjW1voU2q5cDkS0yUhNPhyzWROurevDs1Ql3hdi2i1Zn1wuQ4zPg/UJuGj54f4
cSUxrirEDC3RQrfowVmsPxxNlMl6Z33gNA5FoPbW6pMAr/V9BvR1eCc/1XFPi1tnWHnqgvj1hgDn
l5/hz/9jUXNsl4m1QbzJy+OgbyQbsV1U8mriWBIpT7dFlu/5+uC1+YgbByGpjIWyPUxsxAD2ioLN
aG8Uer2QYma5J9a7VF3XXdGWgiTgUSnICdXdKttBGzT0bdlgkLsFdrrCozAIgcs7thWnB2lG7Heu
REaOL8OKP8ctCK6P9Qq2RKjkFyOJXhlqhBC6a1sO4z5X4vXMdTJO7ktG7Qm6Q53g/9BY63SErERW
NPldD1dhCjXbqtNfHg3uaCtapWy8SyMPsTxu/ixXiB8rh6TuaNDJD7DLtTnRiLAI1lIXUOMMLzDx
jQVI/9P4ANizrizSbQOOA820rxFgne6osw8awPpf9rCpQMzOxEkDwsr04I+mG86XJ+bUrjQCrhxY
4BXtCxgbB+sk9WbDe1KTff7QS1QwOjzf6YR6oSdskXNn85EH5mBo0bYTDxqj7sK7VeyJUeY5EDtc
Cdvt8s3exurpcskW6qdTWegW5ZSxQTczNvCljMHtiCdaDKeq009eYW11JUXKGpnDZzy8ncaLvohQ
RFANpTPPkH11oLcgErNXXoFplVNVsez1sNr42MQ/9jtkBELIT73E0SHVUNZv0LMbTuiYL/PqbQ4o
/vnPPTfnMM4hg2Y5vopURNt3YP1d18+CDVsqC281d7p97d0fV/4KaVh73fNN5068BkcmiS0PE1lV
li/7+4HvT08XE9cP4TdAtCpi17WyrUd7tgypSLYWNAwRjSgnr6WpkBvjWKmP60u6BvcDMRM2FWrz
OHQPHPhQPFk+x6wRSy8j9hDy5fzgrquCxDAm5FmW5uu4FJS9dhl7W7rUkbZnPta9cl3tgZat74MX
p8DWnjkVLwkkHwcmig0tQjUlvJLhLUSgFnApxw0wyMRDippGqo1Ir1LXL+fHjtEqJspNfu8yVNmo
cDOzCAnN3MzVOvgyIG3brZICcuWyYOFGn2kUftqQtV+oECAkeNv4uChAxAmGft4H2Vk7KxgbLteQ
xcpEINjcP44hb9OnUwPI87YqzE3MtvM7FjI0KhnYaGQNyFdM2raXOPHsH6uKwmMfMoWULHKpnR6t
CFMjByG0OD6UdTX0cC+tPoNWkXqz2e1+D34d7OBTIHETZ0j5WZ5anHcqZVC/qZJVVNWujOHm+5o5
mcd11O2elyGWpDKioYEgllXavGuhrStJOC5cPr8Fyke3C/Nll7RevL89GuTE1nbW+YJsTOx5CsoT
bQsogKUbZM137jyO/vQoPz+VNfD0CzYtV3USQRYDxxY65Rs/swxP9ycG4sHIG0xTqHbIdEtfqk7f
9sEOeV0Rni1p4qJxen4Smj8+mPliedsUdNKubnr1+UkZWsbt/wV7I867W6wx0mXtIKO2M8EeVdXe
XNT2VBnTyBHCgoBJdyzUwHxSIfKTHFEkje+N5WbiQLPRwzEMDnaYbJG+IZl5Hgzgzw58nsP4dUEf
HO2ErvYFPK7B4PH54Mt5uH0X9b+FNBogLHRbvTPxol3lYCeFjbcj5+3xHNsjdWzbslfUyvGDv7Ho
aPd0pRNtg66JrzUDoOOeaNkUQqxcvROgT5YfdogvoE3FlPTmTv5eNyI3FmtCdvVelM1MhUpnnveU
y/lMfN0WMdytEbMPCVE0SKjWdAoEzxBtqvtutYatFpp1COznDHtHKmO26gU9QJJaWLNYcRDfFPGB
vD25OC1qfyvgaX7MWfKO7NO7ogEWdoHRQWXoJXzJCn9MZCZbLr0AFMqd2k3qNXX4t47YdjjIMKkR
H/7u2+xFh5oo7FfHkXrstdhxjxefcYIZq54T3l3MXrQZksFnd7cdURPBt4+jEziWEonYC2ui4eet
vgErCplaJChm35znF/6peDrch2N6Nguz+nijTug0Iu6WkvT+m2TsA3vtOnQLEifDgIzirlSaIsFm
7gjZ6QZLixT7XlvS6kVnwZe860Nd857rygJA6cKjCDfxGrMBg2BhAyyjSwEkT2rCE98TOfmyzdO6
bdFqJTxL+Pywb0xHkYAAvJrIM95g+i1xGA8zDsBGSoZcLJJK740lf0Svm582dUBfbBf72SItdGxC
yKDJQXenmTNfCiLJ9G0r/hAWdS1sx7Q//0/+uK2ItI/z3IGaTdhOBjNfEMPnjLTFUHnx8PRb5uOj
TuYgodSNS6RZeZr9MKGRwmFkJOlPVQg7oKSlZr7WhT/HkwTizAZeZz12xhtfUL4PmBFvINiFnZOp
hWn+gltItiETq4ITnLirM22AAH5MXyuzgRXJGYNHFEBhMR47vBNajD8CEDAIoDSOLz4xmSzUN7/O
n8fCwJWta2ynBABXXWzpbYT0I3YIOkNy8kjbPwx2QQaFGEBxs3JkQqSYjkwYFTkaG6927tYWUh4B
R98+zSgNj9ay5GmzPzw2RdjKyB4cRzsdumJp6/ZcpIvp4islCecEaztR3ryCc7kD2kGkoqUBZNWv
mgZpmTvffIQmFWNJgQTO+EZkFJzzDyaExI4pxJkoB7soLNyXdYbPHwzFP5nbUjt3rqQNU2M/5Ihb
prUXBZru0k4O4DsT87M//W1f4p/oxIC3XJpLQVy9G+sTAfv3qpf5+8IVauoMprlMR+XeRCMLUfqx
K/+geL0o6xCyMHpFYBOn0f1UVMgdLhZshH6DdwuxX9eIFajC/X277Z6gAgQBBctHFgst1WFVZEXq
VvpVYFgzg/K57VYKQ/XB/RTZeEAMPxntdQAe3bM4PCpXCZTzScw+xln3raA1x4Y6syDMZ+Px0jwc
ME/KWO3Sfs50+aAksNtcyT6IGtgiGosMjcCVCVOkbrShSPAgW4JM6XCuDHpCpbSGZ5W/Ib3x7bsd
oR7RTbhuocfhDESq4QZWZYv9TgihvwoXGs78Ig4bmMWOhvgOaBZXIHuC12eg7bCLhr0FduX3A/8L
S0h4IAEZkFnUjswjRnelcbzXdi6fhQI4KgH59RdYfBoppRqGrZSu77dXYFy/cNWA7tm6ONSuoYmu
aGEbRaqRaE+3tkZJ5AUeM2T7+KTnHe/ra7PkcYMxtytjkFWYr7dBgAvTgtE+lHmAf9mr62aup2Q8
fZpUdMgHa+Op6dLIHhZ2I+vdA8GsF/bll01OU339ixCqNmZj2M3sdhwR8CyeCkjQOYqR7Gxvl4x/
BAMg1/hrO23rbVHZ8vCK4K8lSANNrSCFCgbe/zsGKPhEw7quDydzovv7wepPIiT1XxZoGdWYRwxm
FCEpLWXijQr+VP++4p56k89Y/KOeKwDlkGE14TFQEUEekPz203m3Ohp4ZfGzb6OECWfW86qblozz
9DkhKdlrrUbr6mH5o2gYH9Xz+LrTr5Z550neBFDIVDjOMAYYjnPSh3xrs69ttcHtnT6yZ4u2xsvi
/yJSXVm6KchlbDqCpmKq3rvgBXFOGK449Bp8Qm62eyx/UzS4/ILzaTaY3roogCToOhFo/Cazsn9x
42VRjuqY1GiO4syhFlw7vv6tlMI5ZhdKHQQM8EHddGMt4aAs9EKoN3k+zNslYEJ/R96Ci92gDsKV
bccW51RUgo+SNJgESho8zJ5f8rzgnVyMFd/e+hA0Mysdh/AKlofA3lov4OOgG5K7+yCiU012zpJs
ZBZUdre2wZbdJTReaaS3+wpsgzT/KdG6wUHoLlIUXTiE823ELKo8+VDtD6r1jzg7d7jbViB5VPKB
U3EZhCFrBXETO4Ag+C9gQiANsowCQBski64BMy0wVmdgYvqVnMEZg3AYQ0NY0TrvuU0wUPthDB7B
2WFW8rHkTA8c0GSEK0Nm+161nzxEyD+o40tEic/lsmIAh61pcWB9+eJHfRjrJIGnrGPPVTI8k7aQ
F1opGWVbEn2FBd+tv30oPSgtDFlnBEu6Olq0MW3BRaO/EkoTvEBHHOaF5EuO7JZd2gSXBaJ5sMmX
7J1d3PEphiRsbTpnnZ2aUr+EClo/KlJugKFBZRsGKlxzn4kNPPFw0q3BzGEgDZUbfvXOQ9qmGHiB
lidhwGWXXKNJEyxeAlzmXDqIZiqCRFrEwxOmlSXVARjHTJzHbN8WS+ynTFGxu/FJtTCOZ4a8d7tS
PSG8uNd+DgHaXwpMc0moDS6TozwKxO1SuQxxIOC2kSa4B50xnJ562HkVYwyKeMvWG+5PaT36mCc0
NjxUxaedvtsPs3Jl5WYUXF8dCxGFiOKv9ytann3ITskRWvNl0KF6YLmbl72ZrdZN5jF2Vqt1uxMG
m4IlujHyYLs6JTei5EtlzhYTn+/AX3R+GMunP/DBcSNMNlvW0S0mgqbpBGk/6ap/tonM6YzfzbK6
JHXk8VXytyxxMl08dua3KQnuELdUlU6z2JAGRU/143i+A1pzTHwbdr34lfiHKJ1oack1l75pcM1N
X5pWeoU2ClFEI8FbbuK9hAA+xYimcE/XpPU2A1Cn5pvAfy+tCtjjLpu5gujkhPVPdFetbEpAUZ8M
aJn2nZ8OiRBiagTdFDfvbcBzY+8/kUAXraBYOWM+Dw6mOgfyGiNWeV2lg5MwF1KXx4xL4OMROSa6
1R9idYKiG5yqLKXbYzJbbeFDcTAJVjhS+NFnFhLIRSIVDddvHRD8vejJHSAtE4kv/tQI2b9QWVcx
jShjY2S9yv3kyA+egXXSJKy8uZu9STMzeNgCIC5QBm6mKl2lyyAV0g1BGHJWxngEPBgNbB+N/jJZ
FlyU5/Xt7/BD1wnEh1k4ocFLAzz0CxFDACsH068zWS+jRKgxge6O2RwGK4KIkXIdwPZ+2oe1RtyF
ASnMPqt/cuvh8QG9Ej/XV1TOq3zwCuaogfjnwKn3hBBCOKQTjyb95uNTXsqWW6XQU4+HeWl4oxK+
cStu8yq+hOeC91FvBaYEzt6GSZwikyjrcmPmBVUiChUHWM2mA4mah+ApXDKmNsMa4mAGnP380HFr
sBz55prytu7kL3xMZYOckwFmq2CXTzaSO9P25utiHAdaVcmYCNlBvSFWXK4r30hIGDslOnq//6WY
TFGRLo1mvHRjRYt4ZOJ2ASiG3okP83Nq29wngh/gMKqO9uHqNn5csSqhdrXTnYkcyV0TEgHEER05
ufmdGmjuD2NGVWvAc54HYFzbj2m7wg/OuwobtmzvU0o/22GP9nDy5ikB31Xx7SamGtVVs7v5bOjL
KucV4xdakihl/eUQG8zLHO4pRv+MJgX4bWS1X+zdsqZo2DsdfvmaiiHJRzVIFYp/C0unR/Cv7RWV
WSrZp1fxf79EsvQyKk7iNMtD/fZ1GjuwzPV9WZ+Y4J1rReNNLLq0L58Brkqwefidl+zSI5z2mWSG
GD0zD4eZEkICiGkRldYF6S92vyAqfIpH28IwcLYuVOZPSqGalncI/HPolKu/FAqYdmhK93eOOFCK
zrKxOhZZHSoBO1imVBDth+LwhkagiuMmVN4xioYH/KErXaYPA8Y2u/nVL6Ay9RJQWpgEZdX2dJNb
MV8FwzGCC3DFw6CDCX5nTmoMMPGmIOyGJ1ScmGyCy1yqF3FK5tRDKqk+sOv2YqkvnbOUU67uSbnN
Sq6jxKE+35Axxcfr2lQXWA4ZL4DMsaxh1E4w5boGO3ccWmp4/AkJh91u6AmYp8y/RzKw0NlfxUcu
cQd/JTgyipt4mIuip0D9Epkz2XfwvdRf9aCSTAkCF7ujRsJuGdP43hPt1VJbdyCsNU8RrEbSsavl
IJtCEgiF0Bw9vXkj+eOk0qTBkrjXw4tsZyvGR80kuaybzI+gUF0i3EA5Vj0JoBNyQwytHBk2rwfs
I+mgC4SxI7mD6itng4JexYOQ5I6u/L1Y3fyg9yxEnRS9p4u5kE16/TG8eSrqhtg+/mfsQKwGTHnM
a7Zg6HXGZH3L9nXSVjpqGeeRVGErWd1zopM9LJJr5jiT45PL+5otA2xk0B9E1h+tr3HiYHHgP5/q
9nrQ7qMECG5HWoDCAlIofJOK2yEpfJ0Hddv0Y/O8Elyk9bm1mjIWc89LarmkkYsqD1JfM4Arjcpf
7G/xY+WgX1GS7tKpQXXwVPP9R25vsgkajBTywqTO14B7QpWRb3+74WJq5sQvztDA2qaL6au3b5Uh
9YUDQRKFOgLAHvniADT6WWFDIc0TVkNCZqplE4azIqVAQJlOn9UBf6IjUUwdzXepP41fBiCY/sn2
xv5afJC1JEzFxEGgwrI4ANvA7BwGHklBerZuq+J26issRrP9bk3jtwhgfm+SHnBvvaW+Uypna+Ah
0uUdT5IR2p6DswHVIs5Ah71zAOs03zC7x+929ZOGxy+ZQ8sIoqfINmpziegqJZQ81e5Rtqyj7DCg
mJyyRFu0iA1iokG9F4RAuh0/Nb6hqyAG/I19AYudqQOGGjAdwpRUrd8nTzESTqMu+DjKc1+x3LQt
Hc6y+a3pF3bzKigb9O85biIfIS61gHu/9LPbCN/T1FWVxkKrHtSf1oerP77ILA0C7zQqcwNKPZ/0
kyAFEZPvhHD/sovLTk5yMnSV1no1pTxKMSVTIhErYfL/Gl8MJd9YtUDmLm3v45MYgWEoCrmxxFU+
2V7OuBeAUp7QGFb+V90CLS4Z3l/XJSmpqeq3YZMiuHG74t8VC6udxFjcyHCJbHSlCBGJhgD3/C39
JhDmXP6XoU8iZXcYEcn9fM+X4i1RIf+RlLxRxmovTlCf6NHx5gCiyitCvkRJRfMgemkzAtt7Q77u
FNC1qQnf5ew4qxuK4GmH94NxEZwaWnOTBYg0WYdqgqXZzHjuEZbBxPltsh4vWdmWM24JYG83vywu
edA1OZaSxMSkFRElX0EtdekyuH9fH7MJIN5eK68HVbv+ZWu+QzOQfpVXn+c8hddLJmETzdt32a9N
fncKa/5io9zkypblzqBzNYJ25UD2UkkNi7kcZPAd3ZWgo4XJCGyZ+JquyoTO73cfaEYbw28XfJMc
LhuydUZbXx5f0YB6QUioPUPOrGS00IAwrB1OXw7P01p4oCg9aPJ7+Dx09kXELEaaNjwmokQXgROK
+RUPYtV21cN6w8V7Y3Y8qsbhPPGtPVusDIKCYTeNK+wHItPgCy7W0tc8Jisogv5yWP3agNyHHlZ7
6GAKqhZASPhSpslItwKJ5oVT3vxtkNGduIQKhvQMpJ2RQE+kNo0q+4shC6RqYROPnOgNpoiEg4be
RPcHFQgJhBpAb0+FqlHcehX1iLY6/CkTQz+NK6HObCryKCEudxADJSIBhl8ukLwb+WVmz/MhHn9f
Tv34oYI2n+yS3igGv0/CRi9s92vRxmWhRJDB2QyrXKqLA8jVBMg/swCciHK9v/nnWX0pjBlyCJEm
xLdpbV9LJRd/K/RcpI5/jH+DoOOLh+w3ze/Zbp/iDEaKm+/NZhjYfzpLbm2olC7yMPgoCbHU2SSy
o3r7wzitEA3EOR0s0I9JGTcVkbCtr3ldbdtNvvYFvsSdVMzqGPF2on+oOHBLxJpE+SEuE9L7mFPa
vRolQChvwFu7b0QppfwRtMzN8HZq9Y7CcGqEZp40QsDPd/e5LHuH0nz8W0sVgVJLNePEdWkb8HWg
CRKcwudmR9V3CBbn9DzO2LpunbXQwNOdqx9L8vGotCM0kebUZYHYaVIsYqaF2xIonSDSZV1p7WsL
mVMp0JIIwhzpOeU6VoLvE3ThEQn88LmajeddHdgE+1nBDf8t+AjFiI1+i/HNivQBbgU8v5spIUxi
tQ24Doye+fSz/A16DzF8660/KvIBN242Oz7FoV8Wfvn46Ca/qShqzf9MuZ8dLGm0YAwjJ24bLyn2
XxHmg++QuZ1JuUaRgj9KRRCE3EZRGCcEslPYYn3piNdEVnNSdz/5rHRFilcvXH3W9KiiYwxWk+L4
h5L0mZy4lGqbhV970EBFvytPQZqFEeS2CaBnx4yiq+W7QQMt39qehUo3k05IfRLTsfTw2hTgYjJN
37Xryd8JMQdi0T3N+xIq307FDhZZQyPNhZlU0RDE8ghIm5OOPdxLYs2uHpOQ+jogKofvUDYQO2nA
WRIsHmUdZeB6eW91zkFj+rcrsVbUDWuHdDtUfVJwkwDbkHE8UwjpJUm3tR/51K2ztZId32/JO9GA
cQdjIc30Iop3MnxtOu9VGw6/S31c7cFmNSlAqOGhsm2jqKHLXrfqLhlDqkAROMCF6IwPbzqQ2lPv
luCuf9/fx2AkSYNSEGIXPSCmypEj6JpRk1r8wYFnQNLlFF5LnCRyJcBee0kp/mj7htqrE+vR6o4i
Ml4HT2eUl2s3OReCdy4TfnZ2y6nmLUIJFO5e/QvKYTp/IVW1f1hmMwyPZNzgWLDnuwLQ731PrUqV
kOyS6dyFe3C/mvRtCiZWhfeBWsIgnt3b27WgAbMP4RJ3TR3+SKK0koyEEWpXDOCZdiLz3WrQdLLt
SA6XiArCRNvU++iC0D3LmDJhO/XXByln6p1F6ZxUxVitUlfiHTfs7snkwO0FfsuGdXxx2cPpFMLh
PnozKZBaGQd0Gt2OYK+17Ea2HTIhkTxK1v0QlrS4LsH9SUV8CfQ5wFHufODRZX+DPxvUwgDtJ1Uc
0kMgrcLelzQHYdNS0gNnu2x13V8l9GMomZAy5P09aDT3+7wVNygP7UrktemYn9DQ68COQEILfXpK
MZHn6Ytt7OptWNW0SZstmzgHGLs5uiKQR1D1xXI6ohI9zr4scjQ4WM/yEvDki3XYGyTegrB2uO84
x0i9mHtpwMoJOCvrpvLYQKyntq9u/wm/DBnbDyWy9XSP4ShCKe+1MRssEg+GWseeaJpg2UJlvJe3
zwENTYVAeG6o55Y6Tbd3A2B4kt0t5NGtt3XhIwmQtECANC24qpZefrGJgTDWIOSMXcHhinS0cC3H
H5qEAVxtNkM9eYVSEsnfOJWUHdUJPyqfj/1Clx12XdXht46MycXtvK9alJ/AZ66vXfLMUf2uUqrx
BsayezQAK4A8v3gORkP2iJwK9ozaNLPsOTFbgcV2vC9SZx7fMshesTOVA6yY4cDBqBzjKSAe7+Z6
fydYRLn77x2zZIs8SpUfv06ThiaQ6IrgZlAQ6wia62gR4i1yTFuv2uBB0qv3s6FGLICiTq79Xu4o
Ng3ovjUXTatfItQlV/IkBMbeTMxyk1EG+g0P1F9wYoi7c/Vljhd6M8PZFW0DrwiaGgov+gLbgbJX
MCMbfIrS87ojKfvfiP5Q0VxaoCi2a0biQfqtDfmzD0VXWzomvDpPngNGvDy1ZZqmnnQyhD3SHJGy
8Ofvp8tgFPgZX+snjEXnUyKt7UMwjGyWQAZGdpIn1wfY0GWVTlv9iajf1tljnT58LgTtyb+o5lYv
fwRk+qqsekJBFuPRJ31WHf/0G/ZYY17StWQ5ui5b2BmWZdBhe+3DeWF7ux7yIFC3gR1w1Jaqu/QK
o2fTmG5f3lgTMKX5X8hg9EnDTmgOKSDMsx77ZlzzYmGIA1iwot/8mSSJJgyd5/BQskENTqs/ZPaW
4YJk1pZ9eiMBX78z7rvPJjPGOa2dUUEyxGduqtR9knffoyz+qpzobMx7GlpAQy1UyFYfYrpxP8nM
xn+fQ1VTTlO7+mMeW7X1j64J0nbFaqDPSU5RlbSEN+pRk9i7DKQA4QmRhGwBFcNQcO8WOUrS7gNl
kBGuat2xCaiiukhzAYjUH3P33IsxhCNTdcpWZ+bYZZHQKBYab3E8YwMHTE7sYZ6HBJ1ZsLjEpQ4J
o2ai3WAdd9nKRBgPgsbf2DkIAw1ks+UdAQ7b3S4u+Z1KrQL55ytSi2azcP3AcvR7PkxrKfXS+klR
Gj4jaKsOmfFWnEHowAxPElHP91JhhdIfl2UEGw4ko3SJNMSH7a1HxywuzFJFFeeTbLu2KltoMGur
nOQBzTcFrohWjjD8YbW5q8H0szpLL+T9jyV0vL+Eu4/xc58rKdGDSjBMCWRkECkGaYi2Rc63ze+X
iSMYKX/mxce7DWcXrc8W8VVkhYosOa2409EJotH6Z8cjfyP/kga4EFB36LHpw4LIYvpocVYwIrXg
SxZQmM7UJf5zu3YrQOR+ns0Ut87xtMmPXihYYQ7iMjuGW9TAm25Fl+U8N2dorsmaE2dAUhoNbsp3
eLj1desHbqis2zJ0QhwUiKlMG2v7C17CTilFzRijs5CMxMTlBBJIdUTy7wZhCdOFcry/ClzcMXZR
rKzh2xNx7x1r17Qaiuo6h0ihbUasluCjjwjzCDenRJf7NQy+k6tNgkDQcrnpkWj2xZtjQBIGA5X4
EJjcFdxdJGR+uJzG4CKUQ8ov9zVTkn6sQEJ5mm0be5dVWW7baQ+3RdiiBbllA7vWGOy1CP/MagCj
CTXBXnQLVobfkcb2I9REFPqgxvy93meacxEy7VJ3j0qDar3m9EncxjiXU64sXi/6huDlh6Fz2dLw
Ow55J59B+O5AEXy35DsZ6dvDc9nsptfgD0ytFaaMYWWfT4Lxv4obWYCzB32YFwUmaY0QkHgmaGPa
MaZs2+ydPzB7cu3735WeqmCxUJFK7BZtIwNPh8BzNf4Kzy0AVtM2ipX92KznRbZ0K297Kf7pKQev
vLxCnuhvMDZjcAzI9j1PY2KVb5zvzPwHglMq2blUHUzdw/Z7QuzwqOnHoaGz4hE1z3omTC6FFRkM
PwTbP2tUBlNuhp9cM2kjXgJ1CrsGXe+o8hFQGrbZw6c5gJaWvNeA4rrkBnpR+tLktyKPcbMFl6Xv
x3bRA7cgX4R+8eFEH/yQZ8/9oIr9WA1Kr+wt+6/B2l0Ypi/0xA5IeWHXWtPJhetFxxmdJhRhsfMY
yZd4OrS1L7emnr+wCzzvCX/gXYubUw3B03+ZwgbdBsYwIEP/COkU+tssUzSiKkIKVOZUS7zxJCKZ
+HOoyB3pWPs2LuA7lwpmLeV+qHtKxdGNsk/bRLCu4ipddOEJ0ARqIEZ0kK3t+i0aimpGC6S6r2LF
3F2hHzzyXvt+laHgmygFgwSfD8YtKaO5kcDyJEwlH6N353oILWF845ljtDiDd0zMLaV9VsKUURHS
dsbuUC5ApUVv2uKVkfjfGWDBMGmjDcOnwXl1u25A8S51rcg21M4wyGTNkX9vU9KuQcBabTS48bvD
Xc42OfuRwbZE8zozyIWXxVK1eWLQSd1rCDljKqDMyf94m/Y9in7N9GDb7207EoZ4lbtICgZxRi22
brsrX9bYe10f2gS7IraAEDwHsg0t6gBK7JQzvOdqAGfccl9CWyu5UI5ooLH7L/GGiyQzjmCrIymO
dI6i3wDZIZh1Nqj8WZfaxRxyQCta/2/B8ROCrnl6jKIOOOveug+dxPmaVbOGeKuToiN54o3bVM5Q
yHDEN/rSaQNYFxx5z2eU745dBEDQ6OP4SB5SPbcMheHvx7cJluHwHnabj3rb1Jtb3yRu7vgHxkLG
OdiFGWvJ/IeBsPz1Sl9Z5Mqu6n30hEPCoODN+jyi5WEP/aAEh3TdaESr9NH6awplfK96sLWPOpSp
R8WFFwJ0JUTo9HAiLI/vSZ5M7LYneyODbr6B2R491YGZoCMgnp9GWw1QhQ6iF4OEwlA78+ymnZZT
MFTIKSxHCCABvJt/HHPq4Y0zTs6o8f/I4mxa57XuZMDj1VdzSPaDuYjhvbK+vg8/lTHYm0fZM4VP
sIe77eaXrLJbLdVQicALeM4vQsMUUSt1USHNLpsYnG4uhdlQ9ymG24hShinohLdUeujp26nzgkZM
xdRjqqCurniT7jZJ16e4ch54dCUKtNdMdEHAxunj88i2MtidBJoVQFsuOQcdjGaZtD9j8MDOv3Mf
cznR+ZC7tLiarCjc7LkQKcHpdzsQoY245clUwiIugDz3gJaBAa58Jj0eb3Jp3QK94wGSkYtrnq9g
/aUZ9vviRmF7JnJiSVj1ChvOup5XDDRW0m4gipw7KaR0Rzstxt1ocn6CwOXTxOqBejHeNUvdzxfm
ht6CSwmAROwx7pbQO1sw0uFcJv6Mvt4G1+mZ3I59cH+VfL2/psf3/IYGE+sIKq+daBMY4+zlec7k
xX4yj5Rrh5khp7209iHBSYPOUM0UAhlRX/VL/yAvUf8yjdwtzwFGOOq4n4pHMe6mHdX9A5XnxPSW
HOU7NNc1SGwL96iyNfkRsgF/hMnuaQEmRIqaoDvnp3Fiq4LN0N5yyzHmnSIEkwXOrgoeow0EeE6e
tynxvICPwGCHqPjFEmsIMEXgblzGuyd/ZoJuXg+EjhCR3bpNMypFp6L5kWUxjLwIxIDuUD4ZzB4n
CdAAkQsPtM5jMAsATv9dEqxrKryUJDG3O2YvqrwTH3cz7EsP32LUMk781Kq43yJMz0jD+E4ZcNLx
D9MdL9aOPJGFKr2HFXg67rlGxjmswKDlGtI28kVieh7IOo9hMSpgh0/G1ZQnq+ouJbq9+Px7kojP
qreEgb3rGEfjFZv9wRdCLpfovIulR6UWutXceYhPjYaBLO+UijNYlhmH9v8N5jgf1XLz6x5NQGqs
sGsPay3VUf5ztvuems0YVAR6cwh21GLah7Dn1c8MSJqk1wJZLPb2lqHXOOmUo2cV0tU6OxpiTXo4
bUjpIMH/2jVaE6IwD9j9hmgmWZm8pXC5wmWb2ZsguUZW+xooI85oSkm7/5LdktgAZSPwZvmzeNIZ
k8kowJtcW1l5unNYEtttdHe5l4zY39HcbdR//VQxP6tohRQgZrmlPGW4LAhH79ld9fzdHFhgRean
GSQhNysj9XqKBsznLhV1wp8TTyy9vv3N3HpgsB267jB/9C1wht+JzZSjJNt3zaMBPU7xBwrX9PVT
iRRl+oontRrYa7FpJYUThIK+buxgkPr2SxAVjuTJXLvEGRGXYH9ZTcwU5lR/VUhbSR2VQuotEJRT
oPiFIhTfYjvgI2x7Ffv/ywhPYGhVRfLBJ6gXKjQt1DiHHMfmiVQuQJm+9JDCtHm1ozcK7qx5MXJP
2jiubJzKH2c8L2G/AlpknTs/hT4/rxWHB9nRJVTjwDiZ70y9/KdmT6opFJ+NqROrrAASf7jT2Pzi
MeES9oOOdme1iT4cT/SnyVwnkfIqP1z8AbquDqBc8xdRz/Rm7UE2vdsokqqGRkiZhLNN9ljcFd9k
s/O6r5sDIkq4YJGc7eP343RTAp5/dOPuhphY8NjqQLIaVpr+mUAV3s2vqaTRGdQ/DSDO7tdn6bNF
iV1NRr3yexyNa38aJlSBCVe44oV1Qc9RigHn3ylgIFpP6MIPAI/1CJByZv95SuMXm9XwfxOm+u5+
Xiw8N62YZ2GrelaHd6JmzKfmW0nSLHVqq3VnESNW6zslNtg9tmHbzGFTLBOc0MZz5gJwQXAQnodB
3rip6MLzNw+DbhUeXcaCwUilmk0T8bpa/41/VsHkLe1onGbTUxS5tBAHcyz5eJ8vNmGpzDmctDnp
bYEFW9BSRiHq3URkKOJlfcVwTTRFzzVLPfwtCRUI02uGzllZDUNLq6k4Q+X7NqU8BRz7TwDboMDf
mQEi3pyt5YVk+5OLgkBOWaYZ7VqvkLYVRo75p9b30p5l3HGTgNYW2AVy/ySTVVJ9PsACjzTQzWcN
y/iLU1PbRj5hq+opXHNnUk9K7ncxuQ3Mr4A2RzewXYU/TXBHJas380tzi3KRvRYtVoUjBqb3KIS6
4IMVbcmG66SgHs5quTrcpSRZILXa1OlRpF8bVYSV9VgKyUUqEOwWWF8XLq9amwxNxNdvzt14qQmO
iqgf9vlNF9j4LxanZa3TVLgWPNGW6QNd4OEP1sa/1o4YbLKYM77Qss1bXXk61y0HhNY6sqn1MPi9
uZ8tnFrFocx9BPHulzDQ/pRWAuuYfU3ZK9BQ+A1bCeT7mDV/zNRI91Hnn3wMgUCRXRvb/DHSROyo
9khDNb7FcMTc6mW6UPlzMqdTQa3LkQSzAOcQ9JPG8NUmHLmODZGq3xnQty5cCU8DptjWEO7Zh2OG
vFFZPbNMoa3r9gPZkzJ1FDlhUBystUTiWSIXwDocfi8DAu/2ybxJjBvplS8X+pcfSJ4B9MoImwx4
YlJO4Ww/PL9g1cP2OhzM/YEsSUTTAIvxzRxtUVIUCsJ5hGO9IkZAMmMMmpUXbqp/ZazO7whK6+Ab
BjgAOfJdAcwEcDFIF2NR9udTeHqVzuDu7qBnwLLLlEpGSdMlG+dSz0nJ0fl3xQkgs57LNc6XYVFS
d0vQqh+TcAz9Qvrgds9+YlsuhloerrM8/VWM8ZJlLrg4T+22S2E/8b6oJlgiaFvd/aNHV0kE642A
GU1B0Xc7eQWH6z3kq051TpjiJPHrCKlqmrXtNzqHfaJt6cCCGAA4M4/J+kw3jbwaqwVnvhd1SxFZ
DrBOwzLDsPsJcQCfUb458b/Y+nac4nz1ZXxZH4X3GlQ2SYS0VOQoxdDS9SUgDIFlql9JAaECOY2c
A5RmngzZBP8elXi0ma+liArd0IbBjtdU15DAo/Tec3sPP4i/cOXiUC8fyuD1cnRmIFPn4FIEcB7W
WxJaRewzpIW5PWWohFvnGV9B3QHhjc6JYhaKItr9K+5BBmESmPhMFMBvXVl3SlYAFyBF3NEL1J1q
8TlBSPXN1grhr7dIUgFuvXUO/eS3pQ3k0HMPQDrbVJ7TTCpmO3TIOfkcIyqlH1ya4IbaZEuOGCcq
FKq7Np5/ustpI1xKbHuUAG2WAK0CgoNzCrYdCuvKqwLC3Shp4ksDBdmCIYrmQ64xywXpZuLy9EJo
BIs9VjXgmFAhhiG+jyoXLJS+OCvRDlhgkWZVUeh/D4WlSHIJcGD3QNqik6ypU/EFE03Z9IR9OsNn
YO30kSCg7A/bZ3wMDe1d3U9HOuBBrRbl/rqf4IZPeFLyNBqS02PYaq1cNV+TtHWxQPLOqnwIxue3
kCQy1FZiiKjbdJwkEmWKJfFVCzE86ne7oPpGWruZjDcEsaWD+zPAhah0XmikBO9pPegcU7gEf2uU
ZOFebYAKkhGcFpGvIfSrmtHcSlzKCQD22lD95SItK16FjEJ5cchoMmnFm+LW5jcC8eAz8oFZSyVR
KVuWQAkbkTizTXM7ECdlyfQvtwdZpOGfO1S0Hnk2S6u/EfoP3EzPF7c0usYAlV9SkDoiTDWBPPCq
aRux/JttkRRwIsC4LarRr0EI9x06dXoYeE1h3Fho5ppS56sin71LoTmTX7o7jjbBGAcExLHAeDwy
hMyaK4UxFWtd4TxclLFnTDruNTGsyK3G+fq9oRbZnlM1imQIt9fFNp4YMuWvWEk/GnFa4rHY+HK2
wXthGVAsoSZhZcK7ucDqTPu60hjtuWY8LMFE06+sae8UI1w28LNI2rYhsb3Xww6tW2fODGo86KYD
/enUMVWRrwOHqESvedBvOii+5F6fD+CAYNV2fR/k6cASuM5uw8uzoHk8j9IbsBY4ATjDv7dPoGp7
1nJJJxUrJorp55OG9BvbdOkD2CyjWv6xNrEU93lUDOsL+cp/tHMcTwOIXk/y4MppZPEM/6KF8vvE
iN1c+4S5zUi+ETCyC3VgVBMvp0CSdpGcTQW7alHhEfeThnEP4FmfHu4nea1gJJbrUd94tXszAaIF
lRBun5MC2gKnDQSkMrKytcs0ZwynSF9F9znoH2CUB33yXkfULBQzkfPv5H51hbTS9nEwz0ZfWY+2
T4ADqMEyfl/SJr+0WqysVo7P9TQYIqlXdNU1DvNOcaB+rKlJuX77bU+3gdvpW7VZcMTAQoPh5+xB
hd0IGbCg7fSvQEt0Qgxr8UzYfv1LEReh3H+uvtd4s0M09N3WCX5NmUlNwhiPCT66H8KaR8ltZ/zu
aHoD4UC33p9gJGsQidCI1TqCp0dMzvEkoxNnvdDFrsTlSyv8FE4wVVwWMlj2aDghkXvOJvDBUA9i
uKBmB8MeDeannRHkhz7oo90ks1B0sMmMVDoqMFlUizRwtKFhsmQmmrgVi+yZCxvYYMTYf4IP6sgz
TSTEFtC8IY1Op6MMTFv1WSufhWsr7dTvkzoQT6pkktE2Tx7sBBEprOC6p81m5oDN9dwFfCcFFUmH
ioTTcQBA0PIjCVWkOoqKKIbRetpkrgsmnFNP5YoP9NF2vCHiP/dVCFqVps5XMA8gLH8QceCuGP3Z
KWoI4QJT2ggXoNVzspU0GsaS7sBUpLvF84oloyUyFGKXoZbXJseRW1E6IkUac5j7trA+3xuafmLy
s/RTZrILMi8+T/JZtW64VXaosbczfBtQDgRxnWkiZZYEVf7f1EPen8pxxEi/dABNsJVZe2b6Zsc2
Lowe7canWmAJRCZQApDWziv5b/B9BaYZdiegNBtKBN0H1E7K3o7jPydX0BkLSHgyyziVpQZYm8gU
mlQG4DH6+cuuzIlILZz7FV9Fqloak2AeT7ZWqXd9xXT1CRl08Hs1jbfxmu4DHCWmY5vWNcIO63mx
WR3WQp0HVUgCLch3wXW3TBgLikBmVGBbSbxT+2kyhLeOASNVSBIq0Nsk75T5DgSLtWd0IPm14cMu
/9+oh8axrG59SFUHPkME8z5NlPmhS42f7OKAmlCmTPG+neclgzquUUiLS4EQAcuvEnI4qpuQRezB
1dHtqgxuZXUZ+wGl9cbDfLgt1SPXvc4qkme5oiikOWi/RtzR+OEtYJlZMtHVrUkprPJCoNR6MgDv
zt9W2zbVXfwTe7dhMa4iZJwDHmmJB2uOchj0WesUOcjYSmiMkPlgXhQL3pUkf8zM6Iw5w18y+XYX
+MfT3BxLHGVp3ZlShk0pejyK604a8hF1Rr9jjqac42ARKlQvnPQ2aGLDgHvhD0ta3qZiuFv9b3jI
VcrQ5tkpGwA84/uTG5wGY9J+XyPKPY7Afsy0q4wRSSVX5cMGtaSPgmvZll/Q5SyeFN0rhvW+3p+u
9vmuFvOGdSpHtmSwzQ/WvADUeQgMxfNGeMbI0BSin8gr2LUtnJgsANLXOnLPHPvNZh2FtZNq52bk
hS5R/s/m235Tes04ZgoMGN232B6RUSWL5xU1151KV1w+ylRq4YC2+/O3dNq66baKi59Hgx0IX0XL
GWzal4zbt4K46M5NZbFQIEJEEl3l0nUQ8ikSiHogThMPxtsXlz0azNh4OFeqXl5sE9+TrvG173GL
2kCy140SrGyxwThFGesLaE4Tlq123+Gy4jwUjXEyrTMirjONOblPeGTJ0qT7ug1ZHs8Hgqi2foVB
mWZAnnmliXMBSCJ9fjREla9t2edVLIzho7UQ/M8nqOC5HebR0ow2mL1m4uw272UMQKoyWGwEJ2Se
gae+HCjnPdtSWxT5dDg5gpNAaI+JBdqjjK+sD03czezw83qrJxnNfgxj+IS4Gi4JtD5rPS+FmhP2
nXe7uZNk9e7UrMdHBCGrlcNS1Z7bFs1SFY9ja7JG3QbjTD75GlYDThAc4g3X9/7j6H3AIlBOWaNc
CqOPMqbYqDBHpE2X+ktayoJwmHMd/1aJXReY52jmsVtxXR8ULWElEiZZ2p/TLuz7V5HYrlYmJZvy
dbN+0XLksMmXsUnN5HFmC1Z8zHGFO3n+xZzgDT9hNj1HOAPvsVy+rnwVpAfOYC8T1dy8qeBO4ywQ
1xaqihqBP5SeLGmDEt1tYAhdwEkcnVyzPMqd7cYdPl9P70F43ZeIJ0BSqJEg6+mmWtbRL7uU6a9b
lTvc4by9jiN2qRgSxzjrgDtnYkhgl01zY9E5I8oL20PT1qESPCeV5wc2F73JI6tIRZ4NeF9MzhTT
6iTlfnFEzRkqSVfwpdOukWN7BtUtDmxoCjk1VsfdOOes8V3vq4XKmB6EjYNuQ0NOIVUpbKsMtK3c
q1VuBxHh38QNCuxp9CmbOmR/McnIkdqgiuujJDNgWEGLJhw3THb6QLLxMh72TzSsIUxFwGxmNw4C
QMcdA8u8uiCcbmbQKfLiVICMLNwkGJS5R4KnnE82D6CwV5phjXEqvcrwCJ3SFOGMwdznX3R50gIl
FTmSGGSl4hsEW8tJbKbJqaR1q/9G+UXFk5xFFqRE0/geux/NClvSokk9phRAr/qFyhPblosZHCDS
HnhakcKkTk4boPo1a7QSHWQcL9ww5yBzUnD4HO74wSnJja0aBLh+VCLAlQLLItShoT5IT5I2wqFQ
kH4Kf52lQINe88i6l5+gN4NB77OgH8LGuowZDA8hSHuAWuLoqsnlrBaEWKOoSIIZAXCj5srkaUvJ
WinQAKPKfgG6XcsC+/hxaABX4dULg8U0ua9jf6kou0YFyPLapHyQ4aSyj8huA6YDoyhiIOYwGry0
/5IyQy0TTtTk8miv3/nKGfWVWlokdLK6H3wYPyHBx0Qy3FRW0TV8gHrK9GDHPhNHcTc+mH28Ahi2
s4ZgCZUtQkRG5Z9HlM2CgmVAIjgZYXlu7/5iI1VlODzsyFCFx2P9kSrsFFsdK5pw+7RHxRq417YW
/mU6t2WtW71yyt/5NoCBqM2WZjy2SMsoIOZmocRce93WVJa8hizyFHyE6z1SIUgGlfnavl8dQ86x
jI/oWMHAV23fcGQM9MqyQ2CDGeP0b6f3RCPn5D/S4VKkVwSMz0noqEIc6UX/hHSenyhBa6vFDI3g
gqvVjhOYe1gTtYTOo1JedsnuaA4OTs/fGL5kXUVjpOTrykpcF3e8gwXWgSoZR/47hZ/PTM3JUMBx
7D+jIHuIyd7Rl3vxDqbio/5bVdh3jo1XbaPzc1KnYzZD93yOR3V/gBA+sYqzOiYD5a3bk5nyuweN
Bz5B+hcz0L1Th+FTfm1DutkVIHoqErKoDEu+EVhVARz0dlUfrvlTbpk1p7TC4TfF095Hg/CbYZ/q
d8yxNmxWq2g7AtaL3HTCDrq+aoOibgTIvERMOMErjvKcrjtLbs2TwXQpesH8nc45pxuntNAvct64
VspY7su113QutuOu9nT7554abqeC4TveYxBNt4rV5zkgdJbHjmYuGT7dWmugmXaShoeX9LdX3wh2
mSX9cSwA9yefFwruPaOwf4LecWpURT32OWCpFb6TfYLGelgbtsUI0Ex+E0nn3X8BMk9NgxxlMtnd
CrhokT0ptJRhD0+Evo0lCSBqBZbdvoDcs4FGbATwDL5RVffvsCJcqGjmGCCfZAHJn0YdPgZhq/T7
qb9d47qhpIJPbx9e74x3qYDIa/vD234+Ujl1RSKk2pQ7WvLFo+AxQ1vv6D2Tp50fLl5yTyLi51yl
EtwwUwSzo2soENVu4W8g50ODzU00Epv8VS8Ggipo2+dddDqV40dLpqn/soLJgqMk93OAb0F4pq6J
zyNyOwhY3nQEwaDOMLEQwGyuy3OLJ+aIerU+MyuvxY7Cesp4TuWvyFR7rTBdMqjGGGPKHJ5pvfOt
cew4UajG0DZYwUBznrm1nG+eNjGdgzfsGLNhhN/UTTvzUvt0vLEZWY+fC+BeF5AuVHx06DAHWE0y
Hrk5SE5TN6I5tegZ8w8o/P9YyJFb0aAe/9yQsPkC8WzNyNM6T49zELWcFaowVCmlZ7u9QLDB/lUK
kv2eecVF4YmvTFicyj5vfPP0kyAKnSY0/GYnbsncD2frbj7hZvGhboA8H/HkqqzVivBuFjOrLAmx
gRNmgAyKcMS3iTD6BuYCxmjQhBEvfXlVgk4JtfXLySmUW2KwHInQ/8/EvKWMj804qZb5bxrcd9f/
a3YXk2/wINJjPdGJnHiQoq1Cdw0xNH1SY3VLsTPVQwwpU0rRk7BaI9SWnD+IA73JQbft33Knw68E
5Vbwtru5rmbpqDSDxrjih+dufVOnx6DBfIVstmJbprIDvsJ8aYC+jZVEfHNSinrkqpZoudTBYNif
kWQdor3uC7VNCKJ3Wu7WUjAaqELf7yh5RGDsIxjVVuMcQZ08RXWv8IwI6wDtcOM7vl1uOGyEtDF6
ensN2lMkim4QmHx53yqczG8HhEPY8kUQlvMQjM2FiDKlIwYWMCG9qxc0wnZTp8ahy2mB6e9n6oe7
mu9AsvAp5NtQ2s49tNUbRIcqVnxHTm/TEPQ+4kUfhfBZtw/afy1XNR/P9sOmYBjazyH2MRr2gdzx
OqiCz3nfWSWvqSEkAiW7xsutIpVdLoM399vfkTseRNWOvuxt0yLEBpNR7GcAp7oIczVLPlzG99va
7i/SLbGHoPrGyIM1VVzTvpClmIrXHPKJcO4b5tomCUsZUQz8yERGAtYtGWmhvW8/dczqb/q0gBp7
h4RzJ5+inA8xc7hnzAtQEsb0BV6Z9vFQpzJfk+rmlyOigW1hs2BJ2JSvbCP+UPBQJf8DriOUXhzz
h6B0ZUECtS4kcQ7taEvLXbcTLBNqRKlWuP6H+qCuU7ipYw8hBMuriCXYMqS2lu6yaZ62X6AoXpDH
mrQIp6P1lw8EVwQl5qKRcfBWRoT4UBBYq1s+A/32Qryplb6fJn5YqoPFE5HATik0KUpI1gJgv1GN
ul24hExPaG/4WTlHb7aUtPtf9LiAheHsBb+Rr15tH7232R86TNn3gvpfs+sJZ3eBWJd5B9GjOmgV
KAApGdzIk6ET0pnKfslycKihyHDA8UPg8i+4p48EuZiufyKVEUjYe/DVRTdE5Fad6Rgl5b2MoEsQ
Mz7bmwKpmTQas+/8CNDAkxSH7rZwnw3Rn5BYP0lR49DU4SQInV+QfYdo5DauLn1mvGjxk6CD9i37
LfaPjgL0V0KxumoTj9DS3HkxG1UCt9tVF1i3n0YYFl15YnsuC15Qp7x67ngoyMRl/4Vg2hbZdw8r
6Ivcr/UT4M6/wkGQ/qHjGwRu1t+bZPmpWDNpLnb0XfmUSWZbpBvNEW2Ab8fdXp7BFVSGcuBApnJ7
wA+6mI7/A7Oe3//Qpiy0GlE0pXB67mxDYRmUwDZt5fwOhCkyviQ8v7tBLoNcFZSDWmY5jHtpB1uu
1wdtmjbvEaWgZfrS7PuRk1eTa1rLFOfs+hCxmMkIv4x3hgiu9Mv6kNUDbmWFSoDJHzopFnkArYEK
UXL6pzROS3kine/sODaBVak++CWCFjemlKFaHxUnoCqQgfrqeAc4utW4l6N+yLtSnS80AdkoXGe6
/5ez7LnvNRi4751gpQmR227E45cjKio0n70bZuvxvgGsZDnGQfbgRmaHCcQH0Z4nClC8dES2FYpp
7lqj8ufmMKMHuRXh8KlBUYMWnIlgeniD8jnNa6pN2Hf+UZquH8xAwpC3iMEmt0gvd2MZecmQwtIa
gNHQ0NvuYfIk6WP7j9aiiNbgJDC4KtEeJUwTiIhygQePSCr+cXRjCfjuN1N9SkwkVLxlGyQmJLSL
primFYRabZUUu5InS5RzGbqR4qaAg/mPSaa7rl9uT4mbED3D17z2AXs+tL2SaTiBV9io4igWJ2nV
vwGAxIEHQqocutaPH8x86b5SLLIMJRMe3diH9hzGqsGWdSqUxdsm+zaBEUWHnoH5L/cz45Flj9KF
Fh6DDxMp2HRn99cf217+nJRCYyQLVhKFvWi7SgN0MTGpOZ9MzIxjWDwPGb3vG49QhaWZQzcBP69+
85eRFjNPZ9F3VH0J6FirYopndqrQItn3OtuFXS6iXIGFnEgfziWjJ2/gH1GPkx66NYO/rjrwacI/
lV8GNGlAppVEmVbqtPnd20+esaRS6MURdGtonZcQBLtkEHtnMRpdsEjYzsUzZu1DDBpNxtT+wBmu
Kf+d0wlHgnGrfa7t1emBwO7tI2h8tVRDAZIa4N3/u+f4NtrN8VJxe24Wjc/3/1Y3JGOzIUtB142/
0Js38IJbq9vzPidr7uRhhCYJ+lmW7rqJeVXRMMeILYH/TiHMwWP2Y0aphXpk0AreUKdJtJTjIaWR
J9DmM2VMG0Sz8rJ/8PDJylzjGH31P7xDpPsYozGZj56aN0Id7X9IZPxCNFphGc71bHM5z2GiyNja
W3GssFnGZQ5ols6tJwmuzxy2lsGnd6P8StfabU+IriR31eUkG9U6thHUtJW/x7//9W6L2LxF67W3
I7YGsCBeWwmg07cxCg8bCtkvCijSZiQRabvEcNpIeMPwR5g1GBlhp4DXIWXFEcCsjwCyFfy7i9JX
eJj/P73vxCVi2q73bPAalzYKKpHcCgGLf/sWvEMsxtK/+BK9BZJ6D/Qe/vBfofGUH6q6BzA+y/K6
orhvYjzvkccWaeMvMH5ILywMXRwW5Va0cWqpYwPQYI+bA/vrImKOS/KrgHOjRMWV+pNecIE9poGk
obVLR8n+JeH/OTWeXXJe3jkzYJA3e0RGfsJHPdbIJ9/cgHxhDd91wfLL/nI+4pVvsvVffq+D3Z5Y
nHXKyPihGzq+6JdDGEyajKO5AEC42AJmiXEQRVE6NUrndT1mxTticSghJBz+ott9loSg50wzlXar
IV9/AZATtZX/w2qNIfVKXXwVM01e0HWbhIJBuu/gjc8D7PxS6ngbf2oVG6YnDUF3/M5aXLWy4OqA
Uj6Kwb7VCvxkB/tPkxqO1wk1iK1j0t+Ny+s2yKOl/fNkkRULzt6pQ0s0pQ+mhAw+KMe+LPbHPxRV
EvwpDt4cZZbqA7U8LduKvv7AGmpNg78indFvBALBEj/xHEHkOO3O/sHjya7aCNlorUHJJbxVTe9o
xg12zroWGsYa/NTvZkLMnwn6HsPvadkHOdXlWHTyqkXll1VZrbiWG5dy14xd3O1XDImHFQVz7SVq
gRJyarFXM7pvxVVGlRBDKHUG5Cs6h4x4bx+iBrmJj2Fg8/vbtYbv3mObsRWKySzrsmqvi4I0vPlB
jee94H6+xz6QMGWKmGb72ZIOO/2xqpgl+iJl2HvfbNx/rAdX9YcdTduDl1acIdVZiTLzaKZk7Q8H
HMNvgLzMu8qQQfiw7LCr/Tnik5l5NOFZcTykXqL6YXwpTghKVqPz9nMY26QH/vDUk2bfdqFj+pM/
dAchr9VFESUvPmycbt7cTGBqfHsq6ZnhHGiPEj07oOV9Hr3jCleFo/I12LN42dEqB2G+ZvPhFw4L
+rfXmbp9BDoknWM7eqU1SU7yMEkJho/LGVR/F+1bxg0u3skmErlp93oCROxhp7jmyT7YeDRAL7xr
ffijnKXZ3Bp16zi3e7LUMJNET4HvvGgmvd1NLYuRQ8RMeTO3Bbkh+RWGSkc6rfbeq6JrxIDdDJYO
Kvc23MXVh+L1AZyQKEmpvqzkflpWqunTXxZ8UbPG96hghd4jdUEeKV92VoJEODzO2d60VYLagO/9
GNBZRcJmp7ae+xOSfrHQfow7fJIBbdM7Tw3ZS3KnZv8l4c1esxSH8/JfBTEH2xw9ryrdhslTxQ+p
RXywNl2KaWydVk4B2EbQmuS3pmNuA+BmFRIoKDyAiO+6nUES1ACtxznS2Ul6phZWaUYy8xsuREmf
sykOLr1V6NXJ3WC39G9Jo0IHcDbEx3qGhp26guiu+iifxFbEgrc68BZ1LUFDd+aUFwNwnEW1cv3p
ZFJyv/hzqqQUFlZTvd+5CLmpio8qOeL5FZhAS765WDt8D27migvxj1AdPs28zf7ZbZuEUZVtFz9H
apBT7iOrgpwUfHrtVdjd1vawZk3GL7ik3c8pU9zQBfATALo2eGoIxn16FVQwK8qYepk7J1mRCwHk
sf/ClU8zVggTb736PcElfl0W3Sy8Y3LtVZKBZzNsn1OM1Q2m2HWf+oJuX354pseEyJwcbJ/TfBMJ
VNBI03zI7w0yiyk7aV4C1PKe69uEC6HpeMBG2gxgF4XiCNhHHCaBnrFDM4hWlKVDzRWbalEHhPpC
EPxO6gIWaHSb5Oulh2o5zVtXndK5q1+ChAmeOAypFuaAdv4j0rH3/TnKp254OOYGaxZilGiOpnHp
l3Ro+unOcVBTDLgphrTT7iutrVEVUrOY1fuittJfhzICuJnJYmXwYAEjlGxvhS8KdJ3dsDrLOrvL
ALbdEDvCFr4gMwQckVe4nYaxuo9u88DmgHkNo3HgNOEKPpKcbGJtKkZEurEkjdj/lWFTn3fPhTCy
J22uAMolmJYX91O5HHaQ/F+IiXl+X1+5q6rxSqOClPZ/rmbm/jLxx2NBfJNn9RbRNIYGynQZNl6M
4eZJVMkPs60VD/PpAKviDffvvDHpSRS3DoEAqNFuHWXLAk2ylOCvUkdWLnNDf4YF4tQr1V5cVBeE
24bI59rmoqsQF+q1OyEQd22rX7K/bLgMBt0eW2K6nbjfdkTnX21a3CX6GrSz9Xksoyzrb1krgLQQ
uvxBJ5flM9eXBNbs8D89GX9Lq4y1CyqZNOQKxPIoYuK4PBqwnJryFWVUJBPpVZ8xQAfgyPcuFIVH
9PrA3MDWWlpPW9ae67lIdYUEA66puMM0++Ky42uh1eslcOazCFG7OkXNqML17ZG8G6yNraapd91q
k9kvXvXYacd+corGON8N9F5TKS1jOf7dIMP5NEGlPxFsGgItr8yQX/6j+REEa8m0XwnbfC9+p+kS
SxoOGE9QfXBor0tHI9funS1EV3ugbJVIz6+9jHOqWCahPwpxXBHNDN7QquGSS6eiiggNa7Bpgmjy
R4A5/sTFlql9izDDP5F+dJImdCIAuWr2ft4MkLmXoIEjD9R0H0oAYCbqbmt/v/pGR78yuLuU1PEl
fcOz8OERjlhGWKIsSDEdI/PTIlngh6SFx1K4qPmBqSAcseM/pmbbdCSMcPPE83axXpFcpccTL7Ke
sgaj6EVdCYguP1tOPFqYAZQt+0nGaAP1IRyGhp6s2ikwlmMJ4nztTYTpvAczjg1FTx69OfHOglWK
R6BLAa9Zs0DOf/+nhiFMSsgjwSzULTwUnwVxarRnROjT6kGV42W6hjLaxrGb9V7boAPxWzLmPZbq
C1cPyTFTCnnQJ6H6eXNasUrUxxcjZk4D0lgm3GzWcdbE4rl75jEkzqrDskdczc/dTvkZYJP/Dyjk
PBwu8jz6VPljIq+Jiui9cXRfRmm10z5+1lYakjMZJelfOpcT+4//nWwp0iyrl55XpySe3nNRUlYN
i17wlrBaId229ryQHSg7P0zw4asQoox+bcHQWSHfMxBQdXwsnHrYrNOiLzVUG61sY7NK1fkYJlKA
PsGgj2zwazL9xiXYonxBy3dP6OBAygbvjLIJ4sRzPWxfF0Vs19+SofjXzkZRDrdixzMGyvF8wH+3
xGyL7LgQ+T5p3QtLDbmvqWtNglmJW18T3EVuS53Vj26NVUREMPqkKxQlGG1/ubcvHOKT0HXMkPUD
dIS79Jds/t+aOYjNxuXXQFF6I4cKjRi0foQ1xcTXK5cCVeVONFCrpQ+VbdAc0yORbt08so0PD+gt
uGHJd3AqUn5ieoV6hwBKq+ZnC/Mc4TGSx+9zQ5XR8QILzU+l64YjDdrxCmtqGU49TLLAVjmViRuV
7LoyK+ezzwj2FSjjyfsM6BTpeGK10hYMiB3YJ56b9GtgFbmy833EM1WA2DaCfYLAntb001sUDuaZ
VfyMoDUmro09PR0YjTRC3Y/EhsD8ovYI9J9M5CWi7XSPZ0hf+pH0Al1TsdCTatUWbLvUHP6k+Er6
BBsrptJGfBY7vwN/0dkv9ArjBMy2XZyuol63WsrCZWkQkJQiyaoP07pqHsgYmIFurD6L4Vvo+boy
pNBHhY/VNWV2X6C/q8dVW3ugHLdqURgm1/NzWthSc5c+ZntgOuSfNpa72F2jJdi4ny6R4XV4TBo8
XxOWyNi2WoGh9zBCLyHPbScCAW1IMF1cbLKT7dFPPB4jko4lkUotugykPSupvy3hOSC25VCnawxf
3ybLBsbidLXZ10C8D6K6jFOvRtwT3DTXpQ4Hh+rWQBtKd6cLuq9mmRdmproWbJNDAWxpoAx0pHSW
By4zUe9LZ5BJyykVPVmo1nHFHcKCnmGmVGmVXInGJqWaJq7ZlW8v91nsY1I6K7hxPu0YK6MpSdvr
O2piu17FiA9SBEeWi9ISnmNs/1tJItXmWkIupNccoR3Btmldo18sOVMp5glmJ5JO/yQkDT9MXS7W
W/NHREc4IEWUHeHyOzoHcEewWiYJ03NhF9b/xrvdYuiqQis0KX6Ju+Fb53KYcNF2DAFtPibFqcT/
1PZb5SKVPmM8F+SLwXJWSW/GYjr68DunVb0EltKZ9tNo4Du1/WFEkVwTA13Rnf/Ybg/+NP5RtShp
gJTo+8kF2FOIOwV5bzoqr+pCnsAToIcQo+ZBfHaHbWehITczlqSzPQWADq4clMIUmpAj2xQzIwxH
WUbhnoUPmUXLNY2xlRNfNd1fWCYYcrrh9kFsC90JVn69Sp5cOFQ9Kzk+BKJSGhRYaR9cReuM9GYN
d8PMC8NEzDhJtWPnE2MXFQZbgk1wArTD1LA511REzdNQ5C88djik5QzWdyrGHbBc27HbrbzDbgWo
AcgElnMXd2K8/lklm8a+rJnLZyKEab/X7M9fCBouAGWOaiQysyqfVfEeawoD9I40giZ33Jrt729N
5i6rrAahqAS1G68LgoGCl3q1pngExJoBn58t/4s+zvgYwRJvqlwpNyIichZVCjmXBnRleSlbezJi
Dfc10EB/Z6ikfssuFDgs84HUEROF4QuyTyLLogPjuD7iZN3X3lDKo7Khg1onJJM/rhdTUAdB2j03
ua8biZMX4MBVf27HURuFy7S3tFO/6EfSiS1p+PPTAMt3grvyrp7JwtXzQTzCqPlJWwwykhfZVc+R
8yNhPq5NYkkhO2b2xdiEeaFYvBRu1PScMYw9643IMlhtfn3iOIvY1p3Mnumi4RUCL6jd0tlIzL4C
XTUUE/j3vswl5DtRrJTuPllva+wsiVddSepASpoAfs6qbP0xYH2PX9SeasYbPSjBdibv5fpu05un
rLD3EKllLZp2xp0XfuzPVyHAiH+nImjZXjaUChtTeb2F4A10CQ3w8JOBGZXnaF1LoonK6BNdYy/e
PBekfcYOcEs/FAf4Fz5twpkWW0M1rgjqAGlcq/EFT8jd0MhZmWK6UOqDC7/a8SYofrZcTxTQtRZR
Zn07KCKEf3xMWw/FhwdtcroXzP6f0TSfYmJsvddzb+eerZRns7atyls3EAHWwYF7l9VywFULag5v
WIa8B7CJAIapifZxp0QtZGJ8k9fSU8C+6auOYDx5fGDQu4eGXxhBjqmZCUr+8/je+gO2YxTkltkd
aBB8tm6GTQKXE6RxiU2uyuVfRG42C5i7A+Hry1c96UKQYw51P8zIkukn8UVmF5x2Oc5YkH55+1eJ
LgIzH3e3QzX8pldv2jOD0ux99W0H1hEwVywxhOOqPZdQjtCQCiBiXk+Oq4SsycweWYTa0ad3N7w8
BPN4OisMjrUTkPQZ9IMEt50nPnAaPweF8qD4i1M8IRxGBdsK0fXZlRSfV1L6rPPsI5K7erJyzNWX
jM8epuNdO/c5kP0a1w7dpIdA+W9id8DmOh+Zj42JF88Jo2ZJsUYsY/6ufyw9+9P3HRLBvE61IOJc
KddOA8gsBnrPMrlVhsl2O4eVpPCdvqvAJNKegc1m5gCSF5bLbYUuVHBPhztIi0se1rnspUsxrtOD
dkluCKxWdS5RjQkFZv34qU9CNUYhPxTfXjSYKzlveVX3IKWxVkgh411L6Hm+Ug4LcV9wYTo6J03v
sXBKLav4Pxv8g3Dyk0d9TGQ4ZX4O+ooQIpfGejTzFGH+j9uIatBwk4VtHEUGvBBya1IAEnNABgUV
ql+1bNJV9GZSoAYUlqF4WORD8d43TCqRM/1RBMw95y5opPuNaTSsyfdCwy2FSjKSEon9t6GnqDTB
rxTdj0gQHNsYRUS6F6Ap1adYMEIwWDDOB1z3NlH0aZJGEdJeB7X4YOULujDtgBL11csVnz3jJeg2
k4+qKOMQjt5eP8OkRGeF0+wzNGACW3kXYc1/gkoJsLyVxtuUWVms6KYcHHEZzkNB36Syq/Rn6hS8
ZXr7HeFBVi4Efa6Di9nBFf2V6RmnbCnYtN4WjltfrCUzfbt4tzVTOWoMNYD1FYF03pCJ2ocSTg6h
kB/X8BAeKfTdwnuuM5+QgnZOwhePvEXXF/jYZNiNFNTWQbw7k9sTGe/KAnAqbHEmUqDcjTMBIWiq
rsttZ6aI9ghLWkjpKWVRqMUQGaLyR+IV21XVho6iZnkUKOS79UZM4PjsG3lm3uVQ3ZhuH9qSSQOB
VIUHEjSFDoQTh7jqE2E9HXbtGwAogSJaFuF9VUvrk2cEPqNIOY193fQuERFBarz5keJBLOXjSxp5
o3afKSYQmcoN6OxszIpQH1FM0NUpDk3J5V/b/zfljhvmFfJv8RGzPrtYvQWiNMgVpPZV33LC4Lmg
9ybqAxZqlkBrixwmVAaMDwiV0D1D900WZqihEfLP+DrfZzG7mxitFpF9B+P1jtcd4+d1LvJWb7Yr
4YkBP/y5fmQY19h/HocQic+r+fSYNp/jYgPTNobE8HqxjFGZ50I2Vc++wZtRbQJeQYhX48TkvTFV
EdzJNXVZRnkR6pIC0QthvQUk1yzVuJ56eCb6+2fMmiEtWV7Ul5/FJN2lw35FNpqGB6dkn6MZb4zz
pYgAQgdOOC/rceaAG/wqmY9X6AOARKXERVNJhz9w7Zo7EONvciMtW471DscM0X+iwENU9f2xafQn
/TYRt3GIx/OTMZWdGVRikKHk/qF0kj97pSxzSyE81Bm58HHVJiHtZEP9LPp6guOtRvmjG4VLbwuz
FpNyB/bYBK9gkGJYkmin2+8ak5PXZfmsR6tJKStysuUBe7oo2rNuPTGe3YbBe4U8l0FctebTS35A
CIuralGQ9lk9y+XGm9NjSzsio8eGImrYV9L/AiizCz3/U0wv9uJS3bQrkLmzIqvLiaMGE4pSvotB
g0vjYNVc2AAN3t8AZQgdBtm/HMd0vg9A6MqLn1O92Wcf+ChQ31O5I+ngF3T63f17ylvE+5bEQCrC
0ujzDH60s52p01Q1uKmpxIfb1iFzesldvyxiov9BOKRc/ME9j+7vb4AFW+BDsLTyGP+Zx5FN2oCm
VLGiYEi6AD0V8uwy775KFH/VALStCvAIrJ33wXj67sC7uQKno2SXjFXpfXpZVn05q1Ujeau2h3WV
5hxFMEkU+xDigNXJ5pYhECLpuG6k1I/2zN2MaTvKga6h3SBZaA9dGCNU+cNRTx//l4PmYOcQiCSz
QnVuHpNeebNSNq3Yo/TTb20hQfNEi8K2cUqlRQ7hCMb1/DBMtvCD385+NQwTPT0DpDxMS3H2rVpO
aW+OvnXxSEBgry54A3CSvAYdZvVFyTBYQ5r7DCEazlaCY3NTA58rwvk8/F216l4j54l/c8bnypyM
Z/CgBMTUs2WiD4I1akwmSml3vKk54KitEUhZrO9nb1bDWQzxosMcCwAEogbeDyMWiSWAQHs8+SIe
8j/YpNj7ulwQ69QXt9csAD1NosQfkJcxNgan2kNoSDn9V9XxrbIgsA2+G50e9T4Vl7qDJqJRt4n6
Ic4s545E0djes+fGZI87Kvrt9XQu6LKuzTGFSa2eAYazRNlYv+FaQmB6Ras0A8GmVJ9yUcrMKfbL
N6od/2rr5NcYaSLAqW+YLWITev4q0QROT9PtMtwdz+JtLuOikDOPwHOjtBSVbXaRqbD1g4yft4En
c16ysGdGiQuyiHSM+T5xLnVAERuObavUuw9tEwDqlmelcauV1hcd+jLVR6RrGkg4++O/uyeWc63e
OdNdKDpZs7YWjymf+MZUWVrepptIS6hug5JrZ1yvpIUiKebxHggzwSbnUTyaw7emWvI/gvGYJnKT
LUIYSqyKzhXB4zUAiK2CCVDPpXmkhNWkrT2gX2icQDpfCo82qI7U+ylThkzYurGXhVP2fsAl8x/6
0/UT5PkH4AbgD9sxLx2xa9GQYWjhKcozgg9K1wd8QvLFxHNST8grofYyK/ufsUVQxbwFzV/+kI6r
fb7xFB6uQasxQWdLjOAQ9xIYcYCAuxM3YsQ0cnWaEmnKFtKJt/uYM8x0Qy7jmaj1+WjbOtI3RZcT
UvtJl66kyXK9J+otYkdFp6xXICV8l5QV1dfCHN6c+ACNJwTqxe0/vO1f+8kYGBsrcBGM5qf6nh2u
AtFg1pwIQBtBOrofoC1rCbYgUetjRlkLMjWgn2jRW8RTc3i6HNJ7bBQ0KOTdan+/EdoamRzAADMW
cw/bo1ek0AUgx9nDLtec0pOrj7Ps3TfQ9Fu2oSX5fYJhLqGOJ8DBeoPlii2/SPx6E49a3/Ym4qdf
bhBmKt6Mz16ulcPa7C1BFw//gIqYNj5brWyEPnklE+pSzQzqQ8XyBlCShIokifEv8PSuTtLV5xxL
aLpTLr71hTLaxulghI7n7j4tGM7VCFZNNLKiyV1sjSFQCDfdzI75xmfWBIGcAclWT/Nmxaw9CkbU
kJOwbChmQ8jTcLFid3AcnlgFyMW3b3RMZ0KcE7t9rBsbLzT/Qo7ONlGcJWT9NtxN67awllCLjehE
fm47jwoJOHKmvCo60NIe4NP0idLNQD5PI9s/05LzF5WjeQAx6y4L1MMLc45fVuU99qQ9AOJ7V9zP
4KqGGN3aUlHk5JaBvJBj9+A7moUrqlYXYI6CJurbQlKZSqsu9bAYsHH8HgKXdIZpTuHpQzYTJsAU
2hSPCrhWO5Alsh4xEOJz4jb46LLGi0oTjvxaBNlwpdSTQaf3ZzNCQvqVRzLvZH0pkIL+u07lrEib
TcQIynTgpevhhw3XnjDT10KGBZc2yB4g/GaWYyDJwKkSM6hx2SE7dJO8H2cEZfVBnWbA1zTAoIet
/uWxwUNrBNsPFDKQfvUFye84saC+hIr+8ASACNMuq7XSDrKEPT0fg/x2SwV733TkdKRbvIgC2cOg
co6XGK/A9ELl7p1JLW8bM5KDI/hnID4WZYsHU5R7iODqkp/HtM9A2UfhuzRkhwlEJ5yqOgFCIG+T
c7uDjIfOQopGoGqJqDyM4fRtVAg7E/tQRrY/uTiEyIMXJWlePvE923z52tYDmK/+TD6FzShiQWOu
dcZyAcNHVJFhZFsQUfXmN/du31ddeBH44E23gPq8Dv9gO06uuCF1kRsHApWDsvSb/EfY8j8b9G2V
1M7/aAkMK+DQRmwOHEThTsEBkBQz+q4qUcUzVs1i9wtZt/DcGgoN2aeIplo4MXQv9kGmIMOEDvOE
Tyc8s+5ZmQzr4A9eDLfqFz+uKhWJBN+v7P77EF2o2qqAhGTWU3/lvrxPR9+ZUaEuFvPzf/i2j/qF
XLnp8+lQTX+jx0N7etbW7PCXSXbQcgrhxzMG/pqrJcdLqzhddt9gfrzJMw6u2dQxT+8F0B3QXwBN
Pd4IqfFkkE8x6ZAWThedrhqZwF5D0rGCNmUZLQ1o/C7eDH1BOSEMhKdQtj71X7M2WxricCenk09u
7qcG8v+hYHEk/IWrdRpcRCpdXxm+DjLLrq/6TD7uKokyWyN8eoo3b3mu1T29lSBlVpyQUZin+R64
lrfRf7nHUQ/lEfcJIJVbu7bQx8E1omRTO60JhI564ZATmslZLsIpVu5l/gJ2PquVC+aqRRzzNX53
/kY5jnz28ABxysgi01oWfzQXDaBiDHhbh6Gk3WrXc/rYBPJravbmPy+1FtkUrvLJ5/uKQ+rxhyoL
EFrkddcdaedvdQvMQj/UIigbtlhAxDq3KNngjT+KQom6jRr+A8++c5jKOn4671We6EGNmxCcJnix
a/jVshg3lyVidLYh5uopZVzEYpFBYgr6cGIQPdS6M9p6yvgtJng+2oWmS29eF5iKvM4lcr+r5tFu
hb8l8BHwfVcGasuFjEHdHp+2SicGQDcKy6zmnFpdMLQ63kluT86Omcm2KCOWfDlCgs5ix8nCf16s
S5Ejbb+rLuPaA6d89CCMOH94G1X9df4bprGLkymFhqG0w50fGDsTSbtmGqU5NDpdnKx9YFQw0/Cv
uY1FNB1mXFvn8innnXwV4aYK2LfSMfy5ng99k3DvUn6y28/VoH9Ibt6q9pr8vRis1FevTOS2LX6G
DzeEsgIz239rQmKlB0X7CEk+wWjgLPtWm9TTZ8UYXD1o38mAU6Fsz3sOCF5I/4j34E7ruaDzxShB
r5czZranIJOszd0JaqAf7mYPDK/Yy4kpuGkTaegLm4eVDgclE0QFNqBkekwmh8UfmFI1epUkury1
2uQCCiLjQTmxGUPYHbXcxlJGXQr6XcWslISyNaioaT/zy3Jb/yNJiFeeZ3lA4WgKmYAaxSNsfcIp
XaEBxv/pSQAVZPEmk31ZWhgkN7egxTr3TgUnQE28zZtrx6HOjScLQhyxxuit0tIDReTsTiVL+W17
bbwYiv0j+1nX1QT89H8dKqHsjaIHT4n48fDst1uxwt5tF9XLPMwrNIiu9vGlVyJkul7awjkfGsDl
AQvca+ktzn01pVW9ESo/CuRCapZ2x8BhsCbolzqRW9KzsW697puVN2Tee+YJNK+HhqFOiVfpvd0u
g6gZLDVBSn3aePXIy7BfS1I5CWuDLooxnRUqFxpM5i2Viv4MQDXKsFjGXsUJQF80GwjUTwcN7jsP
tqV9Y5qigEBFvoAYzJjaU23d7E2hBslqklT79/CnZikXaf3OSaVC1ljdL0EF2vdwfGEH1H8S2eYX
a4PpV+OyGslUpmdf3Mt3BJuOxB1W28kS3sEUNIwV9Qu7eC2TZfqCJmc/dgFoXlcBGIv6Uj8xk684
9Y3/oCX+/jzeSaFhX7kpc9nnRPTwHYw1vt6mY5b2b1xmOrgTNQ21qz1DXhSg0F5munTeKgzI8eHy
0huuWKbE+BLvR5WrKOkRDZA4PVsH9mfDRw07AFm9ygTXyT5FgLncVibSmSWKYOVs0m65K6QMzi/D
egvqiak6fhmjfcxx89B7QSAwToqGpkJgbc6y2DMkQcSXWLS4Vv99JdoiJi+ap0eHwo4++K2shW+C
Cx9TAHcgw62IdT3glwcHYQ6x5wlEzDKVVFdv0aXmqgIbEgN1ZaRaagQp8H7zlQwMVdwgoZ+l9z3w
hyRTubc6pDF+1mppvPxYQpdNHG2kicPgbJZqKp54R90v+Khz5HRWNxv4XJZx8V58A5VYgVGG36nT
o5mGysDUqawmiVZBG4leAolX+doU8EVmKuuNxDQmgG7VnCo3rQhy2VKy/hLl8/1A+9pWpPX2K8xu
oOY1IR4d8P6SuhTLnCfoxYcSu0XBQwd6qkxsbzmCEmuFBkImm6XwqKbaidB1gwXffYWibi3ADEja
PVyfJRkFAZ/+1dVCpXHwDAlA4SBbKySoG4vb+/so5XThIldni6k+R3sO+jEZkse1qgaeLjKxZ4dE
t/CDWmQO95wpRDiW0Oa1cOv9LUo+AzAhEtZDwjkjSVgJNjJskmK+RVRLmCjYCswU2biRcWMc2iMa
VTWaidbmsG7DP1RpTpBolje7waSIgeL6qT7HNGkd26gV/9wkKghzGHPY/8KnH8YMXzS72Rw0f2RX
qtDNeuYBtdMB66yTaGUwNcBVBYhp9g5AoBVmoT9KnkVmxYPw89YYlHjgUC0DYqeV6sUFrsNKqN2p
tEoKY+TY3zI3FiQ3lJnSUdq50sqE+eZjUepOSR8tGI94hzoB4ufv2e0JvH5l0cb+T5eLBhpX/ON9
L+ugPFHmTQQX/fiwhr6pEuHWW6xPKFsZ+f99WaP9rnL5ky8QpCzhIJZ5r8a7yXAwwOZf76ulmVov
Q1eK1M78GxZpdyULb6LDT/TsHOJ+Y3RpDIxdQ74vGjpcOsvF+PTcEQMtn8gPpNkHDSjK5AxhdPVU
nhbS5KMrQZpKcv+ylD1h6x4Xxddz9IGlFq7msUyjh2kFylbMwRpIxSphmIvmtP4nSUEsacG8MdOg
NUhAocu8GDZevDixuLY8ahAwPMAdyW6ATmPcpjmKhBFrLZiFCxv7mSNjPuIVFoqNj+QKVK+Nd5rD
adl6tyvmuBmgkqES6lqFNTL/Hk0hw6uvXMoDJS8s+fKmXFkut2WRhjv4iEv/OQvMImdk4bw9A8JR
5s4Da0sNuB6rrfOvFBV3pthHpvIW9XePrSffUXx9LcP7Eqc6G1AqQtgvQFOos47Dojv7IvJhdUz5
vw4MdHtu8yIdEUYsoUE/rvtpMqRNd5od+s1tGwSQ5YVMSEOoFKZnSKGfuadR11qNGMP8kjBqNTuH
Rc+uNcHrB3PyQJL6kbR6xsAudCVW7VR6pg/bJYVPZ8souMD4r11YX1g9KLpnn/x1UZ7gBF0ed+Lv
DOef916QpkAcAwan95XaFKrrE/JSCSLrc33HzfADvLtE/r0F6+NYWhyCQsy/YSJjP+IGhnxPto9u
3wJZjhKpKZKQG7vVKx/fr35E6kGZpDQ6knVESnNcIGCEuANPhBYmdxcQXPq782BmqRTOlBYUHG0H
M021xxd6FvsdgHKAkn2SLMpr4Pm4LjKEhPvlI48/+5mxYD4EGzYivBWzjgPG3KwAKbrL7McjHAI8
MICeUj9/O+4/kj3zcisOVsbmJlqFMd3/ivLUGDy2jSLqdzgCbF75IwSchKmYlJJOVOQNrg68APl5
88TbTJCHYGEg+pPuBzGLAQufLiGqdZveVOyrCIXAJcblWWA2WAfv2sk/cJEFOFcJg6Vw4eepbBbE
HdFrtg1euM45lTgkAynDkgM2GsLYIGfq52AnLcR1cyIrNucYVmy7xXiQjuT+cF2KO5+elBNMZjH1
KazUVO6zxAjZcqA/bQ3USf3RB8iIrdyHVSZN5zPcGKrOiJoRL74cKZDjybCmhaHtecuhiFa6PhFf
dEgzd3XsUr4fZvaGaUXFA9oOrdLrTtwfIV773u+/OKu8a5EDUoDyJtHGvY+mMFybtYUauHxEGvTW
DKJgL9mzku1VXvfvUzrnKaO/aAGjSTowU+ZEaub2fXAVjj18xHrlWm57I2tiEb96o9/b/s8VG8+t
KG2A7GyuwJ0bjX3T5DDtQDv4Y35dp8PSRuGKrfo+CiS73LtxelPOCp8VrIajUrm6pSoLnyTNI2dk
ylpmjuqsAsEODRqA8UpGmp3UP4FwuIHZXuBoQWsFRgjnVCMvTqXFKi2QBgGeVe/NxZjnm0H9tJTH
4OP2BpktviI6IvHnVJQMA+LnHrliPQ8hDHWei9pv/eVh0dpFEB1KjnBi0BScZh2Xv5/Sj6UWjvrI
XLapzYGlJFnYpWRiVytFsgPQEi+Kq7074TbH6AERYr8LStZjN0Cv1535NLOAEaKtkvfxIJR69gE4
ODjMl2OziMAE+KBVs7hHYRAFcZj0yU/fvDDoPqDKfKyzwyPlW6iAzGPA6j+gkvX8qGcIHi1+oTd8
tvcOMkgDqlkBDWiSbTg05WeV0p6sefSOHmbd+G0wRWv9rWy1PeEYHF5O2ATVJJItlPgXub7OYEkI
lqMIfr2NPcWgMoK6u1ON9CI0kg5fPMInex3eZ3ud8Bb9dmkRIJf+86WyWwO4+Atdez+GJbwGNcNt
avJUrL5PMTnkDCYuHwpHoVTHz2y/x99OaaAsQG3OFM9B3SCNXo04zWBGFIzRrR4l7hkdBFSbJT8J
djGzjv7+CDq6cY12GjsRLvkA57eLaKE06TiQ5Rg2aaUF6meTqnCYZkADLzo0re0ePDC3l9z6cDCN
0069c2Bklu03BeXqx6k2oBYwSN3erxLASUHSt8u8MvUF3TlDFY3NVt62Ry25WDhUBohAsDMwimjd
PGMkLk+mzz/ohwYt/aHKw7d/3PEUxDfhLJkMDml1RfOJoi+LoUhW429Ey97+OW1JXG+Cn0PipQjO
ZMYrORJoDtd71xnpApfuj8oHTMG/21iCYK6zd4lLLBqiLvbfcsfxdHdfaeF86J35H6loZ23sKNwy
kMZsAO4XGr5ozuoNBoeZ41WkslOwSIaTvvLhCFAEBBv4s16zcZpj/Xgd58oqAY63xLENHFb2Azrs
zneEqWme/vLMK+aicZ71P3gFpmp1Fs8ZBLTxP5ZOi8rs8CYvWdHd71G2BdGLpOe0XttmtEz09WzR
sXIfcdia9nJ3TshxPsEY5DnXm3Njuk5ErkChAs3gESiv+0NKdLpYR1RjYjWDBW+T3NzLlhXxHyaD
Hk0uOYa5Ls13pSbJCXnAzO1zn70+7LCuLo4UMSCRVulJdOP8Vl+jdwIhjqmMO/xWCcuHLEAgjlwz
em6/C6KC5j9Pr7hW2ZlOAT5NG9WBBTFqq7i3bKA7HVeWlE9qjcVu9mssOYV8dDoTsb8bEisRt7Jb
FsHw9tu7s3imSxRkhu7rY53uylFsRmy1V2d6oHEVj5vym4ws9OLxh0+05Ape6NjetfeHrpxAC3Mw
+NdgRWIz69nvrkmf0U0jXUDY2kd7oJszeqfbKsvU5m9ywqFNSwcgMmMFgXlKS38qwg+YKqcfyDqH
px0cthx+DbaqI/XZtf5OS3qyfKJDTe31Koqpnqp9J+JYE+y6gYgPsYo+xzPcWo/Ygql074ZQPFN6
Ozc1eL3CP2bE0HvUeVm2bvhuTI/S4viFtWOYhXPjs1O1bAIsWqNyMyYV0Mh6oBheSxU2UyATM8q6
RY/YbCZw7rpQ2JXbg84jLVnj5x14PnIy+1d7XCWK/SH40zMDBiiL1Jx2DKPKJ/2WXJ9Jyfon5O7A
gKWaG3CihiTOcPWjDfZSgOvAfZVQ0FHeN42z8heYOBLQ6sKKsBQD6sa74K9uhkSBhq6alGxJsYKX
j4AVzf2IqVmR51XOo/baDWOpJpBzUEpUp9KghKMMJVd80tQkB1UHfNJxjsnUnCR5Evrx4cPfTdhI
WMgYIJMb6wbtt0QhQlxP9Cv2Tc5kH4ZkMEdJ01X9W2X7nS1XxDfscnkfhd/OENAlwZm61o4cnLuX
78V46z4JhunI94mM4yoN+VMJk+FuTLbg3t2iasFMaVyF9bGAWhfaTAjelmDjwntMLilpEoqVfW+5
xWUO34PaUhyIFSQbd7Z+HZGe8/bXGFN9sOGuY2WMYFRI/2N0lPupcIzgKYt8LkMqdCtVkuHPflBD
ZYN/zLIUspQB5hIZAdysF4ZZD3y8YdRkqeVUyFIZMSWlefalsqgutVRYvZkcTs56wKX0XIT1scZK
4suNU7O6HwvdyZsoVdfPtW/P2GryiZIb8Uk+mfIXPOA/VgtUNyLasZ5DPPksAA5mhny8TkeyX2iD
4s1Q5GNxcnbYHfIGSgXbl79ereXaIO4cBjctJRhXLvtG88/7Hib09IGcEDXz0Dn3JdgEGGbvLWVF
azu7v/UnrFIqTKpn8wZmmcj60GsLqZaEVemthHbQrZGSNgip6O9w7Y7OojmnTRN+O7kkGJHdvN7x
jY27OlKO3BGIHXXLM9pDMfbG60tTyavukaIUJG2wwx57VeVbecuE0wp9NpM0FVlujlfu5s50psAW
KTAXlb8+Tqb5SL1MYvk6YAc4Nwa4md7DFKGbtyWluem/HzWXu/zwJ8lUSeIdKnosbIlmBmMu18g+
xs88AfYVVAnEl/FYUpS/Z0PRIFXT8+PeR4aJJnDU56G8nwTVLV1SRT110kqWkkjv7OV0c9z9jjVQ
NchXL9vIZAQ6IDVtQ8S5uP69mn5Jo5OvzEbM91lQ5lULH/wZbjI5f5OC6biikBaf95fnZJ4qSaEN
wTzXZg8SoS8gGA8u/yLgMsG3Cfvz4CyD5Ok54no9PI5LyDfPdGNfLYp33vjEnViLrG6MnrjF7dJT
lU+ii+/ISbrmxmyn3DSeVHEIaxdH6Yx9mpNFB84Hq694h3fuIG26BGLTl34KxBCg6qF2VhgOdh89
Myip962tAdp5g61e3fuABhTO5Silyz+9L5RB142khQqaq2gfiaBSnC7gzFRFuVlVajYM2wcx/LAK
ZYvFzFWwFHxSNG2haZ3vIQHzfnwER+lDL/JALsdKdXi4L0epEBEQr4L299wgiQY4JVZO3E7816eh
MEz2MSGSuaqKzfXNdeHoQIMxK7x+3V2G4fclOvOiClmWH4XI3tr8XbP5nKqAcUShn3mYiCq7X2Ts
OQ4E//+6wWzje+twYwf2m8Ys/9Y2uj4SjMLvptGWeIYq/rqhTtTcjzHFjhBwpmg555Jo6H3sU9eE
m4doVF0TTNFqIF00VpKW5i7qAxV4HFfJ9couUsgRkaPlFvJTfk7ieBHzoJ6m+/cgEVSSdR7MhgWw
3U4wKWdjaJ/93kj3zpF0w7z8i4rBkgx99AG1rmoAIr9ciJfwZHdEOyBafGTtMMO3myW0zKuo0MIN
fwzeWTh2mSa8KN9Umfd9JE0wY40/5Ns62FkRJB8imnXtUdsDDtTO8NhKOLeofPrtLHc3P8tg0+/6
fW0XwPsBLJBsoRm4suoUGxtwD8CDbTFs6gHRB8ORFZbXmNYFtB7KOLmfyK6AIqAyew5QaOMnEAw6
brcMVWcE0QbsKvBINmR7QsiasHXj9gOJf/8n/HDxEiJ41jMEGv0HpThf8zeMbvSuGwS+NXlhdXjO
0jlnkCBS1ZQUtF5NOl//+46TvJYq+f/RKYCQ5lepS9uQdylO7YdyLtF3r2azo0Zwt86BusvM7a1h
DXCls+xfPoXHGnYof31KavLyRx5coapU9ZlHQoD1hKyNgZUy2RCxoD6SCzmmQ3Bwd5LxRfWRzVdl
LWkUcwXgBtehtAWTQ15c8JrD7k3U0IrtFuRFrjd02xQuPFxyQhv5MLNgWtpHE+zGgV6iTfzI1dDf
GE/4hya0h/DdeLj2tbJ36eOqvdNH5YMmETEQhK8STzv5wnTfR935QWUPbRRByxbgXPZCSwjyqf5j
C84DuSgPz7G20/iFatEiqwPq+nPdinbeGbfsur/G3KymqcGdUTAhHUg4nr7jOOQKlP6y871Hibgt
EzNqfRj0yhrhIF72kLf9w2iJN+FtZil+loY30cEYabu3+Z4OyAM5bcIVig/jxjYmcUsWO4qaQ77p
dnxeVXOtc1fByFe+NeJIHg8IM0Mxu/37tmWap4/E6Av4JjTWsP6i8FjGSTZGL3cCvbhdCWApMux0
Mt06lFHBgPExMU1UrXfV+KbRE3wNjJhCIklv6LjixqGf+pKp4ia6nxtu3ohIz5Ui+pUGk/zR7R4w
AwOR1CWH9H/NTUGSjFNF1rojKpt44NkgZ48Dgfywo+6G8uJxDD66xtBvob+AWhJBagaHuLreP7R+
WIMxq1XlbkH4LLtRPmOK6seWLhw6jLP1bITQKJPCBRxJG4aQqhGKnPmCbP5VtmgG3YXrSZTHV11J
/83D9zVE49ncwBYdBKYWO+aVjBFkkZCgj5r78OBa9sbw626JC2MoFigvD1rvW1Kq3nf2bbUJ37mf
ptsXuU1GUMtdGVQ/mUPLtmcq58F7UTfViFauZr/D+Nk+Ru3HGviS3b3nVZ/DfW97UARXi1AF4lQm
a4AS1kAkjywUgWBs66JvPKb88SRmXcs7gyP0QfaLArIGATYydzxuTfX7I1wb06lHNfNsdURekl4t
1JymaYeivtBanVP5c3tn1JovbqMJGZMiZy9k2K3PyxUuTU/6BhArl5kPXNZIvTskvDeLhIRJevFJ
UtmibleuzkMCCu+7iNysh5srT5F14xTIjPzqP/0v+mmZ73n5tRjPkmZ78WN6yD160Lhowynrty2+
Ym9PclAw0dR8rdrpApb0zJBeouQwVgcMTBb8sNm9DMwZsXWZyzkFPMz123Y1ckEFVH2rOkyCdLZd
4nOSD3xMY0IUpPkmpxQcbOz57dmxR5aXTkjWPnhzM67JTA9l/49sK7ruvEbuUd+GnSGguYDdFtEz
dJ0m7uQeS/DhY1moJqq7ujhr3guXhmP5pK7EKntR1tj+PYzZszVf1EvyuwDIJwrHRyNl8b0zqdsl
IkTknIIjrHsjyM51Bw0rdUsFJupp++8kZb6GEC5l3Rbdg29uK/1VUtZ3YmY4K+WV1UnmeE/K9ST2
I8CRbGBJB8w0VfwzLsofUhKQKVOtVzqZ0+xrGl9h16EdQiYoKlI4rD8Jd7og82QAphD4HRgONMYH
36BFGwSfc/98hcv9ff0iMQ8gJtBOz/dJUuWZ05KCIXgVe6Y1VMCve+P4BqSkJoy8OCTdWpmy77UJ
vOSmahs5/VJdohGbKFrWWvDzY2mVFkXVVUXHpgVKOIBK/fEVHv+NUX1GNzxdDCXSlIyCNaaM+Fzg
eprpFxvp2qkYNw4FbDeisNtT4mhb3LVO5gYv9Qw5Dxymz98V9UNLgzT0PV1l1Vf4LFfXKLQciKRI
DjcCRa+/tccW//bzku/jxgkjvBH5+58Kew5b048D+2b4CCROCfxHfN5j7SPYAV/SsOk+l6l0cLNy
LAleaQTyLnLVbihgqOFqE0wqt6AFIShRw02oOnzIEQ6QElHlkBn3Xqt6dkXZLvP/clxryEzNXQ2y
Rn9u1q2Qkfq78eE5pSZTt4y+jfmx2HUln78VG8JJa2RkmZktJKyXQhOiVXmTOshf6oKNa/yDV++a
xTtJ0O4sI7HHlEcMpJ8TyK2ZcJf1enWdIK+Fsl4kzkKqeFQneh31mk5/eGFpQVIe5xsu/+sgt2YL
R38TXpMc78adVeeuOJMxSuZKmpHIe+S5unq4r150j2CA4gPEg432axKbkIp/hVPrMsuDRTIcMr8Y
t2t1TvtNGvwCIoq9TdWHWUDfx8MetyMKXGzLUefYnt/2OAvfefjJ2YZLGvWkvk5Nm8a8rAfmc1i5
ZdoufuNFnPr3h4NJEVgeK2SMtXGE2Rc0/vphPCQ0ipoTsPfXugqqq6Wumg8Ykdn6sEuZTfwE+J44
h4sk7c5qc3Jq33iffsEs/fZH++M5p7ujv4uF7cCNx9GIX7McmwNySDLriYW3wdfPMgkKZNtbw/sB
M/etGPXezrzTEyYbHO1RpUL07g8W40B+osnSmXZTcNHSh/NCLzhdxrueYarKbah44tTh6Zr/2j/O
mFMx0mX+20Y4Zwsf7yPdRhtExY3rg5jEw/QAYzOqis9gtqJBozJXNrnuZu9faXmGceWy6AmFc2WJ
Q9luSBThtcibcIhpmutnqFmtJoCAZN648DYmI602P3tGBTjyofDt0zaHKdQkujToc8UoDh6oOhVH
SlLr+IZmIoR76HAdYADFJ1ZaWKyGR+HSl55kq4qT0QLSdtzYJiPWNPsHNGwlphZVgm5Hvg+yhxPh
wcIrvd9BHJ80GZi7I+K3bHnCQW1W+7RDYWmg+CR7GrPOV9KiZeT1+9dGUFve9fWgu+Kb+NvTsa+Y
7XNWqTIPSQYG1dvxV5vrL7tjLyqFdPOPaiFGzr8oNavdHt0mYbTbJkgyxb2Ql9uK+bvYzjUImGQg
P6bt/3XInC88fxMgsk/trbLciAHQoSsuoRqfxz7+3Mc77HQqidVrHWyaeD2L6PdATjJpgZCISVv+
XQCKBEzn4oyycMI4MIgGCwhy+UZJIvwwhtbD9riJhenx+rLYTJ4S/vM9J0yK+qzPKBhwdVdWQi69
0Qw1AH66utwqGO6MeTbySJssw0RONPy9uqkgPh+HjHO9J4uhxMynys/KNJP5u4PMRabSygqe9beH
45th1uagOJwv2qMKuu0gmYLZ0PN28pH0hVnNdZCKoQqq6gCnhaTOaq1JLfPRCxVNbLH4k8gEe4RW
v8EIT5SwO6CeJv8d80Lb1TjM/Ebpv5Qk0IdFXC6FuTwwk42ocAgKfBfMBX1+4vViE9SpAoNBy28i
eYlcyn2bTEO+560Ct045oZquw9APB+w9qVcRuVm71pesMSQiVjaWSIcTNiJZzQd7qXeMzvP7mrUB
H9GQNzm2eqK+Tvzfho1UuCu8udDDO9sjx2Q93hCAKwV1ttfHKI3oHViJxXqwA6b1Tj/lG6bPPZU8
O/8OgfiPCFrgf1zRFLAtNKVl+73N8uDGVIohejfIL+1vhmDI09jvd/9nWHlwgFMQvhnfLg/Gwlhk
cr7AM2F9H4tcRTa2xu/ioLOiAfKi3cd5GmhnDsCzdShKdgtvcK8uSAEdb/3YRHPmUbECI0ZtvrjT
lMHoOwao1z1tLBQhfLqwXe6EFKxfcF555bUE4kFT14e/qA/OAwYqp5vOrY8ZwSh3YE4YKKswlqul
hhQ7KVanOxYKBMp6NTLdTuBBS2yBN2RnNSvtQrcaerAKfewZNHZqGIajwWPoWNtMeKdG+7ALs++c
gkGsxM3+gVXN47MztRVu9N/cCv13kTNkt24hd8VUZPK7gNcW3cu/etD1SLfKNFrmQlNuCqEQyPMS
fz9lDQk4oKhbuVPlBD22Ji+XRWW9rKv6FRAgdxJtCd/pTW7WY5GPe8QvsAAE05amZl57XMioWNXs
ULx7U+FcORyA/+uCJVW4DVkHz3phWYltPUKPWoAbu3Q+V6qVX8T8PI4t5neFhfD6aMBrkj9OnXnu
hj0yEBuY/xCSKqYapYj8oMw4I2reZMLLNwlCJRr5C7HOEp0ZRtM4LCgokcyGkpoKybV8GcjSIuYa
Xh8n0+sIl9zKLBtZg2NBFaXbNwKTd7tqfaOznaRXIvjbJZvu1sVlRUsJI+GPqNnOl6KezY1eHsZP
LyJRsbfNAT9NQHGNFG9uvZIhydnDQVJnnW0Vj+4llwz9vc3aq0umZH2yjYkv58F5Nz404huS+pvR
rxBSF8QOtHcGtmjpO2bCU4P/Ao9lZ0KRnN6zfDzW5U5kVLJzEJRRuCkjqOHynR19Bivx/0ZjjK04
H+T1Z+vK0D6KGSa+tCugy4SL3/kcLZCvvXjYrZmhl15/wCQBGeCxVOmaVrLph3pr75kQoAEipIBr
a5e7B49nmTI9fIIIIDm7OhlF/kChXQr+sWpIy4oGsXOohMPHppTF/sxKFgUr1O6mM6qdEYdMJtgE
Asoe5+O4v2zqGemlpODHUV1NcUAAgllNYrJq+t/7MBAjyxJi07M5jV59YLcs2IJb5UeoR145BnQ0
weM8dIycffymk09d/EN/S+PCBVSz16evcqwSJRU1KBwUM0vXIzztn00NJlMS05YECqil9MDRwji7
ObBQ74TQSzrCCmOJvcz35PJsRFul58BMulS0SkAgmDgMIioESl3TEtu9pWOpFvUk122n1HyMp1wC
pRUZW1/hmsznUqc0HB7UR8JWFfggJZR9ApwIbrgUKItd8PfjA4ym96xe7WjtbtmWHMw2KvnnvOrm
o9G1+IbA/UTeSL6g3bdSZxkCU/R0o7cU+lGW9HXuoV/xotTOzfPBCd/gOeKuCyiDY9KgbKq+hutB
Nk7ilIrw7GWsgpisJzw5c/UandQqvis2Be8Ms7Bia79inTPXVirndz+XUEFHeoOW16jlSpL7TP2p
eEREQB23tC5dKHFP6EgeUzACVC216y3zhGfc8De0FuKv9It1+A++E+8z4JRCUJdoobIWbSfqTS6D
HPe/tPApQLkqAih2wSTV5kAqqzjfiRR4OKe9h8S9Ox8mDuOzHcI+NSnDOAESKd6BsRYt5nEkvsck
ZWpEpv+5JR8TcSIW4XIcZ9RTtyXI1ITYP/c7zTq/L0xWofINbtcwAooSzELoGDOkyt2HZVRqX9/f
8HiveoSg1a5skRhx8Q7PCJDCKDUEfVnXi0o9S7L7uGOvBaoyO/yDzRODhGDKIJoR6JilSA8ZQIqF
kkUNQPrAChtJ9Xy13sps6qP9yNS5KMXFwFZoO2gOO7+UXI8cx35GHmV/aKk/jIBoHEptef7vZLYP
riwLmcF6MdoI7+VzkKVi+UgkidcUMwShox/PMFDAXZAWGxTL7NCW8us1oPsluIfpYYWx/F8NMSgS
mHJQvPo7ABhQgkW53iJxOk71eK+UM2QyYSjGHtPBWNSYvclqlKb0jDDxDz+ESnaLCaQ7ElfLtMjn
GrMkDwRKTE3IbgmTqZJnTyBZ4l0sQHaTMdYrMe2rqU/bezRMpTy0a7h2QH+EdIy1HCyIM5B+yBTN
83nRSfMUUaKZei+ZppbsRn/r5hZhuxFNcABupA8Xj0xFZ3MF6Vkk38wLYi0+VdclZzggDVBGWiwm
ehNfa72RWmY7SOvWRFmwGo373VO8b9p9+2ITJkRnV34aLtvKmz/oYR7xoCsg1Gd6EOf2jbb45ulv
LGko/mXT2KyX9oMJfVX6tzoTuAktW4uo5Jbno0EMBO0w9yJ3ijwF64/KPwVVZp1jo1sI6xa4y9Oi
HJD6htfnJDU0O3rkdmmTKunsPDHByfrKkh/TAvQd05H2wvjbcJ7d/Uw1uJOagTCiEBA4iqMpht9z
nDHkwBBEqJPlGxgGorGtVSAj3XldQDnoBwJAVd2bfwiMiwa9CwRzPR1xVIFTxss3o6ZEI2nl+yLr
ZNGGy1zYx7tF7pTvDl0FtMOnlhsDM81tgKpKpZrukwJJ5neCC3u13n/bX+QpT9ANEJvpGcgRHnsV
BZt3gGfJIJLisLxILOAHHKm8PKeCnDRfzr7nlzg5RUbPEqYX4ZbbmuFqxWwPFikAzkg5zROsZteH
QEZgLehSs/Yv46frEo0FIrxOZRB5ZnAdvYpivVSa1fMLc+nnaJRg29O/Y7jB6pt1mSm2T2sJTNxC
VVy5gwfZzMnHnr9cIA2rg7lWpglVN0XKhwcGsV3lC+cHXn8nSRE914rhtBk+7+uVUS4iNBmZZZcp
Wse9GkV9NOxbnWiN+f5reZgOnh3EM/0EnrhACZ0JlRxNW92WMYiQVmx6cRvq4ThsqwKO+Bw/UWjY
qdX3NZv02O9p/Fe+toKUSp5B7YLnfVmoiln7vu0qTQV0DVIG/IIvNRS6T7Pb+XQkKaucjhNUjnyk
WNZWdxAGnhW2pcLOb4to4CTVfQBXrJjbRtPYAcN6TiTBwy2t7i0KZB1WRm4oTo3+mxUIGVhzkBBy
2cHb+8cfk5HCoPxW6vb+2/FVu73PbB/ZlgrIbswBcYi/toOEGD34BUu0vXE2mDzlfSacfB4CZHGb
vAeT2Rp3alCyZPkLj3Uwf349WZ7iMEdYsVCvx+g02kZvMGL1DcrrILOmZw0yrOtrn5T3kYTZq/8/
JeYH1jKZF8TD9zef7AEUT9jzOx1xuwiCVDOUObPpibjFFEzQXiBOVvtDzkIkqm7Si8C4I9CzqOuz
sqw2eMikc8UwTfC7YI1ISwTsmwCmJvwYCjkBC10IRfE64i3fBVidYMBqZHpJdAQPfj7VT5zPZNWz
XpwAe3eGu0jIt1jOu+sGK0ZawSr8e74GaZs591P16warzD9ARfzbT688qlDN0jIGn47llirr9PeR
3ppByOaBq+sTFbjINvW9pgDvcUXMMoeii0M3ytqyFGj5lbtZmOwFZXP56Rn6PLBqOs/FQhtuUeVq
xKFOBFpz5AHVxUZ6p9ziTWTgGFN9GuobEV9OqjrYWK7rcCgrR4G39inVzcGSaEo1u/q5u1Mv8L1a
JAsejhiUkR/YyNKp2TS/SVWe4zkkV0kk9GyPMeyuWXj480jiziHSe4HW00al/EiBd6QVtLRGbBBh
Dbef3uaei8LEm7g/A0Sy4S7wNFLYg3MpIbTyLEbmlnoGptLH2EvFWmkYUxJ2MkyDyhwIAzXShnCl
3T9IFkKIimm9H15cCiNkcM9HvUy9QGvnYqSABf8jm9VLc213hXM81RAeeb7IHiD5t5ZZBSv1hARy
yMFDPI4PZ2AYJ1di70J20zn/vaSc2Qtl0UnIOBqZ8CayXqBoHVxkrXeRJsuCFla0cFhxmSDx+3FR
SXWj8IMA0QrCsAmrX/R74hQLA7mQ8UL8TvbUqtFqTYzJZVnxFeq7SnEE3FoEk+wkH23AhMAoBzy0
iAwpl25GOHt9PQJNmbnLIirXsWU4+RmFg0Kt1m8D5yH5q7HwQnljfOLoAQmW4e4A+Si60x301E2a
2RxP7t3BrdB3e3u9ahd+tS6eKp1Gd2Pb7Qa1XfSF8138CHdhFt7HADRyOhKB/AbOhe+8YuCYeN3s
7ZPzjrzUhohJzLhEcd/3GPe+tuBJdRjS1Q5DxHtCa4f8MJKOKxlQ8XXeIfasVplWPdxFy+RJ5LbS
me7/r506bv12PC1HCDr67fAMR0NLnrot1+MHr9Z8U98NUHbCgM0qx20wELL+1UNzfjkrlFNf/kES
XlQQdEliWFPD7/AzVcva5nK9xkpoAY+IbCVZ12fdc9cE52EKaNepSEDbHoMlL0XZpUF2PYw8ixRA
m+eYawgFauLgg5+RuL8OpFeVQMvLLDvwGlwSjJrMGm3glggs+aFWM4Qujtxke3bcdDyLyLPugqE1
B8uwV/9ylBvPSaLoVnWy8Xl5OKsq3dTsa4voj247iylbdNuwkVwrTlZp6nC5pMa4GmPxwZLtNzr8
hPokb4DMajEhfJ6+HoW553O+bxl933xsNKY7qjKwU0ZHK8URdRwUyv3fTNyduLr5IuZIjNs9bz0o
18+92GKaA1QbLSRGlz34EQgPA5IDOYWtch59gzu7/PSRyGFJmovg50zy5WZxeS6BNspjdu8cDvSJ
rj8Y+WdZ8m4gkDAHjCiYxQglAZSMppTysWoJRZz/eo9hCja9CWPhLFWDCCW7gZXnN8YbuvCN4OMn
2MBOFKqYAybRh6LWwYFxZp6b3k3p+3TPHE1QVvUI2TJcua3UaToIgCW94pe8ErHfypkcye5lpV9n
MKAzIdGeY7dCUqaiWP/Ar0HwxbSHgzo6ApemGZlbFHAZUfTjTzn/IrAJEK+/hFSFrgPnrXWLGukD
Bx7R90RunpxSB7OV+EmR50wBhZkSjeQgzz3sWZgLms3oAqkj2yeUWf8CHDF3Ztm0FGcnfvBW/ZNh
zz8x3NBrtqR83iLOpZAv4NOXc5VHwtyuP02MN94gpimXZwRmh2v4wQ6IH4y4VwaJYY/zq6FDuf3F
WzRbgRpqhgM9wV1p0IvOeFQId8hKcG8D/WU1jqrJ3SIFbZjicCe5Kzri3caYsDqDT7p1G7T/ZEPI
oMRifERfcWytBTSCwazt6nx9qsrShIiZZPxJxicQCclXGVSwuWuqx/LXkqg9Tcr1sCIXkJPK8m7R
1gEXgsuUwl7dV7P7GYnjAY6CJ7pCCBm14DlQp3yZTI5ZnTB7YVCcvZg2oZIyCZYEJ54P4TUwzcSs
4pxm6Z+KkLhBdLY89hwehw8gHZyYW+3kmA5Nuypd2KWT3UXCqS+pIy4MsQwcWQVIzixyxHYKC9V2
Wv8IHTOriuw/wgASdh8QZ9b94PuJ5n/U4D+h0Ho1b4M1UFcgTlBAr4oJ1FmnZ4Kre9RPMm/2kgJU
p5ekOxmzIq5NLg+mSdsVDfvI2OPSMmnSVXXcYnMJ2W2svZboxJ1CL4lq6mw2LWG/5pH4kIZFZJTI
pCjJ+QEdgtgOwl30hI0klEb0YETWZL5CaqOrmhFi37gxTGA5QqSerWUIKCj8G0gRCe4CjwDR8tB0
mn8SojeTKsJx9zy5V/rUm6r95LZzh7WV9UmrKvR+bwROaEu4+1PkARXivcGAW259KyqMg5AY9qAS
oR2nSia5FDQoHhx3WVVUFFs3DaPeMYN/3pLm/+0LKv2yt7R9O+GIK4Rmq2XgV5XLycaHX0XQKdlA
fxGkt53d8NdrP0moGbb8b85Gd1o8PYUT+7yxoRWF/UKfl0xF7zXnSmGB0k6l+aQqlsUAhtdWlvu+
Y1KG2HMV1699YBPfsfaSNJ9CHvr4mKuT8g+UP22q9OtRgC8kqVtZOHn2f46AUFSjrogAmJBpPdkr
MTtmUYo9Q18iEroc7VDeJ/21KRVjDnHhV9ECJaBuq5QexGOoIPDSP5KWcIo+UEaNTh+f5bW/O8pL
vlGrVVTkqjuqYRYoGLXMhSaqHCdangECF+RJkNo2ULqWyz346fOna5ZTmo9Z6CdPRi0B3+RU3oYn
3NwKVpodarOA0ztNiKkcgAwyudjM2YmOQlULLabLcIDLKR4LUxNCXVxyWpYbRVuJd7JwzYIc+Ukg
cbZWHeB13KGEMFwN2P/SUmVggjTIJM9xrrRoObXMqRPylg0mdfrgi0JLIfz2qxk0LAXCiiZ389IZ
jjuqJtSN4ZrARQiln6opkTPHCsrxVGOn6NFbYtrjfykqpbFH8P2JQzUojyNv8DjpNJTeCDv9SKwk
+MY38eO9uqpRrHHqZoMwra4zpOluh+uR7mnnNiN4nqOM1huQKpcK2L2d1S458CyzUgt3M5AY7b3p
YGdL0/OkvhcerbES8eih9bHgOxxbFYaHYzXHCIzCJ+LhDaTWmmO5JujSARMA43uOk0mbEtjn8w/W
5I/7bNw6yCnDg4dJfCg0qtXbJApE4HIfPJMpq4K12ZdPoYkLe72UJ9kbVYS8k07orwF2RtZHFU5L
l01fP0WHDXPgBrbQA0tW42aivMIOLC5WvlQlIjBfSWqx4HBFsDAhFJH/e9Y7vbY5HJVH2YPKHFea
Uutn9+WdYuJHfW05B4dVxxymwoVt289wDHkXTzauzlzstE6vWIk/PYlk++Acgcp3VWu/DTD5ap6c
b3y/uAEX8/sN6VlutHRp/fgw+NfokEAcfn8xkwSJvaY3doEKCTAON5xv0F+EHK2inTDgP1VKezCp
hdmokCax4+yp+s6N5VYac9Q1WTSENTfD/J48faBY/AupxdQF1IcDksE/EJA5HF4ti9kUmGDsnJ9c
n/DtHFPROA25vxwpf7heAqYYrWYA7UiFEDi/ncBXFXOeUiSlQ7lN1We9n1Ur81pgFvkFtrgjgTC9
K4B9ePJtfhSAgv+azOJQneePVv8LPnbdtaHIlZK03qeLkg0O8nTz000PW5br2zzqXdyXPtZndg3e
GogNng/AdT+eRJi1xGY8cseyYDbgqgPPIn1we7s2YdV5c/28yPKedqxKTbHsmm4H5rWyq3DMCpkZ
Gy7Whqs96WNUYrgJTIeaMhqRIm5xoIgq8eK/iS/M5l7y1MemKiwAxkEHL5s6Z2V6a8ilI3nn8YT/
U+umnBYOs0RqesGw5ymQkV46nB2+i0e6afsWAvC2CH8nBA1eF2QvUyeYS4S3rabxARua/u9FvQSt
D5NFZ5LF1WEF+SS6+Wsr4k3dV3QPj/YmdK89ML1Z/IRk3U2DqyqTPEdeOU/B2FTaQi/kZwKyC9ju
vwtod4+MS9Bg5YAhf+7QLPfqlraTB5XKkGpesy5PCczbJLWMooJXLIVlNcdHJzdTnndzzMaLTf5Q
v5UzsqhwdtA+MWIgi/l8H9HdI5bHJZPrHlEhvZRnTfNWZvakEcse5p8kXoL/bQ7RkXRwCTBN6QwR
mMer3/rDFbQIh8SB12+pUYbS3treJwmF91CccV1S1wUxzGI41GQVqkkudxhmLxxvMx1uaUXPbhVT
uCMRO1jykRMziUWwG4080oJTsIEDorqFMV11zfAKODXcbmCbmYWR3trrneK7NcPQQXuZJnFUen2Z
Hua/pSMwgHbmizKRBORJ5+SUnTTr/gKMEQbhbY+LteTQAWABLSiueo63v2MU4N9KglI/6cNVleG/
Qv8GuxVK4IC4OctaqSujguU1jIooAo5r36t4kXKtpmDzMlm5tTrLDiIyguvSG3zMiY83e7OpfEAz
jwvQgIMf+SjcWeKK8eu/EvK4j1df59fOqOxJiHxKGR6q3JrdwbefM6kYtJ+KGDuH8dGQEgFj6bf5
B2K7bLkIBwAuYld8g72B9/By2O2bpMc0TxdMToNQ9Zkdm1q06P2gLcqBSEdb11BnYjb9PvJOw2xS
FAj1xr62sUO1nomzR6WnMP14MGrZsqk4Z+gueupN8djv2XBNsjhbSN+m/XotwW6bC0SKQvdsQhsH
BMhvIEzEXvA/gLZN6OTnR62CmPCCkJ0tQ5o48sr+C6jMAyVlU0UkW0ejp5hOkL2vrMpMf2bo3oKI
4y0Ew2tuAsSvTrG8wa1LoneotaV1+Zey3IVeigFuTNpAMglimccDtOHHFO9r5GywT17ZOSCLbVua
g1zRUrL95aIAk8hhmhGUVTrBSz1Dpdkbek25oZE1mKzXpTeGLiYZx4ycSbhmPBieLTFYN7gO0FfS
F5AX04NY4VrwVkJudB0dmpdI+O/uRtBTRbf8RhpwIBQrVWHr13Ajzpct/P+pH0mDsuQLbJ0EXHDG
KA5unL3LxaXVPDowhmLOGHPFNLft1glgWPzdkLqAuLTx1G4ZHQeGtmYUw0zSqdjkosCgDCeObZ/I
Lh7uljtAUmbQ5VqL2/MPWMxKYRujVXE1j8LmGa4J2XjCRvsrF3+/zVzY4X/lV72yDhcMaSPVohMQ
tesTd+eZypzWlvtRGEwMFdDrRbNNqjQEsVc5cOdTR0fKLXY1won0Q0p3PqdwQxpnn2TuoG2nCu9c
YmyzsEDo8F09cyuJKFIm6SQRipyfpCxREMUw3IR/7HlUgzSkQFdlkla9EhjWwg4hcVRjt4SNZRYA
+Q32D8KowLSsNO2Feo2UD1XJKm80+KRtqxzPX/dwUxiQ/8IOShzBTfU7KyjxcicvqRGe/V2VKlMu
zAlPrKmJ/5XKm0pyTUfVT+5Qi9XfqtSMdm7PC05tMnYVmbaI2w9VJUW+1gLqJdiUy4JXKjdj8E5e
1h9ddHhjqiNU1elBmQaH6UH/QLJqky+FVh2RZHdLO8ZqitW0oZQhbz4+EDDZe+x1iR+lANoiohjE
YtxYApY78Z/oT9PPqGJBBnrZRT5lJCg16kQWiNzQRIzjhbeERxvQNIDIMb0SItST8RrIRl/hICAR
5LwyaZmFwtc/yVb6e0/VuBxcT5kNb3PKCrKh6QN20MvBr1BemOZdG3vgIsi6WlfCgbnIBrqLOFrE
0HU6R0zSer9umVdSb+pjMWXrkGttUF5/b4xlxFtWGcI36XVHUjFqzj6CnkIypt/mNw3eSCYW6Ph7
Kx+uayKem/nEGB9SwhFmoSkoPM9yK3Faa+mFmql60uyULrnlMNB/21n5Wer8j5+7hLPISVw4Gpmp
aOwxP4pMUpLcv8m3xLW8y5oR5nIGHKjpegWZ1GOxfdYwahX6cxZMvSfEdwyu40fyzDW3UspzbJvn
x0t9uqOGl9GToMF/1Liw/kCKfKKiLVeTZJ55RS3RqdVwux9ODs1Pk6+Ic9O3/L95qkrTG1IF9KYB
+BfIBY2BgJ8y77tKEGJAjqNSFwWbrk7fwx3Ssu9GWr9klxrWutYFqgHyFa/cdgQleDjMBOtsG+gC
iZuRArWsNDM/LA01eaSkMplHM0RtmqnjonxukWmPE9+d5+IHdVG5N21O6EhI4rYa2G2TvWx/h7xW
NfMECwamqNvf3QwLhNpyFERsg11+ma0dxvOnAzxqpywviAWuui93QJo8x38u9jPVF9p9dh1ZwwXi
kVKZCqJxYBnkQmm/YnravMlJwEwc0iVFA1/BNa0qiJRy+lVge5n1JE8roY25xH2GjK0+6/aafftX
zieZLFLmQM2jpkc6M5CIHwC2MHlJ6WP91RQwgVr1aJBXzHXG+pkal39SSi4TaMvUVE0Q5vpp1jfH
vnIb95IKV/r+6NaLO7QKXkgzMKeW0gQlUyPx/EsoAapzedsbCzsyomBaftpjlsf8dV6vXzbwKPEx
Le8jXXjS7kG96u+93yNEUS+P+egSYOPmXmRHAvkS9FdaSqgHlnyTpTt1wvi7o1lgm/rY3E4BzZjj
/98v5ujI+WKsKhy3KZzLW3Ma49AQXtnj7mIKF6yQw1ow4w4mH9+TBzfSChbBRmXU1dgMN2sy8bqZ
pDJbPhezqHAkxs//7+Vh3QxILO8fm8NxN3TH6XiTzTmPPNhhP+xbzfHqFB5RJkbShW5qYqpJWPxL
IWKHSMh92G9ISZ7PSQo7IORnvJw+y+LAz6X7+Zqv3A2E85qVV2hl2nONSVwRfYTw9fbMFnjUyCdw
uSwidrVmMc8kQuG5wjXPaoki7SyFS4bL6Y73ugS78ILV4Ml57URWSf6NiFja6YNIAJgWeML+4Pl9
o6gjlPCGYBR7CD/bR5yn/sZfFJszmQSXhhQ+JRxt8x+gnvq5bnoMFPaqfZEeoWPvLoo9RWJcyun/
KIuKUalHqivWbsfaKKIlyemw5jlrXiQ2r+ZuE5Orb0oqSIMX2GTv7ezGzJBUoi/NEwBpJPeJcwkd
LFUK/NQXEai3cVPza884guA91EXa7ouP+kx4D0C/Ti5qKL8VZajmY+aZegAgAyDrFHj8ypPM7d+y
xnYwH5G6rKgWZXxqMctdMb0FozNwnLaspHzrvAXwA9l8TC6Cpp+ut59K/ccR7i7P1wxai/45rcIJ
RxU4/J9rrGU87HcgcR+6shNyUBlc338pUlhMVA9PaiCVZpUYwqWuRC/lZ3y8YCiHSZx0u5BnBGrs
6H9bN7QsQENPtRzaaQyQCrXsrPlTWxgVfrDMM9/y/lEDS5foZLtAFm4+mXMWla7zLhRbHMjQ4uI3
9KQbxNGghpaim8iOLQ3EPgeYWWpBUJ3ozhOyCWowHyDMNeWUbi28H8k4Yid2GzeanHKH0wGWnDQG
gJpFjH3mFeqowGdj4mMgAfCGNg17ydNPfWptxkueTzjGw6sVDQ4u2nj64GH9iGv/eNmX7g+g23Gy
HHNsSJgydjJVGVzsL/QDW27bXYfwI6cn8D3xhn6a6UhyDrRfSckQf7sjYLV4M6dEt5hbqND23j2n
nypM1RzCLM5KHwXabfi2qtFWn6Xrr4s0mieHjBREhrss9fywF6K0pZ35xGkPysm1KwGr9D1Jnn6t
uXKP8lwXfpcrFKvTpn9X2+m2ICet5xaoDxTrmG0d/DL26r4bErkBXdYvkBTt4aiwM4QEFxgbHxg5
wyBubob0W2mM7pe1kqzwPFDI4JMF4RXgJCI/XwenFUjOCzdmkg3Uwqvm+vqaA32h9slx9pP5yNgl
Nc2neG6EI8VytFX134ItY/7oYz9ZM4TA3Rn9Hj4r7NuD2C7Iukp5fwD6dVTN73F+E+FUXT7G82s2
qccZrIwk/c2vysp2dfX8Orh8fbj6WS4W49pe9MnCsy7ygn2J54QiDOez7qOXzsrn7vFC3SGi080E
ukuIeGy7qf7g1z0Cbg6K34vmwQAdv3Ggfx6nbNdLsS6Lx2NIt3bpL7Py89MJFCu6XEDiMTj/VFmk
p/EtFgRikE9FljGxk6NXoNTY1yrm1VboMcNtsdhZOYCVwFAa+hMtFwWp6iH+1VKv4nkJ8CWohYdl
PRVaiGT9nH/3viz39A+KR6uTS1JykVivbzoIcqfNFubdMAA784fnSjL2DwW/skdLg3kASPRfYwJj
MPphy4diXkub2m9hdiQE7bA9fEUsjDXhsyZ4aam706HnZ8/QzY6/dhxnCbHN478jT9lZS5qVDejR
9dJhamMs1irf3qwrHZUcY3s7JomoRkqrJ1luXb3HndDY3eM5S62NBD6gujUtVHvUIFXep49lFw+V
NW0ZlNWgxXJUjEuXbMW8eIWZz1d7FTr2WTu4lbJx2znml+pVBN9+kKsJOiqNjqHdft8azJINhU4E
Ri2FR3RYaTNAW+cz/tzitvaQMIYG+ibQOoionquy4g4e4R2P/zuBEg4vaubHwd1izmVvzrRED/nE
Ea1GK7R/881vWi6RB08rsazUIyOaH0DgRPdXb6/MWjcTLsOaP3dJ9B2lf8M4HegP6GOyrU2EBNkE
rnhXc9jBKvJXe9CBKVMtZ2i4dfa7giRczssD2c06vuESpIp+kVaHD0kiCyggUaHvTK6oW6tAgHb8
C443UIYeMS0XiVv9k7aaC9V2luCoCUsrhx922sDXplvpATjBPoWnRBC9LgkcLuv7XY2cPNbRcwN9
ZNB2qRzwfaQV3sqy47amLwn2ZmEwDE4+UfJutSMXmCEwBQ9lh+IdcLtTnbB0XQCCZG8Ui5akdfH5
LKapedugyPUgVs62LabKymBe9Nn7VcczdF4+v0X+ufqkboqw7TvHwUM9U9a0E5sdCh/Hkh6w0lkZ
qherMFrGUfSFisoack/T0IIbBGhwp3V4CgnvdAn/+Bo05Ut9bhGdPMzF+q/X+02Yp43JdXBPXO2t
Hoci87zYwxRCT5uzPrqCs2Y/9pF/miIB8i6Oh2sd1elqUOa6heG6k63BhtvskQM3bri7nJSTB9qv
2dKHLBbZzVXlU7lIOWe3cH65cEVQnvj2dMMgvmso+UHCC9/RzY034V236m/apzeJRTbIFpv2Vjn1
rtnTYlH8aV5k67xX919DfZUEX9kSZTkaY/WECKJqByjHDtv7cXDYFtChu4UtAifRLW/7nyDZs9Ob
cXxjxgyVfTz5GAH1AW5gPTFQ5bucyJeGGGhUpeSIvJNeJoGh8yiB7r9HX7TYK6/fGR4G30ydEHQD
CwZbdsQIjR6+GJI+PeAA/lwmdrhovCOShpYt9DBUD6cyPSYK2XPiHV0VRNiglMbIQN5Kyt5SA0yN
MbfWxGMMQVtRm7gIOYNbFBnoJXzyQKgcP3v7uBfic7SPSwiYAbk5oigKPlWgOjoNBGLe5w2nLt8W
tc2nS+0LJdhPU7EVPYMSdEsDwzpwtGolSz6Qwk+X/mHTpn+Xlq90aiRrKjgKGgmMnnqwwb3kH1Oa
0iqwhgeDmMgmPuAycngD96jmCedNj5N64t/0Mt7TEZBV0d7VDtrZEehvUJrVWfYbYLRVOIfh1Fu3
0ytcFsDLrIrECdrVLA/UgmKfcnVAaLg/AUXg/Ho69BROChzf7VC8DcmqfbKCVeNcILPrgLjKzv5q
OCF/pwtK9grA6WdW0MztJXwQHGgO5PZ9eulbkrCv0po5aZL9+p5e53OOdlMpukELqGwIMJByL2Q5
54BwdJ6MYx4tyydifXQSECNvjFHYHpYZQGKW0GLxAHgdIMPUTdocTiXy2lUodROFzGpbsOUNHt2s
0l+nqxtUXThUpDIhKlP+KCWrXuKEaLSHGQH/AFSImmXa82gvWERwTjnO+nZ73N6OkCWydsIteD/d
ssiUGVom473sGL9jDDWF9ytHj4h9IqPc2MT08CIh9mjniOW6jZlSd2y9JFakBBfM1gguAmWFeX7D
Q2NDRsj6ynwsLC8IshDuDKXsl79KWfLoFPu0kPg3mpD1XTPWpjL2AffXwv6OuF+pm67CEcKQqCV/
Qjedk9RomEWwHofjcm3tEpn/tbnWfGT1Tj6rxyI78ZDWsFXAw0yMN8FrDgYMRWnvzcOfHo1+UeYY
Hsx/mPIXAub0aEPCa4Dur+EOtcNt+zXt3hnCgZPzs0VKZ6kduAH5evM6MSENXLYC2gEcqlOyy7hd
cv3yhLlW3rfdGfZW5jOX8x74JkEU6nSEDou+QBkwmVPAoaHoOsa9A959GBy9vpRWRGrawhhaG0Zs
6SiiS5f1cXngcABBmcQOVft8Smdb9PivvGDadPTG88v/I9v1txQbfvfT2K+cUCnvG2Hq6iyUkKUu
bqhDPP7Lbqqkt5kFmQYMuLwnrHF0sN8npW+pwCwUpKMdF9X5JH3zM/oPyy+zJd21HZBUqFsB7Aqi
oMFKdwjDNhluyVhP+CY/BMrv/M+D8bZ9HLb5WPw8ca7zyu0ugT/T+hRXEaAIYYcKhny2/z/LSh1C
OgK/NeVvPQINqpWJ0isTKppU331krL0bC2syXedI6eM9SZ+noJvQkzI82nCjI/4+3fjNfohZJ/lG
pypK7HRqAur5ZOYz0Lf5yw2i2FFfb7jaO4ds7IDjMiEXpcOPjfiZ6ZMvpuupGT/maBh5pUUM7v2u
V/IBf3Yct5iUcTYp1ngzeWYisQBvUMmncgL2+RW3LMfQ153zq4Kt52jz//mhUmvxv09+8Ekov9ay
SsMV/QCa8vfRQocsY9snzh9czqJ33fWXFnrzv4MRQwo5DSIyGc8PLXysR0a0O7ueZct3SZvuHQp7
OrJDRTi8jwPK7Su0BmREHVIXMxdXWNO/xBMB04nuwt+pPkEUZG/AfLVfFbq4bAkAAEPLwsImpNGY
q4Zn96TfqZf9XPjcl2BMEs2hRhzgX7SW+hGfsOHjKnFAbH5eKzp7e7qJq+VsdsAeUuOaK15Hdnwg
pbJ2Tgn1oimKmyjaT2JR6suUr44qFJ/wKxJKxpTpym+CMOg33tPLvwO51PDtqsU85XtoXV+549zL
q3kifL9h8nVbN2CZqnYBBDILO/u9vMvlHSQIhKTKmvOMJGXMXCWv6N+M7aE6V+X0QLWySk2WA/rD
qWRCHlfpCFQL+ZULvtr8VOzEUwavs90stMP8zu68VDLUo8gqcdMVloRELzv7bjOD4ZOlAINDdkUv
V8KOqDt20zzLY/qsOa1qnPCQtNKMkEUJ597fhDHs0USE9ldyj46LQ3I+J8AmA47g1PeeE3i7YS9N
VY7dvZkXxxBLiIudmth6DsnHL6YkFgU5nFDTve/Q3/5JXEcQupirWvxmmPQdOjMjwtCTOgAcYBDy
tjF2qhvhUmtHuItsnTSxPYhozo/ysdMwucrUEqxSjzI/JplfjH6qAQ7jy3N7MoSjpZ09KXUTQJ+c
iTpKzzukGsXvFmZ8vSZ1I6NABZYULTYBCM00mbxXJSElfmzkjjudSqtVzOjyj7pg2qSdesk+fE5P
2xLZN3gvv/M910S/q1XdSmkpWhUJCDPyz+UzD+JN97RW6XWQwpPyi7C3xRKtf11Ko+an9O8OZ4ql
KENremNM9Uqbj9ma+C9KDrB8KJcbQg0Ukppwb0di21lnKWKRTWR3mYJ841tPOFm6iEx1N0HrsGCG
GXDjxpResfc3kopzGBmLkeOhR8DzmRDR8V1AEEOqIrLrjCE/cvQj49eL3vx6dzoljWVkxSngcHax
lz+R22OiF0B5CT+nk0Por8BhaCfwJnubC8Q6cm7D5JXswqElRYvRosLOrnyVd1y2lELraRrbedDx
BrznSnZQj4gsrZ0m9q18WjNLKAvZGq2OGI7ZwPUoegWwnfCkMvs9alwrG8xPHGKV2UQAzlqEoDkR
rJjtE15wQlAZaOGAAgGjCKGRAr+3w6xEIthRjIgRBmjJiOr0fJUIg4i8Fmng3WNKUo2hydEzaYWD
PKV6s8+NdwOAmyLbuSFqTaHZJf5uXEMDHBuK7ou99CiR858Tp5DfjEo17965b6EQidEit38rnR9p
c5uixhABCukOf1RXrR3wnNHJbxt9GtEbx/HAWG3f33qv22uwTavRn59o/PWQIeszL2AaySnc7HRU
KAsduTRNRCsqgoybGLfu9M8TVKXlJ7fs+uIvuokTC4ploERGA8x1Tb+pF80SQ/pb9Zo8megTqYkb
KKFwmL3WMJRVf/Vda/8LPXJFLmGAwl2TgBBbhY3Tw8WlcP79050yd2t3ovRraDHm5NjTY/++tNWc
uRMcDTTWr5ur7re/iIY9b2ZtrBc7U0HqekxvvZAgsA7+/3tCqfBMlV/c1kZ/F6CN9CE6j1JzY4vA
tC6aYZwCN+e0uWOpzrYGJltBbyRsXd0KFozZjgGJZ2a8vBjPW/se5Tg54AtBLvIp7NGk9efY7L3I
DBixZqAXZCDpMYfm5ibko6ZVItiGG1Z0lknMn4USU9c8HQ+UfJuqTqkhmtEl9UL1TXxKDIqobFXh
ERo63v0ICsm4Uct60WZkdawsIgJxoaTraiVSxOUdD3keKg9JFjztRRgwDzfE26DOaYAhzmLAkcJN
+6EPBKE+xymYWN4G7umQPP5bNWZJrb5V905L52q13+r5BBfWm2kKm2FJHsFzuuOml5Qnm93EM+QZ
d1cGdsEnkqvyQ3gE7Ueh8lMW0Nh2L0uD4vrwHi4G0tBjQS/iyQK81JOmD1HVhMl7liVJf8O53sNh
ODr9auFieRfbtgvj7dgtP/Kn8T9G45Yhy6AEUNM4knYUpEdia9toG6ClJOf4pOYHqIlaI4ZDUPwT
bMDf87L9Lahkg4siewXyIsI+hSLDTlsqtZ/XNB5wE++dzeEYbQ/9UMl6UuV44TN5DhoD9OMIpspB
UDkzOJjnnBMVo43LtGYDUshgJ1txvnAcebcbqdbMVRV8tlDjtvHSArYgsE1ejbxo9REijokkDN4r
QCjOIB5piMghDV9H9ou0O/qsSzSTqtEw4gQeFnbeN5XMqyh4jhVGpcwV3vUfcGvPv07V3Dbpw/Q6
6nwYMTjp/rPuALSEoxu2/Z9AMBH+PX2urCTzu06Z791pmg9juDDJFUcJjGtn7mq9LzMaeLKieNmk
DJYkLyI3L88moPUrNDZGk7SSNgtH/4M1JKMvYusLolCH/eZKRXQqqJsaXwfq5EXrvqVNxTNxfFEr
bVT9kFaJaGW3uvgqJMca+PV+R3fKXXNiw/IGInfb9/MyRC0R5AtHp4CvCTEqgwpwpSh0ys1N0KvK
LeTjsj3xtucKC+z7+A0NefFix/G/JNSbQikHYSk3e4pkv4shx7C6AlcyRRXDJClCaLEQXXf9QtP1
f7caVl+LIcz1OZsTUM77Yo0AvE0qGEZS/WKHsWUpwgEy+L4et2SP/Vf/N9kT9SugnDmg8jyXnvn+
HgqcCradDGtTLHQgj/NuQyL647MISRycMB3AoH1lYn2h6s4SCW7IwlReBKCdME72Ls0nAM0p1ek0
J5TaW1WNnOxYdsfs+5mkpbueaXJy7DU7CKMMyxaEwg0XSGOpO4AC37l6/dY/MQRv100/4c92DOji
D9vjhYMpsQLEBWW5S50cvf6xEmzAQNoiN1QVX2lydoOeB2HTF6rv+YpJEwVxwP7aXIGS9TAOnfvz
rtmTANLKvaelrGrITFgDSQENjX51bEPv6PuJtZC53zjRY+TeM0Z1DY9fFSGA7xbPIJqHsa9+ezdd
8Q8nJRvc4QOWtql71kxV+YUkvUKoeFC//ykGmPkg119ga00q2++bAEnMg0eFNm7XbFYx/fON5p0v
zLb76ARvpnnBtDJEAItxtnGQwI087fVzHfoMAH/piWrA+SZkjyFUAQeznb/8dPprkEHFYaf+2Nb1
2q27x0e3TX3ZTW2oy2JSr2ePySM+E0KLVL73AqfsHn8v1gbHDlmyXBNqO0JM8SAHNZfDHo8hEDU1
8C6wMVI+6enuY228q8M/Qf1KgbKnO8yXV49gH7E7IRxDK1h2+38+FTmbsQlEYxTWcRp1sjV4VUFl
E44Ow/URt3LMULPyWF9uSUrULURnlLM/CCiRrcdAy4TOAHrJK37+4J9oan7hzY/ljC+Ez92IF+2z
aAhwxSmdPEXYPNf3vHfyO92os5Dq867Qbjiw1BAkIisg1320nuow56KzERCsZ3D8+HU9KgOkbReL
hmmmaXS9ym1jjLCSZ+LagfHUW/10pLOcXdD9fV3sgOr43Po4vBJW03O+SZazuTeqa03sCOE26w4j
vxdVtgkdn9SmGnUbuPF083qZy5/goDFceGma6/ZWQG3TzY0AO7OMF17PKxGZ4LASN9uhDBrfQOyc
fSUYSRLe0Jz82C8fJhGCIGfl2cj6ZRN11yz4xiOk/4w+4vIn5gllDQTzPs6H34bbbnTeD42jLqjU
QgwfuTL7bFkLWKrvvqv/QQnbjDurBSmNAwQIj8LUVwbjqtj2YmH54SFDTWBbuqlJsX+ljQhAERT2
xqQxbL0y1q0IdKYI4qU8BeEKUFRY+ab8bcXuCUhMrnFOsvfkM+VDq7vo6IGtDz5c45ZQFA9Oaxjf
ZwDQ3DB12YT0hrxoQ+mSAeBdoihl6NuQcbsT6HKnSDPo1LUe5skyXwNcm9JE0ziUJ5l5yYNe1FVi
mHAai48gvb1WHdoj/SfOti+O8vHkalFO/Q38s3Ci1WDbb/kR6cu4FkGhOFc+BDUm7VFpZ0Vje63+
wYz9lGKQb+4t3cAuTQP/17cidsy9Fm6QnYMmG/HZuZW86qL2Wk6fqbqJgH1DECibzxT5xk9Kq6NO
Xd7lWhkl7tKWf8IEr65V/AFzlDZD3OZ+XXds8EEnf4XM6BYwX3E36NB6IY74JNLWq5+BdQXh0N3x
qcAvjGp14xB56nRDw2A3mfqdZ+RFwYl9SBq9iiYyoYVqX1wRcgnyHbXnhGl/VMUJmGS+6MhtNP5V
Zr2pAKJGnJJ1X3Za4FR6XiNj4fk+kXc7iTX4uBcNqqJnZJ5HxKX3IcVzquCWaaaLDXYWpJwCLAm7
K6H03CahkVWgKW7n+0qgOaKrQ4RXQx1RjSSmCupDQX9Xshf5BaYiK141R+OdqVUqyX4/p372HDFN
E6W9+EvFjPy8cVbIL23TEeiL2gtxcXBpVtK1gdZ08/WV2QRwwGmvGy0ImW3srGNH+9qgvN2oj5XH
IEnSLRb3vJoa5TONepf5OsoyftlLDk4ktibejU6rwb3UJCh2rc5rp8GWKQIQdd5tHmhKkYzwH+2Y
/Z19QqTdiXpTAJp6hekqzXK/OX/0Xtf9k5FX/IiNRO4KsEglX8jt8A5UA0vskueDSCrRfN27iwmv
tGuJzIBJ2TU8zq/N39Nczq/9j+2G/VvsbMVoaGx0s5nWjVSQaWe0jMKU+G0MUMdflYtDER8vroHG
s+rpynkNX8RA8KxHUUJJlhQssFb8KUOGdNhjPnBopSfoNt2nLHZydLVOYiIXrgET0zBwf79vETIt
W0lqhsCV40khnoI5wRuT86ba64sa4MT5hov7sSPlTU9h3icy/8ldzj+FrJEiqIHbyfOffERAvaLV
5pFQJ5GZDTtI88xFqBqy9c0UwN/wmBycRy8/HIW/nId0BCLmeveQewmasYn1npCRLm40qNe6Bk+8
MzEnaHkjJ8Kpm7AK1sZ3GEHvc84toGiwZqgfLXNKeyo5V7zHUevmSaYKMTR3WOMW1O1Zbap9Rn/f
yQW241ZrlVcJfwIHsT5ykbLSNdl3Dxn4LTc/FG96SWl08glcjukN36LIM+NRbylW7bPTVB0OQqiU
zomdONf3v3bBjHf+Ssqc4Xu4HLs6Q2n3FoZFaK5JJd/EfTOe0PHnrQEVTdmHkgEt98CdwhECFJLD
4fwhhvwB1049VFYtVi6VP03t4WmEvjDwVXgh+7V9JkbxC8DqfgE1rHWaz0dvXrOtV8ZV/X4stPOU
nYDqlWqZutyaYpb9G2vuRaXRDezxiWjJt3+lpvIQGy3qm89hNE1v59ct2JRwwKkIaQ7CxCt18GRt
053smbV0wRC59T6qp9SYev5botqGwlusiHVuMPRidAhUYLGZX8kf64ycqDxC1YYcX87Ny0WrOO1D
BnvqErqq5/wctBb+SliWXt4PHoW2MixxJhWC4CZ1sKT8jwrjXlYFUHQR/Lj1JX3b12no/VPTeYIK
v9wiIw5b+SF1+Wo05I1b8q0L1sTKlJYHWoyQ6GuQzHWxKPXtkNd83oNl/Pg37g6XrG2LocBaGIIE
Ug9/hSV2TwElieTyTFPdqu8kvka9QCeM+Cq7NOVA92Qml3rahzdHC2ODwekw9uvVgGCuVERV1s0q
/gobu1hi2Y8gfls2UUxMKq7N0V3KNnKf26uNgA31yK/owAvZH1cQU/oGb4R4sppIsOE2ep3ToKp7
FXzX7bdk8Ncd8eBSDbPKfzeftbjn+146dIC18qisZ/bbvVUAxtePFpmshtQ6Yjt34B8RiHODIJZR
y3ccX2im0bOinglk0qbNuMM8mYjIwl7CMUkVx3VXBHv7qzoBDtjDSWo8KfF0Yvn0JCUdh64UkwIn
CFvcCzNGsMf11yQIcvoomdCSG/XHVLO8vVzzH4gS++Gicj6DuFda11X0bt+8AGPITlxrA4cy+IeF
2ENTO7MxRJTTlenvzMs2AfhYysvXqIeB0EgrfFulspZFLyl//Qp2u1Iv4U4Y+qEfSWDH7ed2BkUY
nmsw4ojjoPfJpGEP7HP5OQFDEBPwsVjU0GuYh0qa9zA5LndD68M44f53jLn6QK4WbbSue4rfEk+j
czCbqX5p5m+aFngzsP7ad7wihQ70Yg52AGS74nOytnf4L7pXU7abqTo45F390MY6PrIfRCqn1d+M
3UPuczpsrWfbC2EQ2IS8MzFOeURl64wVpyxwOOp9iSo6vA88mRea0bb+nLClKeypOyRzXo3lxhbm
XplXz6k5J5izixOmnbS8VYT8y9O7hHV6IOnt/1VcinbP0MF2e1CwjRWcfH8hsoudmEC6L6eUTMWb
IN47UIC1IWH4HEInPdt0p2Ynuj26ZCtzJ4gnvL2dKMV9G2ZsmDhQfLsiZc5HzInYdhhPzjdEWEck
2wt31bWUaYzvYW+dUHBsE7FjO8RTTOi3TFdv6gvaYrGavtLrwUPX+L6f7OsHR6RLfvmuheuQ4R6P
viwENC6FH6sEdSNW8LdFzoNeSfEeT3t6vg+w4mxilYCGBqTCT+2aIeLXXXPpzqxLs3f+lvrDI8P6
P7bfGJV4ZoCaLGicMb8pLFcTiXQ/4mCGOlQNyIo6xwAr26tbzXDYTrvBjAxUDUpO8/Bpsh+P9T1o
ytdNlxHRJqL1NvcOz2ebXzXvFSx4GXT/Os3bOrMyorG6wh2KFMWbu/yV0fs23akw0Ugs6F+m2UvR
K1iwkJRszenKuJm0hMNP1zSkp9ReW0k5JFtbm4LGQByUfG/ln/DFnPnmJl64MOtPNI4d2rXg1WO1
08EpDHQr5NHC33g9eCBU1b/x/9TUGHl9H8MFONPGoqA8aEhd7EdGTuiporlSNYTajKoTfIz3ud6W
6CHs4Rw5fsdcsULnhoifZNUli0rmbWd/4As7RO7E2PIPopmbKz2X2egxmwSOeg16Ksy7IkllSH24
x8mna3SCZaAGt7biz+fZZBSFflSXJeHy5pFjwphJO44DLwNoyjg2o5Yo0p/WqUbfLpVBOG+WyCd2
g/EnjfNQLr4CHE59XBvgV0m8P92nTRJVmnU/Nj7JG6htQIG0lNP9DAKO6OrNOVCk9vT/o+D1fh9Q
WINFnSMNuGHU/FjflAE5TmTn81yTQMuFn1i6s6hF4oNR+/K+2ZqJ0RtjLg5zW61lVVUI9nh9fvTD
YxdxXbgBPCDwqSkdMd7WBL2UqIf2BGLiT9hsWry1jzOZY23QIbnnqbQY5TYeCbQ1vo+vUM39lwgc
RDdoEOfEhTQyCeEOvKlm+KL69XBysKNnbFDaF7htp5N+UHohlZLi3l5nVRijJKUwKb0vW/afbq8d
WXNGjk2eT3hOMxE7YdOzRU/Ot5UDq3jd26L/l8yp+xs/PXFNQ7bzyxMTzfySr1FcALjKxAZagWqz
5J2NQcdBZctKiXhMmbS6xCjbSqG4VPXxSJkfSJlmlDW879inbmPuF8wMzaYYQIlZ2oRVpqgMMSgA
lSroDfPc+MrTa9Wf9CZgBdG4exsOBOE6iT/qAqyalfZYkECikmxQwVwltmO7vNr8ATF4YNOJ/iFI
Az0SpV/AcgpuKr7fPOo+iTYRGME0Dmt0nHSBUYqAFy+56/WF6oyMky8g5mCFs7FiWZAerM9hvnQT
vi+lh4mHpzx+VngGtuqhqps/rhJkEXwkk7s4pkaFEyFQFZYCoYdVbUc49HJyQQL69ozkj9usvs+q
aVpzVG5GNFwFMsEsFleampcHKgZUnsobrouubVK8sXITPxNB+vkus4sMAlBHcTTDTOD6PUA/ECQB
/SYEy8XAfdNW8M69EPzCOF5ULnJS8GYx5Q/0dLAKTCEtFgGbk+LrJZ4tIxn2l6csnNxm8Gxk3HFt
YW+sDDshfM6Y47S8dS/2tRESfhSJYEJrOcgSduZNniW/2SQT+4Jk/obal9dpNAGhPnHx31S07pUx
3nwdpz9IbJW0BI5aGo6j8cjeGyS5D4End6tsVo9HIe6Nvlg/rWwKajcf9QBST07ycnP9rQidDDVz
XZK8fSNpjfD+UenX1AQZ3W4/0/cAKvFpoounin50kPHYH/ahvtRibDOVa0Lm2FrNNZCvrrGDTkQn
IvkJYQ094mrdpzqIkZp9in2vHvoe4qfNdxU+5PYe2ugx/W3riSRu0NpOhdzZQa+I7x+ztz5OmtGd
jC0fjziUEvPXULrPqF3TrqvTnNHyqTOFkHQEA6lZIxnAMrqf42Vwp1tUWL36dsY0EcpkGbaW2i5l
ciSgO0ySLxbGbPMI7/D9QP5K7BM89L+AyjXYJFd0a7dtfg+139Jdb3dJzGHzS6fWLV88sdA5B0U6
T8iRAm8+muIweGh9WzcghQRKk5XCKs+3DHkDryuMX6tpePaAprFQVHzgiwPGdLnVifS5nT3uHme5
Ua2BcE9Wn9rc6Mqf2QcuGm8lfL9muj4sffwwOIqqK6kYEEtyDVeU+J0XiuNag6OHioBytzvWNBuy
93cy0siIWuHC1wG/wCGulAR5lwJnGr3c9PwuXuEAkSqrUfq+NXRKYCcO6ldgaeS3UaaLBZv8d1BT
hezgMj17M190cDEBgoxB+CKnJKn3qbW5haWtrMjs4OBnNifZEBY0e3ZgOf65qin5DwMJDCCp25TX
CttYsX1p6rCdnGQeuqtjUFY7osS87Jrioa03TuxwCO8WXkH9TzSRRxBL/rOwa8Htgbj0Db/OPA4r
uAxH5w9eObodVqkhVcoyr+K2pXfBWiLZtO4H7cvGzLsNnf7Bz/9AQFRXoNpLLrgRxnlOdaRIJvWs
qP1INXUwbsqqqCrtrl+TqwwS7W+tRTHkHzI37wpFitHzi8OZU5GMPaD8pJDjZJlvKLrEXOWoVNkS
di79b6v0nsG2UT0Ix8hv1cgJ6feM9/mCPwFEiUe/I7MEfj+wqvTTcSxwS6VDuhue1RMmrcfRbMNy
j3g0/mk3M4DIKFQ0GjVMVnA/MqOfcPKyilJTTEpfYE4KewQFTC+Yp9M4PM1zbXEKjRCxFtpGlP9Y
p793fEcWsLaGH6eyzGFkzu5k6EbnDKlm7kaIucoRgjkP8uQ3l6Wh6z1uXkrCKT8SuLF2VLhspXd9
88dGLuR74wvGsqW0m+Y+UWq+gmOypXk8MkZQubEBObyB0qPtGNxzO6ZifJJGemambaQ0sHhvwknW
uA3+fp1cNRjALmgsMiJRgWdL/ITBwNvFrIkLam8u7kk4FpgAvrxF9aTLnK8dGk55qahlR4vFCdNT
63ZmdskW4WsqdtaZtuB1OBheP3j+UsbWW4B4ZgLy4Ypt5zvvOVSjkq40LjrMWfZmZcg6iZygqz80
ZN9CfHIYCzhNE0ebx8t/wAXBN/xvvRQYcW0jwBP/nY9Nsig4UaBhCZWVfPiKF4WPn3Ztzrp0ps7i
tJIbtAtIaV+hLb4fYipTTJmQojupwotY1VxcgjuxXzq2gyDy6W2fyysJ2mIYfVR+lpkObb6KjOw+
2Z7mZuSNj6OXZzGDLTYnk/o2d967h674gMy/AkzTh5jiN/hrWxbi269PHD1SEKIkt4Ut5/Yr4o8L
aUjYJ1M+WHPkBwGcIPjFYgecUVgRUqM29XZSJcv+gKUe65+/HC/LhjaijbOKXvvjdBbU5y7vq/tS
Yd3F37vYxpsfX57/MBxre+ee2iU0QNmUfB627l2Mlb2Qqbmwf4zhOfwH/3Vg7r/2ctfzpRyCvwlP
sy9dpYM9u4TTCAqJilHEzHgC0i1AC7QR44Kg2aBA94HJXiNXmOYBoWkhQ2WHaoxziu9D5UhBT0y/
q26itQZcY8wVZei2sl5yW6HkIfJzrda/NKNnwdnwzkqdt5n5DwNkEdG7HHgc274un6+D2BLH6msM
STGV6g4rio5cYKrlcmTMvdMq4XC6d7YCzMaKZtUorIR6XJbTVEo7+LOheuzb2Tpq841fBgqy+Wsk
vXGJ/gf9MOifPemnEXY/gVK3QC4sfI2VJgxoJRl4xwPWmkfWIzjSPy5vXHRnMRXMvv+jH+af2SHh
5Qb+m/nT3RWJ2qi4Ri9K/OWhMFNt6rrUghAbH0561DODV9GSdoGikcbIqeQDcSZXd1C9gTrODnjg
wTUoL9Xp/rugejOeS2I2335dDFK0kLvqk+w5iO5ZJbPQGjsSQbzDzCjt3HjVJLUuGhWNwu3cDyAY
IX/nG9g0l6iFf6oRjQW6Rwh77Fea+H5y4ZaihEPBRPxYo2hAJm9bFM1QP5aceqsRF9FDdSCue31Q
huhL0CYUXWBAS3+AfNpy5MNn10/f/1C4am1ZkKL9f5VfQC6uuW/11HgW6pdQuMb+KcjRIuIyc2x7
Uh3u8vzTMgjU9E2I9QH2XSSH8gtx7AuydCjVsoK4h1myGEprEH/CSvxI0P55lOc1tIKYOOadZzuv
N5WjMMJwUjP9NNb+ZKg1AQGNwBmPQ/gxoznnEJbhqxP7Ml7S7fLE4c5GCTOiskU3WcOc7tjMPMRP
Z7tfhZKkM+QuHpoE/nV1U3GGpmYadnKgVIJwHflcr4Uoc+xf7f17F4OgoBLej+GH1UyIF8P2bl56
LW7upqdNegIdqki/G8CVAkXIIyC8qDRD/lXC2I2xEOTORPs8WydfEx9b/M23lV94vfi3Yzxc4KVx
tDj12SoSs7LrUEMOwg6hIhZ75nEDFsngODg89skPLVzOakbpJ+tVX54A3pNuSHVoRsUAmGHWrhmn
wUpCEawMGSJooo+Jnz6uyNzIOvMrGCHaPiVNlY8aUhd4efTdwlwPPd4Qtbz4+SE4j/UPFT1NknmX
Gq6LMhTGzOF8jl4aPRsY4tgi6SP9AkxDy8owWewusqsqf3WRQUekqayR2AoIThuRvpLmYK1yc5Ip
bnq3QQjfpwB5pVRz0aFgv4FKWFReiU+KqIh0Gj2Awh6JmDYeB4UFVk4cBIMOWIZiStPEHy1ySPd7
ZQtjoK74LTXqDiwna1FA/5WeRT78uGfxD3xbCR49Y1jtg+Jvuok9wtdeCjOuBjnEH/yjeKHa6fPM
EOit079IHuWaFk4rY1BPM7eFBwZhSQqULF/rfqz0lLiWAea03U9AUY2CNM1F/zEtY8KIQ1fcjeK7
8TNDZ817C/SSXjvkL0G3QPafSwCrx511prN4/dpfQy1SkO8gfxqEObzxiqQc3oOQnTPpcZ+oISvb
DZWmpmCmK6UdQCy0X0GNZSXFVeg2+TgoDVGbUG+UkWculFQ1uKpPjgXW2UuYNnmLPCb2G7ZW/3FK
Kw0MLFO93DEKFPyasaNbwebGCQBnD9n8wN7W0oxvrWUsG49chbVjvjYzGe/r+zpbWoLpsKft4A9N
vzz8w5XCUbdgbPTj8/o66uuqWBQJOQKs6gi7fNmHCJNN2QVcRhxXnz9hx/OUvAzV0EGbmvTKX9vS
1afsir3Xp5RkO4seRV+Va7l/UK+y0UDD6cl0JeWyUmG6QuIPnuPCiaHt6i4X756YtHzS2ZmJI99Y
LYXoLzZ30e7EI/F8dfO8ub/koeFVkDTwlFC7yTF8kWdnYKbfDpTFPcGl0X4TCdk9iT7hnl8NOSpd
rcGInghcHoVJKSSsLDakJcae/UOfsZpPU+1IbaVeoOr6L4/nRCwVhSfBsB77euu9NLdN+tCk1HjH
v9xRbpkz9Uyahu4YGkHlKu+ItqR5nqeZmudlDZ+OGruozbp5AwZoZKeugjTQnWDYMG7/m4agj3ug
Nn1+EIdvXouAxjL7suNhD21r4fxMfu8lZCqkUuAPABdtwF/AVP9uw1zOlJLveYfMrkLRTztrE4Kv
3Lk00ThWzXe9YTCEp4A18onjXz5q342pnk0jFPtqyNClWCn9zze3NEaEChf4mJFSDrKY4ulZjMg/
ASHmUHX+x8SKCETbzLwB3w608SQmgBwnc2xJ2OLgxhKNlAyQ6tSdAB1+Uur0W2DiaY7hf5ry90ks
yQdH3yiuBlsG/N+pvKBOAlaXFxv87nx/uRjbyVaTQkIBuyNcV2PMbyDRQsd3UaInlo1DzuGCK9cB
r35kuQ0Z+6psEBR9f8TZxkdWP5lKXVU/8Yz4Wob2kjZFrknADv8jIXdLFNwcLTMQDHDl49VMZ67y
GkoRWed1ddBIkS+Xs8AqbuQ2/CF+zDIqsX4LN1Ok9cRslmedLoJ0k1VDG+Z00c5Rm9hFWXj25ZKX
0CORD86GWFlb2GO1iqI334Wzns0mkgY8tdR4IKDUyvsq/y0T8wPcY5KniV/qsRfm6ZJ4x1uRooIu
0TKwCD+a/wDBOH+B1sUSLijoS2DezRLe1UWOh+Sz8mPg6GuhKYJaytZUmzNgBYi1DEpFuxQYqO2r
Mk/2rkdSOnB2Yhr++s+r8rnfBpRQU/n6deu2KauWPY4R8IZs4Y9m5Yrjih4BkmlE7oVKE61D/qDP
6GOqlFp+VFRm6L3Z5TC6D8GZLRQqWxzg3yNksB4L0WH4nqs3BquTwkBw+LhbqWdb4a7lDYu+/Sfo
87u0219ifnll44J8jC6jHSP6uOYqA3r/XhflPySkfm8OV2v3sKzZlAjlWOLCHNmPIiyCp7YAKYtS
X0mxUIEMVCixVxz8lbhWOEALIy/QDmsdjlDO/aQ291yBPv+IP8iTVRF1tclXur0Tdz8BAHLFWtpi
JJL/zmk/RzgdcD6Ep2ZaOuJYPtbLGQzDbtiOho3LcvRJha+HKuqgiw4ZHAQWSlruDSjwI2EHXuAo
xakVMQds//xJAtlTMH5NrGHzWL7lZCZGklCYpOefGmU5Hftn3eJRimenpZ6Wq6PIeerO67PZ/O91
dbRUDqErBceRwPyTFjBwS3ahXA4QKGrgG8quMaEESFBX55e0X64pNbXVO+9/J3OWvhhH9PZoOddT
gLeIaXyyiiHIxHVmMGiLsl96ZZkFCXqtQfCVj2H4iNVfqC3lDHV6GVbN4VkKC5mBaFAxWTjwlr0G
9Rlk87GtzrhrYb+5L7N+xeB74TP3UMkLrXaTjUGMo91RYKjspYiCo9N6/butR0WIDahNvBJZBXxC
6E438GTyZMfluVzFyuY5ieQtVMDA+gvoHYQdg94aPvXujxQ8q9eRE+GNd7wBIFEE7qckhb+Xzjyw
y+6wHzverzvEX8WbrVhWJ3pWyPx7YKP2aWZGU57lo9i+JSoAj158RnNUcBTT0Fu/d0ye2xE0rydG
Ik1i9C+nSHGMfiG+/LKcu8iAaqMt13U2YWLXeY5UoGKvdzLGYyqD/n6L3zPDgIfUPMIoWuMtiHvX
Ijyl1DpRfuoIXpaew9Xztvx3xisS07twGxSPrfqWX0smfq5jko06rhXXq3K+unmxhsoZX2mkM5HV
MkaBQd//bZaf6yHrA3ZbxdiF3r0kDS+HZa/EVuKofZhQeXWYQV6DZ6Wb+KnN+qWf9fCzJuklMERW
CsJDYFsg0/lkFfzicmgg7yY8CfCwrkfGwvoGgNFyrSkS6+WaUho9cv1QoLm7d4bRchaW+ZtKyRti
8rKjK9kCVVpuBAa3/fBU6CagM+oFVeShyfWFIvpGEgg/0wodxJkse8ImLDFrCb2VXYyd8jaPC525
1gwWBLVlkgnWss5TDYNEMbW/Ai08ZifWCTlNBON+BlFfN9ttpPZDnF9jG6jsrA8j9ibt00qpq6uM
BP6zYYhFwalYErjW79T5r9vkMTu8E4cntY2Elxf+DDkNZ+yyjxJ/KejKBPpryzOYemzXDaw5tNt6
sOm5Q6SL31v/zpaE3PBRg86hmEphjDErcqT+J9h/lgtbuSHIccRv1CY6AZig6660luWNVIqiW8Q0
gO4QwA1cX8YLkpjHgJqE7Y2MUHZSvn3y6r6bVfOt4Q7F1R3sak/Hq3vjCIORBc1ALBirJcXDNQev
WM6wm5YVwuIRNn6yasAucnxnFwYcTaPXyNxAiArjFu/hUhCse4OsV4r7DKbxmMWvvCrGA2paSJyB
I8Ebb5h57wmu1zflxA/9KkkLeuVL8RjmgoY2yq9w+98P83ztjTfbOorD0Mc0STPckzS7syszD3xQ
lP+0mNnZumC4e7mzJFIr6+V1L/rax01GJBoGLB04c82+nbupWkRsqDXcU0eTf/PhDMU45xx+eJlQ
bPbWw1Qi8gdLt1h6PSQObAV4y0/HKsqCbGiO7g55x0EZLeootTzq8aXV44+qAN3mA1aT+sAMPLAm
QTfuKB9yAT63Hu0c//f3ZaRdQeqVKPAm51k+zJOOFRksR1qzYvZOpicawF6zNw+6CbUe6VM3iZGX
n8eqALhOs5pkjVqA42v+tWfQ3vdSGoWlLpsXDccHWbMfa8slbRHMOAf57qStqUBSm5iiY/S2fdfN
OEMB6TSDQGVPvHs1Jsf/boAmpb4BY14dWkYyleXUC2bCJDOJKeVSnN/ewFrlyn6OlUX6p+U4eo24
gSK7fngJjTEDC9fboVDBKx7NgTHdQreMfsjP50v1wl2XC6cBx6xlseADYLabIq6JvblY8SmmQm6N
JfacJoQcTPdjQFWDwrfjKzV8Lwm6FT5ADF1MU/Iy9N2f5tWB2cqaPq1kODUesGSbGVeeyYxmqfnB
nbX5A3ixcRKgYAreUUhCnKcfNS8ki+hyzNURHMP9zVl4Yd2sjwDGswxPBnyZaYahlWqeR1au0qSK
OpjjPnlryx4B3pS2FKzsaKjm9b2YVCDBISL0/wbFcwWGIrZbp+ulTaDSYyv7RuRrt3Ckxt17T33r
tu1h+4eGRv5MXidw1L8tSlV4GvzNKJ0jpdZ4GLoIwJCpI37IJcqfFk6HEs1vek7qdStypWT/raGl
GfS/fPN94+nUxE5QO//C0yDX4zlRLonB6GhQwYvd3mkNEfhREASNPtQ53gPcFpD7/1HukfdFJEoG
6oatmvxHQ3AN8n93gdPj/X4g16pEqXhJTekqFRnC8oWgvxTtriWmtW0DBEvewq2QIUO13L8gZ2jf
ttWGCcZtdxKHJLzq0uqATMWYQT7QrHiHU1uY6KRST03G2hhiCOHxNJNgk6qQ0xL9dtajhYTxOfp1
UEf9LyHIkiG9CVTpvQ1MNlmN2fK+Et2AMw5U/3g5omFvsVMYJly2xQNHtTX2u8tFYNoOZuEDB0fB
bQffkb0jHgMabyYEJGRAdoD0wx+mRaKcU9oQK5MjfnvymgpUEasXvddVm+A07yi3c++Yjt7YjLZK
9i5sApWUWSwKvbWK15TEKMbHKFix5H5bbae0BMeoar0gY+yrtW1d43tdkBkp9JI84jaiK+90JcwQ
8he88Se3zYhpYYBEhEGAr6YvHevSH/lOquBonj6hj21e6C/MiOn/M0cG9cKQIa8mify3nVDK6Bn2
onaNbKxIwI6V4Ue4NvnId1MkTQIN9kAvTPt8oFshK9P/toZ71ICuJm3p6M6NIbuYYAg/gOzBOTRX
0umOgg4u/jDlnVywdaJs6ANj9fY5DOLUGcpcALZHFURG2OtuP4c5uK/53hb+eHvMs0iq81eNUpec
1AApqSKUQpdSWDREEJCNf05srtDfKDUAdZFKLVFPHtO/84NDGtpP7NYZMdd/va/zQJWnmiX2tOuV
VZj1agm8XFelEJcoLpfsRiIQ41hkc3TWWvaBq+k0Xj89fjl8RkOWcYnVEJz5h7DhocDjkf5fLr9q
IwWzuiZYERD+bTN3+cW20iT00yXdH8MUTenPsy7JRdfdolqqLZ0kBZJbK8z1Wtjfa5H+R7ApedwO
OF+pMnGGcmkALE+YkjOH88C5BnNgGFhSRNi8kHT6ennYdkjiYk073kCKnVg6qJxxAT9jZbDNDUKn
8isT5y51B8V+lpgank8hKMO7yGwcO3MyoNupmUx5QOE207QqDIvDi+BhbhzSicB0ajUPmb9uGy3x
Z7sgSMC3QHCy4D66Hv3KzSbpitpsoM/+DRZl6/GwO4JSe/NMMjTM1+/XoTiJvyg59Y8fL7EahBm+
oS1GGMFUDWUFpYZ2IG6JvNirCL8hyJAnntBrpVqQmb7fosA7EkL5WdgSyGy18rx7oCw9SfFCnS6V
hLb/acxbyIR8d1FHomyePtGFsd7/v6rL+gGUzo5tIWjJvCIgd7+XpFfC9c7hCYsY5lYxpcNNXrRr
YMtYJrJQgtXZX/TlxbKs/nWc72JiAqXUOB9UvpwyatTu1aSfffNHOZ+EWCwx/odFlc1AsC1LQb73
ld2FJeyBwznHVaMJG+WCA90jZa99npUvNHTq8aOzkPSI+PyR+TfVO5IDL4cI1BIpXvPcn9yftUJq
DWUxM7VEkEZ/ycwRxH/VJ9YEDO7/v8veXuHf22hMPHMIyuca0M6sq983Vp9eLiNbtr/HEiLuSzGn
yIzTldf1/Xhr/L4Y1E9+qF6ASk2NnOSIvTtctSFHwaY7ic9poOWJ7LbAJSevBnZAKgHn0kYzXzBT
bUGE0eNwr9kd2yAWrNCDPmrhI41PetVhG4CW9QpbFuXi+hV6HQR7Z3N6vXCmyEvjV6wutFUyYiLp
CB5awAd48AOsc8TuYov3Kj5w2pDkCJVdC6KN56dpf5NFSKcPGGPJMdZzKO1Rh4gsNr2ztgOfQxYd
uEHOK5Ck3H91zW2OMIstuWh/dHdiRTzEwnSrEKDck458n0J1pApWbavjCOSZooi18bp9qvZQNL37
Lv7wlIVsMWPlco+lNh2emOiVgsE9TinYjU8fbLMdTzC4pimA061MgafGDMR3ktQb7AnelZ93D+w7
9v+KJ+juu/b9OGJjYo8Td6X80NjsnFg6XlQhz2W/9AKqhIFZmrgbdjv+uLbOW0jcr7SlE1dBkDaL
fVDKuqGRAetjyrUFmtVk69NcSh50jJTph/PIPESJo9mscvbNKfByrZ2h7LwKVSNb+K/OxBb9XpxU
ljHIuzgBvarJwokuljmHJYS5fpAZmw9i7vFtML0ES6+4pmYFobQu/CgQyXrhWo52eXJ7XZfnrAjr
2JkzaaeuuduPlkNJH1lV5zzi7h+EJDVPoUJ48/RxR2rCnfOekCeP6veBbFl1otUpoA2jWC8c6Fd3
VCR+nqrQOmedvvjsIQfmJH9itk2b9IIuvFpCrCLhyC4aWA4oxMysEfFSWVYI3d2zB10Q7Hy/EK51
3NOoBUPqzEE0jEFw29G0RWIP/PYhtnkU0dRkB4w3Tq/kOrScLVT+G5TYVq7zZgBfwllwpWuSl9GK
EGYIomVCLP/vwQHy6UJZ8C/UXIeQh+KoZCHioVYSXos4Qt/cMSASPW4gCelD56M0j7uyNEnkU92e
Alegr5WLG7zK4YU/9KMaY5lnBUXJbkTi9lUIxP5khUW7l8lCi2ZpxzEtxH3zArwc71mswywaU2Bz
a966vnQ6iu15KheNJf2t1oHtfHxyuKMuKYms4ytrH14FAos64JaXis/PhYkC9wQyryeefk/kGRFE
XPxXmhEq+JL3WiqzWrU5js0Ypvs4k4RglCFd9hc7pTbgfkyb+TRywL4EGUktmcAJO3at3P+XiHaR
5StGW4Lez5KjD7qhUbJs3ftA40S8a2Z9OWI7I2ONJ+wmTJJp21aFWPS9jyTjMsHaeRb1IeGwJwa3
BhASvM1un/4xism3bThsVPoVEfIhwM1OG4yiMXzbEhL4KkqaGjLUjRaxAzuGzox2t9Kfkh7H6ve2
vsR3hPq9CiRHlmPGoMr7QBPBrYwHkCdlCUJrMlsKFYMNHf8r+vg3Mdm8bomFdKGYcAY9QDg4XguC
IrYZiqgfkCOMhK+7oLxHrT1UFZBhk4mxwOoqRaHZaUTIjGbjX179Su8W6UcpyovZX3PnF7/RLZlc
7DX3iwM+S4B2wLReBWEc6nYfPo+HC4IzatF67P5jxN9D6/354tZTZArUPxkaTs6cWpVZh/5gtZg2
5jhOyhEO/6D0WtfaJtWsa+3Y0vzcbTgdto/G+AHcoljx2PdOXpeQz7xeHOjz3SFalQTIsEy+kFYg
EuYgUQSEjbZs2YKYOxHvM61eMH0NkuJH+iQaZnq+m91m/pGV6qiTX08tWSsjAR1uLb1IyvRULyAU
lmuV3NeWPfp7ZgDSD4yvrPuDZhdWcKEkuICal8qDvpCkE5TE4KXE5jSC39zR6HNMqzU+jdHD7wmc
i8WupHJ9lTEGs1t5nP0+BDu5dpa1LCn2c30z9cPE3yElYxo5fAYANk/laW/H6wktTnVfLYxmMRRV
ZKkbkBiD6mAwuAOpqv+GoKC3Kzyl0MxN7a7njwgstwSLON8bTxiQ7dI3PFFBgqsT+PILfqOD9Omg
FWqueG2gdzdWBu6yjEPbYMaFYq1Q39tctll7EZ9Mdj9o+cfIhhW04Q5bv+K6yq0gOKe3+RFNLoy7
LyjOorCMYBcX1PTouOSIvhiQl6lXLk0tojeKeofbfhD4pxvXSivOVcOwmAWYxa0gAc25NGbo+CvY
Yjbrl77Azdjoa4OLiDyMAc22QQHJFTTjr6Em1j3Heivt/3QPbqDEMoUiWXjWt7rVLj0J34ZDvtLI
+wmerkiSd4348IeGJB9c7pIqi26Po8DFWyD+9G9vkPOQYUzEQv4+qK2DWPaXZlFbHNLF12bBUEpE
D6iix0L770DerEZHi3Siif2Zc81XlBn8zeZsixXF2+2DSjyIJbLoXuOeMx/zfmC82IsS5ZEv2fa5
btjJ+SkXjIrYKo5NODxRQTQHmbte8ZAfDNCwggxfxKmUoecK7o5oEDl7iCZ7lqnOSMjzd3KXYwrP
0l6y75iN4KuVcUOfD31AS1QqLxc+gtJnjxPiPsy8XsHQ2rsZ7W8qBCbp2HaAgoOd0CW8OBqCnguA
cC1KBO8g0XHdHG0X3D352vs0v0fmKYdeIkBogB9kXxAnQUqxy9no1Em9whSRM94iocn5Cgdr2kDD
8Uiu9TSpdVE1yYSMxmnWL/PdkvSm64Iu4G+Jti6b6EJ5hJIXE4VQMR/1zdmKFduw5Cwl8aQrmgT3
VGELQSb5IDZnRTJs8U/2rexWIRD37NLxHHFoN1pgT7wPtwWcFJ58N18od+de0Su5nnA68HWVpBSe
L6Gc7Jtb53WUO6rJ41NFbuTJNQ90xz6AFaJ3o/VYuqvKyMJhP+enRKDdYVeqZIwPPJC73cZZundc
ZgxfzvZsS/B4SaeZBSPEQCf2NqAEM60l89vFX59celIgrGcItLYVn9ZK8mG5jY+oUVIsSjK9FacU
JMU9jC/Bc11hH1RFC9EE8I8KyitlVQavDHiMgCaSiMZ2vdhGIaHSHLfHhoRbuHHM01YWMoKiFmgN
KrCiZTrXGJQI9Xwxc5itGYn3KmtJArtdO0nDMHMTlWe0PSfhV1dXR6UolE/+DWpX8Z3JufwOK/20
0+pJC7IscEPdJIIhan0ysGKjVatouT94HNAaJZGYdd9sYuua8Y/5NTBUXkocUwe5eRNTBOMGZczi
+S8P4hkDMkf/xwi0Yc9v5MXSpwKDj617mRhM4VTkWQtY8oTFe92pMEZkQxCChflyTOie0lWbzOxO
zc1siMB0AQOtjAdV3HpcP8NquBO5SNdTy/AoLkF7Udp8OY7Qaqs+3b+d5/+zsTnXKadkyDJEVmG7
FutX0Eo3rc53M8bkMU88t9h/4EU+1p6vd5YMFoH2/rVEPEj4U1xxn4hD2VTnd9D1HR7e0SzhdqO6
k22rHXA8CiHhmfxYeYBuTs7KieD02Gz/Lle/On3sT87JCAbwx2P05xgmFLj3uJm6O1GAVOzSDGKt
iLXC5ecWYMlJ6t8BFR7jkuPJhysjKiywJuIZamYKqQHpCnxD15ICpoirx4qChkRczuzA1UnNv9O4
bIG330LZm0oc9sNBt1c+N/RjiS6dKg8+DeUKE9gfQPjLl6Sx8GMHEPyLwwif45hxgU0R21OAyO/S
HKsG7ZfTrDJ4j6kTmmxZvcaDLsunK7fdois1HmxM9IOwt3rfV+QBr7XiaNOLO4CJA6thWnziRrh+
NN/N+d154XgWW8SKHEb4DC7kfXK4u7iUmBpDeOiy0Hxv7mXTA2RjtYBsNFd9aj5IRdt2STJd0tAt
m1DwMgLWrTxbEomPeOyxHelegr1+klfDkQrmIgAste2cmc5Lo/kGmOtlX//qG3D8IVVwmAHXVkIm
cDfPEH6uem+4FFWEh78Gg8VDxRIbQynvNSqj9XJZQe4xDDrqHDcnqqCKxSrrpGJCo3ZSUjTHet94
VKTNvzlg4JdDI7Fl+pwu9KH0fJKAxYJROp5VJP0cDIwFcjfLHQJ4BwiXj2lxeAbXkvRSUwTbccwx
Cp4UwUzRfWbJnd4IqJfBzKNJJOV/+GWZrsadZdKZhChL2us5IYUcrFqXSOx56gJEkBYLbnyH+J1Q
o37t4YrcQmWxtfiqMB3RwF/VAYzaVtOssR1pSFjXYGTHB9nTFJ+ObI4XiReSDP5kpgXRgCZd/QbT
E6WFY3K9aG37GhqoRCJBy1vZhEJoSL9S165JNIO+prXWzbGQ8tM7SZttvLWANEexL661R9/H2toj
YSe5KxnX735Tb7gMn/mCN0qgTDle3E27FepwBUcq1M5pZ3O5tXCpA9bHNN0DjxPJlw134PBH3UCY
VwnNy8H/BhodgrZncH3t8SO4p61fgguk+Fepn807KM94KdcMYtzVbcH6Om/BvkQnAeYkrFEUPVnE
KjTkwwvF2/lgFV7fBUkowbeOWmOwcOAvy4ks2BBz7yGf+mgktCSwsqX53qepb3NHyh/h+5WuTD35
dwSFxk3QWFWtPvZTBup5Ye+aLi63Iol1QHyynifao6OPJ8QLfnmtaXrh5MbRjgLIAQn5pXzRl0Rn
IJNdelfK0Y2mrEy3RLMMMY90GpzoHrfTCOjEZtzLtBw2kv31xNCKqSECduHOAwbdCaHVajv/lcUP
RuCdETgvk4ZLvhQIh3eh9BdiESF44i6DMhvvdCI2rmnbfqFsqqu8ueijyzLdW2Pp2c6cTAGNOWFv
FA2XbMfK3gLUjogfp/PKaG6NlhzNAWYboDLpxK10oMmkA3QKXvEQjm/LSS0LS4iFF8h2tbQjbHhB
TzlIO3koVJCLbQQtTLk2V1374qwEuDWgXD0Q50EuvUdGCutILtYPNM8O1t1mbkKD2eQPX6539J+b
FPaFXmmbH9Mfi7BA3JBS2vsckOyxcjK2DK6EfHnhefWUziNwKfBmR4XwB84vqXfGup2f1UNTE7Hf
AR+/UtBpDx72s9DAGz9ZUNSAMhDDah9pUM2aG2lPsW5ZrguzZ9xaUHnfvo4LZ1huVEEB/jBEb5oM
l6oKJBxCjjwz6M3atTDssZYJ88U9wifnHdq8gNQVxgfx1PbLFW84OyOQFcn6CHWq/kvdjHPhJl0Q
hwiNzX76i6pEGycj0aUGn4DmStqUPbfReGBQj7fNlXcvKTrzcn8bA0J8oQC5hK7jq9t93ohCPyK3
rvK70mucsE2SOlLWYh9DYl4iWTILsYBjxgnyAVLxxqbcvqLmSe14TI6tziPd02HEL1PMSGw+NfBv
VJikgrDQjvOwdOuECyoEm9ftkUNUhX4fxwv5Xc7n3plAwsala4gMM6dZQ4gUxVlVetwgTf+Zk2Nm
v71JjAtdfyqPaYxsSQRqFYkhULo4cMoaAssFeU1QoexeeER7+sjgAxl3JAJB1Nfhf8io3JgGRMeb
LXeqZPEsdlwvBGLtTpJNS6W0UEgs5EI+dpV2IBuEF8hA3UX5AjmLTwPismciK7yL0ddoNHKpi8Rv
iOQbLsCf847ZBGUoStH4Bv1qbfKpqGWRPz5XPm1bYdlKl50FmJqDUWrugV6QRsLNIt+bQNG7RMmT
eWD3uugRSgkMnber+k/gWIbH+GkbclnITf0FssJH/58ZhLoA3CieL15ffSqtMQizAmrBYMwsMhgg
swBalqDLX9XnJrj0dtBKwtTAT5suk2Yyr+ZR5J2rzVnk+T7a0fa8A0a3jaPGXBxU29F4EtG2S+AS
AF6OnR9exyXKSAUVYTQ7d0CYNf4nVobtv5DPyb5ERmSfEtK31FRUbzaXyFcNUyVUhLZ3TblteWD4
Ao6jMJQDp2tDWaFrsrUMTvLV/UPtU8yAVb7aKjmcDpXjeIAz72uBb+X0dQBz98onbGZOjMEGYre2
RoIJFKTRtcsnv7+A0p9E/oqmLr7UVe67Q1S3QfBphW21NjXK7ZI6g01hThDGJVxZsn0DyM6Bn8ij
XluWp7ZLcgaQqylDedZUH22T3e0E/kTEmcAMcR8U1QMr2JImZoboAQOxJ+OeBmvKMRYceeb3eDYl
Am3oPcWfdU1rR4mECwIOB5d7FrAb0mU3aYoEIDuHiIq9F9I1vhAEIAGaIWerhqgmbvvRoEESz10y
SRV1yuQ8iAagyFJoKX0rMuE+2EJATi291UhlQ5Ewj09lI/VZCjrHz9LNYAV/K3ngUO1ks4vLVwp4
+SmRKThf2wlSehqptl0fN815/9q200DCqdio63qTq+CL03IYUVaiDL0OEiZ1nXlFzCL067PUu3AO
iR+kpCL3cM6R2OrJStr002Ys/c5cqTKQM1h4VF/KODjuwqTatvXA0k5ESBQ6EAmwLTa8uXgzrDGg
Q7qWsKy1sJudbUn3uH4Sk6gR7FvEnSrV0iVCHlPbho6B7zrqzqRMs5YFsSjzl30dMSfTaR3J8Zv2
hioRlny8ztxyVqieaT+3V0GeHWw/MORxOhpFN3NIBIXXHT9csRlziCehNDvwtcAq7OypaLhC0t9A
8QtHaZqvoPF7QS5q0V3O3WfByEwlbYXjB9Cr/GiOEKAdDjw1PtiMI8dkmf2UoMP6p+aAGZZqkXS6
mouGprvr5pmdsvSUYHTH3bCJicd8mzK6zTR0Jy1iUtkOUUAqCdh8BCtxtvUcRnQiwSwHkUEZClGL
by5TC0zPzU2HmQIKr1w8bH3cfI0Vqc0+rdsgOn6CYe8l5i6sF+Q94wSXOTx1aXAF935TtEaYdyTe
HIdZbDmPn/eEnfKew1aqzqY2Be4HPM/GfU6oRC4KZfWBq5O708ajd70FKd6PBYyfp0QGInR8sSDO
b9u+I0QL/t83Sx52KOZf4eBt9JG5BdTXge18nEIjEkBMo5ORocZmqmNtE8P/3ei0HGjHhS20OqRO
nUOsDbjA1TWVryWGbsbIsN2QsgzdCcwkcaZgCkgT8DJ156OdNscgIcQ7zklayvq/LaoQ8rVVemPe
zP/VmaC7IZ8fVDDwxG4hCftVCRphCFc5WIEuNMhXrDxpEsNPfF85aEFGaHPYGcHBeR8INxFzOE0x
2kP4b42EtXitWxgtLXDnu6fbIwwl0LhlDPqeJSzABAVjMbbOvWdZnpybygZP4bbBJdYH4Q1FlDe6
cQujen+eQ0mMcyw6YeCy2CAuB/5czJyIIsY9QnL3Lm2bEyQyobz9CfD+V49hdwpcw/pWoHqvUOU/
WJHoXFLqmImx7dVzQ50iz/V0pYLp7+OSCAxOrNt2MnklUk4Iur9M7Scp0hAu7BJ4k1x09lj3TS3B
HYV0fbJbo5NvUszRhd6oiWFadx824L7i4tka0ipXghgY3nlVJBk9i9SUvhwmKbhUV3P0lPbXTOfT
04PWfmsE0B6Q/LbruVxJz0fK0tFjv0aQViDUAV092uPahl2l3jazSYF8c6VTzGBh1zQrwnzg9B2C
1XoVjVbWWF94MMcbNSgWb6rdNxyV7ox6wSFOmIRDF0mgL5qfk5FkiEsqkHeWNwUIv1rXiR8SiTFp
qARVUNBc7GT9XYOK9J/3QgDGl1sNJ4aPoq8sk9j0+KDk741chkonTjacdwDySEyPbhOr/nKCWkrx
zjixUwWjQIujdpB7cwlz8ZG4QWt46CCoUa5t7eTyJIWB8gUGzop6T4eBJUhVRSAC12UKdQXEqhle
My+NG/an56w6gU5SuVIANO9U1c4DWzln89JKuUrPZSResOh6R5oR++k+7iwCehYAHkl6AdCn2jGB
IODZ0Q1RZrHvCKHzmNUTFaiA6vXFvkvOdwL4HKGdCRP3lT+46z0LxsQZxtuCN7+QEeCNoVZAfJdQ
/TmkcD1XnMB0M2FVk05WcIlFzvBAPxJh0d6JzlsJlxbXWHIIurqEbGazbLGCkyphHdH90pcBA25k
wiSmNKPxZ2kTRjza9e3QVUoRZzqxt4VLe0ANwSXE1732q2HNxaco9WGhKwRAP2w9euBOcb9+Azcg
xaeo2ogyzVUB+TD/bMKdUSIBIvjN+fziIwv95JRFKye2J73HwuW17WvRf4ZD7W0ymyCcM56uPggP
4LwO3WjA/pSXagB7+SBAoB5/TCKBs+lHIJvgPiz1n625gDtBUVTYX749qSr+xj4bH6m0t2P88lDN
Mi7e2tkssTxAJr8PlyfT0ZN4bfsXv0JzU2L/9Ki5r6lrhA+6TpA4pgK7bCKcmvRpnkRYy0wxlIvV
NctAbwJ0w15sfr3+Gud8udqxe0xZLFZUaBVUm2blg3K6JJyzF8TtYBilfOuF5DLsJF1Q5SRro+Cg
7yq+e1xqXvmdwVYvIjwpMt7QGD5PS+soNPNxtUGNMKCWkNGHE4SHFvTZ/g1S1zvkREtlnI+4z+kt
V1ZCYY90i4dz7z19uw1iRUf8c/9SwvaNGdOLWRbJaiZe7Vi3oVzo+BbYM3Twd2XORfl9T+d4DVsB
bGoQxaWP0RzmabAFULObkxckMGT+nmbo21ATyJ8lUD/g4qFH6te3/w36e4M5tYRWWpgjI/wC4jme
agPxafjWlXrw2eL2Il4Kickk01HoexZPxTuilyQRJAZekQ7Jt/5ONnE+L/wHVNfF3lKcM+ZXEoiK
eT+j2njUT7utb8Cn1mZpEiACnBR55mGzMVPKN22iqKcwdRsME6XFfDztKFEmKeVjamvvyAmVuzsT
WOdVTBfbnYzYPYqk+33rbR8TgybA1Ui1kwOElstj6aWQIMvyPbl4ykmHdlTjlN20iRaHQgXBKjLc
E7H2KkXlAXaG7uMHGDe0w2F9EE77g8mCVgXcIn3wmpdrLfOyTKqHgQJJ28obqOipd4EsEfy3CFcn
/JLJHMeoa4hdAMpwiUjL8RREkJEiPPEsjtkj+D9120PTDHU+O/+zfk2c/9jxFMfgFW5wkY/zGbYf
HUly83SZ89ZmoBkMF06Bnw6Gf/A52yHqm+/YzB8eQxBSFklvp5xTa1pxRkZedSy07pIvhaUrk+2q
8OwZgoIsXvynS52VXF4FoNyIol+FAwmjWTYFXaHhNsKmQ7M5LDZd7uc47+aRQYiigKMKREy+xh9d
xav4cdaucpDh0hpeNpx59issuc2OO3J7GoquCH63gWXhHeQ6MPDOorUkakxTxISG8RUFfTRgz/n/
/SlBq36wiYLkdWyVLeApnRht4u0Kw8+yN9tjDroMVIz+PR5fsi0noUQ2+O07qxYOtJHEObslu/W3
eKDsXFykKi8HFwDcfpOg9tbA4n8FhT1L+WebUGm2FVwwLQzAv1ZIH3hZ+QvkOgZU75x1gBATCF9h
2bHflj4pOjEvcRlCWDN7SMHgxO9wTYHBuaUUdVJozy2GWFEZgRs396SRiTYrUKsV3u6nJ7ddLYFY
uYcVfmSw0AIub+u2u8Wco4JsmtqH65RKS7ygMfdn9DFygN5WhAmIpauQ2xjPda6l/eY1O0REo86w
MpDz6ZfIDuxzp8Kx4QJKj0xvsP4RVBOz9IiQhkrVjY89a5DC+lphAxxUE4pUB7tAH+kOES2k632L
h37tLcNjl/kNpQr0s/1zVQ2LAOLYovxzDfRL4IrcI87hmH/0P/OWJxRv+InietrbtrN0Dhc+vHrf
WvHj/rW/UL7Wd0MKHwRzERrOoSlrRH5r/lpyvLzVcfdEgkAEN36FCADopgF/R0z2PBfD+4TbEWdB
Mu7IA4V1SyeakONjRYesZ4o+dIWpk8+WYcn4GgQA/OycJ6YZc2C1rTwQSx8Hk9h7N1f7S+O5tGe/
DBeW7xcMjvVp5RMtAylD6DBfBOpyYIQAJ716xt+mwlDDG14/PIhHlNdBRxe4lrbs7QsfyqZtAt5T
k8qbgbXN54nyPFk5A1Js+gMfE9CmgjLapdQyD61DkEoo8IRqOA/FJMkNjIVy8Ql1NHGuuKAlmm6I
mpIq8HIiYLDVdUFmCoPlBAEoxkL8cjzOt+jaBFO98l3PDgGN7WN9HjREoQIjxqIxto1niY3TG4ea
KBddVZ4dFbLLr13xF6wkhc9iYWQNlMGNTqpvo07ilv0z/D8mMP6ikiRYa6rczuzq+HhNCvlByLZ8
eW8ECtx1BYwp+X0HjP35CvU0B8IBNThEyeaUUOoW8/t/LZh1Ns0HTDr/7Fo7neQZaPtH5YRnk4/U
7bJivIbkXYtRDhMJmH3R6yrcyyC2UPyMUDDH5bcJalv2j9O059NKXEezZeC0fsAcy4Tlq264tn42
ZXuCxl6PGJ2BBMWu+eCvEc7m2jTp/5N/u4xB+gP4BUkeYebxU0oC3O0V2uRdVbE/vk+A4kRMnak8
NFgv28vb1eqj1A4wPAnuhKsvh+GDtmHnZJRKwrC8Z+ruVPlUCzrtgV+vd9huMH5qW8cXRcLndjJY
j4zJTEcj49neNDHQQ3ySGM2Nb54alw0uMg9DN52JJsKqxBMY9SRxbL+KQlBJyaPvc9/KrNXziQRo
0m03fz9mLgHHcm9dtqC4Z4UE8gAoARj3GBO3GYXPafC/qtmGUAqHHm2MDZUSIOAHbWMR9ngNNABq
37DUvbDFoVV+gOYZnMgqBF7jFW7T0MR8/caz0N69oEjkEL7ni6uXy25ZPyzl3m7Sfi2MQeynd651
fMaO+/7ElDzVqdr1LEtt/nOcdN5In7VnxipaXo8AwXThsUtSxOjH5a7rPkmwvKITMmw3px1hNcy1
yrvAltdEzHWIZKpXGiOrD2hbIJ6UTKP4CMkIJ3hLlXyfj+d8wMJGb+H4bax48FASvAYbeFkFFr3i
NFeSWX6zaFmKG3B0gHAVfKdmFsBRPvHkkoBDrNg52oSfIP6SpyOMeCoVslyvBcoSYNdbYFuph8uI
4x3qNM/OEpJATvvtiu7m0FX0ArPM9A0Jl5LZjVBi3eCCS9yCyMOIodMqstHkOK4RpUPQM4ZNovcX
qLz0joRe1KLeoFZMJaBwDezLVlvbGko/oEYQgX5109kZJD3OwYcAwFHYx02CbMywnIYPBSv5r3/J
RMOlqYweCBg909O73zucBFcb4ZaINYhRKBIDYwXFdnSeLChBtQRIL+QwGZiU2PxtMD4b+dI3Zqcm
I79t2U1eMRSeI7iI/nsK8EpmKSuarSzUVlP2lNC72el2SLKLW96DNYOHmTTKqblvfMAg1qOKa0zd
aDlQo7GU7fO+p7gO7Rm82w5szbUSJ5YKM4c89CM1s5VKHcnUaiJCRRdywP9yQIg84LIBLUMNlx+q
ly5EhPkWZq1savpL50bm0il4CpXhhgVlkeQT97ALyLalTwPruGsRz+MigIVhG3zk0TT8r8AlHDeY
s9+TA+yF/bvzaEH4MkoacwrdYXSuBOkonYA5gjbGGiVwv8hTHXclrS6VoWvdvuEe3dCfP1CRh+iN
UHJDEy/Iysp6pQM5FnfZJ9f3yQOVNOuzISOJ1DtN+0xUVEk2UOtgaXHHfwjk/cS+OGhyvZ/O9yGY
dM44w8DEQPv0AdCtR5bMdJp7DLFmCX+i4W7ugTD48doVe3dyQ8o1qEpkXdSWuyXrDQI/2GQ0OeQI
6KQu7+XIw/T4J6KCimasD30WG8ddjJC1f0UGr1yhfX2aHAt2epY7eAshSS/zEWy4JoUvX1MRs5dq
VflytoL2QifdzSvunt6y4qGuACvFjQ9xCwzJEWH2HQtn6cQQu2NzRrBn859Q7f43XTA2kX7YYENf
c8xwKxmjw4M0IWlY/ZP67JMKjNc5nB/+XRNNJ4Mtn1zl+wTWQD8wr/YdXIJlNq4jK66K333TSTJC
EbiCE89SqvCLO96Bf5vv0KiTnGguzz7FrCqQJlrfoAOwDKYlEi8B0xi9eWTIcaydLUF5Y8BHHdoD
zmwi9nIrfhw76AD2rJqgluhVziX4fqXVFbsBhrbVYyw081eEaj+az0+NAc1nwXzXBuGtBBI5HQKh
k9yW7QwlCLOX/xTzLx99tmO6PC4QC61/f3xoafCAmC0bOIEOxfBimtdE/aQ7jVK8TiMPh2VPMdvQ
0CYJLQbYWhCO8rIEL9dk6x52HUAf85ah1iUCojaKuZZo/aYkl/2H6GAOCuwLWJtrP2KbsOjVgS2g
WnNfcwgICat6BkHiBCC044rParlXtHw373w7nkADi1cPdz0EOpcWO3gOf2Lj6H1/v8qy86rX6TlY
7uG1nn88IbmFJ+v1PekzTYC0DtmJncZNWfg/jEgHaEO3s7A3xRsXxmZvr6yXFlYwCKrFa2YWNK/r
U8s1DabHfVNRsUfRwUaDILmF/PUATELWHI57nSCeHNF1AFfNMef6shXJlOsQux6hzYrGixkGOCg0
dXUCRjD89GkfaUg8NkOCb+h63VBwygaTchcDvTzpr9sGrUCX1SC89tnA3oK9zj48eBF9yPvfMJxH
ZNTtgALiJScPaWGzsaR9Nn4NZDvoW5OqbGL0xJswfnpRGh1h5SinabZzuNMcG49orCZCS6xq35Q7
bvAYX7OCyWfWAM301uZ3HG4DspJHzdB2XXcFxCL3blSkBQ9+TjeUX4nUHMgGcClLFXCbSJkyeNj3
zrBuaFaU+9QHh5rQLhw357c+e8hBTZh/azNnzfL5HD1FrNvJJk02oOlWl78cF7AZtskssLljOwtF
azeJEsQrdxaOwKm1wM716V2bfcvBVPJzT8Nb47B25n4vQ1VTgLd+7A9Z37A8ptLQtb2PZioe0YrC
9L/UD8rBwgSprNkHydQaPyNTo3Wdhf7AY0N/bdrfJLu9KQQ7jTpxdOBynyYeQmng2/3JOqodMgqy
GvTvUehCwRBn2ajK834mFgLCZiyaLE30ml2P4TRZ8S7D0elquQzK8Nnz5j4BRYq8dfu836zAWXJ3
wD8Gz56VbWJecutLOTDNS/iIecoGrEJlbaLW8Nn3WnWiYcRjWPG2iMCUjNPYSZ3iioxwh9FRHCwc
xTsXGK1f1SBnUCYageLEDl5fcmTEKqVOW5xiKGLPow2+NnaaCq8ZF4D53ZlhNXJ2XvMFKW8XA6W+
/sJ5RUWIdVekZZszHe5F06dcgX202RXRTPqgfbvWkor0Jfba62JRnP/vZV1DjcGTnyma0BlY0k8b
XBdKncC18krUOd1BCu32pHB2DZLDsdBugEG9F87vlCqcS4GZ0pQFUt/BKSwrQ3+BFfnyAQhpDdck
sz1SIKfdAyhfAsH5JXEWOBYYO5k0pGODUpuhXzdo9gDkqWn6PVxfYz9drg5hwebzOa7fJOL9x7dN
VgMw67j72dHNP+1b5wdajdnqkfAvr8pZnqJk0QS1l0n9cZqWPbqP10qO40ViMRemFyoo1voZxPpQ
CagYhHalvbstdYsQk64U9+I+jNVYZcwWUvl7xuM1MH0Bo2dJ4E+VzvQ0BJHNhTm6o2gtiAgoV5Wy
P8Y2kfz9+S+IIZbcaWbVvXGE5yUs7SWYBsT/H8QQZNotnCS/n1N0a2DDkVqG0xp6FT19XaJcn0pg
iK53EDcqLUPBM0VJl8CLX1jOrDD6b4LKQHICDu+GvivRj03FEG9DsrPlAXMuoQdGBK8kSefJ+2Rn
U8e8JkWg2ak5+IAz1D4n0lBUNUGn2yLO2M4GLyq+QQmT8ajWDgHjZo0SEpP2iZpZNhyAnc68rwGS
AJSar6+EEP/prh91wGFNUSv1ztJSMsXXjxSZDFaZKRhaaucGgQEsgcKA97vRmBeORBcW1dUeteAG
WzMJSizzYcOH7kttCZXq+V9ZQ7chcVFjj7dGr6/3895yTZDgxUnPX3lHuT1EfeCwNUzYWiVYCqwY
2MzfOth9Dv16NOzcxfZaG0FQGZY4w8oTba/1zPR571CtBB0uTnFz0haZ48FFGTu84tbOxZj77QBp
qWvUkW/Z4Yz00ImAVtJyVScNY4W0bH7JUF0KjBfZOBUJrw8Pr8TJTy+g/wou6mX9jtRQ1RfA5xC/
mxJXJdCWF+K5Skh0zro2wgs7crieYQvSdegv7UOoyve0fzbz/K/TdmCHdLCjQ11yAlqNYdThU3Gr
lt4tZRVpH/6jkBt3FbpXitgmP1fzcWcZSd9gl/Xd33qkw6Dzez5uMb+vf8UtKsP7k2MBJu/9Jjvw
iIyAmK5FcZA7kmfWJcZoRwY4f3a/pCgI2sr8rmQXY4wXiGVc0+aRhWhidg0IiAdo1wO+jzcQTH3m
9GpBbUX313Y4CapMRFH641xUbceGbj8NJIGj72gDFvqhWK/WrfNfcQ/x6EB7ga/ahuV/4QZJTd0c
vJyRYLVnCNJQcwz85xG2qtCKAJOILKz9HUSyTq5hH3Wij6I6oTSO/I+eDhI8PiOZomy0v3flY3bN
DU/GL22O0SEqXUdxj7YkN/6CWUSw6kzJI7BvcxObQftfVTd/iE4hM76NrWy1f7I9pdKtT9X5ASiH
gPmyIgrH5cN1P+hRTsGEHwJ2ZnaR5pVwGKXWQZpzBHqrgDtv/hMJFlVN7gLwRTrGdYmwvRtSv0r7
Oz6YFDmM2FABaNP1vWBf2lZOWm1cdMSQQehsMr8rvd2Rnyg6blRJ3Uizji56G6wqNJPuTdvdkf4d
PtQlNahod10w01UFu0UNEE7HX64fXWu3tni/N+Qd7g1YSqiTiTHGJL8EsNeBhCtJO8geTSRrX38p
YQssn0Bi9x9H9rZVwFhjSydNBzOiQaRGU478ngBaWb5ym4Jn0yLMAbAE78V47n8W9tH+NWom2HB6
QWnyihklU8AiRh1mcvd57BnVjFleEyEr62mc/6nFkS+62H2cJDp3YUkQCVBexVyLcAcHj8SKNcrV
e7OCq0NjOzk2cHeNoRawcJhYBX0Zep1kOU4Vk2mbTHgEie0LACVeMrM/MnyfRzpD+HYtpKp8eIhs
spiqVY6/NQl+/qIkSXD7v1yrgagULuR7Hm7ZjQ3XoPrq9mBpPx6RfMvmVGfcU/cNJqu9ok/rCuuy
46jVi6RBFuc/1z6RRiDZjDx9rm47JwB9UWbr09ahIxzZleFwIETbVOT5qCGaGCJ4Imol7ZA1VEZg
1ZgWcXLwBoqVwt6v6JNa/qI6uptuO0H2c0GuL2dhwze5u4cwhLGPaCPLOA7fzNwtC9liC26WdCni
ccaaw4ci7if+gGAv4Cq1A8midDDNTpH00llBRAlko5TPSzc5QzTNTzTJdcV9vLOb693XKy42t2RM
GQVZ1G9a5XefYWRoOoZi4z6cYiktCeO7HHGFp1GjpHJYS48bdj9YKx5tDTsyb2jNNfoguNZlThen
G1GluAthp1QNfjG7LI7KuBCi3GL1VgdY56gq7mtXICONow2MLD5xwHonyJObN4+YL/t/PuU5IoOe
DdyVUVvPkTMhUvUzq8y0s/ngjDXO5hY6/+ugFvZuh3UaEwe4EJ9D5i7d2DeqxaJWnyxaQfdeE3iU
bW4+gFKj2p2uYJc9YztMjE/qSc/ZSqmSYi2mSEyxgVGRHF7D/H2jLI8i6A+GIspT9zL9O8OVk78d
JAUwdcPKSsuSpzCb5F4h89razQaajhWKxD4gJtUaQcaRHUxyzQkS7JYNWeO7sIUk6QchZNfP3Gpy
vATyXBqDNj97/o+QGIIyatCz0lu6keWuyxY0MN/BKT1IddnYn8uWi4v6cAx62STAqbX5yQP5rUjp
T1Q+mR5HzKOHxG56s7MYQkAns4nu8GIlO7uUtYas/MdKTpMahTB8Nz7stzVkD/j4DaqJoopZ69xK
/SDm04fYlAGIyat5dcTDx4ox+1w+63yCkB0XVLT2J5anl4+LSdNBykfqjTtZ9Cjg1JSkyUFV4IWN
BPKOtqoIcdW81lnCPuVdSvdI8OQb5TX4xYZQGKuDvGEdTOeCJVkMUPXiW63pZCl+y6tOXNAob0+A
Nb3oKeDL9WjT1WwvcNNZQmGO31Nf5KJ82IcXRXsb/Xdnz929gokZ1fWUBn1iOtuFrkLpLyW4+GV9
Rd3j9oMi/G0c6AFmMgBy185HvD7itpUfnSj7f/2gZHjmH4o38WDbixcl3vAonmTHpoHGoREUdZd6
0mXxxqI1K2K0D5zOR19EcyMpsqJexd0fGte8YY4q5437LozazQ3kcND4bfSZ85IiIXgSSIYMwXW8
IvEUkfeE+869ZdhiWmdPalKuDWwk0tkTEhYHG9L9QYcXRt3jk82FqVVrZoaDMAgQDH7Yn2mjUOiJ
SxJmpApfw7UYM/F+VZXZLvkybI0ooffkkwPlVdkH8exOVJ9hhyxglFiQRdjZeXXg71c/GkgI33RH
3CcGV+DzmAJNEDt6+Sg+xfmTwZr7PxmIncf6q7DGQJvl7qhfQVRpGcSdQUgK72DytJ9Mik5tc5Hl
oOLx8aMnk0UApOpPNFnZC0ryRH9csCvfWHnwywROLKW3SLjkDwZwITJw8wEhx2Z0Cjrl3ONPdwfq
v4GULaTVL+pNTyVeJtcF9qrWouJ514ZF7yl0PBo4WwWwTGyGqJ3yYBobFL/IrLCx5VBiMdkPbo3k
wXe2E+Zihm13gMbiSXmkKpF48J+R7M0Xv92h/GyACOgsCWJjwFDIz58GWCd+vxh6/coZSJMrrTMq
HKSlQz2GMeqg8fSTtw/npykBa5IQegCzjdAEX8LK5YbXa+xbUlVD3BPBz2kRc5eqJwy+wtERmPnh
EpxufzEMaCyrKpzm22CC/ed2ilqaTPEQcFERV4SDyIwVAofHrcp7jZXQrqwGQ4veqeoyqdmcC8MD
FAWMdrfXaU9TuqoWexw0HXeDhK68Zx9mpgoC5O3aMTXH1wMx49rwyOOJEakFHpFNMGcV4h8O2SDu
/ZRKltVrK0wvC/TtF6naK356+fI3nwTEBJ4g+TVngywQcn2dmBsp1EDVklS5c1VdRP+TSeDhlxzA
XeI1ObLPjjAJtdh6GppJByXIb90Er3sbm/DMHdj8Css0rAAVPB4yOhfSBiH8ZEsOJXs0US2Nrui6
aDNg3fmMBP+T6U5b8aZDv3hYelYWtWZc8uVlOWsYakjWufQXyBC3+epB5PV0xNnQJbceMYrJqHNM
9Rgv/+XFkULKoCykdKHxIyshGbrHxHHQ/la6g1LEevY4DCjdhUw+jRU+CbSqB/XcvUfgZgq+v+Z5
kZzuDkwRHHfYZAQEPIgDDJfGp3jCNlNUE6YmpG1JFQfMlecYetxnIkOYs8UMcSuRRev+kQQ5AB4Y
TT8Y4S7Vqd0aLjH41uj2baToIGn2dXawVoIIL5OT4wY9fAaHSNX+sHuANSi98AVO00s2uZcgqahd
sPB3fMqALyAmH/NQIMh6ts9gbcrE/9HewJmYt9w2LSjXmA0Mi5qg8QRBGkUqow3LOuU1GK4OcB7C
ATuyE0GR7b3cMKNemMHlE9aNugeizA/UTW2Zbdza5SExqf0k419ToSX6JYuMNX1k4QA6qjfCPgzr
m2Bvb24R9x5en2e8UvNMavZMphw+Lx12Kk1h4OZkm3eeHvlCzqS3MZlhgN2CVpzcg2aKwyKuJXNn
hJsbHsUo5+Dxt/ehT6e9Zmbg6y6z9NbrmINLK3PnAOxJATzfzO2FK6Af8B8mU721SK9ht/tjMnPW
9x/WLwD1Vm5jqCCXGrJ/GXm5wdrB149xuWZtCv1b0sQwGd2izUqUamVdS4juB1zvdS2bChAXRzhA
nltzeDkPE8zXozaMrmfWXxgJ66uMtoVrLojxn+qee0poVJTjQOPm6KzLSN3u03vo30be1Q7lm1p3
D7kC+hj+xnGpKG6WbK99bgfNEqM5Hc3P6R05LscRY+jPWUT4ZoeMsWrPVQAUyWuZrymcER4d+7nL
t5M0xCbt3VIjSFTkmSjqrrx2bDA0De3By9o1kMbLAPPDZNqPcspB75BHRIgkKWJ01s4yCnZ1Onv5
iSQlWssgIGOsWgYpWgJFtbYLwWGbfLvdgt+PDlHnHv2IvsEp2La+7xaJER2g4kGeA0efBOckv3C5
ZkxWcBwQmS5M924UYx4InV+p6Wgy2TqTEeDjTN1AuG7uWrOOqlaF0oKnXI+m5mFm2FlGe3He3ayl
IiRdRkaTewte842oOESqCn9NRAjXL73FOhzhGHAq2heRV8OaDDDJlSwvuA8acUXgg/2t2TyLZJiY
891qAEPIoTQGrrNxnfQE39i9lND/gfu82Ea0S1smAyszUhoc9zZP4zrcRouS32RSS/3K6ddq3BVj
pMsci0LYheppPayGFRC59vUmXv72p8dLxiaJN/spMaYEQBDr5Oj0daxFPUYW78XGfGj77z8VbeG5
jFnSLc2eMldRNOxLxEH45YpFY8JxRQ+fEwP0n6wAP/+UEome3QfguThHXNG19aQA43F34zpYmz0D
NXWXd+28zzLEbc/sP0hFJTcDOoIxMKUcV3RYiFLE07bfP6V31f5tqu4Pv0+ST3ghR46PR0HYi2wF
1Hgz8/i5+Xm56aVMWQ3EA6P66oa6up0+vHx1nxIergX2oEhjFIU5z7+Fzwg/p8+07PkbmGZTs/uO
8vZhDCMjcA8YnEnkWhYg/vLxUAsKDWQ9SZnGAicnSJKwPxMXLxxT9pKz4TtgfWWdhmpmGWoxGYA5
GhKU3bAwh3lzshBj86MFTfM+HpwlcZDwjoMmbh0y2wrCI31O0EkvqPlS7HzHMruGnspNRym8GoBy
D5yHmrIN+GnDApSfLzDAT83Seo46JBp7AEmRWMcx6L+vZYkU7W7ZlGhiyZPS3EJ4XM4iAzY2/yIq
UEOQHxgxp49KiVgjohxm7rawxoFR7HOKo47D0MHiyI3W3istoEqo9m28Mx6wiXFkFnljNOYrsyO9
74dlao7HWsyPZM5AcDvaPJ34wp3D2+HnS4kyD63BVaLjdfTfJBMG4CJILAW6tPDOsYWPvlRkvEh7
PTR6qj4zFxGhspjWO3OKETrlVSZgN8x12rDa1wUugHUTjWbrpJNMasdhDAcVr9BOTHYL9WwOkMIt
iNUpUPBKHYiyBGmGJjleVrjXHm+NPvbDI8ZdnxldYB7hxfoMM6Qy5Oo15jWHu7UwZsNwQavV1Bv2
ZtHhh5mbi3ANMaducpW6ZGPK/lCJn1m1LYDyl3dunW1bA+kjKOxPD7GQ2qS77ONEVHF7XF4Z+Crx
owrIZgB9sbAFfRYIQP8GPgn6+agRXXrWCWdTr14LuxK6GYsg82Tt+QX/iN44xsuOYJyO24B3Adnh
IUEwxBkOolIphYAIxRRtUYbfhAHxXmBFGDsn0cmEvskgzvi4wtAqisn9qKJvsHdnrM6GqRv3bXUP
prLVgGv5VNdfY4yDkhwGBJ1swMJS/4Gvz++GpCkOMf4aEi2LAb4QGefqGzL4seUrXlNUBFAg55SX
UEoK1Od0shtauFMuDAWOUI/I3NKk+kLT5gETsW+jiwGVK7gmQWKSIo8A72QarvA74aBlBVXi/+ou
FMvI77BP7ZWin2gmOo/rAdzUdEm15EPs49Zc51eBD6W31P5Af0x5Nj3JxwTox6em4DW2/jx0cjoD
MpIjyiWMKOttiti0PYRyrcAcszIRh7D5nL2TiVbwPnoWFg6506zCqFLOJE3g9oh3Ws/ZRy2zgP/+
pzxp0cPmO32ZNNCl1QCE41JICGI7iCGsOFmItfHCpzikEk+aWnamTdTKXKlM1Kik6eJ7oafQ/94G
ftgw8HYJSlt9DoU4eu1OPkvVlqglFmd7SkUAbN6pgqA9osQwwjrl+T2HhpYV6B20wVUcKMuNxbi6
YSjT1Avs0E2cMBMOKN+uO5n7x5G26gEOBEQiBZbHtrdWCS1JaHhUCCF0V6snh3Uft+5jW25p6YDq
g/tfbMeNWgUMSmwAlurTFa2vt+Nk9UChqWsZ45KhL4yKT+sTlr3LN/6d1R5C3bKJzF5Ka+GjoGFK
2tLyHw27NqULU3kWkZBu/AFhclnj9sYlSSSAu1sKTe6xiRbQ3OSX/VHsJEq8+H61aS1EHk26qWDE
DCUuTzSFoV8KOOLlZGzg1AtdPjEzNpZeTjuAQiwkNBZPf4R0NaKJvCI8v82f9mhBts0voo4sRTmu
9G9uDDoLkEuOJbLLjmfWQaBT/bx4YuwWtYGKlTS0zhMxw9sRNiUfvUzWRmhYs/WF8qaFh2t/GPnS
E0IjKplEHmWq+BELCcRflVvT3LiiIjBlMfTVIVza8RsWeQqtID0++sIRG8WCF+o7aLC+Tnh1mWsy
wZiRlNbf9PWKcipUhqAhy1P/mDAoHuNTO91hA+Trtlbd2ep7hBY6Z7tn9MKZh+voZ12cjtO7Tig1
8JBA9eKDs/eIBbgLAnMqvuWY3DggzIkD0ohqJeniIopiF44L9HGfgsMAgIXTml+kqwJxdDEiS8gA
EDzD7Dqi+f4nPv+cjURyRCoVzXWSwuh0gN2AYDJ5JemRfuwm2lhkWWXq5PDpIJ9jUo38McIwKDaN
07wELKXD7cjo1Y1etGc7w9N/dVr275urxZtB42+yRylRehCW6S/1+5FDJRKjmePfii2QNd/XxeEl
cAIPP1XvoL7UmoERrJucTR16Sn+zM+Vko2H6sGCFFNLCa5fMb/8LXddN0zWZavjK1r2IRtmuSQKJ
2rwOQuKYTKX2iLiwHG6SXSN/zJ9bITH+fX9qZRCBKvTLLDY1yO+j8kqYV44BinuV3EuG2lwO9noq
CDbrNgs67PH79YAUCO9+aQS9dfThKBuKyQqxnaA44xJui67t5q4KE4nJtoIo/pAUbgXyu5yKd8/X
+47iWp3j5Op78+GNeXWEk35eLxAT91N0NOP3S7iGkbRnpy/dypUfG4KwF2NGEQ48kn/86owwp58K
bovLWlMWQTVlpQgCnrrevKeMbwoNVCtwY1IHBlJqLAuZ8uhonCCFffz8n5yht3CKaNgYue8Yuzga
ztapXQSlqX64kbanQlmVFpeNCtfDjlrW2mVk2vlYeHGTNFAqrnyc+SCZdf0NtQbgJ+mxeP8QwPUF
ebK87dhr7IRm0ZrNm1P0BvkPGO4abQdSAQtAp01/CkaUE4cYZ3ZO+1K9RMVXnk+Y0dl3YE3rjxnm
5A2fjwYJuYCgY5/3AhxSBZcRGgSUeErLtI3AJcxisnqupeyQzOWi/c0XvSMJNlzH+LVNQNbdbHwh
ZmnYb/akk9l2AA8UrsR5g7Q+bLBOTLaq9OOszt/sE3E8sE7E21a+wAFQNOfTPIvWooX+t0IG8JJg
JPHy4xA9jxqN5CRxZYZGMjylwiHokBf9mMsFnqdMC4ofSxbTwsjcAwC2+CSwUfcOnCzO3rtYU7cl
rduIz7Rzvdiq0uLYsf+cw/gjBBkun1942bTpGsVOWZHiQ8LWzWO3v0AjG00G2zxZrm300oKCNPF+
6YudMsBW/ru6KdEgUe6Ts8UTGU3dGQulDCON46DLgMbyJ9+AVhHRk/Qd8t+l4Elu2cJzz4J7ET02
wc1prhc5fJni4GhU1ujhYtJSguufqqYxOPd4m6rFPQNQb/GaYDsLvZ23iknwVYf4Qjr+1s0RWiBN
0Dmdc3y33Dzt98lFD1KkuDAjeS1fU1iSWHRFuFpzICPiCV0oQcAD40C/qUVyTmVCKDFxxNoj4tI/
QbMY6nlUnCvxfyf0Scvi7E5mc7TYqpWO66T8QI5hU9cZhQ6+l9xD1oFIIAFR+LvwNjlxuTMLJq7w
Yo0QKmkPUSb80ibKSFg8X5u0Ey//gC8RALzWdt28/crMN08qAWEkPpmmSkASFlbzJC7TYyyqPZWR
JhfBcvtnst2Cnn9m7PeMsg++mrrI2m7+SSqslZ9c7aK6YHr4RlNcsOqp0Z1d0PBI3gzs50fNakKs
F8gsMe18d59Ym9gVWCwH6VrrRBubqK509x4HxNyTZ787pP9XKYPnsDT/Cob+s6esm+DigZtoi1Kt
1zjJOc9LmOP98nFhwWV5hCFeabMuWTKTKaQi5qVSDXz539RRA3L+xKQ/cekLUF8FK8CSyTGy/C/f
vDb2rKz7Rhkp/LKo41TuWTglc8MyTJFYOr4oLzg3N7bcePEsnjshRMJo0uVDb2jb2oaT5h2G+1v5
G1xYebS9woBE51DEt5DVBYZP9aG8hrD6auDst6EGCjG0lLdxnTBNces2D95J9gZwCbm7VFZRHTkI
50uQBAKQz0mR/7p5NELC5GdtdSwhxG+9RsNP+MHEq7qonkuR/jlEJ/HlGeMVTiemNOXIDbdaZ8wX
EDGA9BVU/NWO+FklW5EuinjaYmQ7o2Q9dvRcEIW3qA5UDDm0cfH4OV8GF2X3H+sYweDIpFK3DAMY
PB67dofXqDrwnjKwHlkUCAW++FyuEHo5e9ZmV7H7H50Dt9hPou8E339baObR/mFYvL4WKvyTEV2F
m3N+2iYJqRzgAHoHI3lT5BzI37sOAJEuxcO/n0WHoxcoCr6ijKo60ZBM4vBd3NuvoewN0b8R9m2j
AcLPSwYnt92d+fe+S1lo4gDBcNxOXy3B9PUiXx06iZqPjvZVncMUgdbnH9ziyIxl/bEEbknbQBcY
hTxZJU/Cj8VAN7MlFC+r82a7Ov9s4T5mHbiW13rxCdPAzDD18PyHumVcXu8oNyjFoFhoUhbSk+78
VSX3PIgDA62WwADliXnP5Cs5l7qs2yI9zOcmHSkvZTBYe7i7t47Xu6dDyvOs4cffsXC9IbpMyKgn
Z7EGB3QEi2SdBfZ/CFjaBb8jlgUMo/QJ/eyUQ5hCxtsCi7Ben/KMN1P48cS/MKzoGVb/moupCKf0
F14tb6AR2kQ+Ovsi8qtGomxZBfDddG6zcoyTEhYMx8RbvdRHBAZ4lrnttBzFjgIXSLxaVQoZtjyw
Qesrl0qHFW3pDQZC8xYepOq4eBWnthAxVvECMYGrWJw6y/aBmbbfjKyMxUFHQOsAeRXqqwcCIyhh
F7jLiYJRAY3nYa44hd/A8sJEG/9eTlXP4vsyoJ2LpiAgeuVB5ryi5EaWOUFMJ/3PkXQFRrDrjDJD
Yc1mOeSxu2fAgnhf80I5W6mnGQDddhGDqrjiyYNiNykZ5PUq69KyFVayCziUTiTxR+zImBIO2N00
tzCmjUecFzia8aWXxiS9UO+3wjuHNiGTKk4WBLUKOFFp0oBYFPkyoog3VjB07+PL4taANdPy8VtR
oRlRJreaLW7xAzgNJnfkL8LlLbUHPlYZzv4cHQuAqKjHK/BLsFyiI8Pz80fP0G1xs+WwLGytwRbl
Ko3xw+g3YOsjGF2Xm0Ya0TpCMiU6h0x4Yrb6UAE83D8vOQH+VNGzUntSQTiP5iqwHEjSWcszVYVV
ZlhBny4v3Lz2M2RunHnqpPr7xl9NgMelBuLTGvvivcw98OQnGRXt1jtOLzTQWpPNEVifmKCaY9Kq
8/WatLpxPCemkmIykvF98zlXn2NO9jPzJimCkK7hNifw5tDIQza5OTWlSYcj9ESvK/bjPIH1E8Qv
ZyYj/QD+++5cqDw6YchOQCabzSEvklX1C7NFWcVJhuTk7Aa5F03Rns06aKwpMkObXzHd3Y9DS+8T
hR95NY0A0N9CnQ/nHktp1uwFgzk3/fE1KyY2n4VqXkosBZFU6Isfllq4wgqBsaSWYkmuxRYwXajW
wus1pbKDb/ICoI0eEdgnKOGRxQTcP6QdgehCeNATeqeNU6w5j5JaV75sYKepQHRdJOjzK2FeHRCX
dEtmL0YUDd1LSsAptRJKPf3azUCwP+nMIwBRRxKTtzI4+I/Y2VGTNLKp9vCwNlXoqslxuMNe/Q6M
7ESg3cHhGr9cC7e3cYLuYGPIRAoo/5RLawkmQxVFyxfrqkmT+r+iYNmCjP6ruuLDR/hWfPjkvVA8
zJBoDuuXVJRSIwOXVZaV7n7aLaytk5dfLPdatbC5CUCWQWTaE7t8FqX1nLTHcgSwW477gSIRcjVq
bMfxxE/OhGIHIe9jJbhjXoQ58e9gB5SR37ghK0JCHWm0zvmxY7qB9r5w6cEw10X7yzYukQn/lgTF
eMTiKmp72zW3OmEL3aTgURRPreFuMLoPBVKkwArOugmi/CVgsUNEiw8BgThIR62dogpXIa+rZLBL
lZjZxXYeUg3XZOb0FLnd4cV80uc2vM4feapez2zY131GGjd8wsShYoU3nxS0SlnAsrfP8G3k71dE
tRH5sByARdmCeJrytvmncQUFHGAAvjKY/SW4pUk6ln0yaTieeT94Fy1bnKGezhfRhURwDX9wJkm8
fB9kq6W0FnGCK0rZBcEk1yqpTLf7/OJL2O97UzM5taG9phqYFkuBfihSJZYgdIbB+NnRCCQftDNj
SkXQHKwBkwUxor++SAWccqA5IrvHeR0XI2SEdykYdKk64rjDxe1Sd99ONzePoGQ/X1kDb/khdfNU
SsU79DYIY6R/qS6Yw9CAkcnNqZRCnwUwzmOCiiedZBT0pds1oyHAjSeJAup53HN77wR1vMl/257+
df3CbtKpkPOQ4tXf+bvGz+d9Mfpfj4SpP+H4UYvaekhMIRN+h2u2M6pbvUlOoHXid1R3VehEIzfh
9hq9rqc+vKT/mVC4d1OSSi3oaSkfq7aSLCY7U66tB0uQV34K7oHuHVYI8rhe7jarG9xIhR2PKBjT
xzJIE2MsHVG32g4gOftGuJAM/wOT8l7K1FpNy3cFd6lVrqjlF4f/DdVXR6xDbG2rAccqPTSlAjD3
jm4fTmoJDDbL0CR7bcumofdn8swGTC66pTHnxHx+MsmiYrdvlnItwv2CHyC6nYMCA0HAP5Ry+Sgr
KT+Ic9zbtA4PRGhFA0qTJQSq/HC8KiFIvBKK8Nj3ko6tpsKcRM/uGXjN5MWPAGc9sjMHB1q+Azim
FNfa8y4XxZcxFcmzkXU/6GgGvRpIHaCG6yeEWjIaplJBO0x48OyhJWSM7htzUv5hPoE0pZj3ErFb
OhysiCGVEwlOqIBMjpqvNDdJe52b+0vZ3u24uwqVARMzHImufzVmnGk+9dbxdiP9IGuZCrHt1yIc
U/pVloA/dHK9RC1y7iDHdC7yfjM/XwzCRz7UlodPoyROvZuRiq/NJRUFcUFl05QQMrOPK8JvKcZM
tK4vSEvfoXIbNeOgr4+lCfjDOnY/Yhvq3hJu9WLG6vqFSEcJOX0//jIaJA2sanlq/pcBVhcnLNQF
KZ5QV/s0Wf/7l8GD0CNker1kAtBgEN+II806xt+xuEtJZqHBll/+LSbS3EYPJB3yGs6kNJ5AgNbC
5+E9sH3soM9INMLYAT83vDYFwSSFMC2Taa3XwHV9csNI5CfHA1lzBaErpWhY1qlOe3VXoSDxnrmC
a7UapWIAOUthbOX64RnZygdnsCe1LcFaEmgbrcsf1tXi94Ccva5/mmufsqijkhsYGJkWszTZawEt
GstYip2d8enS/SYO2l6na4s/d2/RLklEqemuwsaiOZSk4CgNfFWMevcH+84FGNW5j3zVJinw5N7y
1CFIMAlwC0r1BsR27ZCM4+6cERlgXyGrFDvcj2sZ9ksWQssLRnHaHvFm0H/EtaLpJFE6ZeSi2KH6
Nh02KJ+lX96w1X5PlOhg7imxCEin1K2cHR8dvEGrKiYCvbMcNIJO7oNHS5AgUZUaBJJKRWp+5e+z
mkS7pm5sj1iN+bFr0OvbvM7e4z5iYzTecJtnyMqu+hcmu2c0yenT2oVtnObuhMp4OAjPChiFOKw+
m9/O2f+MH3IAEoeRIhWmjNvUCJYKhtLjfvbrfHeRR1Zd1ECuZ1ggE7WGTq/Q0KQfBq5Lu/GI2ikx
kiwJQTO7vy0hPPN+n1pgaGLFAS53SRedOWOgsa7ZaHHI08fHTNoFC8j9PV9L6dFuqP4jkSsO5RTd
CqQCfFAAX9XmEVHSLml3Dc6gT8cQLIDLOXKN/uGoeiUtq1Bk3YOKS3Q8koFRdxfs8e+ajnnQCYv0
GJBeOK8w9PpfN58hPBm4O3aATagXH3OoboJFwNBII7bRbjJbTcnJCJXhuqNHhrGwAm9dE0aSex7p
23tGn5Vf3Dat6xttdwmwUAMOeiykNBSIXnAIWnVaxIDjE1TlCmC1OmkE87nFwVWcr4Z09bj/9KrY
43a/kSdeQx/xxkPJ6b4K87yG1tIZjnmA72oJ1+hSi1AhFMLXTa6Ik3SHmfVWU154PeQ9gcziNEcr
KYGJ5bByfkKpT+7OyXvAb0nVC0ncuckIQ67ukL1Nkp++p+vKe8RRTL2ogUIo7P5pBdRnRAfhUTzd
CGnC0fWsuDU14ou72u1iQ6Pae1ObSkJy8axhZwuCcuKrAfbUse82GCA+P4rTQMqItiwMzyVZ6Cwv
0D4/NtGkN21zbVSmOLeOqJUYUiKcLpS9r7sVXGGB/sCBvysvicV97subEQRAwvPleYI/eCVgSdtd
6k0IthjOPsEXfhey7DYfuO2hJtKi4W+SgBOwud14JL0wjavCe7F4oRPbV8GDSI3sSwA72wJTnbwJ
dgjrgOZH/lTchOsdXy0lnOw7hltRFVrl/RhsbdyTXc8qXM3hIte7fuZpa8b7Th/Qa/0GZJJ4nJ37
Ocizrdt7dygA6bsqmim0N4ZRpgbhi/iHi97cNQ8uhcWkUyff5tLHExu/GbGEGlOMD2UsGDGmN5Y4
ewJnr3Cvw+JpCLfsWFUkfv7Xb0amQW4VIT1z1Xg4TW9suR2h0LdQVVtbU/9hM4eLgXTrRqd/Ilmj
9s0XV8wwox6N7iliSrL81QtdfMhfxX3n8wt8CL/vhGW1g6AS9B0oG1jL0ViKM5kSM3ai9YwpJf0l
R8iCV3MRF82gMc4Np9aR54gmf7csswETgTdeME7uyfPpxhguM/OBL1OkuIiT6sxHcIod97wzqSl6
mAveDCprFQAuwtvVmtu8uAxKTFEgMi/tT3Sg5Tw3V9J/UcHgzBnYZqAINUHr2l0f7FttwKx+8NWE
Vpjo1gbBSbo0Ngdn5Y+U03o4RhxSJhSGuzRjsaX7Qog59qINlokb3I0BjJ/cVmkYuyyhC/c0J2oX
XsLukMVj0dfd5SCpISTEyqLgLembkf10WmfbIPR6DVh1gIrxejKboC7B+7iT7NaWvG/zKyZqdjuD
AdHN1g4QpsZU8kpr2/Xatdz/IP1LlPtwb7Mh47kNYAvaZ6AZP++WrF5gWM4l8TsZEjQY1AlVx1iK
P643mm6cN6p7U59eYpdWSojoXcYAEkci5jnSx554INmWI53O+unrfu5CbOI75pk/5oF7+mtoaLze
QRz3hhtgkafct+2ijV/vexx1xNrZq+NqgjvFCdlPx7MHSo1i+Jbuhe6IPCpL172rrv1n6R5UedfH
SvFfe3kGicUs68NyKeQmoibm+3QsOQmyAxqpcRQGXJc1fwOz8S7M1CZ+M39HSJFOY828Q4iLGcJn
b17qTOnZ4/VKsLes3WmsqkvMl84+Hr+teFOHi7IF3C35ZHMIdxv6eu8raOJk7z3+V95cV8ehV04R
VF2jqsXbxpMpR5C05h5fH7q2AKRl8tHt5fBME3ds3Y767tXaTZu0uxvGCL1Y4VNYVR0UboyGsOYL
3LshmPsKcWWK9ZfYpDv9uzOyRz22aD32YqABBW60Hkl4+CXY/5k1AEYd1lAAlRBLicGNpYtmnqC6
yG6jecBmJzrPBATjI6EmdqDna4DYD8L5j0Okq/MRFPcUIcZGX/yIOgj3y/soPdK4kLT32kl2Dw6e
n+SI3OMtqji2kqUPvtZIO4sRoNXOlrMIbokCSIsaU27EXB1Ji0svT9cjwAvsS98eTlfKkjyTuJGM
HQBuYypa1Sodyt0TOTXrAWZMMUUsqj4X786Isj7Oyozl2hjf5jirO/bGYeUjy4v0/UjPSteQmKbD
u39kNTAH2Ar7eLpwUw+7LOVcqNPiG+2nvQZP1AL1tLxLJA7PlLP6ks5E+0Y46J6NmPvqd0p/CM0/
421YI1PTUbCSIlHJzSREy+yrP7xP/YU4KofEplg/lP5KWI0YDDG45tY183hIHe3y2cdDHs78xtHF
kYS5wjY7uBKtx6fiNqN1qjSClnwKRmEpSDJ80ruUfA9JBJ7NFkO2e+0I5HwOw3Y7nZVvGlewEFI6
5SzYAiz/avhiFPwx+7nLAX7RPe4IdkDz8BhYHQLMlmihAL5iGhj5wnZSBdxuuxMao6EsDQl8xN/v
E3QTh1otP6Oxl381Ya1aJBRkbTS81lLDGsmcwTnA6pQHfyMn/vQCqTnrjmGbrbsx97g7IsAAno5P
H894V4iFIDzwca2ShALcKbJCQqRNkh7sNVMW9GaXNvhdgWkYbg2bMC74rZobiAG498a884Iy9nFw
IwNot3p10n1itsSElRl3G/qPf2lsyQCLrixfklVCrdgiYnfwgtrkndVs2QqsSdNuTBbhWlmVcJcs
X37q99cwg/DC8u1sSNI+eENMXWfEVzOks4G5zBjZ4hE+MS7ZjgayqhCxogOIzHeX810cVLnc+Jni
qvuCvkGkycqUg+HuC6lmGd+ApEAuyHqdQXeOn2M4y+uBps8o1F6RQ4qwg1fg5K/iSn2x8PaJsdDW
1pNV7QjwGhplRVBvomIf7MiWHFBDvhQ3EEG1mLwUn/RGFSr31QuIlmfnCnsGsURkxbjy/5Ftadm5
HxwQ/WM9lHJjGIa7EMpK9GG9TQ1huziz97+jUtT+Czw+9ULNANHHEi0wdJuK1bdcvJh9ue4nrt/O
zDOx4NXJppSb2VmYUs5xm8F0ts8E8zophBJSPF410r4jWyYYlQaIgJVww87mQQv8ecsT2B9gAsvG
PcysVGpuTZVXr9tXd/FgecJi/VPp7Hzzxye4OtUkQsRT2hvsA84oZ90EKGIVdGHFqfiXoEiNRvPM
tD9Hz1Baqc+gmu51HABDc/2Z1o365ooq2jDbGn0nK1vqrA9+HVxv1jH7urfOI13FahcF9AIoxghK
VaO84fjVOsKgjkLWfzYqAGNzp09k3rCpM7gKgPFg0THrhPvsNA+ciKfAKaN1QaGZ3PQDb2XFnEq7
wzHYHmZCbXXo7v9su8UI5uOeqIL+MJWqXXuRBNnoep+nX8XMLRMqg6Jq1ho7CkBsChSItYTlzpoN
x44BHgg7WGMp/vnYjVNUkk7Pcyykx4d38l5ObypzeB/koCNMV4UMDUw9JUfDvVbIID1ESz0ICK5r
yBAzV/RVTeR/Zcnkszq9yfqGSbDHTClIrR5d2l/YZmikMq88mWxcbFEQmCrPi104c6OmT+QRKe6p
4JO8eqKl3v+zhdDAUIIRnam7gGCzeegr8/GW8DKacA5GmCrVcc381BwfGAeewsFxC325LdpfdeGe
iApqP5uv3EdgcFGUAuHtm8NGFd9hEVxI/844zM8cXy73CongSQX3CvX/Y61ia6n8tTgWESiDTPnm
m/hFGGb2ypzSFgyHDqhP8Ob1o/IpQNBXLZU8Cr19K2qYi8UZ01bzAC2jaMQHNQPOqA4tF2EznA8y
nhl0Y6MsT2WtmHyYCkWCoMmZ7EEyqPhmrc5ot+m+t6QfdUVmlOr2Hy1YngFZcx2atmAxLmPyAjVp
qJW+bfCrVAo4JWbVih3ivzOAUUE8EDbM6HMJ7sF2wH2GEx1OQHbuAqASrakfPIfIIUg5hYR+EMj4
IcFis3ADTv9r0eFAzrXPQxqVGWtDAVcBNe7nxoTM+/m+Iiaau9sSTzPc0k/Vsf5PMuRds/D/l3zb
nSTeoC6T1fd0ZOKqMeDDP2hDGAivhFrIHn1JbXSfqxjzhoBvGBMWlw/Q59DcsCDc3++PtC7SE/Fz
0cr065Ph7PtOdVZbkrUY55PD8FCzLB6X9e5Kab/3ZFvgMM06c0nXwmIUoHW/fGZLYm4D+mEg5GqF
voDT9UzuO7iu8xiWsOkuQa2pIeFHy+aSf95u+MoYa4sIuRsjjLQxMuA1IePP065l74pZ53xEv097
yFLLPqmKwF97RM/q75FCCvN/TdFHrNpLKzmI4Fg2D+6DYCg5dNzD+UEYDMryi17dYknPEiSMMOW9
v449qaIZx+5m9aar8anKPuLENQKhBeOiuPoLt9hiRvr/OgV89d+TyEqyUN4b9+XwAj/wqC6G5fZL
p7F+KRHPEXPLLzOuP7s8+PIP/XSRDy3jx5fL15ZG3RljXuZ4i191TJ58TZVrF9GMH1AhiAWBmZ1c
zNW3WRbO4vkZoBjVRzwJyN2ybejzJ7x3uX85wuJeAdQgVp7NM5M8D8omSfO3sT+zQiJKrso6dA6E
j3LwRSQMgatKYRFA/DG7+wAeQiUaaxpUz1TtatwyQ+ciAEpvmmA8AqIxueyUy++v4q83yJqjJV/R
7qOgoe1PZOQaxyUyGis9pmyzYtVdTfLw/2XZ9xuV9avHz/wPgP+bLDRVMZcZSy4H1EqPHT54T0Js
WSaL/m336c9rjSRtK+WtjA20E7k73CYz9DrFl6ziXWwLmz33CiKfMe/7GuqeBEm1IFWXWe+oneL1
3e7jQYhk/Ax6b/TYh0BWvDienA7GMvfev/USmLWz2cQb34tL9+iln16+vAe3HscPQaAcSDBHa8PL
E33Cu+N1GLtVfizFI5071XA+vgUA5llp15xwWnggdvQ63X75HJUEZ5YK1JBeE/RD623r6Wnt87gi
TTcmbSZfzeHqBcO6FKU45fyDxmm4psVFH35nzKI58NPebj0CoKuShShWVlLo75wKksPxJRfFE2/q
ERwSZiNIqnWM1yDaEcLC5TPH552HYPb9V/IJSZ4v+1knODiD2mBBC5825QkyaSvdDcnKY0ky5Qwm
GAY1hNSXBgCnfYiPo4Swk4vo5xPKbrevF5EwQXBsL9iSoVqjWdhvTAf58Hr4VG/D2m19RBfjq4x3
zfi2Ta4dz/vSJVS2lRy4WZRemMIAOnjmk9Oaa3siyXlHjDsXQK5NOKjE/pGEH6DbhgAKxnsSzVJf
jo8WUielTjOyoe8STIFK+SHJR9W1GvOjs5qJvJpUtztrhOaT0n7uPN3lVx5PqywKW3crTRTS1lUN
r6lSBqmIMvAr+QE7vJpea/lC/55gizXB105kJj9aroUkEfYn+zXitUURkBU5T0D0NQaCcZ847wSD
QxKd/DF7Qqk+cuJSKm3jnUtOx0C8yXkwS0odXrnRifJ0eA9hdbumlHjFt6zhicmYPOwbNzlZ5Bdd
9VsSWsRkmqWlDkgsD6rWFQ0SKdfpYwU4i4lpuYOgd8cLHlrKDzA2zr3P5VXken2dOFwHrAf083zH
ZgLq+ymPepHn3Qhb2AVip7QipalsWgKbwLGmQF5wnVmYbxf78xM+fOjbQHLKrm0Ef21d6KUp9vP6
osNSsTz/jDrqN9b9GXGjr17QdvaFHIjlSV26SCXS5++FrrzM38n28Tnm8JgPNEZ7Qf/k4eULMXBW
+v+9/Wf/XUrH/Olaulg5CBnXDYXd32EwDxwvMXGrK6uqwsljQTkaQm8kkITU41i6FRdxoma7tya+
GrbCPucjd2TuXn7h8bBEz75Q7IAiBPbRbiRAOY2ATX8QNBMJk9eQBIQ2b8qKuUiOfMAgxcl//ra9
t0i0x4NRicKJ8+S4K4GjGnAcjCGe3pVoa611D/HZH5hfUCpQ5CDI/xF8uvsx3ZVQAB0pApX2GYDq
GlBlosFoSrlapeXXNLeaDuTstjEbQEPc/84C+xP7TAhmJfArlxMMqAN0TbR2lZgN6cAkMIo5N2ZC
/jDSwAzTk0YclV0W8Q3gXU+amDHeVSiLqZq9M5a/nyUlgSoRpIPBYQn1oz+ZYsQC4wVI3xWOUTO9
ZTnQY130TH/lKf5yjKSGXlb6+n3BWOXvVVzIQdin08+JXeOGvKGUE9boz0sbDddA53B+sLkwGiyk
wFfkMpIYeL/9WyZDkwOlMTobFMag+HdGAbt9BLYDO95scVrVHFc5+u4UHmzVgFq2Sey8fJ61uXXM
vz4P4RDoMzsIukSgs6H+hrwVJCENfV0DD2gHxyttj+RjkL/YhtUdzurnAwALyUbeCVJhqw5bhP+S
SN299eVwEdrQx9i4rnf5oN6XKpk3KEhO5nO1vD4ZJNP/Hl+pJf6Jj31D9KJDyYkwVThOqznpMYMv
c8yIhL1BTcMMGcFnPINuO2Irippb7MuiOo//5LpF1mEmeuqGg5lf5s2T9nfR2P50A8RXyaxGgCv5
X3QuBtBDGEg3tK9lilcYpM4CB/sha2E9/h8gsffhF9F8f3JTZX/Z98b6gJwolo6B4Ubq2e6EHgKi
L8fbfJZ0YaYoeITBokBIYCtorDM3YkZObiBa2IxXqy7eGDBhwUJgFBXlS3YPGAh/8HImpTu2uyfx
z1YXyJD/yLZ+sTA1bkfk0X8zX32ij3oy+U94MOH+SvDMp6MaMO2o24XTpAYDQVa9ej7MwJY7U4WZ
awBf3I1iQLUBEJLj5MnOzgOkO3QOsF1CR1ALvbVeaWeDKFAsx1kboicqGx6xzmcVexLaK5oimruo
29AhLAP0unKyQYEDlDvuThX5Fs8Q/HE1c2WJmr+YnEKcgpVRs5l6NuaZJk6Gz35FaSH6cxHO4WNT
zPSYAnUTef/3rTrEHoe+Hwr5p+mzCBlczskgLjgZIQvifyRM3TTeMynKqU77lpRuyoaXcYP5F1cw
/JRoW5bXqK7gEe1DWWtQXmJ9r5Qw84+6AFfXrSkBjsn5vVHN+CIuM666XDPIHIZGtMeqDh1JtCBj
ZwEYq3xbOxBo1S2S9litIoYdTZz3ukkCosYsJiL0CDNz9rKoRuKawApxo6wdFW6DIf5JlKBDS1X9
S0Mx8cuNCWuZqRSGKWbJBNDeSsXe3CLZGv9VZ9ojwYTdu6Vv9PyLaepr189TxnKoEYGFQYJbIMrl
ryXFZGsFm+QWWCE3Us9/VZzL72Dcqj9ecA9vuxL1FS7goJiCIX1ABt5CkCfQ6BiYgBJmZplSw5Ek
aaqgZraHo8qeZSCEMcm2aR0oQwha1vlV95kOUVZvl3TtAeJ0t3cQkcQneRSu7ZSNPOaPDWSrRdmR
QeXK5wq11u49hedPcMTbnRezNjdLWyHiyrj9CmBN4QfXy6tv9k50uDuFlf7H8Ne3zAeuS9jxKKXr
xwmlkfRckkTuEV0+DHcCTab+gN5hnueKZiwYmoIHWQ3qcLJcv+mhDWaW4JBNRdxV7ePzEoz1HUIf
7kHCtq35G0VGSCGBCZR+ik0uXNiJ5oKEalsfnWCSV4F4qPdRIYJdQDNJnDUKQR58bvzw1ykC2TcP
HX+r0vtXUpGj/z2/hiwcahoEdzHoYdUOcRMkKmsdPYDp4Q6XCyNbqG3hR0O9XfAGqwU8Xe6G8AX9
/B+JHWC0yTodzM3IZbCLc2QWVKkFb/X6GVVOsZY6LTzSM1gvXFJhK+nD8zmzrAWJp9+J85A5NxnF
JIyQ30N+eJmDV4q8mznYs/pkoaVo3aN0EkN/sTsKeIou/MKMJGy0jbdj4DpFkyatiyzKHK/zZzqH
U9qajQNr2Gq0/EC39SPwviqZcX1lMeJp1AQuQ9GSo96GPXHtGtiiBHozBFmukHxFFUr99VGYqfDf
AcOIIg11pB9sy5yai+6tUMQ254kgDqhaGdOKzj8f2PqgG9ZMivqH2nW7RK82SaKvJgMPWyh3KPGU
LXkQI4V6/vZQsqPa1PLu0NY4JnjxuQGPxrv/1EzzjfQY/5mnafeiGautXkHTRqTT8w9hIsazEe3Y
6YH02t6W6eklYDFZ+JJmyZCj33l21zbgN7ItR0bxWZGKFYwsBUF0z585nDA1QnmxgpbJ9/62/A20
pKA6YzqalfpWx2N6g5E0tuVGBRjfO8vKhdvbLuSX3DbSwyJIn0p2qGY3l0woo1U6ZX+fC6co0O3r
fgFTlXCnwiUY0VUPGs2JUhtfneYn63QvYsDFsplcb1Ut2djCN/Kt5GLR8kfKYp0652ipYjXVK1Gv
uYCWPuIjW17l6HYNrbrmTaiL2joCMr8cPZhT1NjaskV5Ejl6yaQFJ2WVVgR4YFrLVlxVQMU/+YIP
4mp+c36vXVmZOt3zbTUfosBxl2EjyeyPxMblYL7SuePqfgSSeAXJ5vaLLSUgECFyg4UY7fEza1y+
BJiG8GJnd8EBisB4lpFNWmI7zpmd+JjpBj8NI3xmkaBSlkfQhXIkA34lH8411jYKVAlubHDOGoo+
zuY5lkWoP9QsEpAtlBb8KPIOtP/JyWgv6EK3knvP+7qjSLvzXJKglT5zZHx/5YOwFd2rQI5R5b3q
vR1zg2+bl3sTFHxWmtpwadKuGmXrQT325jOPwyk5cexObyn/lFZSPUCxHDIL/nAmvhoW/ptrYCP1
KcLGGTNff9R5yDorsSManBkay5zScOJMr6dtUOuB5tuefiTE0D6qprZ02gk0E0vaEg6iORmPHn/l
+K/J7yDwxmPkKvDB5A8bjj1uGPFqPs8V6f6U2jaUwEPKZVnWtb6hf+YHSefi93+KYk4GOtDK0KJe
Yo5JqhhrVnBkONXkV5RHpeVBJcDIu/myZIW1Q4wqxZD2XkCp0Uje2Fkw7snjraRepJUvuN80tprW
H1IL32XARxJk3p3inbOqY44/rUIT6NWwxmMtqk73hfUvCVz1n/CEBQ+Vtqs0Xyts2Dha2yBTIXFY
CmEcaTnvcjbI1dDwS4OamarmkSQ7Ly+TR0globb/KwV1ukj2fI+WQ/yVHCe5YhPNEioroysHB/0V
f7ljk3sVVIeLHa9dc42j76kBXuGVUvnNueSYhomvor/dq+kgwNQsdkHfM5wUZN0eiNGGFnhiW7kX
RMLssONe3OzuNW3Nscu8r3e2EayMN/Yk3l+C48CkY9D1L5ChzRC7LUxPC0xWDyI+lT3mzAokZsBV
RzaWupxvNgclkvSQ+27Hacz8uuVROhRW7R1ukyHeXlahqMCmLcZH/NtBrzyL/X+ZS+279LDwzibY
AjOL2Pvuk3rynmLn4COD2IXRDAWue8+opmK8MPkrzVKjW/pughzsJp4R+lz7TzkLYhm+vVhde4dE
nAl6d0i73jjVWFk0FJLgaUzTR/IVRDry3H35EOVWXXF6eo3RMNjItWk/YAHXaQZUNLftjngw6Wpj
bUhZYIQ3r+l+/5kUWXWOWMw3lXNt7apxHndpDAYGfEl6v73uS0vdK2rdGDp0qD8/ecu+k6GAIgHI
8HxqRNZjtFeIGWb39hx/6qsu6S92dmB5Ip67jXvhXx1Y9nLYuwPSx3/vFOfE+l8N47Uxdc5g9OST
o5yvurJ48MpMZdTtY/TFxAcpKlSv8SjQBXeVlAKIKwcjvP4aCe/7atmLbOjmA0eb/WGL/rKR5EVM
w554u6ONoD9gib+ZRuyeiYpq+KZNywojiIy0MnTfz/SHU4SdLUou/EsAxyi7WXQF0yqSaQUh+y94
h/DPakVaPPrh3jfugyato67x6vnwjntxs+6TWdANu13USmKXmXBXnAj0FprZgBHd8/MpdItJf2NB
YTMcSjjzJZeCbwUJvsZ57/yqzztTGrhSbG+iIvxKhE61nC7qUxbHxZzMCyiCP5EWkdKUFIr/yhPB
M2KDYI9F3MP/21XnxCOlKxpkmzraW1A9WgSYoF7uDasrr7VmKRvwGKlNFeeD0KFRtAE0fejivrCI
+y/fd/JXMDRdRvstX8sdC5B2OOVhGlPwkHlGcp7zEz8E1509exI1JNylzNBxHnWBJ4xiSxXhP/eF
/S7KpjJJOvceowBkoNKptgsqz6VkmuVxQ07ZM3biIUtjl4a+7qwCMbN97LdwRXKZLtQ5KTOk+nF7
CnTGwurB+nsXBRkedQmjOs9MJ7340qRaTrWdiO/14WI6+UQ1XTcR9IxjRNYfwRThVEWZb8g/h3dd
irooaGLuqqkqV0SvVPUK714nMU9yZv65s8NPhtQBmDo56L2w2FK/jFfWEe8J8oMAcV/y7yp40J2O
VapV4OS3H6S6JXPmKdFaHM0hmAizwrwQam9AWmiEORalQjeT1O67Ggux1i+vkug8qNuYlbMifH/2
TDUQ6L/l0Nabhm5esp5Sfi3nQi7nGnRfq9L0i+h25kLtQxYSSGwLt0qJvuJwehezincsG/LRTO4d
WizWScen3oaAzNG8/xVEwFIKnC15Ic7C3f9JJpthydKie9biJi5cW0QPjoeySnGRejv87hXGkOhe
JG547SLxbS2lqH85GdqAoM1E5aPip+lwToHmXl9lx2ZFbdQlIdcK6VTSZ4RuA2wFWrr+ewwDzCmR
Qwzc6+CC0nl87v7aNl/dXTGW3bMdU/yntdjogdySRH/MWdexa4TGKJfJeo6G+ejy9O5Cxl3NFDOT
+gUjAJ+Ah5pMEsp4fLo/jfUXBGUsev2R/Q2JMS2WJZ/QWh0LuS+oaozt3whrzrYVNmzyfsH7zTHC
Wozj9fSIVT1+woSSbGg9SRGoCNsdqhOxKrYNrFVghrlMMS8zoNb0SnPCRmrnUYkxBWgUjwAWQ0ET
2k+f6okzJCH6rGL9A6T306whtLo0umz953g7rxEWydmOZMvLQnF1giUZCBHUXlop2aEPjfNGphsC
+skjvySQPlOpYI5NAtKCgMFZtgtHDMyCGAeGU6SX6+qc2DWubmkAJWhkkm4DG7cWsHnzDlBF2cS2
jmQrbROS8QU65TQ9B9vAn2lW1M2yVgZ80CmAb/wsBUfENObINuTsGfnFwKigGP2mVNGapamFYtO0
vPFxWUzZWErMeUwRHqzZc2u4VwlyQzqpJzscMNTJ7U0RJMADX03Y+3Zpfrv9GEFO1sNnqHOKfyAa
dqUFFyM9mCjkm1FI329bsSwYAeySW4X62wFKzcBjJ7VrAzNrytwlGgoqc2Vm8cADc9XqW3qYpoQw
0QViRPJaMO7PNpPOffQet9hOj5/JNHVzKGc3rw+HGwk+H6riPvrk9+Ve3qSDJdBw+NXXAa6gEp9k
9JKNW5cITzJ7jq9eLGCgy1ebq3G3dnVdoTYEUgqfSpSDgkBvzaVax99QcYIdqVmfmKkF6Kc9KhtD
jhaDxg1kalFEL2vX2gHVmw5dOa1DaIcJcRYkrqd241S4rlANav2GJAe0F/EKsVxYIc8ce09ZPuaP
zkjUFWBZ+tdvRbjyo0YnoXQWGhz/gGmnKrtYhmdj/S6t4JQpKhuguZRwKkirc743yHhkXO7o4lpf
Hnqy+B+RH3AnQQqsy3RP7Wj+2CORhtFVh1lFVHYwePmlK0/O/sl6RAWnbnIO47vJGWQWcnThSLjm
oVVgJPvifbzz14sTHMlcLXlqlDH6j/Tkmk4IOzc6nSa1B09DO5ENeYIB3mMG//ugKaK8L4BpYicL
0G5n82NWvWq0adieVJanzqWBaYqYh4zMSBtyryyhkkJ7a7nKJCH4PmFeTF1lBj7Ixs6yT1K0blN9
WkZ7D007psLw4OJ59UYsaCTlnXWyf6Tlgtztc4yqvUoOwX6XLRIn9cQ69OvmuecWgTI+8SieRr2j
tucVST+QTku9EQnvgoCL/9b5x1gMNI4O4pTobBmxp61RYsygFTC+3gGyYTHn4erchWim7w1/6I9V
XfcbFivNTYyLVWcgN1+UL7Qm7wQVphhUtqdXXy17GfG6b+af4RYSMrt/5LJJN2bPuFQ+OxAChtks
o0BAVvVJ6p2JFUnmfQUpQDhPakb5KrT1olFfMkqRGTqm6nTFFkMUG3VzfXN1qdQufT/dZL3u1xRF
oQShVRI/8jR4aY6/9QvsyWW7P2wP939k4IYcW/kINtwjEU5yEMsjjyQrIDhFrcsS9cOaOZoUOXm7
1CMe2r8A3fk3fk4ts/emuMHz8zODhZpBYs7ax7Tvsigw8bRT2+nDF48QCzOAW+ZebhUgvJRmvEnC
BCw2yK7MdqzACFAEZM3BYaGUcKsC0wwMK2gSXHgXPxvtXn2EHViiBxUKldiS/DJXxESuhgWWN9J1
50QqgVkL4EK4+Fn0I2xeKiUok3VPz4V4Ka/4YvMW3NgQuVLrZAQyscROmWO7fL4jy+ll+Su8RJ5O
YzxERVn3/W/gCsg8MJHVbWeakT5ol21/Mj98bWqpxIl7n2JZrxiUuMQK6xzjOccUsaGVnpg+IOyz
m7ZrGn5Y4pcAHF3JQOq8jhOjksWEVjru+zEYTJvAUSKbVDhRt7lOpYfbuHe8mHn5+TouYQ/rJVYH
FVvkn6GJ8NZBjeBOomclN4ikYc8cml0GN6mZgKTxFSvrDHw6OZI48PVmE6EvKfpmYTasFqhTqXaQ
eG28u5q/RK0OiS13QxK8U0a+Z1bHskwDPxCQnLjTsceLfvjGN59Mtxgx+tzvLqbUWJO/oKy8lL2g
a/nOqxRcKezq1vHwAzErrmRY+4rI/eLqCeZTKN/tIAdT5l4YCpB4C1T2JKh1Lbs6/D6t/u8Y1Jj5
rLBsWixORU/lD+ss36Mz2A+CKWJgULkpsyXL4xMlP+khmxlL4czGCUzHXtfgkugRODGyMiMG/s4t
g4YOC8kcOhGCCsqIQHAEl7ItF34j+eGSyNwknPmliYVxT58emz26Jh3GJhBHGFmzOXMk1BJEN78G
1+ervRbgMSnnLB+6oF2+TteNQZBxReTYbnFZDG6lr8iOJgLdf4a9Sk7uGnr14mLsgpH5fN6NkUw/
WAEjVPjyoVBSfrvI4yZOChLimt1lZ47I78MmEdAerNIj++sglTq8ha16RHjctdrdhi5njKvRj3om
kon3M021qTqm3j/1GLUcz+XqzdzY4DXeM5yggXqED250coxu3+P1qubtEl6c3EQA6o5rMIkHXWeH
wu3EpE+zPw8Gm3BF826hp5eopckT+s5KQOiV40SeXLPa7h+IMSWxExKa57dEkiMaeym/VNJ1MArd
dH7IKSEY3mlG0FZsVutihWb5eS08fBQ1A3MgKTwhbnxoU2lxCmHCshUoRgyv+K1alIl9NcmhRQ/Q
DUcEmmXhVRvw+dHjbsrbn7dODr+z1fDqZnXTZhflIOXqHnvitUzj39pww6ijY84wxroqHk1aDvU1
4CHHXlUUNju/Eaty+bMKsitNB/zMeoNxCIjbfLidznfWwnel4sX40rtEb/UTstiKlv51xqHOVK5k
QfKkn73fYy7d+dNrnHuAtw5DB8cbwQqC//FAG1dyIMEu+ZU77x0K2X+5J5zJrkUFewi02Lh1sXF7
ePN0ZVk0lRnC+u5Ai1II3zL6NwQQl8mA4SkbxYsi2WqEo/0K4fvGFxRnqvHPyrPsPWjMGPdhCrCK
i5Ud8E27/DKCLOAxpteytuC9h+dmoUJQ6NfL+GeJQqi6V/pMroZMaIkX5Hp95tgNLMjv+A1tHPWa
n3iYupLITn639FSTpAqPRrZvKhIEgdwkSPJGDVr7rFlPzdHR1xleoHjdl5CYv7Rq7UbNTDKunjPO
i1+/DWDsEWLCAZ06tg4uuSqJ5cguAybr0QU5Im3mtc0m9Sd6hc6/G8/t5llNxNwf6D1CBnIzeHd4
tNSBADp3N+Oror8KzCXyJKTTlPu3giOQh3qhzBYIE0tPB5XbM1AkDOyqbV5Oouh20CQc7OnII+t6
9jxtxuJj0ShwGx+ekiEnaP4uezmDNBTEocb7xXemSBuQTmV8BdgEZY5rFcSxg3B9TTPriqwe8fGa
7VnQmtMOxINvFqPAL0GtKqFEbdIizGSdnSDzUJw0Vl8WYMZBV56iW4iBfxYmZi+G3klK067HiNQk
ydgDS1V6oq5c4kw7/u1nOYC/rtAx/osRQLN7oXDADTuU1yZJ5UMZDnAdNVSblHAfYGst1K0it3aR
asZsm1vvw1AacGuDVxOxt9bB7VdATC5dffPbR+y8w8a8nfzFpvLCE+mnSDTatMdcaMC5hmBSoAl3
MSJ7icOwGwAMZw9qVkROA4gXu53cOHE/2HKQCoWRJM4YDyNoxbUJ1kNbe0Rpto37FAQ6foXx9Lui
nF68vkZVMs13mDz4imEhVK1ueEX9+jqyONgxTiMPFMFCP+nXdPXMbPbYucd3sH9JGpPIdCjujXjo
j9sEeNVzFs9SpbahVMqf7PZVqlWUQWg2gPRPisOG5q7S2TqbKUFoXMCwk8mOnNZ0GXcaqbR7iXrv
WqxST7Y/1Hrhnpn51OdbqG2LLFem7Y6QvzXkIMkmYDf5tcxMyYWvZ579/Ew1pYMVJ4ChdWzYiN2I
T6BfYdFfz0N2dMDCvig7whpYgd8nGt87CZDvKOVNU8ORGXhuZtb6t1n0ZxELvfmmmrPUBz6TRJYL
Q4fNmiL794P3L9FeK9NRINjBJMSkzrvcbUNrCtvW7SS9sLLnhF513EZlDQJ1EqgKjcbBwtPIh5lX
Ei4ow2XjC8vdkca6v8NTTQyIQ6QOgJldRvINgroNN09AhvHeiOJEN6s+kOmQmNYS96WPetjwLjBZ
/UxYbGKPCZCfSZ8juamyh+fHfQfHTbfUrLfTpkcHIi/tlGBR9LNAENTD3GJeLpuXnDc7nV3UNvT9
NzZUuKHVvm+4OJzQMLnrHkAu4HnHDR+D9i1ipkZlPTASvfX3+nCqHaG5ve5fQzWM/HWZyjc2YXAH
hl9fbM5eppRDQpvcdzJg6CIWYRAHE7TophgOFn6a6eSM6mC+vvi+0i2b8kmAKJod5gdFporDOtQG
yiD1eeGm5+4XxX8HYtYMg9HduC/O3F6IiWKMpt93iwPFumL/1hiKy9PLjnvRgBN8XCYR2iXalZ/i
V1hoFWzSY7uIrl8F61epGJhI03BlDHIOoWvNstp5fYI7AryTuTy/YtsDqtUZPCWH03dswSWZ4CYC
QOFcfr8cSYhPZGPAuzVdTMLjXLMpA1rfxgHc88GriWwzQuhzmuu28WxxlXECiQvu0aJse56Zvwu9
kxNlz0IIXbYx+S08Uf0UcoRNvxtKQyYZj5NdBCSyWXFCqR9O3jHFcZp02nKjVBn+tkSX7qJIbS8w
6QtN/uSVHDUHgAne8xIC/iPQ4Ph1RRTnhIdeMiiHkD4rQ4gDzeYBcv+VbRD/yhKQsUSiPyT9w8zq
4E5XMzLSLAejD/f7rWKt4pc/YxgolK3riP3bsUw/8XIZnWtvfDSq9RCoCCFWTuSB0zXzuZdM54eg
i5aqpOs2AF8FluswXsefbDPM8eBKplrUgdgwMNqBhJ5UNdpfVYpjnKix1NT9kQvqBtGOU7MtU/E5
mSOQXuzga+Mw+tCU5rqIRlwMPxA/zrtho0FfrXdoGtRu0fMuqMNdhPguePgmNQF3uLb2nUDrCurX
lFz0A0EKX3wq7ktd0FVbZu2fAr4axHsisGYa2nTMbPJu8hy88tBS/mgYi2M1S08Y5QcqnSbvhVoL
5hpGFRX4Rmicwp49CXuYuob5nlefWd+UoZMUFptjGLDsK4fh4CVf2OQVGYN5TdaOOtKdAx2o45m1
EPxtF8/ClxqRZu/tNoc540VCKnJP020oz26Dri9uCgFy0FZrJCTRHsBkrjPNrrKRESw7IOedQPPJ
W9McW6xMctRPNpVJU00gedJsZf8AYjJz2cq20dKPFN0prRbuM9rE9yHlBUNnSdZ6MdVIFQFRefxw
2vd3NSQJeiGkNUbp+bIvMBLYHxuZlKvpawqDTQFz9uBB2P9r6b3KJFmSRDyUfQ0QnaLtMc6j78B8
Rowo022EwJJjrP6UZFgANmOqPQbE55DaR2vGC5fjQmiPFf/COrT0eORDFn6lS/Xp9N0qh6T1vMFv
Tc4lANKiq3p1zYfQPLPelDZ13cdW09kIGBt2ETAkomCQoN7TcvWstt/pAFFGdfqOgTqaRi3gdNx4
pM1OSdYlVhZVoU3FE2rjdRjABoQnjpAEF00oDwg/HMTOEfqDgkPeKC9gnMXy5WKgVphnjurUSqA4
pFeziMcLq2BEC83A5CW7N10MVPe6uGPadtyeKEkSP478uR6YqM/tU4f4OurIKMYb4fj3wyGLA9wm
ODztvAW2wY9qWFG8J4ZBzDJd4G5b1+lKwtbNHdK+OZJ0RLYcy5+nAIdNos7oE/K0yaD9afs2VAzt
ikxJhffqXzHIICqdO66LnVAprQ1IMCd2+X8pCOX6U5k+OhWmmn/WkmekRQ51TBakCzPUfWomFm/h
mC69llIeXJEtFsjrJheftbNefkNQVz+SG8DzSX876UZrNFAzcmf2TxzK1XDQF/WoVQ4wy89+EEnF
7m6UyQExG5OTbj9gEbpCkjahH3MtuiC/vnMfgZho6pIsLMCVWDb/SloJaLm4Zpz77e/C5WvNQm/F
ObEnHbd2GJIMsw98VvK3XLvSxDucaK+Jj3S7jH+P+487zmCPh9nrvrKRfwA8fOHBaUuvpIIW8wSx
TWGYJ/MOLx57HrxTBkwrY1zSmN2iK8Dm2K1V38ittNUxBpLltSPx4KlZYIZtZu4XIfWmCNe52eHW
+TGXx6pLkY0/NL6HX/Et304Zh+Vr+9LpFV3lIF0L/e4CeZnWA/EnH2RroZYRokcaNeqd9fLQ4FLM
MsoAPKX0jajRMxyDa1SQAGojZ3RvkQSWgh0oIOj+kceQVPvOegqgTOdlHWoC0MXDMYrvlg+BsCfM
FiLVJs1x5Fjl8sVzgT76FGclmBvsVtrQiezB1TLfPKI1HBvsysA5B10BS7FkxLq2c6NWm+F2eLxe
h/WIjoajgY82ix6zkr3Gq39vOBtV0nPFLjAkWAxwMislkWeCyU8LF8pLu0JWsYozXaRkFH6oJ1qU
yPtt0soK//W5CAuDu/s/PSgISDwFilVC5jQzQuxT+7xQyT64CuwQ0VtyZoa9YawTLUGpHG99zmbb
6XqR5nsyNpFNOrLVQUNSoMGOM62v7vzdyMb/V1JRKL2vOhJSWzkekWIpggBq4ctPESO+YcF9bGLu
v7AuSjXSDhf3z8ZKd6bSdwrl4KTNfzRCbYZn2qb1zVKb91JRB65YEj6aOeOrTb0yy0BVAcWH8hJQ
wxhFEKb/x8g+D+WBbNwxaQ9VV3o1cYUfcFBm9Ijn/OwUtn15469sd8tyxSGIQB61oD8R6xvPrhgc
478rimdITjP6E/xxFcrzRyN7I83uxNkCTgkQzbE1o3MXM8xGsX5HAGN5i4CJy3gGDqJ7B8XXbxoP
r6FRFzLEJeTrtIsHIw9WK1qyPconFC32TRgnGan8UTNqykSqwtSzYlwpQ82zJCxT2rklP6MVFC8n
568YyIVARPBxMZ5Yt1CXf9fPcs4XegfOYlUnxSOgYq8aqZ9Uo4fjDNFBBNJ5ID710ruXph/UVbg2
MXSCaewRj6C/N0385btin66KNM/ujgW4GHsTj2b0RdSeLDG4Kdm8f2NHg7RE3OenxKhAInBkNZB/
O0AcCU5MeYCz1sRXSy3t2H4wfrfcFd4MStwhesw6blCQzOwjG+qRLBMvqpiiPjdTSHMkIpHQv7iY
Fbn5DtAVd8J0+tAXxTN8Cz/zx5hXTaFfhkN9vX1+G/RwvwIDC/ItMoe/9dC3eWNTpnkOcpQikari
aYZCTUu1ww11/4chWBFUoPWpmRUWpEpZNtYNoywvaVYayRg4+8nADMtIYEXmGTYTNlFUwwXMJ0UQ
Qnf8gzm2dGt6ccVG1QfMs/mAiwUfZCDee9s5bUbCoN0fr1Q4Zkt7AzxqowCySGk5KQzq3AM6Cb7A
AC0IW4f7stsbrTQC6xzR/PCgtAtDVDn2AQ+lDyH/hEj057dld+ROO3n7YXKmOCsS37NVJbOtlZYl
Dd7XaPkXxfO36/WlJQ7LuHPt4/ivrztI6jlh71/Z2ExbnKePitoE0Xjrr8XFSLBwLpMcFGVQAwEf
8pPEOg9RD8pv5lVGBwqNCDuOZNcfZp4EMfGdorJ1HTLPEkoqVB1zhrWMLR4CIkXGwlqqUuaVz9zv
7PgXLQkNkl5mUTN4CXN3Hf1Aep1q5UTmc4LETOIsWJu189SrZMHadfqzyBkO+TPMcHgPuyiZe4/6
amIIBHpIu8lm0mbs8s1Y1HO1x4qEWhRKC6DwweGqRzlanRaGpznBC71SL0VqZxOJZlT76ITJD0t+
WliOygTB6h0hZRblR15WuDetTVUdgiB5tCXvVri7zV57PlWv7eQIOB535VASahqLlakJrLjbZXlo
yVlqlz+lH20qcRnLTONkm4orlxH18VkVrMeGEyPSCj9OXJcz/XWrPLxShMl5QuXtYQ+EpEwbyDYQ
CJbJ0UUkUZN/PwYbzj4BulGThyGD72kGNK7jKDTYUPiICEmkFq3NZEtoQIQvh0Jy2zapON8bFO0U
0Ic+Lo7blGyO+B2d76aDhdD/6enXkl52qKTwVb0l3JSMz9mYgXysuddL310yJvJZ0hAFAb/qbXBX
vMAfImpcEMVIlIY5NR5nfCi0r0FGtyRFhDahor5hsUhMfspVEt9Eg0qR/wjIohmWdDhMq/rqYNBa
gPMPFdFWOGRNZ3zxe2cePXp7AxR2+lhbfmXrTzLTUNZ9WpyOKMnOaWQCUJWaTNmYfhmmgE4TYWEa
epiduJdb+ai/38Vf2rWUcfBBb73A3GoV3+v7TG4Cr2cTJc5jjNk9mMIB/y80jYmchi24QB5U2wgf
lwerbzWwZDnEqONG+NOWSvAQX0+1dbz2QaCVTG0XE89A9EpWAd7o9U44wJtQ090KqASKHBELnCUo
GreZ5D4+opCcZAa9NpINrledIuzurc1v+VN+AVOdDL1lzbBmidQUXBG4yZ9nilcuFWPs3Z/ThUZV
PG35ioeIBkFAtoXRO1SSChzH4gAOyXfvTeLM/GZLulmiyei03uZKF+9LRAf5w6sipfqfTyMwnMzs
rPKpXYRbQ/V4TmbFoU8Hle5DYYyhBaRD/eKtNROfmNWJPlD9AJlwv7GHzt2qYHvPxXwVCkpKQ1l7
coWcR441vcnXatmxT5ohpQpSbfzEId09W/cpSlkaFg8plFxMqrYCQ+I+BEGF3tbPLZab3vi+xVUx
DaTfZSVJfhtWxqJ864jXDyj8qcPrVfsL/kPxlmuOKyMgnRvBkoNhwNUUwjixqDpkl81N3kfCHEva
izWg+9TRS24eyujqnaicdBsyLZJgUxQc6uCPmoXGmF7XeVxhORJugP6FiuJngnCHUBolZvc9+c3r
yLce4kLkZ6sNuOAR56ziuSs+bPyNNZzRBX0DB/J7AMJOT8WJnXqAlNWCe0hXarEteCGsVOg6HIzs
uZWpQUs1eTcc9maU0YolW+RjXHR+GOu0cwR+hFG2xwO6j83Sy2oe2DNcjObUnwclnVXHyx6hKOm7
5tTC/AI8E42FoN0TJ9tIjD39xcQEc8lnxfQtdY6Fd4D3837VYtK7ny2xJ5ehYXysfTsXQrXHIT9D
KexcLZEFpweUH3+0QRTtFv3/VcU1LkWtZ4/HYtqWP00gOQI9A5l+hmuqgwCb7nG4n58CPoI4UBR1
Ud3uQbdaCGamC8Yu3JwB+tlOMl5D634VQ4N6oJlcI621Z4SknTDSfWKqBJhM7eHKaWEq6gD+QrDO
G0NJfDBvRsKeIppVlVUHn8wFEh/Cp0qabUfze4drDybhZOHlc382MJU69QKcJJQk9lhED/GWige+
IYRy2eUWgUUznHRC9H6wX+dXum0pe7UU5mQ3X3ID7/rQlbvhHilUcHJvzSE4wscfHd7c/MXXbm3y
L49Yga/iz8BRnay71IUwCMRGp8ZUBHwNcQVqOALL/v5ZTpMz1Ynk6ShXeBWmXLjpjwsxUlVpBczr
VYo8/6JMtMxqapB9dIxRVQfo/tlJvlCFxLNWRU1pe/iCGZpYzd482hlG7bepZFAjgsIm0ClPKj/g
Oo3ckKuv9zjBEo/sZeefIQA8bMl8MYItK9kuD2Uti6SPF1eRH7+48sichEG8EpWCeUMjmZOAzGBi
9/WPAwOoV1m//VlmQ1cNkubFfvCyrwRQ/BhiIli4i0ekbaQKowEn0RtBayad+1ys2eweyypDnPQT
QNbdYY6gi3UqcYu55iX2AA9si9jk05s8l9gOn9b9NHmZfKSGmxcD2NLz//kid32TQH9whSE3qt9J
5N24c4vV2CRrz4XQhbT6YpIlCFxgKFRzZaH7NtbUoLdlvN01RRFvPfl5DOcY+c2Gjw7dBs3DRiw8
9P9c6KzMYIB3Uj7hoTwxugNUR3bwHrMzQ7Ff+HaW/TPc3YYPp3z1C9m0allQRZDeaePBLJ6xIjX+
hRpd8rvZxn9RukGd5bP4t7BARgOqL7DONjy2eJsjb88S0OIZYdmFUgYaukI3C02w5dayDgAvOHlU
yVXj/wbflcO/hLpS0SJdalLyhopQBS2GqvfjVRPjIt1j/+jA7G5FWOA/PrSPfwIFsrFUGklXu5pv
kRF5uW4xM2DjQ94PRTgOkwFDsy3/w9V8TO45wgda8fo/uglMrLiuJEKBXwJy8LkF2M5cbAst3w+Q
zNX38FaC3CMny1ksMXMwkgYC8wwhzwwSHmSr99H7a4RWfsV8jAk73d+79U8523r0tHK+7U7SPgM6
1TH8B9eVC0tR88GBBLHej3Myeasl6RmtPkRwPP4pLkcGw3cehznldt536aIANKjnX8iYAdDEd5a3
mzsfCnmi2QSnna/zmzLYr2epP+aGS+/M9tNCyFfXEd3ABHETsI6sOUQi5hAShL3HDDTpOhDRXxSn
5AJY8lVwAcYp3AhKHivwIyYDwTDeTn2NR5nO85JATUtwG58DJWsQP9yiLlMKUCN6wgI4ueGwGDkH
JnjjjaHkRKm9qh3lpFUBAbJg0aOukIAZwqVZHmQ+ejFqwJ3Z2c+edCbQsIPPEEciBAjUZpASbLXL
iiVR3hEZhYLtcdLmnGi7YXiz45AxAxMRkD3K9WDfV3sYgKZBFScA0AWTQHcXknRY8G8me6Ocp6OR
JHUKhDH8lG8HMO2oCsT6bwiScpyDC0VNyX4wopwdJjRz0GLPLZjMYTgf6dfAZRxWNOYmY3pEiAsq
InTPu0f2Q/y6vimz+7PCAlM8pyfj2GsvckuNI6/OdmTXBRV8QEDd6pmsuy+PBEwPQXDCekgu0U2Y
Sy3CPugTS0z+8IO6gNs2UujkivrEhFnhY5USW2idRdVmA99unR9BPGMilTvStsgoHTgErsZfA3J2
3eavB27wqWyhKvAYdE/HBfNF/0SSRsp5olS6m4CsGEM2YJdyVV3rA33FgCsyMpJuT7eiFLDKjIpO
zsIU54orNSHMRJCYqsRLv2UvjD24TDnew+ukUCtxMSEeDB3xN+WbfsfeqNHjJQulxDKcQcO4igqV
uz3kNxPKRRy9/Jyvat1AdMMwEJ72HwwjMHWhMbij5ZfDCGb+s5b5E30t9aakjwLlJxw+22Snp5y6
dWs4+Sa0pVlup0Hpai6/BiCsVm9Vm0eytjJzWrMwF8+fCPgQwIth5pwMCZuOunI9Ig6oQ2XDiP6m
1x0NHACSPLppz8wa3ugpI7QpdVw1KyL6maD2b1emHgRIWfiIvgtnMKcbOHS9+K6mTjoVSMQEbRAz
2lhlkiOnH5YIhMxdTbU1vZv9zFOcEahxGngYf1nR83GIIeClI8C1E2h9M0cXMZe8idhOrOk+MO4J
h/6iJSloPGEIizzogwnwdiGBveLcSL+yQfVBaKw3o/g0OIPWfT/hl0GGxNfJXq2MiBmSGmQx7McK
CvTxExNjlgYqWrgN4RG2s9wZVJBibKhgyoEATh6fNrfPIRycs6xTRZnnF2saBdUmOb6dK6X30a/N
xqRckHBPCOnY0olQ7Gr1Urgt7/Vii8OgTesj56gdcNeP/cc8HWd6ldrpXxPsbJ2GDRe1QG33TCjt
eCBPxB+F4dEK04fuEnTPIt5TPtflhXBVe0PXGDp8N5SfZ1DzQwkhdLTUs9rzmiepdE8uzXklOkSw
pk0xuveLQLVZlgz412C2DNCrokFJqbrJbsqLbcYZpgVgl5PAPKumBnpxFmV8eDmVvF7WEg4z6dlJ
BQZwKpx9a2/7tIumulhZhfH3hllat5jA33Q2Aigr6I4RyT33LEIgFtdHOngrofo5HOp8msTmZqnq
MwGpTe7q7KU0koOqGv4bwAS3yqel9OpOfLn+nuEWKq/QNHbfTRf3dgkZUonu34W3DkQ3s7pbQsbq
QnDDhUwA5hdtNJTn7XeTzfVtRGYy1MgNWp1pEbcUnhkGldpx+MRDNNIhhbF9nDI+geKVOV2alQNt
X2bjQyDqWG4MkjgLhUpj+AEiAWXarGCF5cbQDw2AyRln/lYVQzyts753ukwcCYIv3apK+A9mBbEl
mQANkrsRgkxXkk15UCo1AB2DGmjVrc54m0OGdmnRGl2D5l4tl71Q728tLQw56PD9OTMQJwACq0ww
ZTrrV0puaww1n4q3xnbzLfTPdq1+aSdIYbZgkmu0KIYufECX7JrdYwkd0FMupBFem65eOGkVk6TR
QxtZqw90OxroohZFw193nEqwFK9Wi/M1ozEpsA1t+7BYpYKGuq/gVdZmfym7izqCpjPXp4CK/mwM
DIfXZS2UXqcPvlGCa841eyX9MotTA/alJ1GW+ucsLir5jAbaTgWmcgk8UNwwHLikOLA6gRq95Tg0
HYFDbn9uXXIjAE5h9b77QkEVVTvZbIXn6tXKdsetLNEviCNIHSX3CfZGrBQKLJVAhPnaEW/q6TMX
gDs9IqUsOZkO/IWAbXQyYYFYIYKeu3DJuwNmEpp5hmO1WyykPNu5GwoMpZig1SG/tBw1Aazlj15n
T5FsNDNa85AVUaWxXSkT2q1Zv4eJar7nBpEyvwTabJf3X9W4CxPoRhYXPTNBwI5yadcneG5iqDWC
hY0n2r979vExcmTRTj4HHqMdW1bK/DBTVS28xwM2ySRxOEYmdYdgynCBWbRfnHMPOGNXpjqgw+yB
F7O44LcY70E5MkkC32hxSXsHlcDYVBEor+EPOVPWBcK6diyviOu8N6gQlYU2oi5JtxEsmqHg2GXM
SCr/e3Lmp+YatnfM0Sq66Dv6B/L8dKVV1S0ov7859tNKhj7/GvhJCe+CJuCS5J987Bhx26b+a6QO
Q1m5Qwr+F51dAEBkv8s/FNWgPaKj4M/6by5VUxeBQdgVQ6uR3kbb6+9svcLxA0SfHlw1D8D9xyEj
EC0GFCFrRoGPdc68mCiKfI9fu733J7Pjji0uhty9AUlCWCWHcWVaL6KX9I5x9jSn4DZKvP9rtfCp
HYofKufLyDPfMmIVePjud3W/AEB1QNpKWoGp2BwdqEFcGXHTcbqnL+LemXf0+/hapnM6NUgIiZeL
zWdpyofGw73h2H0Fo2IDzS4PlUAH5X3IcCrFPs/q8N7ydEIpFEeSoksVjkdBA0RqT92W7hlUsOvO
5DK2aNW2jz6VdXDQGj0sZh+aq68B9+WNad8D+/aX6xNGtKl0OTe74yYZFtXIU0qpj/IGVDJJRckr
ry6icspHRYUAYiLNazanQHYhWnorICbjnefKcW3AuTK7k62D6EaGMeiBQWX7qD2DyzAstJiU+OAt
OEW4HovP1vv0zD2BGfHM46mVDt6m0aYkt8x0ZTl+qLdS/2vD4L9mn34L0lJt/0K2QcNQtK+w1LDf
ee4iNRgD7ZAyMkJu9LznBgiwfKH+Ynf4V72mqO2I41nC9VElc0C1zBB1GK0oiv0dPRfB8yC7Bf7g
qPD9S8mf7C7v6bWyodcLGOZLgThWZcbeOCsPPoRrhRxE8dIO4ogmEkzpGEOWgFUdp+47lwp2Cdyw
sCqqIQQ2Aywfn71QrOKONN73AZ+zHdapZSgbTexiuiyBsyEWIa6vOI7CatnRahlEDZujgaz83I6v
VTc8rDGObv7TZqwRLw2C1ISZ+3Qm45E8bJnZCtmlMkbUiSWAX2pa9ycBSZXAmjK5mRUPs8vPBGO+
l6aQsTTju5qzvh2eBpU7o9ERRY/wZ6L8YAqoResSWswSHPwBVZeFAC0fEa/SlZiMWjxwnE1ESa6O
HZvgEzRpxZLBClLKjIBbpkqf2VahISQPrgwoVw105iEX8Ftnr27OvDhPrhCS0MqZa1ymXu8jflFA
yIRZW/LyqgZ96K+8+Zu8jl8xO3caqxLNuxCHYXz0isvRq+48XeG1Br46w7r5FYKjtuQ3fWloxVVu
WWbuKL8R8OpG13HoZKGihcc0tt5udilnOgKvl7w9uKx0gkOkFIy43+TqxWsJnqRK5WYIrQB9d78A
PfzhZMKZ+IO8WtAODn0pWe8Q6wpr1atErSDdrzeOr+8W9Cp8g0vIHmuGhYLlBBHvcE3ramiC7kv6
kz8GSWHepjW87HhmGAJc+CLepOVfvo3CLHJnIJGtsCZzbruWWFoTuJ2Lo9o1sqYmEbcYOtEEFvui
TcRWZRoorrS5W7CWeuG6gQFDsYoj031h9TEeA63yid5jFYuJHwr6dfh0EW5qht/Oe9VRm4LvMTyf
IWSnx1A5fLBy3Sb4RQXFfmuGNfswsGqMdblPkncIlLETCH56Pbte7WvIAgFZkX5MaYaR9zguwSQ5
FGKq30wyx3AKvi1alJAFvggDnILaUYIw50XUdPjjb3SM+CBmchvPaqMAKMMjKckfWlpbRPk5i9rg
sH8l51cO0yY2UtbKKYZxm1yBrcZLplt0GNC+NjCvLQG7Netek3yGGDkY/xQ/xxL4U6XYYibVDD/g
ben4ISuKnLslv1Ycxcee9vGVeJYSyaxvLLcSUPyf7Q9lyX4QTS4ymvMlZdkjzbzOj8+d0ghQyI5B
GELBw8xGN0ki69jUnTFAGYCSXw2lz4LA6N+whucO5mXVyNhFrcURNGZrN10pJwCudHOuR13QFDg9
FznGyQiIUKt4ClYbl95CROMWjnC9diIVAGQ1j6NHZcN+CTk/rThixijXBC7aJ1vkfjyPbQQO89mX
HzcncqfxuiCdrnBNk6IGZbTHiMdPYC3zCNv5/UNN3n/UppnTRms8h/zZrU/tb5BBoG/iI8Dp3LAw
y9VGHjj9XKXxbcze6EYO8wD4hMzFBo0G8bM/DdZUhMwANuMfQQq+vKYKu4/wBN/TkekgFN8ciVhk
nkJqkGl6YGyEG4dfzjM8Mu60Qi33kEzvSFctEFqISV+evcfo1orRbKYCKcUdXkZFropKeRrq7bc9
xJuxB36BYrbE2b/q78RAW1c00WwqtIg89hr5DrIgzeqKW1vn9fFYhCDsfMxNlvspVsaoFpTczzRl
INMLh6Nz8q5V8FhtKGz0Eb0n0LWz54GUpwzGzb4IkLLX9cfPEAs1ry/kR/3MegFX4V647xIAFqSl
+Dqs0e3BO0LK9XTyFXp9MHXJgX/AQpaSg+/+8raFwUlP33aGSHxDb9MhMtO/OX8Wvm/JFCxIL15L
yeGgd0XFSGR/d8VftNNBCRJp0mLFhFeMGfcSJ+da2Jxn3h9ZR7+KPHhUvO6ALLt4gH4QIVvTD86J
Ia+ZlpiIv1P10vX/sHyzGCrYQNoY6DH2xyUcRqpyWkdnMlduSU9wgGa5QJ1zU2EqpnJfkyPeKrlW
bshCGxgptIqRvDHQo2LVt8trRmrgbPG0xu7e+UoI9kWUeWnxUV29mxU3W4CgXGe36Hks8NWaV0M7
tOmDmRal1EJ+DdE/VAL+X8psY/ucvRvAVf1zVkRSSJLO9lNHuguDuTQkGqfWsj9oKfF5AgNvExWQ
CimWGZT7TL+D5xSpXEXuJz1iCucrJCka+4LI2Fw0CjMrlxAOYhpthQ1ypZabRc3juB+p6XVDqhJQ
ZUOXh/4mNDbqol27xL36zdo69vX39v1+iarKBfu7xLX6gAOH7Wwg8iRPfxIY9UhhMctw7YDlugcB
F/7owUwza2BpA1s+TFRJKh9DKnR8x4bpsAnWR5dff4yrLMRhHhUISJZUoGXzc62o9gbhZId5k6xN
WrZsrLD9bq/A+Zfr8UQdpnkWJY4pBSknVfJ3lFhxSbCVwx3irxn7uiEJ3SOzG3vyfc2ZL6wmagLI
colyirr/6pvXLpsaEMkqIB81DWaYUkqudV6fJCf1af/myU6Ugw0thGNudx4u+PxCgTQ1vR4hlA1T
212vfYWKiJyfknNaCFe1F2nPt9P6MX+XfrwWMXW03gW4XUB9JeoB+klykXBJorctZjE8M0dOWCtP
oyGzHMuQUtcMw8FTKuUaUdNc8Pi7pOuUCVQ9kjHPaliHwq1DORqrD40gojhC9cT8OuujBhxhP8lF
0kYe2KS1O37GY1No7WG75mMdq7mpZqdo5WVebn/kAIealLjyiodwKYeQg5a5TMlpgRPtG1pQO7ok
U1S0+qiVn4BDmKtQydZAzwqvRTpHVqZokLDUtErTTIc0azEUNypP7NV0F/RKOXUBabQ0XoLme96I
oWWYfv0CHVYMleXiMp7fhdT3zvJtg5A9/cBLlUs97q1lfy9yJk0lMktTS0TcndqkaC1rvpc8L01g
bKyF5hwRtvTBrLIRt5SVDJ6jDpLtLjFqNuoMBCd5Lnnec32CGgfI7Bxmk1qLo5EfJjttJ8VSJPod
DqDflRJWRFsCWAPs9qt7FsZhNT+/eF/dtPukqBRFWBavYIIUKwznCMz+3aH71fotaDwOhqjbpVVU
0cs9KKcspC6ZMYEFuo46ypGJVlopdEC1p73ZqVF3h0M2wVJwN7h3oWxJ4jEV0xO7Q9SHk/Mcevkv
dUuhPazrKbNZNgLCTm+KlQa9FA6IW7Chm0II66kOc2zWUavQ0imHqrUaHCTPseQGZ0lMumbgzw7y
T6pYbPjJFxUMTKSPHYmx/Xrw6wL1p4lOxOgxcbuNGYwNu0rzNdJ59WDeKOMP/heINIpCMtFv2Gyz
tG++QovRa0utVz4j4iN/x19Irf4GaxRmsJrkKiVFgLuN79N9tFlyZ1+otl04o0227uGAY8PNTZKb
KOxn4b3GPrVlw1boWIPmngb4jE/VOreNPH7IDVSiBE372ZrhxEGExdsM26rBmVb0UIuw72v2bP2M
pVtCxfxZ7ZZ6f9OKd8m17eqwYD11EKhe9sYZEgyX4JyqK3ld4ZBW6ycWb9ymdYDHm7pKhcrmJxzm
tCklXvaMOCTcpRu02e6DVAqjzPnF5k4PhI2EvSINBJ+av1411YFOF7X2xAesCt/MayI4DTalQjLI
IMIyrurT/TKA3Dmt5fhtx0rYwyMZn/dvPlINULtWUzrzH4uSxvWoN/bFjFiduDZr88jmIR3S8EWm
r3rPYpjA7S16pYze9q0gQg+yqbp7HXSEGEeDDE7QlyUNwzCT2xY/N30IFj1g/FKwnGYreuXb8Fkh
LPGEHyvUbsBD7rKHHi/CDErlG7dcEwLMm/5ALGUaZsRKcn0x5FojKnywgI94yqs3KC8x1E/ns9Ru
G/wvto8JExZEYQJ3HXwIXLJpOc1FGoU0ZW+sotrxlDSl2RO7e1QJwkRwKWeVCIOK0KpPcU4yeTEZ
+6473ft/gLFnAvRGu8IloyZmC2+ovlEBblIocr6fjJL+5uycgTWKxC06HKuoIRQnFpJR3GzgcUEL
hnq/R54cjaKx+SxAaxPQiUAPfn3x8CFuZBQ3pXyRQyb0WkWiKAfe12nYx2zXXmxpOJl+8xiwH1g5
H/oa12WReHQvEYMB0yqficj4dpAjitBGmYVQzYBghvY+mqoFkWdcPczH+FR2ZImBaNyFUAr6ZLcx
hRAgU4a9BGOGk1tXS5Th1pLP21v57m6eIub2y7/KhTVYhsuTl0o5HVxK2oysz7v1kEDpa+Of52tw
Fr154EuUzge2GIDdqonxeyvqqloZT6IDogniiW4DT8dCmXfrE3vscTJQ0Gj2UG+xNFrfuRn+ppb+
wI8Hu0gqZRV1kkuvR2ANAcCK7s4X+tpkcWClR1/jjAEzF8BaID+iUIeDadZ5d62IU8+JCLN09vM/
Vn2hkS0+QlUlu/ilu4fsHfBf+e8rGwTmGAIMXfrO+VJxbgs0r8G+SzIZ58jgRmOm6TylBczsJrYa
dPLQI+v4J8Aew/gRUdter6JIdLYRd3LpRxWG6AgQFkhTdmKEWK44zBrGNOZouXsE4MsyoU1oQcvp
dUhiM9zEZVYUQgZxMP8zDErlmcJIdBP8v4jwArpx6QbPQehrxQJgeZHLN5E/1QYHHQEPaiDWyWkK
MMcaTw5iqDXALjw/myJriwi44zFYOzvSHAfwqg7GMI4MPKEEpEeS62ayqvxSs1E8uBNivaRMChcz
QzcJcOgko9kwHUJPdedHz4PnEpchQKqkeu4onkcFqQ7W0IMJaK6AhQb9saqfuKrBUVxsDQQwag4G
z8jhb4tmMzFU8WXxOp7yLJRwijdB4ROsVDVpvQRvftOvbF3/uEC6qjABI4v9rA/qIS/qss4XQ2hr
0k9ffht1lux1oEg0+UjfKYAKQSOPVz5b7trb6rPO3zpGvDnWfbJV0S34/b/YG6qGzgopxDQ7zvSG
esSWpjD8t0Zkgmi5q8ldgbthwnYw/0mgM01wukotYqq4ChSYiuvs1/ayi70ycX7ngaVKKPuBfLxg
CeogdlBeyc5Mb4t72HQAZdaG3iuV+7m0uOGd7cKWKju8qJqLWzTvkOCEik9dm8xWDzrJP47HQp4C
Arvi1XVsJiWDi2PYXcAsfN0tYy7NFcMmSCa6TFGd6+hW1qTriFKPWNLgWhuLRyYpFZMnyQj3CTTD
5Dmsuay4vqCUQsN1q7It4C+tZobTxIFIBiy2jZajWK/YQ9N8TbFWaQLZA5aKWDGWLgJaDrwxX3St
kyvT4gAsQUGV/l+mag0/3X1F9Wi4o+Frp47CRfbtw5J8p2Q2ZQEUmjBa1iQbWmIXsFFvWaGdFJyM
R9oJsnXDn3NCGx2j/3Okf2MktmYOMnakI5erPjqYBovwvUcc8cBwwpPTLdXLO8Hx2zr6+nBIMRSB
zDEij2T3rghPwj8+6OFyaEW2c8c0YiV7TqALQ8mODgCDUnZ2a6K9QfXlARrXjyXixShV0KapE1DZ
tlZTSQnWzbZKqtbgLGuYWVycB8lzYZodvmYKLBPNPn5wEEi1mltrCMFrmq3+sCfUHt097FX8nWbx
b87IeqYNCmn7u76gPPZ5W7kqDi0ShnPMVdzQf1gHLvnbhMYcSj5VW4EfmbAXMaxwFdy09WzyQV9l
2MYeTOGfK7SQo+isx3RZm/dLIKDIww9x7MHVAHDGO0fKRZcg8Q8Vm25KHmCT/9HXx0fsr/GtGs5L
SMxD+9aqnsZj6bvCVn79qVjnRs0NVgMD8MV5pCHQKytYwTxIQFa0/YLF+Ee+BQyFjbJqLsZVkJeO
w398PmvYPnHzg5wAH3w1lfZXyyb4zWfQhV87Q75xifUDgfQCtuVI2PpcK6+s11C2oS1k27UMZMPi
agMDixBSIokGTbchFStHAUQjc2Rf4ClEE5Qo/qf7bUeSRKb+ORfDHP9hk5h3vxe3QqZvFiE2L5v/
69bcFvPfR05s0siAqjzeDDDGi5bZxO1FT1+16yrPLWagBI/RFRSAaRPb74YPnlr4q+k8PC8vGeeN
6ziWaAUZ50uFjuOsT/6Y/X0xYruJqGy4YmxQuSO8QxHCdvB5u1w35QZ4mboFtEWTgmShFVlgLI89
W4EjuTC0wy/hprrBlizSiO1NGkKmyQs+pAYipis5lbk7iJmb6Z9JxaD7MEbPW1AyIjv6YewjON4c
uViKqWDTuB2h+mXFr3YVNaAVbGeiJMSID0KKjy8BbuoYNYhtXfbdbFLHvsgANsmayam/szGAG50Q
61VrfewMmqLKczP3rrBoflnbQtgbybBX0s17YGCJBMNpDlwTxGGnAUVshPZ+G6+3wJ/TqGabmOWv
29Aeh5AGwAmyU/5SkFmY5f+8sYABceDlhJlNb7FzvJUsi6Fj1E120N2ddMervAfS1lDitLqrZH6D
t1fw7REDkbNTklO6r3C6LNxfqlDWtfqOKeJDqXxuKC2gHixNq8+PwtW+dfbze8iatZAkRpSu8Amx
zE8FU65aGeRA/Wmyskyzvr9hmYhiCIZ4Zd5Jdpc3h7BTWIMKjIyNwmItsRL0+yvLSsDdytByRUBW
vYN5V46Mh6/rfRb7obZCQFXxcqIBLgxes/cnin/gvpWQi4jTcl1yg7iimAxfwNyXypdDqtseLIP8
dgIiDLJGAsbyx56h4TnEmG4RvRaGT2JKmqeaYH2F5VbA8/v53zHWgArnxsHneVHC7j/sNOLI7Iuu
oX+ZL/+kwZwjjlppFRgmbN7DqSJ7jeZ22oJzE80pkjhD9Ecl4XBjg/UfAcwsyfhPr+wM9ZEfzY0j
4o+ajyy+VloHH2EZDwHUfNHGbsX9wcB7heUgpgT7A5mnYVIez/Ddvc1MmD8bai4J5rINTP9srtaa
j7oxueoKIXUnSUYioCa+gmFq7cVINiy3x2vGEo/1WzQxYNvM2iCG6TrPTJwTc6sXj3yWAqx2hsZo
s/cCUi7wfa44qyDoy8hzU3aV6isGF3fnAeCHb7KsAYT8WGyskfw67xzoyQr529St3ppeXTY3dE4L
TZXRGnfl6hcZmCuM5kkWU55/kv8syTYtdjK0sVoPaIK2rvvewzyW7Stst7sq+rk27W19k7b/JmA4
VkVx5bORXM44qj2CHhRp2EV1AlRvjpBYyU8KKuJE2WD4cIw/dTIOKGgG7nymqjYCWFQX80AMAPsF
Qy8gLN09Vbze/u4CgEmUuOwS6jZ3FgiRDhS0RJ2myWi5aoaf87cZs33Kh5GwEYZT5NlhdRHaNhIO
ivaqqFWn1izo8sA63cSB6eEDusEFIZjxPrqWhS+kYXljce0IAFF6HSBcCL/FNfX3HY/YbZgc17kR
h4D1m+Kkco722e+IyQaqWh4qCN9O2L23m1ag/hKU6kUTIJfXgWAW+CRve19b+LFUJrE51LoPhjhE
oQ6/J1PvHPnHtmyiM27aD0GsNNyl76cRKZ31pgLS3mr6F6NfXU4ZOjqYCkPoRxNJA9gsJ6cKVSMx
+fEhXKX+sp5YZ1HIy1ggN16stPxyJy/WWIHPPw9IyAletUivJG/4gfWuOnPo3qpNEDcVvXrPIF9F
f22jcDRJyykBBTupM++D84xBEgC95+YE4I5PpRjxSu/4mKVhRf0BVuJUULozAMZED/D8yrlm8Wlf
6IRrnG3TzylOsWjdPADlYiCKbTbwqcIUaISyuGC3XaQShBrn025Yo1p7JnmTJS30Gb+YkhWlW2XT
0D/yU39sjJGMANIRdzNHqx6b4ZSOAYvzmS7e2d7S4VlqOsEOr5wmph0iuczERhdI9AN6Sh2AoN5a
CXWRGuLIDl3dHFOOcMwHJJZvG6us/c8a4oPPz2hebUnt2vLQCZa1GBkI889f59bjLuTnIWN14RSA
qUVfwlSsGJTfHtz1mUWvnSKqdaonILyM7hhd4tgNf7hVyOYcR+qEKogpC0oiaHnabvHNg2sOmQ9L
lFLLm93LV3ZSUIoWVuzqphSfR7fA/Ndb77e7D1rIj2/6eWs13EEbf4/l1xe2M7D7MPasPbSgcsjV
ZSVywK1wz4zRKSXdktyGkp72NDUBJZ/tRsX62ykxYN7v/npF65hxFNiUC/rm+wEeOXGNU8wkWSHc
nJ4SnX3wgWaAowSJ84WEsJkN7FS5fgxQ3yZUppcKJp+aHbcR7/ax+rzFjyI5OG1W58h1itMAvOCz
a/aEwvncp/sqcdHOaoQHET6sssygebQz1X37Qtt20FS/cJAkVihRwBsJYmgGa9cOJ3IHupRH6DLE
FA5q6tNDe+GQh8fc1sJtElsvG7c5cwd0xxUyNs9tISm/zcWV7jRXI84ipKayzZ9mSfK9VIYV9g7u
cVZGew024HRgXYu9fGKZyaha10wWa7PTOT+XfBK3XGQ8gL2KXmCsR+mDnU6IwyW4Xj1JrEIruFFB
cXVUbR81H/7ja1b83EyKIJnXFfPHkV/9f3zaxndeli5KuPdS2ovQaG2sS4srkphiAw+/lmp/KjNV
Qbp63OIcMP/TrqcoszqtzPNj5gdpY+zPb/zCKeRHtp3ZD9xj6001hP4TLVgem2BPXI7FJm4mObVE
qoEDFbhFOGvcCHnFkXU3cPZBtQlA5qrXkTlU9k/nhORJ7LZaiwITG9uyWNeI1J3OFJ2kI+K9IZCi
asstJYPi01vdDkP32VoBkMqvHJRtz9LIFxckiU6u5uAjFsoyQnMDmPzg9lsN1/JVcPZkbsdJNsGP
aaD3qogtXs/JbncrNQILFJ+Ba4l/h5zClkpyOXhHpwf2npcovnq/4KTu0u2kNMPsisQ75yr/5YIH
gXXxNqjqPgkXcb6C07Wjamo1rLH3PzrBwOFzoX++9//viy///dWekVKaazKuNhJEI4xjdhxkhhUV
4bYkXoRmZ+IHUTY9XxqZWUYMsMpW2TxCEdyxtTX+9nbGjT2fuo01uWfK8B/OtB/ftPdr4ZMj/0UL
aQUiyvfHIsifNH6MZp5bW8mBgrWnWrB33fHuGuSM6xs/PEwrVG2I11YjpLJHsvBzdR1CTS6ELp7u
nSmN75UXg4pjzDEYVwORYviD2B1qz2ljjvRFBUNGQz8dWuQ2LdCQsQ9Yco9DBbOrGqfcuH3Zf/g6
l3tOXeQNOHJSg1dXm8XzNjkRLO0Y+SDGQfHNj7/siqGeK9sRU2CF43oGHJc16q93KRmnn49h8ObZ
lD79Jdx2fVtRyDs27HfXVoWrq6DSkrHUzsEd5tFPUxOeIaI2cdNdUH9INZtX6Od6DNt8436KzQVu
TYOFsTloMlgs8AePSdrLoLSHYDHNk6bDgvcQz1mc/4sWXNIyqUz/3cC47ZQ2pXdfIYfQIrCJ795X
gk9Eg8bm5tDi7OpfXNMT42cIgToldHFth/fqb6DPgKatXbmCw2+iLNaQZgBzlu9dFLw7ZwtUJ9En
OtzsEC1QQ54NYq7nH0Ozsr/an8PjxTauPo74d5Y/XH7kV1Q+iOssy6/Ee6ksPLYRKfyEkygdrqtr
IkbIaD8u+gsl7m9akBkqjGMep+UyD90iInnHL2eWpRAnn/A0GUJjpmbZ4wfdl3e+gUQW7S7mkBqT
o6/u9dccGjo06SmYX9dMlKkZhAZTkHJ5OJhjefESGMiymiyKkM6AyjpicyDIK8V26bJvGpEzXI07
oippf9cEWSY33pQmiTwCqO4b9ZbJ9rR14xhoEeiqYaRNEh/LzgCzLOXbhO4mQNP9mdaMKr6vE0KH
4K7hW5XpoyLGKV4sKUDv0htpNqb87LV/74zBc4dvdn8gG0mqo/cs1Ld6r8SzY5EpHnmemqBCSy+D
A2xR0gpwEmv9PnyOeTnTHXYNhGFwdc+f0ONebb7UexzcpAo15rwZdhqs32ok/3n2Wr9iMONdCDIQ
iVZvTBKxiMnn+ckp668BKHc6aTQlIY6kbhNYB/DGk/35WsOd0IwOMptPObw5DafIBpWC/ABF9LHg
L3W8LoGDpHJEAGJZ8KM0dTNR2wDmIbFJxF82noexvdocGeWgBF3Oa8hhA9lPiQi87el0j8pApK5l
U3/B6A7uUCHJD1J52bB47demd90y6Znuj0KHrNVvOx64n5AHbTzFvmp8nbhw2NZ6ieavWiyM30+s
SQcBi1GyZicSrhkBD6O5fQezVCWLiKIbdxFPHp/GouP1rPrG9j6iROjrWm4TrK+jldAFQZDw30+X
/J4PSp1395JEwz3eYX30odv/4IwDCFJKAiqMkyr75SOjx6FqyaJYBAVDQOqT4pfdCuKOEbiCUNVi
ph8gSXGPynNcyJxHgwhAk3//R0pcDvcJSxmDjFEtmfLwwcA+W74i8zvW5mJHfQGTUzExZL0ereaG
Hokcw2s6VbC1ieiG6DYZbbOkuDo7sD0F3iSmnO5uEYXPhk3xnpGQePsBCNUiQCPvFw5p9Is7mmX6
GVT6FlNAznvmHVE7mYJXYMNKlh9Wk2wZy847bAs2L5jCxAFBcrY6dne9Tr59oNunkWguY8OcXGGo
ZwqVgJzEyqmNv/ANBv58Iji5X8wKFSfwXOkX4n3sc1AMbPHWUBXWinRto5Kvit5Ql8jsMzMS7vDJ
RaWCiX+TwtgPA1qbT0SwEoV1hHzBH82ZGY99LUFv3uFQUCO1X9lnrNozyZ96+v0Jw69n2a3o3vr6
lQC+Bw3PP8SvNzIe6kgJqqfwUNV3QZGB7cK9a3+UGEcsIOJkr39XuAlQKJPksalRKmB3TEynnpxq
Gp975nypaQLgpros6c2qGMtRjdHel9u4U+BL92a/Iuel8rAs+3QJbILqZFfhwk0ISrFDf347zRUt
3h+qasN7d1mu7ZKOFmkfBQ8MK2bTjosGyq2oehEoDeAY9Jf0VhfEA3W3XbDnjtXr6kgmNqdKSfgY
NfT5U4rM+0FnZkQjOFxJQeTteqt5glgiQK19/DGxc6DXqPkvqNSQjmFZYBd0w/DwfJs30lVBrI+P
Wx9V9i+HwqnkzW+FJ9511XKP/1pHsV33sBBH3NmrybpoS9szCcesjbDw0m2xxVJDu8PgvRri+eFF
ZpY63H1z1jCRVtfKUZdoneVUft/FXAURhxplFyvL2+JMve+s4Z5ArgNyseRxRsPq94EVrCCcLAtE
TYcm61SWa7Chq36zQMqq2WrGp5AYxWEZJUytk5sX63+9scchARrQADRX8+RqzhRTaavdCUmg5sZ8
INpHg/VmeShsPh90QeuOi1iBTK7U78ozCUFlk+Hr4yWmOxAYmQPbIw+FHg6pC21UnVGfaSz0glLa
ppfDemGjFdSe2zeGY1drCMesTpsO4uh+S6WB6bliWrCS+G8p7JhPIsAdnKpHEbREvruGfKfm3AbA
c/SN5zUjjZU4P3We/OqGJAoIfYq6pKqzzQ/mqq+Txabc8h67JqawtDod4EOZTo0NJe5QlBsMkcFV
5iMb+txlyACzbVW/BekSfah1fNBExAWGdFpkalNZdYk7ikU6RTUStXef3CFI1RsrnQ/fCZ1K+otI
BDsqvpeCYuaOIQLc3DHXaqFPZoO8RGXNUhKj95x/724c432CvGAohWwEMN+8i6h6MbhQpIU3EsOF
/i5i1r0hWaFkP8/wiNH1ghBieISVT3ghFyxnmwUokX9uT5Gp3EYvNHg622eVq3W1gTF38mxVqoft
4Uo9a7kIreaCstWYzpWfHfa77iWamT2X4bsx6cmEhjntAMpLOK5vEHESyKZIYN1jGTK4uMfjkc/7
dd/QhfpFdwIPBkzOG9yS8p3RT5pT0PbcQU48qNCV185bAC3GAhKsY6Ul7eZ5BcA1RPEX9hPEMFdi
fme9/KsNtR053/vJiZTE22MgnSwXoa8izKnVWAw418y9ZpuHpkxiPUsUzHeM9c4+Yd+DP/Zgj1hQ
ttS6my5MfEUKqYuZFFeVaDukULcguSrOUgb6V3XV8484V1sq4/9ZTlq+Xag+Do3f8fgjx+dTf5WE
48g9E6S49mXdmnmcGsIeXya2Icdhg/t7QsFBjhcEuGAWvilb0ULpz6biYAon4CpDoWy+A9SOqWJD
j65IUXh0yxlGLlpAH0SkflQYnK/b7fDBfrMAvfqr+6J7cMFs/6wWYZX1KeKj4kztG/+2m0Li89Dw
XSmVpLc3VqgSVfrfZHyEXeWD3VcZqXTkeJ++IGJZHi272JPXOAyZs8V9Kq46lPK04BDCR1XOUkOz
Lqd1T2ZjjG44tgaAYa9ZS9iXUJG+GqQKrZcVBQLXssNq/+B8a58yxQ25SFNmVtAORNuMU1DwE5pQ
ZU8Oi2eAzFKY2XlbS0P/Vun7LeMPB4NwqrEZMhkYjdv/RoGTI28Gj2rbwnNQRbWwAYmXLhLxvtt5
VG3TUXc0WtanFWUTvpQFWtmkRuO2BL+s59VGlpVVp12mimblCsU9OkU348r/8hCEzdGWMftwjpdB
Pc0xP4UUJSOm1W/MdpkZdtQelHnIKOYDnvFL0i1dua78mZE2u9RmEFTmBSowYFFMgCymzE6gawBf
N7CVD9ueVmUet3JNxAKdenbQdsx3aim711+LnkRPJMJTrQzf0iQOwEwo/H5gm1mBIpsyCc5gzWLk
Uu3djDfiAAeJVFXYbTBz7aSS5A9DmDgpXEFtqP05LjW96HM+ZURC8XBfRCtLg+YVX1UwTQc/udDb
Fvnneo1Ou47sEVG69A7rCwGY5J3uW8WUcAybUPxE9GWUTCgV1mi/Aa+48MVELQ23Hy5u1+EBEsa6
oRcAOw4sQEWMZpqnGqaDgQ3iHyCAv/soZLCCY2XnCPOXfQSXDuKvhNDaAgO0BV12Dyli5MxdJ3Pb
TnR1K4yiZs5Q9sZVGaikAfNqGfgHII3cm/IwRBpIHMayc1wVISyWF43PY3JiUuJ2ozi5C40iDLa6
ovtNwC05v+zBSQdlJIwWlk22nbmE04r3H4rzpYdO+1SvqZlwhThwBq2cOUj7XmAsOtHsiiah8B0a
zUQS4D3nzoMo05kVoyvbZ3w4hFvlHp2NimQFT7ItyH+fhArgOR9+/EQkbvs9kKnbPiNB62qAF+2o
NK6dOrDMKS1zNDziLbAehFMWSa/qPS6l+x8jqgYhUlnbER1NHF4C7wKJoGGp/Wx/pbkslRu2IsxA
VVdpqnGqLu/oR+R6N7pI4ChzvjPrY/0gSRDqiJLOmlNlqmKsmRrq0PLYXl9Uc+gr0CgV9jhWcWyO
fDonEWdtyvb9SGhxxcUG+EEhmBBWJOKnm6Md+PORLAOAf7AaT+MaM1LdKUItWnWbyA/lg2Skr8dl
IDM/TSZlMj5o9/ibPPkMfpg474SwGhgjgOE1J6/5GCs2RIYHWjufMmblItAqLV+Aev9kaPMBHtgB
lLrYqkL+PEkcb10iuEt0MliOr+bKRPGguzgH56L/hc5dEltvjmGrDWgWDYDr8iBR2LENeJuQ5RMq
r8x7fkw7a1DJVYf6bV9bVnZUt8JbqPZm1zoPCJjTQ2zAkaWIsI2XU/R+STKX7gt6KFcwL6Oat0n/
JNXCLFiky4WIhCKWziZZJapYQ2B0++5gQKxcl7Vft1baN1+OzfjZ1IPw8517IgtD0SOZHKs3qp4Y
43seHq5cZYDT3nK1ak2fsPmvveIhGx3lqilG/6sckE1IL0x03zkJyrvhesxRE/KhpPXEJzUtbZTl
AQNxpazfSaIsA6HAvnoUzqwO0K9ydRRItLjsDcCWxzNZrVjyWSdx5g83/5g/mR9ZSbNO7AnUgnHI
ZPeAYtSZjgwZ6rnZNUl6YJPXBCfH7ZgHm8F/rAtMQ6e7WY7Bq+WyDtIcsp2ye4gurPt6uUZLNk4w
jYJBSZwq/TOQxpejbL0mjxoFimt0jsgxETuHYgwozscO3qERMbmFkrQGLMGYiwYGN7k8ez7Dhppw
r1ydRxUxvkkgiK5/rnBblrF7eQwr1KIn6r8s+0i7derYBzdMrB9csK0EeIy5PxWIV//xu1uLy6h1
val+3wDiCLSJPeSiKqAylzWX2W4gh6UwRKQghpi8jKuz+uYgI9/tPWu72ofd0iwGWYXnR2r8iRtJ
HS7VSoHl/t69eT9POn/t6E8hSENMPQtt6DZglWRKT3nemitRZfM1Hm4r+0m4DiQK9OQo3xZv+3G3
GHzx0bi6yKoHDqXF/Z3ncZlYK5BLzspeIsq90FgQmG/Pjdcf3vn9+SKeMZe6Kb/QztGOFIrPxXin
OWuYHaItzW3EllJM9swjdWEXPzKDoFOO++UlO1HL19phzY8UPvnULQYG/fgr0k/xYqVeM9ZiyvG8
T6DLqlZG2q1u5m4xb0NktP+IbhE8qRba6jQewU+Zt6qvwPvtkUNxCn81SZYsqFjgkyAxC6NVFRxB
uP0bkee8o8JlI64kXHG5DZH8YQMSkQ/9NooBrLIoztID2LY4D2S5gKQYOKzzAo0rJG9z/Pm9PzHr
1fL8IkLPBxKXSW5Pa3ARct7+r2dWjl7nH4VADs/Bp8pNT2GuUv47t6KiP1RGhIotC7GQpKc6f1dj
o6VXEriRUWfASeyx6zNOcxtj9v+GYqdxEptbmmy0xyMtqKyrt0wZgKQwajS6ycV4kwtPTV5rTYJj
RBgbz+jkbDh2IYA83INOukoZ8gcn+0BGl2StAP+MRfDBBQoaxQ/dngrdF3WzR8bgmILb8cuqW3SX
LdMTNEs6C/WuCqcIvYzjKrcrFdLbrEOGwzbckQ1HN2epT+2pDsXig6HP/OGjpF8O2ahzTGeioxsT
6BcMpJ/LACADIo7SN9xCuHr/5x99YYpRnbYkSxRW1IkqmU+X+lrm9XtV45v8+FZMpS8Ctxs9bTwq
ygCYyE2eEQL2pGSUxgr0g7iI7EKmi0FgDhzS0fEEHwWjpqMVVFKOivnzBizGJPuGB1R8vmLpaukt
VG42TS62Nwt4/o3Lq/1j4qV+uQv4wFSZ41yfkbpeHlxiu9w3ijk6wIRPi17dDA+m1YkLMLkWCLjv
Dww3e+/XJvsjwM6Vk89XU1lOfawwjKCDvbRBEEpBg634FWYA6RYhd3RHH8nZb0aC+fL13PAUD0wF
CxlM4dJXvNJ0NPZ3DWNzRbTGclvs/DpipCQx4UVASuFuqxQLAFxO8Bupa7vtARVMxMmM5BS+V0vu
KwnNcM8cvWRfEOUUVBR7ezTedPJ8a0Nd3qZzDr1I9RSR/8+mgdwzo8HdAPvQI+RoK2np2f3PPpv/
blD9Sw5T7v+JkExUAhnpFtaGGA4dd+AqDT39xDNgJpwLg1rVzHjKBjwOoC7mGGF1Cj1FDKZUm5U7
23q0LRnb+y/jHDuLb1z0EyG+wcksNH3117DuvDHVVaFl7WERrbi5zNgffWBEc4VdTFsj2jUjj7dV
ZPQ+yqwkeQmE/iINtTen8lpgN9Ho0qlFSC3u35IZeu4Sv2V/+5cSqxBAUhsu1/F3YFRDQq06FoTo
IRsQq5TVJfy3HAh23R08t7gVfg9JqRddgtCKZ/+1GYn536ANjMkM0BRlNC9F4tZ6ff/t7t20v2V+
1kOfNbUAGOr2ibs/mU2Mia3nUVsLJFG1rhVo6Ag5ils9pu/9vvla7M3ltkC/QH1eIXQB+84sA+lW
FQZYuHWf1rPGMwJyFlqeD+Uzq8Szph0Qkkq9xXhxY+WYWzL71dA+BrVnvT9AiPIsRQYIFZB1YLrr
jVpHalsxBxSDWgmuLFspYr8BxB2YWcFXkr5i7gvMLouXN6R/nuuJY+iH2QdE1tLL7AHcmAfzLX1d
K7pxL6PMwzzlw2oI8/lmhy1UQGxSolOtvq8CmPwzp7Pe+OgZ+wMxQMwfv3h05bEoUUhBLOkMQXUJ
UwSEo9s7R3PEXM0I3tlb2MtTwueqsDQcTupTfRDJ11r2ADfeeSsfBeqPDxkYhiWMPKfoG3xEW9fC
xhz7R9QJL41FiIhUuWEpeYOgbe3IhQ65j9U5Skdk3pGgkXumG+qv+7/iAOfBkMkIZ1mtoaUP/I+z
LSz6QvHjXyJO6XleIm/k4YQUtQp+R4ELNg2fvgIswT1bmuHY7Pk7yPGt0nMYIWltuyBvrOUso4LN
mdyopRZsBxFWT0CxakbYU2tdWTBdh/MzeP42sjAb47odQySmvSy4IPNUwlvXKYVrKAnsuaMjmR4Y
BJfdThEr+u0FIg8NzyRsNRqvp/ipHz23gc4+Ti6578KUp0DCnStcMVQPJ4PqcNVsnw7Zr45GJIlK
I+qNsjPHG7J/sjxviXrRPKo0bY64IMAW0xGY5ezdfZeTsV7e5K+IZW8KnsB0IPmJVk2VYjkLlQ71
MYCEFDJw+aCEdFeZsZ3/erBO2Qj9hKP56LIqZwOOC3WxvguPte+OSvsIWY+YF05vW+VuLWYCHaYv
fBFSukyq64TsqhPxsM7I0KdEy1S/UwjspQpbC2OyDWVgX+88U0jkkcJOiMmyVxLZ3abD8YHVBnQI
B5IGD9wDmhoeWK5iOq7Pa+5YCUfRLirlkVLuKMyH5GteWqnh2yPKkw8i8ch1mSeAbu4HilgE5mKn
ktQU1BNZibfAVdrhQfjW/ujDF0UOu1oyqYrKdzxWTwY+NUWNk3Wsir8zP8/MW84CLw86UjJ6krNx
nykIBpkfsYD6rbXORgGcQyhvPSDQ7PTebMs7fdgDV0BV3Sp0AN0+eV8Hk8sO+UuMAWYW0QPu4ySh
3k5IpY0C59pbFnbCsX66uNxaqu1hIpmLtFcG/fY/GdJfMh/yJD3sSnlndVktn66KX2yMpZQh+ZXi
x76wbgS7OCMYvYTSp52nSExwb9Ujta3vclCtTwuLIA+2DfsHU8Ei733CxD+PC+/sjlZa3godTQrs
iMoJJBDuLGsuoxRzQHEpqSCScP37PPtsbkM28sDajPVbaSFChqyG4mDkAC38A/Y8JDhU93+u6Zb1
ToJhdejrjcJduWUBy/Y3BoncEYSJU9Y85fE/rT73lL7FyLLH5eFoLOzJdcrFI+GdF2q91rrSKMRb
IQpX935QV74ssfvThqQOjphzCEZ1oBQeP7LKO4YyNXs4a2jXJZUw296T2yfdYs1KEGwCYuMDifkl
qZxjOSYlCky0o3328j1XRm+K/kPBaSlVL8SuLzpC/Bngw/T3i5Oh4I8QlhcU20/8AbvXNSK5D24u
UB6500VExYKYZq/2i3HMuLb0xU2xWI0Nm4JMpEjNLxOj6UyonGisaKtOheI+4H6S6+PX1WssoQ4s
HB4kj5L+yGI9jej2kA2loBMW/qScS1Nlj2LP+rkl9RvosEpMeQBa7cAamijGRVi7db2YpsGdNV5R
mPdKKi5qLQG0Pvei3hX/sY5o30SQfDSlav2LluKoBJrJn2Q3c2/0pyg5jqVaV5qO1w/wpsugCoy1
lK2epdD8HyyJ+G3KqOsQ14CvlIQBOxd2ntQSnzU6B7ToXO5snfEeAqBnxVpfK/D5DAuPgZ+I+ZCi
5gaBueCROfC/YzzxS/1A/UjuWjoY7s0LVUY43oTFXFM6AP8/jGPn5VrnlIyP2l2aEX8eYchb6uk0
e3FVLCCf1movOMXRNnK+E5U0/BAL4u1BjWxKnYAMz9s6OVRY7hb78ioApAfT3VggpNRkT1kCn1Bi
4b1ZOi11bcVzIay89nOKo2EaFNHDZDJAiT8k1WLe/7vek2lMuI/Oqozyw5bBpiZvJn9C0teaeKxD
UMYtBynM+hrKumIxzAh10v0quoNG2mi8IygKFMslN7WqbKG8ditRJ4toSCcRV6VSdgSSqT+GliFW
c//dTJ0eXfZZTEcz5WitiBvzHrat3uc85IuV7+gvhfFaLbB5vaHEb0E7MF+Mq0ynM9NYpd7jT/dP
5GNLjrQbcQMOOVpCNTN9ITW2o2o9IbZE7CYgSE6tP4itUSzkkS6svwCB8IsUNpF0kd5f6ow1Awnr
0s1SBy+g57GIFFcgZ3EXetL/oCi0lozdTAkBxbUDuiTDtvyz2f1/HeRFZWozAVPewmIehEJHB+AW
hMR9xNHieybg5pwJRzC3c61c76nWR/tGaijEJovN44/VMu1DvKxWQx02jKSHcVBRULbe6U4CyBY3
iCXDtywJYJyzQ8DFawGMxyy6pCaSVQ9v3BBYY46aPtY5sNeyrab+xDx8BeNB16ttO9Pl1FgO4y1h
qkSm8/Ce7FNMLe8NXbtbwEemb+HSIreb7L9Usi6FvQJvqs9UHSuAz1jpMjvuwaplCUTVCV6uLXTC
TeE4uxSJehzO9nQqrcTnVYxUVPOZlHxWdrogvQdLNp+Iszsh7dqfnq2qu87jrKotx0I8dwIIwtYk
VRLTDwzHXfLwSK4n7zZzsZKSkyxxn8NJeciYjCPotX3zxyK1LvTZOTo9m4ji1ZnhaK44+8+0oyiP
c80BjL6mig/xWthU7UbAXSyrhxMM9YyYyngom3IYIBqtMPeanBCOk34u9qjobZuy08Zy6DijRUpD
SvcQt6zCGrJmEyAdc3h/M6EViqxUOVKIWql3sthU6NVX6c2kz+YYpxeURAP3jJ/BOvqtOMoVYA59
xJuvQv3eBZCtQdrU3INBeeOy57RLblDI0zhzvJtxFDfAQ+diC45R/oU+wzBF5GtrkxBogEbgc/jv
MZQy8FziO9cdxIjcM39YtPfofi/tyJ48bxbtTzrajxcIF50/B5eQGmsQTyy0FDbR8YEOQDV81Dno
hpcaYz0Jjrb+0bI0nKXnymrwuXsNDTGzDZnA1CS1jUMkuOFXxrR8UiElvsWdVvDp3Qvpl5NUsVwf
dAmNNlIHfd5lVQQGnxOoXLOctWGaHzHspApPjj7MRwzt/ZaLz3SGhMN6w6IE3GIu0gOqfQAiuWfQ
T8fY8nz11KJ2a2DlbDG2O8I0QhNaLXdBrOL5yMUHatsdvwPQz/rrRhREMx5deLGhgZnuicg24Pei
ATpQVKuyj4Owqr9zeoZ6dh39q3JJsRzq0ndFGW2z0RGR1p4ktOsGyji1h1gXRL3Q25H8a+KTzowo
Dw42jC1kRa5gdOG8VofDDY5KCktgz7XZSKKX9noQPaoHi+F9P97et2F2e7N6ggO6xsPFVfIAUwgh
0ozt65UUWoxLmNG7mROrIRrc8pc6sKSjBVNVzDkh76zDY31t92btl4Dbnoz2QQB3mjYaelqUvV7P
tJA12qYnDr2CUb4grjtrgbusybRLtnw2Rc5j+XDotPbJ172GlrbwD76sgJthgW85zwvCXaJrJAhI
mLHD9IqrsL/ChqcsOHQHFKufjUGx5MNHxGHsmT3BmHqJbMaC9mCENtYmY3LZ59XkqxnCCKwZmczK
c+Rohzu9h3BJ/G88ghHZOs4c/JHfiU7jSNnoWSq0H7xfBQOxW08xJUeVaIoizs2qtzsSjN6Dld4Q
TQWSjRtprul0USjrqDQIqgL1GWKtIC5a4IOcQkK5U0i5bkKX84tJbkiRfPJlxnmVx8KKSRO49yhb
Z7e8bOPMMwZYQB/md2AHAvwW5J6jAMgNtJEfq/JXKWm58ApVaKsjKtGfks0sHnNjrsEVrbzE7Ere
GA64Y2vWDGkeAhvxC1hb/vYRsjTDjs9RI2nPARf3sn7BgBAttYKVzxDKK85GXYRWgUMQJNfpwOLC
ogPldwFcjnuHS5xsqagK1d6xyOuzKchjq9nS6plYjQoMYIlXu4adrmo+XhovhInCNHgKn8pZcwXH
8uG7wo1JFtSG+qW/601i+yp4XQhPK/E1+LtNR4j0PzI7/YX3FcPyK+L5XyOxNs/BVc1/w2m9isq6
iqjltJIpu7o0k9GbgktddbSqeQh07ZCIZr2XHZKBAtecE0RhoPJoGfSlHsL5iIut+U58Q1CCbqlp
X6as5i6XjfuwI9Nmd2qMZS80ob/1tubJEWI4toSsfzsfLnHa7VgmO8mprXabOc4FcJaw1IGPD4Qw
xnGkumrmqr/jPzdH3suQGxu2HI+d9GNYPfk9XzW3/XIbDVw9w5jLUip4Y1RJCQlUguk7gKNTVtUc
gGvSH5xfz9bq4p0sr/K3dNjNiLjrvhtWoAdbA6lsl2OMEC8LYbuMWOI+WMjYlCW/hhswh7WO9sXo
hHzP+XVNpvykj5mrpNk9U6ztby3//rlrUKp9NiyDzs9HqfmK9+pFO/NGH+hEsJD2Q3v0179Uz/aM
0WniUJwLTYK+YFmnggvoSiOI7mt4Ecqgm1CoNBA496jFvqdtwnyCcfNnEUkFQbF26kqwHZci6VTI
CuUQrQF4ni+g0U2LtLZ5cH+hVjCH2U9QAxI0prgEeeUtYY7Wpfg+WxZsFTEgw4IQw5pOqWMUHYth
2JXYPQMczeBFaQehwPUxpWbousYYU1CoJil6K4N9C0VQoTjRofAKmT18jmP0TtlykdZP4ZEJT4Ws
9Y52hatWGDo7OZfYj7G/gLH6EH5ZmpQEAe/xM2h8/BndIw6XhPxopTxl8hUDl+9tMvtA7M/WXi6E
mbhAoi6TIlpZX8COgRsSr6pchTwsX9n73WjGnMrgqKvR2Z0JZ+bkECrDLFO0LN+9x4xMXjNwlM8V
xvgsxwhHZAcUoud1f/cY4lefI0uXUiRPXaJfJRClE+4JJ4Hn78i4lLDoy73x2CSgrK71zM4T4U2p
tN/TqYUkmqPjck8FLvNcGBMWfUtD67w8PZ8Lr+CpeBH8nWUdBFESC6z4UikFwX0DA3SO7WXYS7DL
aclTunMzqzXeo3QqQCW9jAaMG6ni3zEpJVKsqXFvJzYrDqA1etqNkDX1B7EK4O6gL0f0eq5qrmk4
Nbbi+akAi4BaEeYLt4TdnK56lBcsL8nqQZ6w+r4JoN5dhFA3k9AE7JYb3JqG/L2aiteJUeUai0sY
ucZxj9g59j+F+wvYb1wIEP7boJ6aCej6Lfrtw2lEfY8k9HRqJnIpLKtpHc4OKUlrI1U3r+xrKy+r
cUoLbylQ+gTFU0jLeIBxTYiqrH9mAjF6j9LFjXXd98xYzSd0Ml8uh2p2W0/Fdtqmyt6ZxQ5rNHi9
+lB5lzy49hf+YrfxQsHNIQ87m/vFCrSb+znHAn2CJyWAQBJrdZcmc5EWcxTL+7NolfBHD3hJOwCw
Lc4cvqR4VhHdHYSpUxOoEBsIHpIaFyuGlXAuK6qj4RU89UngPnd0uVrk88Nkjd7lU45166qwSSP2
081sjAz1f6YJsqQt6U8rZRYQC5Ngadzr43xk5GlG1N5hTLdBs4BPgLmp1MeTr1hfX1SvJ5Ef7TdQ
CL8l3nhSf9ozBo/hAxJy/yTeI+sigeGYZ6f/TnEMb4U6qWZmPe3v2MLO79jlBmVQUo/VdL0kb5wq
n/6bdgr2pLSZjIuB8WR9vnhTygQQecR8RJeap8hjwDaAbNX7PzN7Cv8Go2qmnqDZEvlk0ey0HG8t
lIie8kJPbLBnUfasoN9a9h78P/z8k/GmVRp0xOAUNDduopEHSzDA4ZaYdOnsBQpoVtMaNosZUiZl
UByz6RRUHlj76R79EJJNInBstiYW2u7yvgklvflk5FhWis6dM2HjDnU2Mew3AeJSx0IvDQ8e+L5l
SZSSUkHko0pH0mvg/zFwVeTkjdqXwjZtal3TP6HftZtw2MxWtSxq02U9VCkj5cLz2MpV+4APHvG1
RCtm1LwzJ6aBL6fwrKw21KWPRbnNRJtKv0Z3guZLfULBnsZ+OuA4abtrxBxIKcwWqEgNhCIJyPLi
D9Y5JaERged6feVFc2wpSojD4cKVUshFHW7bGV4FERE+To7+1TGG+9AUehTrfaawQ618lfDoY7K1
fhGT52DGn/LshSa5KMwU5xnr0v3hGN+btsTUdVDFEb1snoR2Bq+9uUqU+c3Z+gZJ0+PHZcEoMJFe
moUdQ3fUpP90r/tOzRNvHCMsKeJPCbnnzlhJiVmxSf2Cqiwv3prKkpw97TXPafln/VXRcNM8meDO
8R5WeUgWt4Ez3F1JmjjLwh81u2WfKwf7IPuudqWjdJYhfXR375WP4s4n2NjfeeuAXW3Pdz14gKAe
KHGIt3iNzkDHDtwE5apQ7TWmCwn2QnJhfq2Xbcy2uUGyonm0gq1mky/eaqQfVm2YtuDqWfJS4859
JutdafcxZoL57HywdkhVGcUWpTva/RA6vurPTIstfAYasHUyVOOGQN1rMmZAm8bqCQ9Ssq7DjY5i
yR63DQCrx0h4sNOrRDAWprmPui3DnWi2Qq2StF7hNRCV/+DROfxEVfn9jxXzPGV0yqxeJpfMdaW6
RG1XtkQxqfSdzGHKnHJTMs0gNf0A7ogshvb/SoUdMNJAz6nauYWmcFSYejGWgny8LxmJxX9B3lue
GRr2zrCwNyuqKR6Oxla6p7yvSQj5t2/u38fl4MNMSooPy7Soi16dIiPARoXo/zZHNE7+zKZm0wbo
dcCly4yAcADHncRWdM+g7r4fqtm+YBXf3etrDNesty4NvaTl68QIm6/on1S72IO1c8BF/X13R+cF
Vab4NrxAXt9Un8ydpM5lDvepDa2uf8jnJGXgyewjWsJDvVqrtM0usp38AjAuvOrzXIQSrBDGrfzk
/MxbMFF/A6eFjBvzJH53I0Q8OkgqTeOgI/2HorS1O4ByMYNKQb1LNr/nlJ79nsBwPmbICC37lccY
yFUlXt2FpHvwi6SznQHDzgpOR8zh738MgvftTJXJTZBoeQrJl7WRT3Hi7P95e1q1S89vDyJUc8EF
9IffkcStYXmRDMW+J9FLKWdB/NOtbVLPplzrJaq1oUXDlBzGu79aphScSXMORGTNice6BZitELFl
OqqA9xeiS14WobrycOmxLlwOn8YAYvwwCvyRCybJo/PPS8Wo0QbBUmZtdgX1Hqp2oyf5O33aguha
WHr9rF+1KxI26tQztIwP2UjYNkrrOMa7hgU2ozrrK3WeiUqnyqZ+jN46FjcohGQTyGGEIxb4wuIf
w4b22naNTVreRPcuFFHeIzP1HWoqdP9ECiKOKN4cUx6agbXm0owhIhvULtO8u1FvaZB+qqj3sgM1
LR+j+tqaZ+5lZv8J50HWiw5DPShjauF8gVRcyLK7Dam4Lm4wDxL9jRd7JtGsgwe6JoDhJwbV2aUv
pqvOwB3R8hPxn8vkBnLnutXEBsqobOjTfJs4XJFWwB8pUSssb0vppYkrAVHKeTe0ljE7D4r5EGwP
ifzn/NZVp99LuoCgsHl8WRWZBAdRGnyXGtwn1+RKRue4iu/Fgrx9H/jZcnoBuXT+ih47wTrZx2Ud
/mnyfa+KPe8Ayw2F56qrFs4itLoK/ol1gCFv2fZH2IS5eeshS1+qs6ICVdIy7hMmZHElMQROmAuU
uFb2hOvqqyb5tI0erlK0cqA6NFmbgITWDInVdztDMQ7GKd1j1MDZWINtsvVPbCCZdK43a9M40sc/
HJGbA9TC7UH4jrGjM29UnQiQXnnTOHAYQKBpt8V/7nfWVg5hR0vN7ERaIDVvz1AxBrV15rTLUv3F
fRpNyBHYeo9GTjbOKV4SGROqtYMGKy9ECRptYpgeWUnoIjTqBc5a2vnky1oz6DKRZ0BvQUpFuQW3
LbnyQhHkd3rQ3GFWPOJFO7PmSUIDozeTv2HP0464qVMsBhmgntg2zVVJMQMUbmFZEhw5kpk/x4ok
H/L6a4UUGWv/fIKKG4yTIpGqo6ounjoc6QsIVt76zW3GR/qyDYNXyCGyUiAwJwyszhtmjP8lQb7z
Dvkh+7YnnBT3hPQXi7UykD8CtBuQpJa1eLBpsIywzJ3dv/LDZA1NMIdcz1bgfyvr/TNeYknNC7o4
t9Hppjc0Ltx3qDorpq9STlGT0XwV8Iz0+wyNtbPv6K40pFyxfhWxenkxdYoQjPFwVG5/xC5kjpGK
q8hAJfrPzLUw/K79I52LBVRe4lZwbn5V1pLjNJfbtVP2dNuWR5Ip3UWCwgCfKxwL0c4eKoy0nBsB
HI2GYfDQr/E3+artKBHjVKem2/zLSDilRDLueYhXx5ddPl8263ja7UhkWoZi3gB/h698PR1WhbXD
c3AN4z+VCSXvjhHoEqdmFoZ6AHBpJh2n6oj8NONprElajmD+KBq7C/D/MOIDM+njbYTMlFv9n62K
Dznk53ld/GrzTBQIib5DZuAQI6sDLwETVbAMCTV2ilrEgMuNXrIVRrqZm53bBrag5WCAJdyUsMkv
zeZeoQlwHj2JOZB2w1hkvv5ZpPrlTPO4hG6fQkEFn2BieYxZTZJTy6sDxkMNzcOIVrR+gKFTlgh7
IBSd7oYJL3sebwTO6VHuMQr4Rv5xUqJtlrmESQfxyVAguCX7/YeX/c+Il65w+0Kye4betgbmnulE
BBttYgnMW8mdiR16TFH7rHrnUGSThyK/SwDAigCfmcjK7QZsBaNOUP4zUAScXSltxOhOcc2P/3cS
VKJJIw6kncTMAOqhIhFQCew+qd6vtHv0h60j90lnfluTL7dhzzVbswOEAnD0tjgrD4crT7yBBhvY
WxeG1KZ9NN+csqm60ecGFQ24E+BWtNxUpDytjVaZ4QzLKFS+PZMSN7jlnClO5sllFixE6jwGCRli
blwAn/9hTPUnFWxWZVeVCZoI3Sa3EKD6a0v9VnUZRLD4vzKKDDVa9FoNssSRL2QvvUyCDoXutfqG
8EHXS9shloJ4ztOPZoEd2Vqjx7JMpJBh30a/Ywmt7676yQNgaABK4p6e0UwA5RxL2yfSfwjIrkwh
17JUf9RqyrmVaXkagXxaRxjb+jlSt+xCNFaujfK3ejo500j5bZSgQElKxchysMOM2CzqZOQYzDN3
GrJdanstGMp6ISZwJYUwpf4pcZ2etwb6twbh9G3c+tfklbwYsPX9lvNS1upoJEP4iQ/fgXeeTqW5
tw1jynoAgxh5jUp5Sul5wf0TcH1z32Q8tpZ8g7GvrAt/x0U8shvzl1tV2c4PxTZ+64jQJ67BeUxZ
07suEBVe26Zlz4fQ0MF1mwrs1ZbwJr/18TMRBGwLGRlaotWBHk3viOCBV9ztQQQyG/vTK1+7fFV/
1d54Bw4PFjM3dtUngvkgDkGt8ZcrHc0x1YMHMGnRYV2X5OCTYxDQANDA9GRQYYW4CZll6+K4x6N7
Pa1X5t1AxBDvs3v5yZR5hOBHs93PrzB/heVotdTD5nuM4TzzwSsfCpuQS0BVklfigKtBgoSvizyj
2okJ0VNd1eO5ogMbwc0E4zb+QZErp/hyUPFsuWWJy8DqMIAXB49k+rqSkMds8S9rNKPGqChVBdp6
kEA87M/fBBKiQjqlD09ggfcSVMH/JovDR5jWIJ+clTNlYrjygKxBBSsLimRS8B2yP2N+yF+iHFTk
a2ZUpllDFIqo8UaP0YTCCCVh/R+W7rNvMGTTgqBuVBeG7PUi6WGnamxzWQ2MjKS4NkopibHazQIw
RxZR3kv0NB3OMTp/0Ksd9+wFqAPQZMYdO9BXRQkmyyEPhrfLzZuVMZIqBHI9846kRcyhhXdPowym
Q5254pmE7MBwtgUFLSj5pT3WTxsCsD0WfEqjrkrzSrvar0OWshdTkJnEv5L7zQ7vCDjoyUu5bepk
ByUbrPlv5T9OMgpO9vk2WAhEKhL/x5JGbKTj0kYrdmeEUTXzRehcUyVRy3oCICYQCMN9rzc4K8Lr
KGst53Rk0rLejAOqFHJShYxtouFblmUkazgqAPXs9Mf8NPpWpy/S+nPXVsAx14/op+9yCiqXp9wN
oghaZdqKIqXM/f6qUJk3okvpBAzV7Bd44TyjxGAn6SQlj/K5m2DpdBn6qEvb2lcVyMyhLnFK5s/k
vGooAvTZ1Lgp/rIuQnPLB3hPqctN5JHzNsxGkwuzFJTxXKkpVincrugjjxrEjCaVDnbl61O3935L
LPAslLEaxsWmCRNvEa6rOP14zCMKN72gKa6WX/37QhyzmI0zRVgznUIqP9y67C0dvaeCz3FuwvFi
+QGPz6wPjNe8dCEGZlOxpekFZD0z2z44x8VM/zZzPb7p9ilGG9K9Vkc/ajaCOApcVO6OR8Mkg3W0
QAF6mz7NHArPVUqLOtd1ICYU2IQ0tRerOpYRI3ef80ZwJuLCSnbGy804i5w99doE+zw6ePE9dvYs
r/Xxs9IFU0cTJ49yXKV7rIBoj734Ic2aJ41ttTHf95Rrv2JZxjc9phq3wEEJkuHY3BxMUtmHrN9B
sgIBPkJsBLd0vLfdADx+cM27Ge5BT/kVPCnIGNEpbdVTaf/D4kQl27xB8bV2PkxImX94G5fvLVhz
bJ245HBupKWkhEc6VSygxlKiZ62S+WzEdY7UTADsk0LPll/7sEWrmGlF0z8/bOvTR87S0igYKAhu
MPTXv/hC+xGJcfOSppIxiQPYNnwrVEPJ7nHyspHWeCPdVz8TzltdN5LhK8/XDYFM/XDVe9CRNf0C
4upzuHWpQYaXcWjEg42YXVCCBxHR549GeEFHEfUOFN9lhgxVU9ucRqls7qOjqZbdTyV+vz1h1tNI
hXxBIUZnUhzcKtUct/8we8lJKPHs+PsdnXziLUCiAt06kWamg42//rUbZb7HwvxeMDOy3ElqAWxa
F6/xUpaWVk5FORXISMqcelJLPPRf54G8YpdKwH9CZFs/h4OJ9Wv5mV1oPd9rPKE7APVK21M6vvK1
Tb0EP7XBOw+3Sdh4rx2/pHYYVplGWg9Plxj3WdpRuavJct28nM48tMt7eH4RixLdfLmEeFyboT7J
cxD8OFgDH9toazrxbYdlzpf2Uj47g7pWlsbzEGMxb1ZpvZ7loeFTyj2SObU+FLBWzWEaoZHLsfVU
b2Nv1P2QeSG62so93/2lFokZFn3jKeqd491kcDThU2XQzzWvR67bNgQdNfESsli0xCsNYOJA0NGI
IDbv8LjJ7KASEbptMND12GnvaXiHNlb1qSUx28lACUfBzfqOJzM3CyhCqbZgD6MEdJlrdh/Mh5LW
TYH6YeVDGIwG5J6gpE3aUEQRptaetjK7iOOTbwRsSE18B5LZQbnSzImafZTKCfPUti0a5R+EW6Dp
bzEk2I8mBNNZaVzMdRN/nFEgbABeSV9KtMhVyJ3uSAj+cLjXHoKj115mAF7tW56h2WzTQzEgzXr+
C8nCecTB/5hnT57LQpA6dAb7DwfaB9Ha2z3jT3cnu4uNDisPGPSY9svn41jFCYJjcqAztEKjaB2j
BhbSilNf3pnUPHPOWooYmWrZ7F7PPOLGSngQsGtuvNM/dYBq/HAtaR60YTwveVlTrIjKubEe1SMC
ZsHgvzYXJBDIF51SR9JJ3cEyRKVwlYKeMhA0e0u9ncTVCKjUN+0v7zcyg+OC1GdhQcwt14L7q/2H
PgqK9Qc4ITZE3p4StYf6PMKZuV4ox2KgI9ieCLUUKXdBgGhm2EHvhg990TuR2/KZ8LOFIPN5WERl
n+z3kcwrpVAAK1PdzVYlqylHjjlR32vUHQd0zMacrbKw6FDydCRNtXb2m7Ebvb0DAd7MRSbx3hMH
cWU4k1x61ph8MLffBeJxS/GisDIJOk4l2PldT+YX44EclE3NAWOvqBt6bgpEOZ8Vl9mT6ZsJm0QQ
O3M8OMjjGvwAyag9/Wx2jfkb5sJZnR92Tg1G/E6gAnH6fHzWUxJLq4ROuiNh0XJOOwTF0zk28mJb
W17uBhois8/Z6s/TGn33dD54gbJXP0tPTuqHVzN/ItUBHVMhM7t2wWToToKBI24jEAPbHZkntCIL
vI13jkYMlNhNCmxUGnJfmxpEtVSUT40qEKqL87kdFLWMd4vB0W7wATiSvMh+Bx5jePYhwPawfu/f
GV5tliLqOSb33VXRcC7siuPHiqNHwuevU28b4A0b/Go9VsXGCm1RsHgUVoOnLT2402292tLHyI52
xrauiPain8H3qrlBCu1avLjeY8mRX0cy1FO8bEXBreYBkWk9nKc/N0eDzIQ04uBdlp2+Rsja+5GM
YrmKZf6ITxg4FcnqPsZmcO2bF7uJuJcEFr7lH9Dv5Kz/3vxIgtJDixGmZhakttT4ptsKoIItMVXn
eaQjJxN/iQaeG2AUsjvCOebs88LOpFjLDkcQmk4ZGmiamRFE0Br1P49zoxeSiRow0IIVQM53CK1t
7T87WHRWcUzPc9iZ2rvvieqv2fpfwlgknPcqBWphcaujDw66s7wnhKsjyy1DkAuxvuQ3cE/1aS4j
Syk4lNTsA00kbWTOL9DocJqOGuLDZt70Rli5ZP7YOSK1FX+IOZMrHYjzt3At/fqT8Siwn7DPVc+Y
ENlWNEGCwieg1TK9m8L8dpuWAVHYzbygLABWPrz09Uv4LWKbJYYuc4V3gYue1NNBrbOFaA23D9yp
78/IVs9CBQls2g+mAjpzsglfq/OGnVw38brwjm0yVZrYGzriyYdNQdsg64vtDX7QNFNRWksaSc0T
+x90Qi0q3PuLYTGO6eLKF8m+0uS8m0mosisS+ZoB3Vc/OwkMYdhw7wZtk8rXJHr8hXDJn/nqLqkI
undndZEYWV/mwserH+JibUGNMdEwBbLlP0gKnw1xe1Fy6jptY2n8T/MxH2VcZ+RsJHFRUcrp7rHo
DRkOlBm62T8y7xshOdn6+A/1Oi0Bn4+xekOdXOltyXx6NSVIM+4d2QylqTYihXuvzHf8gR3q4DmJ
EM5LZ3TfKLUrRR5WejOKaTa5C0vu1LrSA5LwRPMIDJ1Yp955qTXK6aSTxGve+KycBUgX8VoUtO2X
20T3Tb6NJ6FWYMOMEOlnWZPpcp39LZdOAzancQAAoy6nONSQENyGFlFEmUDb3knVsOr9l1WzwYVu
RWNjiFidTuXUeDA2vRtwhqR0T+98ZBz5HoieV1ArRDFO5fqID/ayifXwRkQ7T+uFd69pqxKAF2kD
D9P6WHTH8OO/tGvjEGrnfbHfmyzOm6oZUNb2q/9JFjLN7bk7vBTGRuFkB1ngcVwQdJcc8dakJQGB
+UOovT6mBmH1FzGXSjQ9IRKkXKjrzB5Fh7nN4+8LuFdYwUo9TF/WMYuDF5fggGDiacw+NQpoIlCZ
WtcS8nzcvjWDXzIMX18L+RQtk84wTn2aylykNQWDLURshXwRfYh8/13HPf+irUiOyxZQQpiAK8SO
NYS3UknyDejDJd21U7BXw9OxgbskggFzAlp0bFotxIRIG7h0Ctl4S0YzPm4jLzNU8SXq4UOjF8ef
HRdCd8lE1du/WXO0XCERhxNW4Qj1A+yuxlvR6GNfLKdyXV667nUexehMk4GmxIu4SErz2U2GkEVv
e3nt93WhK7Mqkhc4ZY4Xhh8j2OFtMI2B8PNyCsMYZe8Q7f1uy2wuj4+qbsk9AK1PFgfo2YpgnMGF
44/hhkjaP4vQ1EPkEmi5VD/E55bOGmFl7niu4QslPs9EsXTSnh9G0RV5R5pWT776CeEciSZitJgK
hIGN2pFv8nlGrYNi8c91h4Ua6NgRacyI43a6vIG/c8fZD+mwMfYy8RTKu5fO6leigKcKk0N8NiX/
RHlNB68A4xnFf2u1UMEj8geXIsUW66juTPpVIXfh1M23D0FTefS6zb1/wv6RsjSITSsPPFTOkYKo
JX7I4yGuDr1FcYWIfpp9Atyx/RTEmKcxBt8lIWzQP9WJX+wW3Cp0UP9BgOgWK79S2tCyX110PwXh
Wro5R2kzeJnHHJIjkn+UNMFkuFBA5GVvRRU81fR79JrGvHNM1OC+r4tj/s/sdkIOY4BRQA9Gn6A4
pAFng5843i9qbycsxoMam/Sls2Wa1cwc0ndROjRn3Odvginzd4l+zfNE12qFKbi6EZahsR042zMp
tC5OcARy5hKI8GuUSNhCeXYTdCaROXBuDNuPEBbZUFQtMEzN1Sfqsu6TdMlXeYhmmNge3PstpSHu
sLfKDSMzwFqP20dgmFY3DBiBUDDm+ULs3Uk/NBgo+AsHauKxdbhUUDsVBVLntcdquM4E0weZOFt5
q7751YIj065qnpXNpk6ZFAlqkJY0t1Kmdm9eJEgTrH9QesQ3dinDt2LeQtIWiWmpiO69MhfkxyXD
uy+fpRJDvEbUlOpxQZrJPicTklsarTvfWV/M5c6s1bJiPkgy2/goUGydxnk4m88fJQt/xRtV7G16
z8oonUfMVomxwFgQfiqpZjjSTCdz9Dsk4Bi6t9wXVa2CIQPzacp7N8+qy1fb/ES6Pa+SB+bgZQKS
v/Jfdlcsl/2WnVn9aaHfJmIVETXkGTt9l/U5R4kyT25cfktUXwaW4NA3Hi6y5uEkFmV9wwSySnG9
yZP8r7G7s4jNWCDoAEy76uWyjGEHvsnSfpvc/DDo3rVP1akQP8mwNo9KakUefrNfFRzVp8H9c9BK
r9HGfSitT4b8LX73T1RzpDU5dNt+4W2TRmhTVhV5SYTy6cfOWEPsMnyFkQ1dIqJ8QjpPAyJAL9In
xjNsVzdp5kkVz49PhJB4ck//6+/hV0L5vxsXkgXlYMajluWE0PNvxiHdA/S7hJGUUBoxNJbmleVt
IrTMJVBBulV/F7HNBf3krIvI7FolyI90/l3Dm6IVRfea0FYVkiEnBxfANvht5EZG5xCEtdkIDYJr
kmDe7gJ675Hp5T+bOsZpzBNbijn0aLcUqZqZEvml+Pg8iYDv4FGnHRKmKKD3dRpfwNasFNNx2yIn
7iY1UgwtRFbFlYAu2plHjgC62BEM/SMfKaZBQa6+WgmxmK3e0kOzgI1m5NYjzeLXyUBoFe4lVAWS
zptrpg0EPLJaNJRs3qgP58ga3GmKerFIHu0RwTZwc2L848F2v85g184xKt+w+6dmJ7mg2WNOXEdK
1yKaDefoK3Ij4jX5IIA6gPoiVYXorlvd2w9mUOxW6ngSbn5ybOyRNkxQMuCV4m+X5kmHrTbloCII
wiaTW9dx51huoScl76RqDwhqtGPGaEqWmNYz1IUyuUAZUxHDQk1Sb8KE+wv5tEoLYi37gcofZAbF
p9VE8avO+YCZQ4S3+HZktFR4sW/Ne6ODPlV4/GvhZ7FpCK1+ZfJ0r//mprEVkxSjT9CTfONQJ7LZ
h1evtr61Zebff6O+yYoe3pE2H6Gieajw+BbB1m8+h6Huo6Z/RnJkxeRWXUdqYknaI7PqCpGtKfv/
660S/UXE9p+DNbGLxc2CK5YqHByPYzM6FCkfs11WX5k6fePdW4rfhUW827oSt8J6KUDeQh7yUyU5
ZWQjS/Z5pZs20+VusC3WmOlPUHjgf6XFkaQ99XfGASfCjMITedcq2G1x6LFDf6C2rOUv0FdzgaR9
VZdDxYsZJg6ZClxDCEGTb/cYDaj6sx43+iRUGP1duyDWENgOyLUr26iARSee0f/kKVgUpjLQOjGf
HtT7RPbtThNEp9k0yAobI0Anm+9EGRBwzMsfWlTkxZqgP1+2jyzxk+t82JyuUjPsG9Erbz0xIwkt
9iidRvUeZ2vy+rZl8RWJfKPzCs60BWH98UVBt3QlyStthPX6rqiJn8DaOs6FdaumELR8meUgH7cY
qy0KjoVbnoSjONjzodLA1xAuvvQrx+yiZrO0gnLnXQXtNhCgYBPoGdXe6zuPbcB3S8arya2PEAuV
sc+gmyMqONhHqsb+HgvfgP6MqfKszm/Tk/YTQ48TCPzp28SBfWuapEddHa69B1pS6rDlT8Yr3SBj
NbulVtxYD1COypHG3ta/IhbHz9H7VbK7F3Rb24jweSg18YLwr+ZydHxgZCP+IHsMYrWjVEIiBtse
ftsLk3L44XfFvH/00sKjeHYSY8dAzDj+bARAkwS4ep+ueH4Td1O0endwRaaBV9Os7omCP0cTXagp
4BZOWX71F6GoJMQLSpK6jRzc5lx8vboMtKRA5gF4x3w3j3YnsxdtVuKkEAV/RLhAG5VDH/az/cJ3
HH64QpjPBl7lYOAlbWjd+hXdJzHeLwU4HEIx0xiHkWxw7OfoMt8+3j8zKBz6CvVZ3ofSSr/qZcQE
wQ9Rmp9CjF+xdm1bXKQaiaAe8tI/Ymco6bmw8pjKSHFTTld0wM2BpnXVBWfQI0oOEXgsJCsFJN/l
fys5cctEigEzWwJyzNYpz7xup4mqIgYfMLUnCNY53YPcuP5GbIfnOtwgP8uABN/PdrOAGkKRLszQ
L43SfVr0jNJ0HfbG0Kcj13xwKp3oz+WadnPtT7pGiiLRJKYWquc77p+ibS8P79bL4v4bXgGe+ZWv
J0NaTM7msCP7blAN+4Y/cgUj+H2TOM4daHmJbyU0UvoX7a5MjQXYHYnsr2AxmxRVzaK/R4A/qpEh
F91v3CG6kQJ6djHNB+y3yM8NrNMc4FaWFAQyDwX3ICtU/JQH38CSMBRj8XGCXdyZINPCarRRDBGU
yjp1T+aL7gQn9BB20srNTKZd4EvpDHi+pVe9/v6HNRdoLBxOb3kziy1hFq+nePy1p6SiVdlF+7iq
4EY/RwVTo8hYkU+6LmakmUmmC+/cu+czvhFKV4mJjvl7s9vzxD8zGPJaMzsEf/FdPUFOgD4Hlf4E
XN2iWCeaK+vrY1wdQjqdzBqsRRyhJ2gDuDeXhPe6NNxKB91CkQw4ziRdnvVMQqL96Q6OyxpSi1ee
246Y19NKfW87IFBiWtTFBZuxDuKHIPrD5y0uE9zpHIZQ995z46GubMr/UgBBChcV86dOyczPIlxC
eSPshXwnDUGCocmEt/LErmLQVA2rsJp8PqF1rZ6oEmx21XKji7+GolzbNTOW8Thw67Cz/EJ1//vc
X91A+HNuVjn0DK739XJ2XqxjR+hLvRk7DMOguyVAR4p2bVfL/h6+GPFm+Gd5eeK7ShyunX3P7qWq
kGW9RAG2QKjPaoFFYPSKQGObyvz1Rdl44vof0sKmvIbVsy1xPcw5hslywLPWMfZFABuhk2EhSUdi
vnKH2SBMix5hCzaCZ7EpnHnqJx3fS3EAhjuk4jmlPEePVZdiPR/g68V0z4B/G4cEUOsd3Pw0MJ7y
RkbX7XzZC2q2qWkrHU0ePdHRp13OSIFt5CUl5p45kwWL5HvhvfZhs5q+nAF5k7UnPsnr9J+yCNRY
mHVP8KT7+2jQP4Lp8npDP1o5AkAM3tPWQfVQMQyFyY4TquKjCgIak5UCCbNNTCKfaK1eCtYAQXZo
K34KkOhW4bSNCTKsbmPtNyAuCjXvL5ObD0U5SfKXPw7imSxM3xfDZ5WZt3xDDG+GqMRT+/j0cezN
actvWtTLsYMvRbwLb0SWl5ej4RFa8ObKxWp+Fi62NP5FyFyzplViDjeI3rkeiYEAg0+ohpcAfeUw
fqxrTg7XIpKe+wZ3WtudyUanqEBSUDVXRp3WJByg45gNcBP8KbhMWFXP/Loj5IhGRAOceQGNyuP6
LtJTaXZa1MwEdGiFELQ4EJLFJ+am+Z9PaAgPShBjobWK4aP+kAkmlq9EgNbWq7qhOcriIQ/S113y
W5yVSuQXy++cIsRZueoAR15ys2RCBMIvAD9rafvtD10SBr4EqtdmLS7E/wO68t5KG+mV8/wq14nO
lOqAyrVM2XuZ+BOPCau4WEjkQpIKD6ludwKorEEY7s72WWdFiiWPupSZfJ+lpfyvsGdX1AoyJRdc
wfzQi4JsjxgM6vZrhaZNsa1wfSbymKSMv/bc1maulbdRjuuSt5cEQK5WcG2E4BtAqOznLVIs88gE
YNCsYpnR+jhuN4kEKQKdEsOR4+i2PkJsFJXnaCq91jjBWjtvT5HRGDyFq1BXMYEu1ncaR9PJJmuv
p+dqe0YvbmJxHrpD4sEOsVEdbVT8TK5+SFWLIikqV8eExe9fBnJKFXshiBy88h9TkyTJgxBoyc9I
r3oEokq1qpO170Hwd+VRvBO5W6U2Ija/4U94xPQd4tfsofUc7qyJgsLillK8ZiqX5noI5Ht5mygs
r9lrwuI17GqT5Qg3hENEClna+ZGF6FAFY/Rjd6LfYvivt+VTxEPpL4EA06LUoumynxRtiv7gtK5U
rFdwIVPbzTEPm9odTBqwQ2RmTSNj+r3/W3XjMC3Vefdv9t4bWzNidWULHV21Vfl016cmCge38QXd
Kq6rwEh9U645hBPJ0fh5GeOyW/uA0+7rzD97STxaLAPWn5a5bC6rUr4BfXxsJC0U9m8YU3iXPNrZ
0x/zS736ReUH7ofgFi1QG4DHOQa+Xy8HkdVta9OI19P8+dJRSsjbX2fqj/qHgGUzq85GgsCekNhg
UwRm/sJMcGKcM/NVgrWK8AwxQBcLVDVk07CX1frk8yC/0XHn0kPfTZxDZyJ/QxwCrV+nYYkUSfzD
nbH4KfGIERNpcyM0EafRZpQUQqslsJUMRUG6KT8vcmyCn0E7TtJJJ8bm16PoWJhte5aIfZphf4dV
nLGY4Or94CWvmew2xiqRPjZP0eHhcfoBWwq/GY4v1dCniDzW3De4NMRSPX/v78rgOqHf8L+7TIrk
Yg4VUK3XZDyxg3FsSIuWunmSLCVkFaytQWrZWbyLvelwRXB3KEXNyjapL8C6PDpheKyiVL05RDAO
4sLt2poPL9eu+/j3DfpGhNpQESe0lSULZnuGNlzqDnFvs4zGzIXzoJWSslYx53Xp2x3mWznxgaxt
9rzlSfGLm0zLd1Xdh331kXMZ6dbr6Q+z0Xbpwgv6pGBKasVdvMLHgSRnA03/Gv5fXQpLMuGV/ups
UzEnKnLWQrQ+i3Mki3vD2Kz+VesdadvZX7gBg7D2Zr4t6dvtCWHCLU4QbVOYqoYuUTM6cJbcG/uz
NfuBxPzapeI+6a0i5uAKgeTIFKgn5HtC0htrpjjZ1jJvRRUXw56r/6AcigGFcXhN1H6Y31fErbi7
g2dxipO77gmviWFgqGabPDV8WtDyn1KvnTK0Dk3Q93Dz0qOLR+vXhVyPrZn8Rn0gfcuWF4G+0FUS
iPutRtOJeoHFANLizb2aRh5bVFOok2Zmap1sROCBt+rBoG0jNSA55uf10Qa8h9VRTaD/qDCT72k8
DT9fPHYXLRyga+S3S8TKR0LJmbq0kqe4LH15xRBkm5V2PfLEVopBLV4/esUXVgSmx90A3ZohzlCi
CKktlvVqDdvzgYi98lUrMUBT3vyEsbaHTFqu6qCHInj1qY8ag7FfFYDj4eXKjrEJFuxjEFfLyEHJ
pMhDuTJIe1aq8QR0Tmmfx+2K5PfIJ9vhsMJavg8ouGqCBHwWIh3V1XgOL5E51hQpQZSKww6wTE9r
Ff0XFIBEFP4mH0dWewPyhPtdQAAZ1u7LqsBRtZf+G8xJRf22oo9FeRnCZ9FX0RlywONaMCN/INDN
y6YKKme6NnyIIgapL/MF0118XG44uvwfdUBnQsPrIrt0sisXb2KA4zwRuYOfzlbHYnQJ6MiJ/075
JzWmOab8oPRRakinoXEXRWV9M5GQdPSCnXCOl+rC6gY0cs5jlYqKxNXjCp0pgESjRa7czXp57CRs
h+xbjzWqqV09mhNfQu7UiQNH/8Dr2hn34MF4PUg6ZINUxOJ4TjmHFGx6RgqRYVsta0q38/msalzm
0OkxoUo/fzJho/b5j/jvkMRT2oVC41VPW7AGpFNJwqnBA1TMB14N5Eo/VS3Bcp/NjnYgw4d73WKn
8FitJGEnP7OIAZZAV9rkSvhNBh6tOGVOemhRQNK792uJwg1b0mi2+dAFHxbQ0SSAIiwKX5VGz4uS
rQO6yS73LM7E26EtXQZmvlj88WYzBHWNP/6OnQp+hlk88Z03WgZuaQML0JaPjtXzUyrHWbnqc1Mc
1wyAG/u+XrQhOr1ljZBd1mZHULzj/K3dkNSDmdPlNitJgfXmzwrrAoEpyZv+gCgLapzcikKLJJv/
bkC4JBfBgQQ17ybN/MjxC4HuqfTjXZOrimXvWQQuBHJDM1tXh36QhgXHNHkbLYfCzNpj/pR6T5WA
bbR3BUy+Uk8d3kGvocR8+G/bJgDjDxnuL41Duf6Wvb02lnxPPLNrGqm+E5x3G+Ck2jtHUqjhbGOh
4phptsewCOUzpSQkuGlli6g1ipvXzVY3ilr2UOHav076Ph2wZdregPGGc+rYuyP+q5DxxEIaK0Bd
0fPM+LCRSn4l2zJq+DQf7SvS5C6gGRf1gnag/2pPxwi5hYe1OTQN1UI7co7DOuqF8qUdgBE3hi5T
mz1cGhDO7x2lAuPbvcvfBEXJcISEJOUoigZuFV9WtYIWPa6OxNVlWk7tqaxHsMrgvD50PXPYIJJz
SnOmUtv3ZHf2mEg4R9doS9Gpww0o74d6TP/PWzU9Tsz4ilmJOQY6C7NCe1/Az2NwhIUij0P7aD3S
zguB495E1Q3h0z/rZP9rIYDYcgMMxwfPX+e3ITpoSPChQ2dycZS1l+H4XY95P11RMl4LAfdJHOs6
KX9VUy88P85tNVOj4BZPDwjLkbU0PQtg6MLwm42nSn5vAy/RH68yJPBHwuKeBeGOBxVboW81QP0+
1LtTC2u030nCLgreXarJQr3uAOQisJzyd5NGfUVbA8FpTuDjF5SMAbNm2GX1BUJmMXZNH9ETZHT6
r92GA4o0gucnkUI9iDyAi3BobT6+VB9N5soNR7F5Cz1TbAAbEBi/lqXnxeYCEY0FzEWTpD5Xy9Ox
IgN2/JOh9qgzZUrp8/MMkqHxE8k6OnBMXUIBU3vB59zjsPMi12vDSCYCqPaWqwOA+l7PKcn4de5H
dUImIoRQE4JW8BGQb690gJxblnZ+XfcDTgB9l4ABK5aE40nRGoYt1CH5/JMoqrHsglAZzbzbq0ge
HG3LByafD0mOAxNyOwHPg18Cp95MXIwQElw2b0UG4yGg4PfPxsDy/zbiOBNMwjGD7CTeqZ7PZxCG
3mV18u/K1V/v/gOAm7sgHeA7SG6HhbbQ6C7HSNOBowNnzKh0sjPufceoOsrtFRT46R7ZMxJ8BymN
zGGq352hG4ppW0llXk5j5V0rEevUuA3Bcn59OgkLSdNzGK3bu0YOuMWCgR7U4bLKOLqtwoj+Rf8R
s9FIi6Xpnujpkxrj7359o/Fp8Gimdewy+WokwMOKWG8T3Gg5uLDjAdQOEdrt7RWGOPa9fy1L5M17
7wGaA6+EblnxXjkZ8v9cbzcLLFqsU5vXkxB3IP1P3WIn4EAEz+YN5DqvTHFxOySHSnoAY8zEiG/f
VdhErnQyOzwFfUt25lMRp/4jULrlksGszxgPMUYdYz8wNbSqNrTbK5AMVU2jRakWerjsV9mPxbsz
CQKtBZfogkLjDDIAfSkRugjBxbLfekWbo+Ize/onuti3s3QN4Eu4Yx1/qZHeSkZoXPzxmU11dUaX
rbRajS6Z3/3mTd7L5YQgbcpP7XoHR8lg6AXhDBBXq7qORPAOgQtIbpba92KXXi5GSY1ody9n6XnV
lInX6juDzdEkH7E896AKCwF+IS3V5NcmQh0/fBFPijL6z99zZVW4uNL+YbcODKtCsqBm4weaSwWr
S6qW8ydPxkpDUgB0R0BfcPuzSznUHsSmnkXoTkVVD74k3VtkM3ShM3fdQaTONxMqjMGjKNZVI1iI
Rhu3iY2SYoYrU/QXfn4pAH16J4UdwxDEf8Nj38bQE3umi+YfqJWlbsRDgmAWY/7Tgl8/GEWa5QzX
99xtEhtfw1+axz+WOwOrvKX+29kP1wx2sh7bjWWMOwKiOJzFtbhU5JBcuihkl/veau6ygMyZHfQu
9xpaIC4iTD6VsdfQCcd1y7YBduu9n7bEL43YZcgR8tKiaOPCCxSl+UUg64KlVQUCE/p+buOdyAlx
MQTW/qRj0RYQPyzq4UdxRznmCb3MAvxj/o9t4+d5uZsSNZrKrAEe3ievYWe6JhapWEUYn4tepRga
itQGVK37fYiJl0MxfnQGb1uw30uZ/Dy2Iuqoxw267gsdbyWSdMH+CRlDBL+PazMb4CHBOxE+ijjR
kUu8rGnHi1Xo3r1rGU5km0H1LKaCPDP3mDm4+paR/EWEHNEIKnAy42CnzEi8/OipfEBdxH1DKUBU
TVvrxYHOmfpS5sen/g0czMbyG8oWGsyIcmdHbgzqRoArRBl7pS+PQoJ50dGS/3ElmHIcGjl+QWAl
pNlwfd0knMb3GmYtUhiWJYNy+KOyxbOmkkmjXabE8o2DvVdRkBKJpEhlMtH+MMf5hvCwUbMfCnCG
Ki8ZHo6PJDQ90vMgC5ORjouISd/u25cN/jQKqmA/kfsCH6eZFm8knMdCdOl4mlhg5ASK1YaNn2Ux
imLCNUmlHUrWWoneNwP2w+QVhqTUFWxt9UJRKTaoRHMKk9vFTKfHf+KDk3aqZjmh2GP7HRzi+L9c
rRY9LOBDPWkqR8LkwKx4pbdr6AhuGtbamY5hINFmN3RhlGcnN5aldm4j5QH5vL1j06Ns65D3MXkp
JD63MVv1vxcYBuWcctzpCqvkhTAYAWo6ku1gXSGZgtgjWfWOL4zjS+Wz0kE/2Wxemtwg5dQupOog
doEvLPIopSLburSL5GdY0a1qmZbyj4dGZHp5f3nzZQoVSET73FZh2RgXqrDYjNth7dQbunc+e7uF
0rTQ86alvIkb32w7Qi6ldHjop5sUkBsj4IAfIdT7EzKoy0xBFU9ePOJvk0BmkrCzwqXyu3Spc+20
NtB1kwSx1K4NUzI32UFjVZK1BbdPgyu3DNEWsEVlMHO/n0+1SLMh52MaBQ+9KTBgK1+yc34Vau6B
hj1WbCUIx1QFU3QAXZDgBUZwTSQkPfmlfpFJWFcPXCbjPEJTw3+r4RdCWkN/fhqTdwDNVb5oBJxe
ZPhdV4aPKlezPajPydcpsMSphrNfdarGgXoJxszqCn5AgjtxYbmpmu+H6MvEfF6qeemny4Y/ukcF
dwVntwhy5Gc2SZOKqjiulAiRGw+BHqNLqnRpaQez9Eo9/k3zf3lkSwLoZvhRq71B85KHXxt4OIoV
EpAV1oio7RnYvN/Y94nftb24HlyIlfDFec/N44yyGVE+Cy2jXEc93+SbEomYy5sWarvRIM9By8K0
5cLTjYQuhaYerJ00kUmjUCniH6FTb6nVW9M/0WQa/T6/WbtPJNfpuTKx3pLXsh+91bLjvIMYYg2g
mwYn7yGytCIqaxpqJJ0hCy97LJhEBmtkCSknJic4UfuhfspWPINQ2oyAiaD4VPNiVFlczA4klLTp
NJTfr9X++Qw6x3ezLb1ts2VY2V9sxaIIuz6I2phNJ8EDOM+d/akrMfVkYjFKtVhiFFhLdljy3XJA
sq2SLaRlXgG5VaLoIR19h5h6YQeZ1YFlXbbfFx7arZBoE5vBV0h+zQ/+bYozQudHJy+/gOmCzSy+
ZrWZzfUrUiZRGAh6Muz0th8kSR4J3eAmlTLY09rwQwErgUNKoE5pdOXYESxyUDHz0UdL6qYKSagS
+YCSTW3UoVlbyYxaXKU6mIup2lqZrCOfJ7+pFGPQXdMpmdKHp1OEcJw9QIRoNAjcq4X/hs+eUeTX
l5Z87AI4WyyRU8ULM4BmaoFV8gG5cKuA/nVxV2WuM1GvvezL0LD3HSh4FlP6Vk3fXSz/Pnf3FHyw
ZjEBiJnnpiGb4rP18WH8hZyz6OmEZHW3hCb0dB4vZMD222OB7kl7U/uGQJ0lapxZvkuu0MwQaSb0
DT8EY5vkfT9i/rVmgfWk8l7uU0wYG2Uh5NT+XUrdaCRgl2daSL/wnvycGf5/GhobMz5YcMmflFQm
D1KfoQ8H8HLvTd3jc9C1akn3fSU3eBchra7IIYNPFR5HYvyAROmgQMxUESO5rRn5B4jsEGZMeCtI
pEfR5L41rSlmIRL1uBAR8RqFbRl+/0wlgQYnfGsA525s9rAgxu4q6imFe1VH9THtHUFYWBXGE0Iv
refOHmpKIovxkrRkpMlYnXuvKbzqHzg8x9pkRAmosQuzLIlWp4hmXdOwimetO/7cezDfRi78b/wH
fGjQoDFvMc5OmLV3E9eOup0OLpas26Ms1IAJbLX6fn/XMu8u+q7g3puvk7DDP3ERxCaJlR6QY+1E
jHPiTkvg9njF+WfV+1q/mUH/mUYrS3/BOXw7U0JN8eQZjgTgcJOzNSwZVyZCfwVXzocBvm25ScnS
WzieE2+DPaBvfObjcmOBpz9GxqzNmOjcGhPGyKG+Qhp56Dxri2Ki05P/4U9KdntZ1jP8aMdw2n6G
BJ0k7Z8irZZ+xh4C2E/CaYXdy23xmCJLD6YlDn2sZr5BAOICtouW4cJ17Qob2nj34RVZFOBFpG/w
BztTGjJRdwwkKO/dfNPfojHVuABHPpMp/00GMWNvebCbcmjMbWFzt7OtylL/q60PxlUP0f2Uz+2B
ypc2lx7T6xu7kIom55MZ7MuUgl2M3ksztg4QesaG/817cCVKFi72oRhXWcnLFEpHs+quySi3CGy8
eOrXqSLMv4iNMZFo5jwVl7nLg7PmXujalzBMg3nFl9VqG00eM2a6Ykgc1StUdjk/JK+vnDCHCP2T
WMS4H5AXrseG2FwWuDTz55bLLiC0/J8eEI/bXLIB8QP2sYBNc8UI2uyK0/QKhhyx9psTkM4BV6sr
nCzfGUpZgJfgP+EvcGM32nyti7okkO/eVrkVj0x2mVc5Z0G8CRFr8/ZpYPjZZvQ4hN1FwAxPgytJ
WG+Bs/6PtFUNcdxqLOgwgVoXsvTurS9RiFieWbAwUZg4hE7jHAEqD0T5Ua3rWlcxWqBHKqK6pAqh
KEyPzo4ubCvy7hMf/Kru+HIbTo9P7yTCJS9AqG1pJwYkkOcFnpLuFeDwwzheZacxU9Dw/nJdK2PQ
IopnZ3MBVBy2EY7U0Eiy/WFdP90YfvJzMOk03oweT/SEBhINb72BBhHmLWobRfSqnBXWYiSzYoGq
hWhRHGpJCcZ1WK0mZJnRO75iJiLYcA4xKTm+j+l0XnQ7tyIg5VT6ACtSJF2OTfo2QWqOEOmsof3g
/O+LWQv39kwFRqUTb6MbnR8OqEV3zcs+YwzQh25HZzmIQRNk4DrSbuuRL/b1aupnQWwCA1CC4hyd
fsNotcrfTwVtQJKDi3iaxHB8ZlAAgRScWbpocFUMBemfjOjyfe0d+ygLsJlslYGysovxFvvtVYEM
hLWREAGbe+bgvDsg9end9Y1iocIfiHodbvyyZ7X8J5nROmj7LIoysxQEEkbTYj3O2db1mDLLNz3s
nJ8vcvkLvazJ4jZtYx1tIsNxi6tJ2G4wFV0JnrcIpGAFaUbV8y0/KR1vealXlsAsZ4ef77iw0BIc
sGCvMVUYAn+jaE0GCl4E8VSsiKD3F5/5WoR30c4Cf5D2vuWS0lzkImcwPp8L34PnAhSufD88tKCu
E2gN4S66zNQdXUisznU4bE6iqWcyVshZ7o8LZqhC8OFAAFbTMPjTgS18z7Oin+TgB1LsySglitVC
3zAqBh73/WMgf4nsK2Dys7geZR8dtm4gPs2XspJ+U1y9TZu1lAVECqrrsT1lxp+tP1E+qq96vYL8
i2JACgpk12zeDOBkVe6iaEVNiW/JFAoJaRHfHn8YBPeNZFI2pTrPGaWSrEqgKrQ7DRlV7NtwyIop
K1ijAgaauMHJJZoIsyzZ7q1GvbvGwViURbBK91FpLAPpNpO1j56uNBteVYAldCA/+ih17djfRJ0Y
8Ox7ODjDNt5Yqpm/HalkrH4duSTwIZrq34Q9HP8TVBNZsPZKnk022xvFdc5INC/PPj1U0qevhB7W
rSqp7BpG9t6bXiGswCk5NFJm8SmdVhJsC9R9fpEa4riUeQGNxyveE8eJ3tH0/iLHrRyY4ZjFglMq
hjsj0gzZseOQ0q23vRV3oFBbCuEdYcmfSP+lsb04D8JgtRW7MkCykrV+TY1i3uEBb9qq03sIcEKf
ek0eekyMf8W0H2h3wFRrh7in+LsUq3ttNNTb+g44NJyDxx2vNbEx3iyfEXQDiVBqzD2uFudS2kbT
0p8MbCnQMHaEWRD21GZmwE7VsuHJs0ZferokM/Kuuq3nPz0KoKNJVo57f43HKKfAlBuBBoa8qvMY
6f5upKS+qcdQRgKYY+TLZi+B/ubdh154MyGtxEDTF/0ilk8JpNJbH5nXM9A8K933m+DDwWJBnXH7
O5a+ouatBo8Nafr2VteGON1nHNzFS212Zla7A6Lgtul56vqVFiaUScLu8w22FHpkX3K93wbcNJsy
cbYj/ElMVIJFsIbLVwRfZuHOracOW+lenEetfLmNzqdVfdReJiXldexgSAfZnhfzh9yIq8tBRZ3T
rjrTOWt4p5jxNOTpQ2UYEs5bnBU2wTqCoJGOEJArVWGvKW7637LKgAaB5FF/NamX+lgDGMsTe7BZ
/HKWtbvGpjYu2MxlMpwX0TISJkXfuZEGzkd7n5iiBnQHLHMdZeXkgNSn/MBNimb9LQYQ465PAUkX
N4gPRaMzPLR9OFBYlEPb30Gi8QGGidwEA3wHDdi+4ek7ZBh7USzmLXvy6yHrRuLHSxtQUqm8g+eh
t3izhI7Qa9zG6OPC00b5J4mNnFVLkhFn4iMdN0guFSRdphWQOgblR69ugdIG8bTpNMcvmy3++yYY
zJaRESfgyVoYa/BaOy1sPx0G14iVNv9Ww9pE8TfaDbz1kzqhRuh80yqV+GLvqnWveoimpW1oSs8z
Us7oRMocj68KEJZKeMIXKMQtcFftR9jVUwSyMNvsa8mh+mlQ0pGW5lElbQR96JaJKvPBdSTKRS6A
LD0YctaTWUymwbUd2Gn7XYum6F2A11gLhDIMPLeboZZ2V5Fxp65Eg3yFZgHrpAY8u6wc/3D65Jf2
tJNExvRXOkDSXKK0Dkn70fN4f0U8f8DDxdGRoKsNX1MlwUjCeDv2MGG22w+hp+roGD4zxsxHucK0
yIeFYyZtIm7uHp4N18dZgXCb1r8nenAdDrqYELcnksD4oLwqwM6WQHtJ2aMHuSz9wknvqkxUpGvK
xhEyYQPbaEd7aAtvsB1BlVKJI3eA/ebRCA9uI9dWrUsi+oRtdcNejoWlvmVEEgoXBCQh0FmENAeX
rYlvQhze0EPH9JjHyB980PVM0hUMBCwWhESW5KoP7dtcID+IA3/Yw0pFVE75T7iIB8pGVPRD8Vkv
ycj6AdpksYwney/09z2xSI1Yim9hEIN5zu2QhpP3VifLLwPrRrsLyBJmc6x5cLkD6CuxcCCcvPHA
270FTUfm5nTTIaXkjqLGpPBDGQ+jlCMlqb6O3xk6jFUcOVhFIXMAT272DFSi3vfVqOwS2vDg/5pg
5F46A6cU+N3Wr4NTQDjSB0/twapobLOJyDrZUv9lUnAQvvLRq8CUdHPBt2kUjLsPTK9yOFjgInIB
Fv7FAwPJ3sYS8P9pE9fXsBQtL+lLbNLLReJqahfT+IZMVqJ1pFheE/h0nmTYSFY8zZP5YXdnd7IO
tYEOiPac1h604u/KTF9QtFVXVEt0QOTSOf7RUcdOaE20xfWvEQM6BrDD6DLldNcmopGh9AtSbLI7
KbsRDYI3LNrfbxxtlmfDhFa+P12UWAlQer4RnJqFBh+gvyyFgR5Xe0ciosmycQi14TXjBeT2NxMm
J5ejZPiccE77fy94Ed8r5ny72VhUSRIitXQnNEvOYpxVBB0FLFlJY3VXYgaIemiE6JFt0KViWRWr
Cr+Jq8fZxCmUmNZUxMeBar/92Z9o/6UDVPuJoW3jWqXKQ2q3mpNjkhVkClLzg29Aq9Na2C02nfx7
1c7QCGLaI79fO6NlJF8XyjvFHN1IjEToCKcJPhdfMpJQaPEnVGCwpiKuhJ8C648pPocapC/6Syoz
zualhMVtyZkExNrPpNt3CQoLoqZszZi/wOACY1Irq8WFej1Zf3+qA1SgwjrGpta2NFSXOomGq62D
zKdOeYpbbogrh+x7+MXh4IeLnd+5r8YPeXpQD39SQTHdiKn7u9vfRYpYvsenT/LxxxpwVVgJPN7b
JnVppbzSq5BB0Q8fZfsfiuyvP3qIudBrYfAG5B9iSfiNc/Y7D6qwqdbacxMK59JCVZLCsCIeIsX0
8GjfQqAuZufsoPjico8EnJyD10r8oX+JBBQoJGM+IhLXrwhc6LfD3mI2a9CXpRmDtcoFGDBN4IiZ
jUz957zzZpswArphozrLVEpHRHLCygd72hkZ7FSAf9xSuNfRFjPvcU+9UvWTJbMp2seupZ7f/M+e
GvIzXr17LwM9gpyE6lY6RgJu8AUH4PXcO3Fr9VDaoqXeWDFPbLAmpCTGDGed69keab4LuKLRDZ9T
fdsemqudzOS9NyFiPwYctjkHcuz6rbpBfHi3VW2RkGebFW5vZmSiFpCOzYZnJLbAmJJkIOcRnHpj
t/IQ6zfUKMQEZt7OWkLE9LaEMy9owi3jxdeDucbP7wGQOV6MSbUcZXYKbBDfSl/YbIcIQaZpqcsq
2Ju6hQwj+yECYdjuRmMZ/A+XmLw4Qb2becluithuyqRWFK0P5G7LI1GBC2OjvJCJMH9akaGQtq+x
x7wHp9tALR2sRvBEloJvdirTZMQNrVVwUy1Ao+d8v8EzqhOwxkdm1aUeppnZJCIkrF+Hr34jOk2d
2hSZ5J8W6mvBfD0AcXceSZaghz/onG0nuvOZiI4wakXYwGTz4LU5L1z+2pfZ6Uvz3UaTlqMb+puZ
fSlnJVeedQ2YuIxGIGhQALnlYlol3yw8Qd8pr+tP1r0vLT9PkSAQvzs6JlhBMYSBzhTLIF7xfZun
GDY8qConU+m+VP/FvRIQe9LIKKlrm08b+qS8SfWTa9+0enTbSG8XxZGvRt171nkNVrw+NHA+pKn9
KiV/77MMry/j6Sdl84vKlO7edarqtTSOsf8tS2zi3SuUoVknfBW6z85ngBSj+6CgPKJRIWruQ8Vc
fJQXQKO1AVWJCo6OjkybyA3nBvaXMARywWvDnYN6KaTwJswoLhCsmCNKQDEL+aEszLFSzMORU4An
2bxU7EOofrROMh7er1R/RdGZjpzL4Zms9P03fKTa3VtD4sBhlCRIVWyGvUrSN65nigXkTX2pEjzY
THEBMvl5f9CU0m7+97cG+4tmyQDZ+xA8cpzqkBA5ZHuZ9lQA/NMpXOxp2T4qIiZYDQ/5QsvBjkrw
MGLalq82lep84mhzVj15eyNO9Qnje8y51MMYD8BjEwNbbGhMxh5WPfpx7rT3VGXtTSDrwAJiu+QV
W/0TsBoF2p+bhITL0UhAPx6TYFeE3I/LJLPMhZhtOwlKkfCe7ikuU4qcMBFEDSJKy3BuC5SGK+9I
HD35LyrSELxYtKAdwBAgZXZRn9NY61FtuubyK5r6M5r5aWuGbo0zrg7RKmHRuXFU3bS0r+1bdPAW
hIJcBiQ526zPXPqFG2SNv5C8wVRQky/vDXeTGualruIYEnm/HE51Cqw2mNAmjEQ7iY717aW28qCv
NMOHLhlrn6n4TjQsw/dkrGJfWIbw1GaV2zAnLrQyEf+aZ+yoynoWlDE5psmEUoTMxsq8jgbAhiB4
UKy6uNFDxh8RYQEGcHLUEVsNznWY2jCzDrk/HwMZ+1667Gu0LfU3C0x1WbdF55WprgR8wwFkksO/
oUCsHOiThwTSj4iD5vod40nM3Br/zMxqcI2sNHNpqFocCy8Hunuj2eB2QtMZoDK9xZykI8LvpVPk
5noh4powsI8GXwPLv1EkJCB2/DXx5f7IkqIcgy/aV4mll3wWCQTYaBIbKnoGZJGebp0Re6snAfD+
0TO7fzRqmvjbY+MvDY7auoLWzUY9uU2whUGmcnJ5c5R5l9bOwR4pCQHXoYGco5/oMWUdcBHI1Dbh
wAAuSwGnt95CGikhss+edrYI8Ct2UaKqiUC2RD77naRsGmmiCos2iezvOgCpmZHM8I5b7lpP8AF7
4b+Jq3AvgfmQn056rTAhN4ch0nc2rCzfwVCkiWARfX6XMQkdJAueEW9qpCG48mO14gXOIVsIbsF9
m6wjq7UQ2+n1nn4YfvyraYb42XEjO4EAsCjSGIlE5erJb3Nd0WgDk8SF311rnfz8FhwN3cg4Untk
fIdgzweVu+/jz+18ECJGHLGzwDedxjmcL3kQSRhNNHyRIyI9qmernCllaA5u06oF+4PvK3irvJ64
5kLOOXCd6ZiwV/QbZw67Dau7rIGYnN2XbNR9mdtTl+LVGOjuco1VOLsFCt3QcPsgDBikiSXi8dBo
Qec6yjhAAYmZtxJ892kfPsEMdgXf5nLOvKffq8lK+fxzEdpjhlfr5d0Pb0kBoRHzfRnc+fplufTX
KxBmCALkiuMP3dzdI/p8cMHtgzeqNXZ6pd6Ys2dgmRTDUtkEKQ1/q3R97+iREvCZbvTpm8cTeVP7
6l6UtdCEWmQyYhr3DMc1B8L/+l37MhsowEld3o67VdMKjgOau4GQCc3PU8dvrLh8w8N0TIUtOOZD
6gdsYzfPWG6gn0tjL8qGWTCM+6EMmDmgPYc6WE7qo9xDMiUaKTJI+eN+KSKzDanGKSzNugUdp5Q/
c2bptcO5Bp6E9dVVSFQzQ9ONSAdyPEPLIx2wxkRRPkoJ0RyklayASF68bEzR5OicP1zCZ3h+ZYEj
bQIvwnPqhrtbSGexIeaYNjbSiF/y/I3juXVeHC/ExiF/ZnW49riOzghpb8v5fbCKbY8w1C9fL4/5
WHwyl263xUADv3DfgZVCFvZMkWwv2s2NqPLTNG5BDkPx+uoJEFOKLaDVRBWG8Yv+FBCtfqSo6cs6
a5XnAlmcfcvNx7Gsi3cpxJPhf5ZHySvND03lkpw+2eSsSLezSooNjoJ6hqlMDJhIk/hs+/V9WqNl
WPjBF48RuWlzNaSLSiTGNAMF+6U7/GSMi4TCaS52VafVjsuaWt/GcyXP4huW2k8uQGZHLiLqMd/y
ARBMLGtGVXLxfuVqKF/25nSeudodnvGPyS7dRSh/cM/LkCYKUmpSwfXDcovF+tgolgkgSMxBjHgs
7CxH9vKsQm8SpkqeO+22HMv29LkIurhkO9yS+HOwwQ4LOQ0eQiaujskr5aNSr5eQaGuwPyKH07Lt
m24mIEI1q6lrTT62DHA5xCYMpXP9aTC1hyqSOLAeYL8oL5uZiAVkoE14ISSa35zI5t0GwdsLiazV
SC/z2jM/2WMz0syTMbJk6R6tTpA1TmHj/YF8rVWSfwug9CnDxVP4IwFlxKeF8FIY6UbSCkOGp0Hk
WKaJY3s5Dp9Bw5Y/oICEZe0w9GYZHsXEf29pBCe6HNBLRDR0+LOVaq/PLhxafXOKSWKanQDNVTWK
46/KhxpysRECSrJfjxG6DNEDNFAw3spyzPdMFtt4RNjOhHvehu/fKr7O4qVtuWSeDE5VWg7CBOOe
9/b4MxKNhseYzI8i9y8oPmvSScwLQSmNDUlea75XxZb9LDNL+Y4O78okmu6o2fcdgJNCTI0ICVPM
0R//Cob7BAeUpU8V4kO/UUlQ/zn8SUkvZp79k6qGIDqhQ/gvlnzpO10KmbIcCJvpRgWCg1h3DAHC
hpWJsR1wVEvwdYezp8lRhVZHMeCUO0xIggQSHrt5ntEsgOGw3v3Ok/sVpiWUxy78W6mxj0sbLaqR
bQXDmWTZJE/2jSfo3Il/KmjlPzZqHVaFJKgZ3Eri/FZ4g2pgIkhE62gfjC/TqC9STfl5BLNC23Jg
zShbV/P8qnPR0PCBZjk52IVAcJEJNL1kGuIrrmE5sK6EiixSiG963kLDrEkQ8iG9OVIYfNPL00Hp
3IATGU98NKRUgHpK9aICiKlTP7xaFf0dqIl+jzWygxm1K8yYJDHcoPlzP5FVMZGK4xfKAjm17/BJ
3hU8slwTlr9zxtKokaws9qiCHRzUi6PvUePtyM3/vEXZon86WJjcvp5FSNWxmsAdJQkxJRey3wZu
JEvMNogLBV0ZdCXyURX69QEcNOknlkldIWDt9f12e9GDIWD7vmVPqCXYmTQf8PVN9AxP/hfSWnoL
+Q7NAkfuqVPohczmjAgDghpL3dJLIh1b7hh+EUnn0wPiuLtfC5Mt/AUU0qGLYY26/MxtRUTfoVyQ
O0IeDK9HlKD/QaW3CVhR0oiadnwASEl3iOrCxtr574FEoa3MwZGllUJr1eDbOObigW1ixneD9oKu
K5HxjyHybiw71GywtJdjhfqSErBs00flg3z11yOjpNyfzd6m26rcMRWsB67pFjILBZQa1H9JLxcE
ScBEmIiOn6BLsQ4Do6wu0p43iiwURqs4s/pb4AMbOppquG85PJ08zA1SaSba3rCtxeDQXr8yuT0l
cnplzmKYZuGlABjvYJONnnetk4f4/sRLsQG4MQztgcj599WKBOQSiIyoHqbhig3u3V4YmpTJzNmI
a5uOzLUBkQxkMRr5IP/mIEKzaCM8fg+r7UtXOgPMrCtqIh7JSmJ3vkPs6VS1l40L8YXftJMPW8kP
kReVRBHiUBOFKqudgC4ChGxZnzE2kX0mT22UwWv7Ujo30hExCcRVnJEJgpQ8fBdlK0AIjtMIeV8g
A6rFcj9fm6oYOLNEkdeipXdflBWsv4GOffXm7Xas4vxg7qshjw4sV0zImQxrzVxpSolz0piMQPGB
qwDqI7tD+qn3Vua51g3rhhyQEKXMl2AslWRb86+jIyYbMrgHAOjJOgWk1enTU32JYVSEYR3i8+7a
0ov4XLmQ2LlhbuDD63LSvSeU3/ExQvO1oWEVWmL1o3E86IST84LulzI4TjmdrjbTjYXOflHJo+MM
cVRooukcvszitJ+g+Hb4uVmVqSoJafPAn9b+oLYcJXyItGJAhRC3J/c57MG4n+EHROD0rDcOPTZZ
op9w8erRAzHjPxa2drUFO/xQ/OeoxILatRNhpqAVgqC62DoBr3Cnw5LB9otiS+d/ldhWwFK1HnkZ
uCo6cNGvMEoV4uWWn7E7O5f5aIJVXkjyIp7cdgi2iwmwellI+H2yGlQ08BDUFV1dVxqTE+Umz70o
Ijr6eJw9tOJGM9YLXekWSesUwhSmOkNC4x9dFR9U5x5P7Wer0T4cfTrXCXQLBk8nzdf2+9sPE+Oz
enr/BU9gguSPQQZXmNOjiY5WM8RR/TpreqpF6WEP3DHAgAX6HJhk8rc4mpNacuxJRaKmx6W2BKul
aFrlxAx3EBjqRUC31skteG2lKOg35EsWpyDe33gpu2UNL0wy+ivbHa21Mtta2MEtJpOhZMYaYXvf
o36jvaegJynDMJGyw8EZXUPRzovHUAd/eQWLI0phO7uuNE/W9qohAsg4YC8ehIDA/lwLuXT6CbM1
gFrFav2dg2ekMQyJLnlEr3srqZaE+4EwaQaz42sYvy1+bMJ63l9x7N7tMW11T4KWM3xmbgL5eR8S
9QPX3MnqbV5esVGrKvIEvMsvfWIMq8D22EcNRP1/jRSU+DCZCHNHDddrm+Y3Kv3Q83VJ/9zJrOj3
8GlZnGPwBR1mR00XqxgxM5RKep6UDOKQZHlO4qeQDPU0Z/ANUx2i9fLLoKfVPw2XrNsTlhZEbr2p
yyu8PWNzEjMLSx7yjb5GZuZDw1P3PlU9xfsHXoPl3q+AZNlfSJk+NL9knoN8N/lXGVWBBH6oVyYu
Jtoz2nHipPDcEud8J0e4E7zUfkJ3A5qIBfCnMv0bvbFqxHXuX0+Ql5I9ZihSymmq8fXIA9yBSLUG
88QRN5LVw4d8jtvLzP3y7zIDyPOcGHQ3IIKlvCVkhJJMi33FC0QXz6U/TlClWpq5IC1fxb+zxeLq
VEWmxDcT2Reg1mtrlVVcgpWfhrg16jo6q89Yzgy6o9cCd+SmcE8cMF1Q10bhfsLNymgTzn3nz413
hWPu/LJZdgDEQnZ3PgdEIbhMKtCeeM0V7eqf0lZ3TZcsQYkAW0v4CR2IDOQv7AMqCALyeumwi7Ta
niDLnvoMr2c3CXjlpBuq6Ak5buBKf3F06B66Ic6DFOgTEBVPoYim9H+0KgzHVFI3JurImig9hFph
xpO9JAh6GOxdrMXOpf8d1KGp4pUlpIpV5SztN/fG8r8F71Vi+VPT5CTZWKMrc/DHtZANU47EqnFS
nynvpZpfk9seLb9a0ycfu7xk9OZx+7l8y8yJZEfGVCJ5mAaF7ZThJhlWktBp8SHSdz+vrc2ECppI
8o4cckJhTR6os5m3pbctxbMvIv+N3h9pRT1W/UCmwJ6vSoBSkYpO6wWvYGtS4CFFtDbJfsky578g
y5735Ju4l8VrNYBHBhVBFiBDhAaZJ65E+n6koY3P15hlCqGu8QsYE9tk4cOmQfIm2P/9hdjbOolc
weR4Ku8+q3qfrS065Qai+p9RwNd84R+9lgU5uHgFxME1TReTcCtZACWnoBty4OcRUYxIojNcyEZ7
LyuihifyJMX6Q24CdHFtl7NrNjCIxUCLmj6ygkpNTpe9aIzxJ2QPXq3E/mvGoBmAluY40mDzTRtd
FtOjs48Wtuh1V8msH1GESGZ6/5/rtW8NeBrOVkrF36aXtHAzIYf2yRWCfanmfLHwe2t3uYe9w/7M
f6FHB4n/rIbFpRwF+nuE28glHjSTa7ju/kQbOYbAUBCxcr27kidu3UlTPvfjbmfj4EPQXEVuquy4
PExbMJqPYP7fJ/FX4wBSeFDy6Kggbkh+nl/NSscNYU8GFKY/jRMJVRr6oL1F4mKzgwu64qPqzKUo
9gTzWNweY6Ps5V6pHwZJayrwn6S7JIG1tRoKmy5KI+J+v5rtJsF8kZN/gQVruGW3uGKu7IvXW6Ou
7Up2iDQastXZw8nRNjhddUglsF5Y08PMnQB/Kkkl9nQuGYR4j9aHnK5gRmgnSBsgl0KPDVirRTbi
F/KE/UEl2kLcRYuiz1U8z+Cr4nXhooXDLa+FyUqpHdzjS+z8hCXHedeBYAVClyNsptt2xSCKu8FB
ryvJL2ToHbVngY1Wyu5cgNJu2XWIf3qecKecBT0TL/Dj+u3WpElNs9NyBv8Wu099g+i6ysLBdWn/
nDujIraBpBynvLJUtJKasclNYzpidc7B68x03HCVUwu7rY5Gxsq/wvyNlZUAYVfvij+m
`protect end_protected
