`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gBBqHtY3Bunn5h37HpCTrctVa1SkpXy7VKKB+BLoIpekT1JpAEXVRxCRFlXm11bUuVEv/j3pO5ho
t9pTutZSCA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rT5AuEipXCjHo8d7Uq82KPZlLJRMWXHoM2CEgdCzb72AUhqeRT1qBpZCSEtuISLEowB+OqwVoPB3
zybnMbwQb0oxhzcN21zHYr3IRmDn/uWaTM/MMZ/bnwJHAXofyVKi6nJ1ZcQvvuVCoGL8KZKn2sQY
BUZNn2IeXewaklPHIeQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ddHO5ZrB/psVOnMQtFAGp/GctaRakAwKZKpb8fZB+TnHO79YBQYZi/vlr7RpKlgamWNfGsIyviHi
4DIn7nUd5XwZ9QHp06khu4m91TFepB2UCDybY/E+nqujVmmRIT1MbkiDUkGmGhdlaRTui9BlBtE3
0V8M0AdcuyXLUOGcPYN1g/l0n3iEvu3eoNOYYP/kCy9cKfwaeQHNoZehf77AMdR1pfynz4YwSujK
w1CXonssc2+GvTDEUoLQ4/Q8xeAeoZGD3iG6YPZW5ScawzhsAidgis6DgRGKTAhRGMtozCJRfR8G
WFjtcUsenGju3BFqb5waLMbDwCr9/0sFXCYQWQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hcWMtjkawP0pEAeHRPrwjlkoAY/aJ/OE55+xUYc5sOa68hwNrmj1qF2ncvb087ShjKLuEH0jfkUo
QzvhJlOJJxno7QOxZuWkvY91+e5UQOL+2j631nFnpoZE+MloH4Mb5itp/2QKWciAqiwm0+YgSi7a
rgZJsggXf51kL5HqrmJUBWR7819hS9n/qP5XtJ8y7FDBu4ElmV5DY2JVmGTJzFc00gGCP6g5ZCbZ
x2WaYEa9rwkMAMQIYDPF0j3AzZOJf9BZ7TUjt58OKt3LANApygtniZkFFlRSo2PBSQ3No628n+ht
7Do7iCucrGBsrniezp+n7TPQFoCS/PsKj/0Zag==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M9pROQR4pNGukvruDI+JPpAyg6zBwqv+kvFvbZWk7i0NekZFvWp7FY0oY1eWZ+XxMsuNHPA2Plg7
MH+MJl6VkCL/cJ2+knD2NcU1AoFbgFqErwcWRYVepmitEaQCaZwfy82Wax6bBGqHKP4X1cQ96V7q
2rHMe6dFzQ6sbZJDGr0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YmZTg65xAenvz/Kb7OqoEnjCRgOo02BX9BzONEy+LExgkp5FbIUmzte7VnUBMqyOfrjbhR1gwsSC
E7jpY1rpbjcIx+SqgamXNDfuW0JF0+C1zkLYSPYugbcrMUXpChGH7bk6WesFdUAwr/Ktyh+Urq7s
BsO32fxnO0rZxYMJ2voFB2hV9nZov8aL7baRr4ZUYDmQxS/z1gPpjxqoqa1AuT1OEpW954ozW8uP
b9TWRqViZmVvgktghhAp5Woa6dttGplqCv+T/yd6WcKv8U+Pc0RzryU8NUKwL/WxrBgu7Ba2LvO7
g/WeYyKq+hYf3O4ZtyuIDfGHBhcpqCUnRRVPSg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XSieXGZEsQhOJ2iwjK7eXEWDvgXxCQanpoMe8ioBhtE8cJi/QGFtNn5ZnII+9PCK7NrWxywdcuIa
c1zWLFnxppl000eGkfeyNxHN6jZL2+ZFu/PdSDS9iHl/x8HlFh40DjlqTkoxZLUs12OKV6MsJbnz
eVDzsmiGuMCtnR1GD1O/ajyP4J0vmVDwGm5WTY8NXRuJODjlsSgGP9qnxTANsE2CJUW/5VjwahFd
lnQc7QKxVYFfivRIxRpjMPi+njmOySEXEEwVklTwOXobxyeOZ6mOeReGoAhbJivQnsxe34MignfB
cR9hfUmEkcVU0Td9FY8BgXjUjjeywjJrKoW+WA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KmpD3XZFpLe8+sD1iGwEup6bfACKiedaS21mQM1V5CyQMjx/p/K/npJNenB77Gsv031GbqLJWf5V
fbT6GSFj7BtI+Zci6hRlAkvZnNNqCaWgoXdIoDE+CXp0KnBn5CaDdAN7GUQ8EPx3UkZWDjZ95/80
Pd8OG/SZdQpnjtHOs6dZDthcXgcestj5Jl3/O0O4nevBH+OB7KqzA8UymTcf2NHBnCx2s6nfDbW2
C9LgfejwT0EL1/dR0i/f3AwiIwwTCQAXxFiE5IaoctK3kg/KtdmAblRzXI6FOvwjGAZLCzA5JXkw
Nd/EAOBJn0Rk095M3rpMJruHjbzpAn3t/WzMzQ==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C+FB8r/tMxRA/SU4aH6F/elCSsnz+M7jAys/z8YFGgwvumpGQFigA0D8dS8S5DvMgxfak7tlkOE4
LEte3Em4KJ2VUGOWsRCSJjerMYy7DlhPZEE2q4yhdU7fz4hQsYWnnuuHt+uEzyFMESj5KBVKmURm
a054fsL6z4UkeMEwHG17eluOnEb+vJWan2hnHekSxUgqYY2FX3PUgRSO47TX4qQiQa4pdDxOB9Nb
dtmBxXkxa1ey15e+nNZf7ZKQin3MH0JTFjnbz4n0D/ERFnXqnTG4Z2M6RKyohLnj0TyxBL4Psmgb
cJ53Tx7rODwX3skEPgU3YIBRbnoh03Sc5Fr2cg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
oqrjYA03Dpn6UrG6nwymuQ7cbYEL7RazMOBaQaZuLQG721ZukT6Lapjs1uaioob3cqUzCVZOAksg
MqBLIjbB8iS/VZpvM8Dg4mXDt9rJE4Xqbl4B8vp9BTsrgvCqF37VFqlT6L08AhFcqlIYdqpRR7gt
FGWWjnIBZ1QHxOhuRIxy7nXnWAP25RpmkmIQ367kikuJPjyK+L44yqh1x54bD8qM/Lya5Da8hzjr
/LEFm4qmRAkhyoJQSydYYW+oAnR2LbfK8St3EOYYiR1j7fUbYA5UM10hVMMBnUWKzATSukqX0wvG
rs3YdSHhadbV9BYXKyW4xQ3lMFjDXCS0AbAZOYJZIHxmebTDGOA4LX48xCssHC7d5ahlypdYPKfd
Q2PyIcQ3JVPOxI6ljgGZNnoGrl7XOkPte4nx16aYyWRXgyWMUwlyGhzg6mHIRdiLxVoc5rHid1ZD
XLGZvMmtdgma94XkHsP+SCOPv0b+/F3UshOtNmQCcwhbLVi4UmgRNhPJppvGO9gnIUgwz17s6ZVJ
GGGnW+cWJm9GUy2RS9dRFJYbMleoQ+q9/EZSc7rNAcs52TJvXAqKbovUsSInzEspQvxcwHJBcnRn
nT5A7h0qHt7dW3HWRiIFCDLobH/hW+NphMD6JlRy1LXTWkd0WCWSxFJhshDYAY7/p34sLvNEXvpk
pO3BLrRX5C23MHa5zKHDgvO6dFM0Qhyju6MB6RDhrjgJyRhnvFuBLUUFRs6lWdSIebbYkOe2z6se
QAq4AH0VioXsG3bcOuRUljuiRX2yl7nb4uUnjSaKw9lmhQAbHdX4eYRITlca+fk5BCFdhyJ95mbw
05gP8zQyNHcZG0YzMEPpAA0WLfluSRw5+uO+gSOHHWVmLuCGaU2tMEU8cLJ7UYr8AVZhYLoo7xPD
RyMv0YM6Je8K+UWwwXcBrZemfKCyCf9xbHGCXZgBy9OEQCpvvWOtUcmYaMdkiujgYSS/e4q+HAZp
lPgZnFl02YEODS+rkwpFC47DIlnyRAi034HtE9n4pqjJOzy2YuTr8PUMDGft/k6wRclKlnxd78Wj
xFly+YRjSccmpHz48q+PFkDc21mEM/gpKpX6eIpFTQnsdQPaIaOMl/uHQRqrD6LAqQlhjRU/b5lU
AnOIg9Mo6SeO0LrkxbWtOoZp7kd6d/z36jNNGecyZpzVaVrNfsok28mzcGpjzLmz9zUciT3oIHFv
kCmWMcWjMULGbKbh2/7tv+Jcp8d/PW2NsodBZJB/9yRkogAWn7bqGH4JXHzmunhkmanyuo1BiKQi
gFChsQqIrZCrtNxlP7DPXVD8cCW2FKI+n2LgDEPhDICbSUfvEGfX/WsX4XwDrHy99U2GEPEepfWs
CX8ZwciHIIPru4fXHvw2ukyhx103vrsxXdxWofz+gPYVj1ZZMqxu/OPnSOfvu7nskKuPQulDHw6W
aMHZKKjdKY1Hlt1W3tBEIXYWbobsDr1B+brwA9s72mrMHzofQmKWssD17BRmI+p4LzDXRtA8/rPB
AswPvA1CEqaa/Citfh0tWhgSpHJDILR8rtQb3V6EOe7IKA4D1gDUJfFcYwS2q3YfY5Zpaer9yt5c
D+lM8/mSRLX/zYnkrpVTDNqwPDubwlgQMsxYa28Hpw2zH2bTJ3OSbm7dBW+Yi9O0XXy41pQAANYm
19BvUVPEQNdjQ7uSg+eRAz5q6LdMJpuzq7IypYwPJO3Z46w96zxZi1uVfYT1HFD7C1QDfaghooKQ
ZS0BVsz+MjPqvN6UbuM7Rcr2rC014hRN5dd+zYHYfDhecyJoGDLNKm6gQfwq/drnuRdZMo7fsOsg
OfvDFQdL9ljkxFyYmkwHYbXPEB28KjMv7W65qJVaeR39rfw12Os4UvXNJ1BUJfCXlUSuxlgHEJhH
Bqmkfh28FT3jjsz+52ZIfXr9wTe6RWkQlEm511A1V+MB9AduvfwkWDKLNWcXdkQAWkRVcOCFXr2q
nu1FbOoHG8c2lEXMt3z9gJTIbk0FZr//nNzswn+f+3Stbs5AOHG3C8TEdAl/2jraKuzyuI1r3DHH
SSo6miZSMTWTzgqeREva0PWIMsIPh8PGREWMv0XFPJXRV2wrXcoHpUQoW273sorZi6hBbr0Qk+Lz
7XLnnSgErAn/iSuiP/7alTNMrkolX90ckJMOhTe3xTUfJr1zg2cE5fYpyT08tKbxIH+K/f7Jtep2
M82MZGCP+C5UvnO7+x+sphqa2vU4OW4+LgCE+s4dYoeGPoqYhCbTd9qj4T9/iPGJLWn54LN7zm/t
gxQhT7MwX6wBl9YWw9sr+8yX974oD+4cvU3NWEHSjANVtBa1zs8TY9L5+xIw16q7Idt1D9jfMmnT
EhbtasWWIzJGOABDKWxYZhtj//gGO03wu00SSczS/visq7WpaGfWg1CgLQSYApFkcmNXVw6LaatI
fl+ZN+p7ee2vDI8rb0CLhgNl7hWzq45pQcHUNKQILfyhWcIMV7PVUyq0lCe2DtTjlJs/rI3ZHprx
3i+SbwKVp0I7R9o3v8RJpItQj6+ZqI7PawkfYXag4VXoLWjzFYP0gR7PISiZDwqfQ77hSxasJzno
BRUoDrFV1a3JpHamh2UfXpyJkTHd5+16WfV+07LEW8g16q2S55GxBLVjN8WJFYSXMOYqzKj03v+k
LFj4cFL9YQ53y73A8AL/VhbrXiGV9k/Xps+0ddHQUzH4y+zm5619Dup6SSLC3LxwqNfxi9U0hwxv
80ZMra1e3UbfEbnJH3kOQfwGeV5nlzWYcl/XFrWCzZssDR1oJ66/C9Cd2ooDfEHX9q6wkVHm/z8o
4+WEYZmguardc7XnSKtm1Avb718l9jlRgmq1bbgKimwVkRF9akAthjy0OgY0xVQpOBb+V4HGJY2m
S4myc6e901WJlgpo88mK1V0ZxXqoNY2iBKZR+e9Cmckj0HHYFlRlhCO9cJ9tG6WqCuj01eYwwiN6
KjgScnAVHSIlXlVuWw5RACkiRhUQRXn7DnQSmE3kbkA0WTBaU0yl9cMpYnN1M6lrLMZ9c3AOCX2A
445NfyBvNEA/KCBjjO+jCU6kBIHsRZ9xVs7WtJGgXjqp/45BN74o2qjpnbJGiIkVz61YDiX2/Y5+
xIZpYQdfCkH2YZCJjldNeQURWujXcDOIN4WNwL18RnIoTm/NqfX1CSoUKN+pFcL0Y5ctpd7y/3ge
b/wMTcHWN81udex3xqSBIFGLVNoABGNH6LN1P12qO0aKIzPPjjdbptrfSgkIeZ3yKebfn3cHNSA9
lcd4Vpck5nqMyyk8Zit5EQfBT7LP5PbbYI8kbCHAZIkxKAyU6VWBMoCCtF1+Nj+U5qgNRwMezRhz
Qzv4ApbuyujLSQ0PtHAVi3aNzuImVQk2wC63Q4avICzEGnwY4u8F+X1ldU1dU9S+Meh6VWT1EVDw
H3PLlsv61a+YdYxfzSk/WCP5ixb07WKxFQtfqeWEOwODXPBl0sPKgUVYDhBjvg7gIDj+Ix/N0zW2
2VgcDNcGVonoITfx/UrRStnxwSSl16jZIhIoluM16xm5MH2qSwguP/m/XEOyrWSkbaH0crw5P/m6
BMpKwDxTflfy/mZCBrZ821VxsskLcWvlUDSbsX9zDxHvsEqk5eTIbwuYHRx1JmxIz7uP2XRPVHx+
Y84oBtzA0wrGGFQlY226+ut/G9ZulH2JWgrlQR17mEMmIg8EkLfAnRn4+L15Ie7AXB6zkKN0bpf/
8QsnGNvd4r5cfC3GCHcBTasbQMB5Q4eTXHu1A8zHlu7TbiIuG0otSZHL8LRdDhCfz89RPDch/iKE
F2GO9I2DmsPxHDwJr8c+kyjvhhC4p0hM20/7SOYO4BCDY2aioihU4Z+ytVydpN2iM4i/T9ck11Lg
vmxDp481oGKV4ae4oBh79VQdaYutcm8C5nCj3Q7gvk98tUBBCQfV2iZ34aC7S7ABo71OFJuYp508
Ary2UvAt0l42Ad8R07F9VL3aIqi0w4uumwG8NwkFxsu4Qz75ceaNe/qcpKFZNJvYgJHrEYPLqz5L
p8oFqOuGyHnMno/E16Eu0XcMeJEvj3IK6E19A3wKXwkkeFeRvgC4flLMXYf0vHQnKR1ehdYYbpqr
tAuAna2ixTeujYetqxBDLxVpprqYE0DfnAxjiqRNZ6IyK0lBNui+8z/UEX9ru5uFEeBnNHWZOtGC
OecgUuM/EGQ8pCgaUIoR/9QfmP47rCPvzK5t/ZiBt89Ga++4dV7MVS9DsnMIAP37gJ356oWCMx2W
TwZ8rJ2vnxlGrcZp1eYCOU8AsEwQrQjzxEl9VPkefeQhaT/WjjBpEHPNsYF+/PO9LtRmmXDuNZyH
WActNoQP2hZXzX5+mgXFFr49fZ1HqIA33sjX7B1KVnseMEv7VRxfU1M0cdClQz9OxOW+DrmVDN31
M0lA4oYDgFjEYIrMAvk3zN4RDGMPX91I/Yt2jse3k/3rdoSG1ZB/bANjXRHlqmy9yuOwGAnwrYQ3
WweaWrUMufuqQb8d8G0vDHv517T64+Tu8+r0OWNvgN8OckHDvVya5Knq0O7E7U0ZeBJpW2Ub/Vq/
jvLucOR8jXAbYzNbmohKL1B4tCL2sw9fZE4wk8nxtH0XDCxwL4ptXbyn5ooNYwqaKMNsLvBYckZ3
rhsNq86mkUXJg9zJtMww07xg1f46tWT1KvrXE8PssepXAfzu4cDPM+CcD9nUcbmVa05+sNsMVgrO
dttRwY9ubdBb46AyN0NqXlpiLiabqDKSAczefxjD9/fpqgCqU52rZogHNVMfTHnMeVu3dWCcZ8tC
n+1Q+CrCf5UO4OYAG6A/j7z0Hsg5SIOuQ+hNv96dBp3gj0lR3OHGu5gj3LEdytNzMGd7YCqn/h4y
shBi0mP2MMfWxnvSt6zPv0JiW6DbhPFJxgWvlwozw1GQqXcF/WAZrCCuRICDJgmeffiFvA6n3Rea
3HADB0VFkKiE5F5pQirmf1ZYn2MrpjILWT6dho+4/7Bie51UtW1MyeYv6mpXwvclcxtAIJkbpC3E
M6vA9leGUI3P0zouQuHTQgYjouRwSGGZtl1xupiawa2h5dFl9pUwbnKE2ftecUEkEd6ZvPxRAag4
u4CSYp+WgZtkuIvhqS9hWht7/3QuZEJcNTvfU8s3dCw2tqovwCJHRC4sc0s13fdgsiLJEWXIzfWz
MRFctqJpxmh2lPRMsjLQszZphof08+6YcgHDptMc9uQyX7AoGOySLXl5qlw1CR6RlhRLbtbTfeTd
cIdzpO//30doUD8kZAD5Vy8w8wXDV/5Ijr+vN9QRqXq7xIMkZUalVf5MpGYCenNfWDwYFgiwUfuu
o2BejRidzCqNlIHTqF7LXAVns3ewz24v9lirKpHotcsuBlo6B42qRxaU1NTj7x50R90GIaqXI7cg
miKRKFGtrJmYoujSoqAYZZwE6gPvkW5F5fOfJA6xy8lAk5bXPL48lo3GV/iArRfI5rLnYdhjYbqJ
r/c8sj9PnWuNjjBr8cfSvCM+unmTkD9DVcejdnyn56Wh9MhfoMtvk3OdG4MwQWwt7OeGrfoxYM8Y
Jqedj76kxNptCzGZagLer9OU7FQKMxyAxDRL7sw96z8YW/WrJuzviqAHIf931aDcP5zw9M+a/GhU
xQroQzaNTBmTD0Z2STuXIwv/lzjEdquNfNK6Lpf6YLQ19aWZxMkcDEJTQ4LrJI4opiq0Ie23UVDT
la5HY1l20ThG+etuABYIxqOLEKfn8+tlIn00L7a76VdZbSaTxufeXH/b6Rj1TD9JEBLwbZkaZaA4
RWzMaQnkJQ93jbE/+AqkilwLCRLmjjkMUNSw/5gpQ85rnX4YCxO+McgS5b4NEsyFHTa+VIqbysWG
ab5eOciSE5LKxgDnqY3Vl/tgvSZsPrsqtSrG39aLGBmNjUdr+74BLyr1gM+IzgiBRY2F+tqwtg3D
4K9ioWmQXa6qL8W3vSwH87mNwM0q5DJLALFa93Y8W4F7rVsNxGS3Y7wY0YbtiLaD2ellmytjMo9Q
wFagaKA33RpE0OOn1Dz3Mndsv+4T0OctPwNnOXBQA1AdyrZNpiKLUxe+7Ull9RXFHPZHSdIATtHc
w+dJjP4XjZh5mgG/6oHLQpg7Z+YaCP9scVxKbGGpJEKEk0PIznozrBTfkyAF7ww0inmtua9ZW6Zn
0bbeqBn2Fo4tG0c1OMk/phUjjIWM1x/6H/oG9kPJwaNAsM/ZmlWZ1V6FLrcJgb8fLZZOfm4dJQk1
EUcbiM3/hmiyS6JH4dDC02kK81ZyG2OE2jPW7y9oqJqHAmq4HOao9G4IQTAEQs1L0BLsC7FFs3Ee
HSNiJNoDHC52tZrfHKcBDxj7/CDAJIBu3iBN5TIAw4J+kMxoBbdtY7tCKue+wByOTBYbiKk6yvHQ
8f+VxOL1G8sz/gN+rAGWj/EwhkK7BRfusKEzBhCJRhAOf6AQ3iRNpnM+2X2fXW4obeCUvQsEChvS
aU+oi6SpP7qr++xqMSVQQor5M8gDFRMXrbvvsO/AfSxFW+DT3nNA6vC5GP9g/sreZ5o2utsCzADj
H5xDnNQi+Ey86eFQp5GUyk3iS+kVW6c5jK0rvoKj2Si20R+EdFFJZI486L1zDbOuXBWY1Hv/sCvv
NbQmN7UuGfOKJMrWuTiMXnNGxxEHk28Nird5SX3/lThr26lG/TPxi4mf+ZBMxvVjtYqedTH7MhwH
mbKcBU7kTnx4r7CTeLlpjcLtzWrbM9viyycusOKYZ8QAQC/1F86iqwWDTuDaN5Mp4P6TO1+YZMQX
6g6rChO5X2IBAMwUPcwC9izIevIm0HtcugzJ5uFFlhITo+1EDZZj6ycegWXxMeIwQn9nkY91NC6K
s+LhbB7ni1eic7l6JeKx2gZ9+hC8/dYRSYHDOugrUiblNsVfz6qWpM0zk/Giynlv+1RUWLnSJEOz
kyG+EFH/MU9NuIsu2yGU5Umfyg17DH5ZlOQQuq6aFboI+ZWC9wJ7B1nfU56czDgrUfZ5VtDy6BAU
FsgeEsHCd+1xvPc0XqkNdbSXuPgRcnGdCe+azAjJ4oLW0m8KxoioF8DmvuxnV6eJk/YQntQSztQY
mbbDsdNHCY0qANxBlBdn2N66L/jhAotVV+OgsySArkMkwsD5VIVn+SnibcF3chTgKu5np8YVvFCk
EAsHBwIGnENJS1tdoRotTs3wJdEOJm0y4OjdT6Z29AbhveYPxFoILx8AG0RaE05WQVj6sQuGTKYE
DoXdi5rX5eh9TwpGS91rUTm6A7pKt9u0Xbqppqy994+Xo43hF1AnDetD10FvVvUE7y4hYRhgZ7za
F4lUIVoXa/LoeHj8HzAG4rBWXtmP2hMMJRpBbcmZ5/rErd9KDiTWqY0Bg2chfBKga+SLzQzRIPAt
KtbApBmanlNAwifEFR14TMgekXO+FkRosnFPFHTMRSqqqlFZd04VoDw2vTgeufhiBttukWeYn7Xq
FBW4UlbKbTQOh4V7NfdRHLX1IRrD94Wbp1aP6gO1sPg2GvumyX3XRyEmjcy9e5wmwj0XNIg36j3e
mlfazuspb/t7agtIIvpZqokT/zNpXmNAPvJ3sQ9qSd6B6XlHUdHGQYfsTM9CVeozeE3Emdu5LqsF
7x5R7lMu78qkV2w14HnC6OZb23L74iMjepH4XAXMyLutwTzxIX53xlv69dAwXOwp37lJcfSCSQcj
uLcAFYoM9uyImlcADN/rYECqih0RCbb7oEP5xte+BDuK4VDIe6TFJ7Mfuix8SKQYQQxgfGgsZRV3
/jFL+nuiJLySMb7TRDKCiqBRcguGpJheJxlJNAEfd2iqz80uTXu/0uXIpsYwdo+jNlIYSRgj7qkL
OT3ArtM0h92Av23/ajLeabNCIPw0T9Syh/mzn8wlBdSiOyIn/B2KZMnazjjgsHLkYiLdfo5V63l1
mkOR4ZVKKrrp2rdwVufI+pX0ueub1X/Zwem4E3sydIw0KBV5Wz96PpgGlH/GME+u2x82BKJeuD3x
R2kd0MH7UlQE1yvGDAigNpkldyRsB8mYlqOUQ3Cs13iUXpkmzLwZZFT8Wpblwf+Jt7F928wxSqPN
POOITUUQTliaTFHgHyJdqcsM7e5MoIR1Iv/xvzKLwc7Rpm6+LDgiY6mm+gmB9esuqcFtVuRWPRaG
pvMNMCgrG3d1b0Y/hOp4r4KkOfmHgRw/fi2FxcxRIKdYFw8eKaxFtQ2cNh4cmMQplcOjPdQk5Ww0
LUeW4NOPulspzQG2KkreCpMDJ/o7AClkdwfbkReNdzH8tsJsozu0S4KJ3N6AIAT1KNLU6MrUkbR6
JgDJnUhPNnSKxAPHhSuAGMWbvtguSQPJvdLznBrXY0IwP9RnH/3UDO+XgyMUYoMBKYoBEQRrrszz
hSrU1g5ZuRj6jLSBJ+gjaMIJyUnDAaluMMjvsX1/1tvweIfigJupeQl95oSCE9yg+2p5W4qz+WGd
XPMDHNF1tG4YxRHTkeqwvb87uH7jDwVx8/hfeRc3XRyaP5I1faABWda3DxduHDvy9PJv5v7U0tF/
KP+mXpbzNwAhvz2j/hG7ESj48KOSUnvwj8+Og1OoiMlZFxjm0oqlBlDVFs+mJrVnMaEkt8Yag+cZ
ssbmEECH0R5pSM3yexfPH2cDof+8EYcLH2yyBzt4PkloLXRz7x1c0Fe2lVpyxglof0C4gLs8tInm
QvU7fk+txdVanN135RQ1uY2/5J+BtKUD+TNGLL8MCM+EVJpu7kM5l8mDRUElRthLGRkJkKRZCFpG
uyBFbNa/+6AMyCNL6A+y7sNauAZVztoA/vrZOnit/tK7lxCu5IIn1gkTleiEYJkigsfmnW7t/42s
MRo5UMEVEDjPttFRE2/DShiqxO4B728gJ7P10GR4C8bs+c8b0MJCEQlavw6kYK4YWm9G46GIaagf
UO0kRfonEvBySp6d/jUWHaKmHEdve0nuG+LbBy4k8+BlFjoMrpRTKCsc2HDJD91s9mg1SVDMRpwh
KUaOuHg7P/Cp2YCtBBQoMBqSrFtbCMuQMk5joDHop2KjI3MxonLNWT3kmB6u1PDaejPjTyjbOJR9
h7xzPxFrSXin6SOEJpdYC6NR7YzKJRPWM5G8qEL5JHqaM4eqLqBR9fDC9lk7Ssk1qkH1IW0U/9Cq
LHHR+Ho6Z7546ge8JKpTTlTg8zHYk0viGs788X5sCkla86gxARG59xvEbKlCgVJ4RDqXm05t7ksq
2ybw3z61PnP95VOBYG4d3jQkKK3uxwJ8n2GW0KQiwJkJS2zO1OMoHor4wP2LAV+25zHaOuIgF2Hw
cTemopIh+K0yoCAhr+ysJ1RJVLtAR6gxIc2oXctz5Z5rrY3LnUyHJ8v37RNgMlEXkMIWjKDYmXGn
W3OXSqC1YXZYFFyeNCDfyCKIthDesCu9wT2ZyNWjIGpZvA6WzqRYfBwAQc95IkMaFoISj3Zw2bAC
ohTdlulEil7tY2jrHEGUScbTw9+KySBKHGajebBqXT+gyfqrF2JfoXerLW8O1Xg9h/nfZ6wZKYco
Moc9GI3B8woqEuRcIbocjTlWpJFrNvGu/7iu7MH6DhMUdVoEV4ChbxHSE5cC+HV+EM9bd9iglV7E
Z4W15tJB2ktJcw6QF2tOA6+RKCHa/xWC16HvI68GVSfTte1ywhpOREr3dBwpyBEZvpnLiNA6gSfv
T2IDnxkp4q7frTOC2aKlsr5LWXHQd4We+LKShKvvhWEQ+EUMJs5sN6acnCdEYLtobFLZNxmSkexa
7gS26uIhPoF8Ejo9to+7ZBZX5iMuc4Lx+r0ah5ZC0O7tWHHGafe0r3Ezj2mkPVxVyQJU0N9eYn0l
oBg5nPN3Y83SFy7X7UULWbIpC0w4zQNWYuTe+ZkmYxm0cTWxxGM5YIUizAiDezQy16rxUXOux8JA
FVbO3Aa4QW19xFIfVmIkPWnyv9JNkBR3If3SarHNjYnO0IvZ+M7eJASNpogMDP5BQFCdgKH9muNh
DxqbPrKwVAMwCE7JGIqqtKCb4Uc+56V2C6d6pL5W9CawZYFUREMSBTJt7tumtUn6swwccOooatfe
rwo/vwnESD+Ip4fk5IkKJR4aq8aLVo9XbwMHNDDshcDLAc25cu2sFQ6j+d97p7dd4aos8d9sx35B
nOlQweHk6DJM+lbQ4Oi0S1ty/07gyZ7eAf67e26Vx5tG6Knel0EWr0OPL2OTBDoSK4mXRbwaTh3k
HOKIodo3rOBfUMENNzVtO3PPY4ulubS/Vnqi+w/2r/cFi6hE3WpYfFM+c3DKJvIrUwst4sTPVuzF
AJzvBjnFonPCOj7YkOV1pxK3VgsZVaz/lg+HOIN1e6OmvAEy6fGx1H5pIqA/vuuTaaciQHQT7eOK
rgHunQ8u3YJkVJwrD+EL7gUdGAqeTqI2BAGrQix1FVrnuXsDWHHYaqrJxP5vmVrGMmmr3d+1uL+e
4Tx3xw8HynF+E7V9WBUpCrDkyhF1l2VoNEP7Bsplr/EAIJ5SYBUbcu/RMsueB6qc9qktimJ1sgJR
Yrs56mD3V2CSo7LuywdULPAngT7ZikAfb6dL6vaQ0rC3p+6cBx67TNYy4vQYAso3NsuaqJbVTylb
JJ//t/6O/HLiVxOn7cHzqZcModNwNWWWJtXRmgR8GHLh17SLKM2TmBaBLEsqoLvYnsKz4jmCEDqH
8l+1Ph7mV2+uPbVNLn+sR9xrMe0FV9iwH47BCEnHjENZbCUTcsEVWBdBo3pDngLdAfxVpSxjBQCa
0OV2Ceg8oWp4XSX9zHoxOqj1oZOupnIBIyCGUzK+YikodeQu4lVJCdqSS70INoMHlcZUHte9VOTC
7Alp66s8yKQJ5XvZXxM20Ng1g9Sy5qu9hzRBBj//Jca32IXPkyxCwZKVO/RhijrrKrC0e84NhBVp
gbROfgLru9s82lxbWVkygFnTEyPtwJnZpEug7o8zaIiQSwXG3HZY207E6RbgExCHqoilqeLErkZn
oGbLwhkRk4cumjWIGOJ1wMA2y7eW/DuqbeO+zxm1bzmONZBXxKKANQ3mo2gwv2thdemE83i2VtIz
IRwWcWwMyv3RShLacwEMYsvBVtIKDrDOD7tlgv3X+7bZTfBdRHr76TUTnsRz535CWe9rhBOGRLlO
UF2rrviVmuuFeOpsmQS/NzmD+fov1nS0Lv+XUNj9OBfa1YqDyyBeH7HgyDa8K99kKfWktBQQZeiK
PlGKMPKQ6Si6Fc4U865IA2oATFvCxsQkI5jFKGKbv9TAFn7TWO6NSSefxKcF1ACdU79QR1pGWYip
5TjvZLM3FzKr440BSAPVReoORZuSxLTnGXm6wjU7/tyzsFT32tMgDrcJa6QOR0/qEoYshAHre3SF
G28qsx5h7A04HSuJEmBxIX1MZQsO8SPU7hGjfdn6UGcJhpggb2LNypZxzuntgTtkYM+51/freOaM
I+FnDouuH9nhN54Wjdifd/wHrEUGsEB9H5w7Ta4uso7GYeczEmxy23U2PQKYqyUeAmkT0dfVqwYa
LNbkuiuPod96OTf4rgWBkl6eZ6sSbhbKIw0VbuQegdru0pZYBuBdLIxrT7UIWDk3DEJtWuYkrf/t
BwTYtO2KTmcqXdRJgrDG4VKFC0CvdUfu18cLVfJ9kH0b7qVgVlMkOF4Sn6mU7C8E6A2GengWMMBj
FH7UR/FaygfNSiuf28XWWRw6Iyor+jyetjkJt8FYmqM9qRWGMEhV+oquAxHM1oRXsI0N54ENraBz
PJmQ1UCSVBL8Rf5i0MeTndYDCZOzfIHXglRWjeyK28eB1cQM0EzHAa5bCHJdQcEDMWv7dWg54YTY
HLN97Ky4B6k22AU1qdf5IPZ/8C2TyaiThVClmlTvKeV+xmYKxqbu4IoPHpO9n9okiIMM3wu5ekUy
fU2wnwzP9gp4y2kH92JvnJaPGgIc5AbnkCDME6iRZljHbMmWzKYMZWuy4Pm6ViddvBP4NaFILMg4
uFPeaO5gLiGPln9+uATuBre+BYnBF99XSUWtHyBFTl6Ca/oON5vwIH/o+bXmtT6jhtCRjiuw1/FD
38CXjNjMMxX4cgpFDoo0rKUSQM3LayKpGeYBVlXFEAhTAk8ADv9FPKY58KqsGRpg/YtgvS3PU60m
JiK5hJRRnUdomtv9XZPy9nIXdpPPPqs0z/Tq1oU6SJ9vZGQnjpvVD/2+BMnCrZ51Z2wEbGVkIEoh
ZMoqN39z0omCt0l6s6P+VxGNKakUAIaZo8/3TG3ktMfAmrp6XtAg5J591ki5+lGqMikBL6PVjl1Q
oNdsDfXoIWl9YH0HGd+R5+11Xp+MfxnLLMDpRdQ/96ZCAawRONu5W1o84KNQj1ippDQZ24AsUWAS
kDzT/UqHnhPZIDAoueiOMkp3WuprzZZB5CvUOsQyL4Q3UzOsvHnhse+o0eQiseEpTn+LFaF8irVK
EcqkXTPYP9Pu9qOERVcKpQCviZre0Dqi46zWMi9V1ic3bnkphjuE99lgwV6AzfcGXaFdOCq9dVd0
+FQBJP2YgQ98sx7ARWZIr5rMVkRaV+VsIyAkviFgF/bfa+Xxy3YgWr8KM5KWrKqwFgq49VyIx8L7
DZfsg6E8L6K66eQaAWDgVNaTHY5ci0PVjC7dGb9+ojWvWYPRe+/gwy2PbafdRGOMfA5Ky3a+aiN0
2QPffDl3xfK4NJENyo9ZCKFxUeuQUaFYwnFHH/l8YhCNippzkSiMW1uOfRIlWSYZslub2xa2odi1
+lWUMX0VJRj6RQU5BKt31rs8/xYhDGpVGSBYt9GXs5owCb/e/1MD+SNLMEiWoOvPeTBmFarw5/bm
7arammZT+KE+YDYOYC5OpFZz4p9CJZ3oos896su+PXIl4OGwvFJnNUvBA7K4MCQaqL2UP64brchU
95UFjeQd1qSEMtZU5f6mewqLzqyinOVataGoBONhsRSV+SeC0+YYrwPsRKVT0vOR0Oos7Gl0FJar
KBPVWt+o0IHWTXBXRoSF0wMTaQdKgNMeVkPHpzP8pOhNHrO2KkNTIbqfv6YTokrRCh90OcORr6Cy
uyVB1EfIRJTqYwCdPxuUGRsaG+p1mD2vt4UMjiyPgIdVfZMr27wNZRQsfZLRx5cYm+c8oe4gD06U
fdZaEINsUeawqJi0aYI/j0MVFi6qvqaUPi+IlO7xIpgNQqzo72ySUuV6Eq98iMJWLRpbLGGatu/U
xiTgesDJi1yLyvm0xy360+OOUUpbg7hISObdtpAhXgDimzGk6Lw09j5YwL4t4do+WyTEvYFmsVp2
fGDL/U5P4r+qhpxbtSCJ823EIkrDC1ptd7wtGI58oA6ZjDRf5LLaqPSyO/V7GycjXrEc46jqkIPX
db3Vlj6HR/13dLHJhRJA5HRQxgaYX/GiRBID43gs8uTcCbDQhaBGOD9O6dwjsYFNgkyh/OZ3RlFT
eiU2Rc07WKK24fIdhThyeB5MLIxDny31/DnaZB/swHKWlqphURPbMVvunf5WcQvW+a9/k+OLho5d
Eb1Nw+fSMq8JkE6UHNfSnT08Z38oU9fJepxB0RPBHXUxZjXZZd+BEe+yk77Ztu55GdfGpHyntNHK
FJUaRVNCjsd5zWZ17DkizUAfeGY/rKLZ4BGrRatge57wHC/Ufu36m9os7mWG3B5P02MSy67PJynR
HqDr4WvI9bwA1B3LmEJZrLGBqulPWvjPzd0VEglCJ+mf6wKW110ITnx05OO79PjAP1YOhTGoZHUk
hz2GpJEOXRI7x2CGMVStzTDUyGnFr85Oj/qNqsIbmx4Uq0zLXwtVW6Ot8MjbU9VVk7KHSLaTgjdH
HIXoReXYRAxZdrjQbgG1cCTZg00algfpTof+Ml9tOfCBteqSLp7+CA2XLCfXuZFV8HgqXlbxV4lf
Hod72axwSs1ZJbH8pxfUbMR02orgm25/WvcESLSvVM0E5gaRdCiuoB4NHE2Hc7yLrH1N6/vpOfiG
EJp9p+raRlDzUpRJUZPpkZXKFX1llUm+PF0069sGWBowfMO/EJL2ZFDtDlmM1MHoM72DY9dHpk1E
6cT16sZvhIfKiFhBjp5RNUBFL5U7aNhkRECbBv4KALxvDjmx0rJ/BZHzqUvkeuLD5aswuEQ0SqRF
zPib+bO2pGKaSY+QuCOBoqg4jrK89QYqVBC132abrmfBTtHTpY1+2DWNqvVVlz0Y06syUUAzIqP6
bT6fEPF1Ip7T5lN+5qfe1Crz9v0tPBk9JLVgWv6OjBx8Kwt+84eYn8vgJLSmbsq03oYDmc5zCqg+
z3C8syq7Vn1VsYW13ZnSWXRvLYUxLoo2HnU2hHWWUV8XPnNjNi86VFOeiGjfRlq+YDcID/zTPxcF
gPIbaagMwIgL8oyoPGNTXaStNJsKQmaDFaAbr/0gcAwtGTdE2G5hM8xC+OJeCAicdrj9JcjSGHnY
p6Uabv96yWNIQuhb8FrjQNX53j0/T+M4mPceHGIRI3qstobSIii4v2gi2LyGVMAn5SkcK29eFm+X
McuobWysviiuXCwmNtj0lCtCjZrhHSdI62HBmgsX7TBEz8o4ipY5Bl9qlGio0kM739f2TKtmP2FW
IsCW9pXm1+0YUJITYB01ioq+zqlWZMFoLumlKHXYXxVfUvN5mFHaqI038QMwj6n3YYJlDl6Eqniy
NmJk5YkNnm8EJrk32S3if3l3LpAN7Pk4wh9Qvv3Wze4pPD2QPKcKrun6GlofCFMovPQUBtmr7qsk
LYI1jd0uhuiNrhZYoV2HBT0v+k6ZT6EZrIn/AhpJVSSRPbZ/5t6c7MsMQ7PGPX7I/GjTvu3UjuWi
lIRVXlVg6O0//OMEV5q0DK8MV1zazTVSqg7F/7T2BAXaYuxuy9495t12Yb21ZSGidVstH8zaDoCo
BYc1ykzZQSBjbl4m9TPbOrs6FGzTVOiXRqsSPhtUfYsmDLmx41i0Zx02eXmQBY1tZsP7VwDck7c2
Y3EMcgcDBZAnKgoWvXsss/muxzRQ/aY78BmyEpL+7mUBH0TS/dxo1GEpK+Ryt8hyASC6Ys5hCd1T
b20tXw5Lolzb3TCPzQVWYkIcxqHLqVCbNtZldHsMJA12mwb8A/XTCozJDIGMQmgxYUyc1m7kHiG3
ibO3hPZZKDjbpgAv3spAbc8/8lJRYUOqC8sEkg4UIGTvohhQkx7ZDaN+qig7tfyv6uiG912wVFMt
ARu59QGcKJ2JsqAJqjot/3wj8C6ZIhcWAdlIiVNQIdxO6LIK/BS7ZF6eYocZQM1uBKtxnqy+OIrC
bfJdq5yrW/9nLmZoVuobx6idqmOV/guiwLv+r24OM/n96RZzvQxZE75cUKfe85yquGHBtupxWVYD
sOzSdBoLD0Kw9IqVWgLTqfbft9suoKnq6vB69ryWc2JQo6vZU9bWWsLyqtOruuvASzgzaxVYFg+T
PSgNaY3In3Ld+/4cE94AEO6/nAaa15rHXWgWRHUuCYpukFr5Xi1VBwPqpwcPCwfWNjZl5rWFS6Xo
JdM+QE0fjSUBrgQTwo9PxL+cI+4FYJv7HTWlhO65t1s7UF/psKL4G3lSSS/uFsFJ5zMbFBmHo4Bo
vh/V6u3+p7mLMBXGgNymwoQ1YQBrbkzoGULeNeS1UF84s7kZh36KnWGHk35mk5kKdzgkoeHgiVb/
NpvaELXjuJWxyfw3dIB551C3It5bGo6H4BBFBMFkj83otqvuDhFJTO88SvfGgM6Vs3r6rjlAqVrw
/AUOLOeczsV5P8pqjHNFwlNDMpvZz3b+aTfkbmre8HNP6rhcelQsacCTKjmEQE7AVIqrOFr11u66
TzlPvJhYFAsulTriYzzimCqnWbuVwY4VHOE9R9PmKk1jTp0k5E/YeSzwqaQzthWldUCIVr2D5aXz
HddoLP8v3l1AtNz03CFrtp6lbxWgURsaJJevH4s4P0nTlu4lz/WJb2/2JZEqOLxmGH4mImD5aGE9
yw2j3B1aYF/qvVQLMMITjI8Lp2Et4veGArBZiva+noiD5AELgLTw280kK/rbRTeQfRsG3OFTZTQM
pHyGpTuAVrsAXPX0LTFEbIXF9i0cmDmCqOyunWt31extAtf9Eb/rhf8PZfe4OuRt5ZduLiUiIxYx
+xUDKa1zuqyxL1NGDIUf1rf7OdyLAuALC+Tc2McDCUApUVNQgchRZS7DHcUDGZOg+D10UeDgJNF9
jeG2zQ0W+TeWR3YA6NajqupoxKiDQCiSavO4zb/f1n4k9y7jHebQlRyr18z1/IDALEVhOVMrGUmV
sp7Kl+hs8FX1dW110MDicGHc4H+sH3QUXn/EOdHrnje1P+4XoW/slW7qMiJF5v2g/lMZ7eYLe+r5
Ct5xaIOi5jA5pzKwopzEKjdOHsmWt6TALN0pFovPfgAhh7A/TIVLL/zqE1dE8+fqTSjsGTlFy7zG
L/ggQrnQUXOxhjyBboowIVwTzdpqs0GzqBMVcGb+XxrfxwhwdXlahz0rvibguaVJrQ24TPSxfg4o
NECTIbHBXe7PaXGEzPzWl9SpsQy87NOYUAtw25O2588iCkPO5q70MUlco1gLPfsRFr4cZpzyM1s4
aR5Z6Q+Dxd4HssDRXZpGNvlhOzvgXeNvZVC10GbrM/TgNSWPlzlV0FmCsOLfH2BfdMOwfVMH8pSz
X6pr2epleVnltqbr3GOXv3mGeaFTeahUIZhMiV+JFzHQfIPwzbBmzp+hOmz7LEp7Mnv5qbK+I/eb
b90ug4z3QxHyAwAV13r0lWFSNMVwN3KTXCfzrXaejT1m/B/OIuszBQP03i8sjBaOUv1P8Krd4ZL5
PyA+oNUfIVEL6QxFO1wrn+LUvJIxxnNsaOS0vIWH2GWnBPapP2C8k261Hc2Bh4+dV83TQO3Haihq
4EVYbSqTI358b0fUeJdUOnnHVEYCgCsaCpNN+ERTpegjLKAL53Ce5HWdrrDL9VIv09AMubQO3Q8m
9WV1fx1P0uLK1P+3bdFL1zF+oAXHnWUDcNcUYmB2VIo6SVVQhcvXfRxHpliWdFkA9z3jGOa4UIRH
rosSl4LuZBFbBrJeMy8Q55Xkb1pUCpG8A6AU2lZAqTahlEfi2LDpjx4EE8KhMurT+kEeNLFEyWKs
xJWpDIRsNfS14GdOlYFEFVys6R40vFp21EATS7yIzcvbtSdsQLrRN59ibjBz3I6JTAcP+l3z7PMg
4QS05WhIBjbHm/I7yHyASt6Vz0qSuHXCRXr3PhGnHcNdcBkDsUzsVn4RPmF7JTyuKM0gFtuzHaHF
/OcYVOym8pHJoGU3GA1sMucCFsOgrLVwSBrmZAG3A/7iLb9EiiDm9tEofo9kuAjRzbwDxvpu+P+r
o1avYe99H2JQTXdmaJwyAjYnLuBxVzHdvHHo1IpEV4GTLeVYZ0CTv7rc9l9oTMxCZpfAcdYMi5vU
2C2D9VxpvQGKhqHdE3pSiNHmC7utWOkmlqORMVEkZ81oeIlwneh50kxwLlKZHmLmPa/zdS/spiKh
AW85AUpEljHTPElmTfan0A42Kafu9vH98jmN3PiPR4nduF8fVOjZBuAR6HePOjW9Y30Ep2vVxGVK
mDKDKzXAkOnmD7deBh+KZpU1PUN/lkYkVoHWvtbq4kKSPqptlHbbPkMLjLivuX22mITKmM+x7lZX
q5IoAuaEGMPRq/o//pKZL1wMh+7yb/Sm9SP5cw+QltW4GGb4db4O3MfN8SpDJbvvK1qf+tk00mRG
vt9TCXgvqFtNUImMuI2bkwM7C5cTAJYv2OA2O+9JpRQNs683iDxGGAOhzUJKqhCZztPA5D75CElQ
peJgptXrHZLHdItU7fnDFMpS5ln5BbGuLp5QI1Tj2H5tsLAdbKG5EUUqc2OmQNqliR5tQc76f6Pz
MnStWanKt2U+neQbXkfemJO1muIXAx6pL7lQBL0ASltbBXoVbIWh8ehMwqtsBIWMhuLg4+YaBcIo
bw5G06WgIVpjHf2t8KagZ2fH2LQFM68slanFy9yVxFK6q99ttSuMTs4Pv6+3Ob6sA9/5H2ulMrVv
+g1BZAwDaQiwYApT5TBwVSbTYoqQdtRW+645fg3DhYQadTYNbO7sGw6Bl6wGPknCyckFTaEeaAp4
kJIaCoIwBcIAjSFYAaVf8lXXruJWhUUSKUkSzRmOLSe856A5Cm341Uj/SFa66Hhbe8AfsPTRYrWp
lyBvb4v04X7iRlmN3vsdLXJibHGpHGbNtcAj2T4H6e6SygZMjeiLhyOxFlAk8+dLwXivUHWiT57F
5SShL5xeKcTEpV4k/YxYiinYJC4+kel0OtrGsLVjgXWQSZLHn319vpTruEJKs51FaEvy8LuoKnc4
ClWyxyF2zVgJXCBL4H0DQMuK/3xvUrLdUdQcMN1DU0aTN7qjVdESLIIbBXe4pfOvUbJhKe99VEOZ
JUItRTTRRfPmiXJskGTCcJvT5ZT1dCC++dsZ5/NtJlhGXmNzTeFbwgzgbBt86HjkjtVMmqJpJzsQ
Scls2QC2TQ78J7ruEevZhszTrpw2pzN/6kb91tdnT1U/l797R+SSlTY8aEuBXntFhtmgjdqMcmpc
8fAIo5ERdx2rf6HJNOtwvY82u2LqTkzaUbj0SkXXc/WXp1mmsixrybbNTK1UFsWNUP3IvPX7YNI6
M1bVXGhB3hDilDZV4oCrTEyCj8NkHS7324NvpWfJP5d2d2LEYIXKkB63i/Z8S/E5zm4nPHLXPwT3
EAhejyNKpL5j6uyz50mzVovL34EswB+DkDYLkgbj3GVd9lHZ4D5XyVwCBGXcUp1qwW2TjIokMUyd
YBL0CoEQdQVbfCDuqi3VXySnOnIip05QlXKnPSBrQ4Q+43B1Xp4qlqWYgNARUSBMFqfOlLdh77hv
xBIzLXnpPVt5WvXKUAYbom9sdkrvan5RmBaLuWVCip4umV7P2peRbW9b14zsfhMccw0k46N1X4Nj
dX0zMobbcHaTSO5GAZF/1UigktShXSDaMo15Iy/lCCpqRdLh99UTEXbXxu6T8Fr47APkr3ZPFiPU
lB4YmBd2X2nwKd15Z2Lky5QktmpMe2mRN6u6ZxktBp55TQy0KkTYcHlUcgJsnXod3lEe1K5qg8+U
4h+RzvykPbUOvelHHD4vU/SvczkRTs5M3R5d2aYUzTVFA2MVSNZP8v33jLhKixAXvKPDK9IKep3w
DwYb9iP2VMkTUW80sUIPWHjISRFSn0+yMbY1ngjDr2H+fwRU2xk/bVG2+LDIzFFpgZ+Lb7lIzdsF
3NXtpiTkLQhSM0xps1ZPHpYFsRbDN4MAyAvlTxyz6Na58U6U9MUzbs8DchNE08+ciFOdSpaXkZwL
8xLuVMzmHvGi2JRxghduZc+vXnDun963NcDNUTGQcRW+JPFEWaKmrp/dabS1uKHI1+rNDA2IeBRU
qGddMMPYnnLL86PD1fslZn+2t/EXsr4VaLn4fKgDW1L0ZP90WeIA0XHgSoOTazatkab93VALE6hH
hzu5VveocculbNwFGg9Ntmw19pjI0oF8WgKOKVQCx72SdSYPdrKs7tCga5wxHRlRfITIBEn4Hb/M
0tcKXaGxnbaD5ScDTJJp/+gOp5Vcsdwi9mdwMRuVyOnhAEcfHK2LcQ2DdGg6M0HcC6O7em0AExUA
0ya/mbuwxqPLl4+zvJakhTG8fF5qrhj46CBK/rvP607eDL7ffzSpS5yfIaBYgNcFUoMcCvOTS1qI
v6Ux8N8ZBNmBLbpa/ED121DV6hpO6V2fVRwaZzBbRw6t1SA7POXcDJRK8iTthskmEIk3kWO21U34
MPyQxOXo5K6/3YtI+H6I1vy2Tkdr4a3n1MrCnGj/MMpgacP6aGYf3Jv9a+Jsl95WEBFne1yArJH/
EJYelBlJVNd9e8x5hnpwNkrcGotOHmc4UmtEfOMMJfC3TbrK0fhdHqt7se/U6O8FXP+qsFQNGdTk
j7jqnb8XQChREGgQogID2QBwUqYkyUByvSCjdN0bME7Kt1AOIhypDn4OA5mwz5z0GL9sH5ScPPC2
h7FOD7ArbLyAZlYf/X27Wnt7DvNCJ3IURO6GKgQ3yrHnaEHbBnv+5i46g4YxzxLkWFzid9xxLBh0
cO5A/u3exKIS33SSxgAQJCFXLQXlqn+XVelv/t5fnNdpU0qt8v2Voj8Ka5nEotle7Z1dcnrFWKFj
wbqKFm3myzckilE7pEEsLcObuWsfPNS8Fu023NEA865dIXGJkoIYfGSO+kXamg6ZjylctYevEm4S
SCDMpHrnn1lqY9qs/zatI+FpDGR7CmMLV6MMq2zmypiQ/Ipb+wAW+CltKOLjvKb659ua/4vtZ2uj
0jbJ/rPpQ5TgObd7ERvjZmOKDkC+8qpK1ylKtLbmpe/VxF6Rsf1eSWcyBy+pufnZfs108pjRHX91
/nknWyQtwvCgREjm98/7DGmrxp15gfEiYs+4VbGp21azZ6Cx4USof8Xkd5qnAYxu/lPRqiRsJREX
q4tFU5pcDZNoj2GLYvWvE9A6VNaVQV2pQYluwbmxOTkDP7xjeW+YF3pqWF9JWV5UxrlSVErGetyU
4NoP3dpoaJLFVgtMpczECEJ59wB0mhpPxAlVwzxhpRndZXWnbKbSVZeU4qUz25qrzp3HmmbgNqd4
92dCceg8We4jp6Cgj1yid9I7/Go1LF5eKmyyhL4ya6i7ArPkZyKC412Ux4mUxO565eaZ0PoCt6wx
UZRky+79RevTQ59/SYKKNUWca1hm7k8ImX1EUsoAimMF2dktd42x9G7Sol+q3CY8/RNmpXkQUCLo
noWgU06qQOBQ7B3Tbm6GXtBPC4F2LrnbegxBkuobVQrtisMElNhdj467OjwlHO7TVuvkEw0IwRTR
KOuFNfuLoZbBIJfhpf+1DiBytFXIy7fNcikzNTpmYgzkWLvm1v6fFvUlCyz2ew6a8/golhjwQtsJ
fg2FNmSMsv/YxkMRTTIs4Ml4CUEyDCEaR1sKA/a5LJaNOASsGmMP4qJ4Mk0djAmj1VPAsEIpfIHz
Fuy5UABZR3HTEfvNWvz7ShhQ3115xSSuVKMnGtBsmSiJLqX7orGMuWpRsaGEYxreJobXYWjo0V+T
YNF5pMoEUFVS977t1NVfB6h9Dfpoem2oq4dH65YfGejGT2BaoBUo3vnkX7z2ElnIUjp0DDSItcQp
KfsHK1YVxbQfAStLFwtEvTo4cO7kio+8e1ewStEXWoOk2yxI0w133dXjl5H3JDjhB5fBX2GAP6GN
vBxwUnbveWzAcb8Pwr4HU6ay84wuAT9YKw499qCahD03PlM4RrzjmnlLKK9iXpWpdqYABDQQQLct
Fkb77yRkJfmMTPH1Rea8nW/9JBE5GOWXN5ZyzK87JqQGgMeG3Xy4OUdymInyEhp9f9ZSD3pcSj1Z
G/6USLfB1tTlWttW4GifhRSaZmALh31erwcXvSo9WmCszn2h1IIwBHDmSV1rilHk1iZMoRzecamV
qqU9XKLeNygVZAHmrGTuARbGj++7mIm4Ts6OWF7E+TpB5BYozGskB84xILH9qCeCoAuf9xZEv2uz
qI+PVusM+YzeKh/0D/Sf1S6NQkN+VWuE2kK2EWJrmJODe/FX+3Bt7YrJZ+MEm/BNOxprkoyi/aYW
khYgBmW7LN6cIzjkJ480n0gvvS5UmuNO7saNUGJUVVhDB/t6l/73+ZAEF3jzVCDxHPTEQ4K3hQGp
i6fF0RBbACvI4m7OsQ8IhwGV9Wf6OAv9wljJFb7DWeQpCgc1dCCIu1y892trrzG4l1z8k1XHBOf2
Euym/NuA/4a7iEZbfIKVC9B4e4+MAwy+JxyoDfniIkVc1Qloe0hLG5Qfma0YKrJlsxN4T1dKIiHu
pFPYdlk2mMQpXtt//CmCEbuhF1/Cbj58ONK0NySW+b/+f/zNOusQ9kGApwC0EjR85V+oEvO8fbEl
Y0fycO3sJMoEzLBtZs8vXegS+9/kPcK5cIqg90NK2F2Sbk9PyMRTjlw75yzKujZJ5TpjmDs3x5nv
xByYqyxHZGatAhcL40WYH3fp4qGRDC15J0zXOQSmlLB2JkI654RiO9bRrOloRtAWqsapvEeNxlYA
0K4SZff0jdhWkeKhIquINYriMZ0ieMKKVdcMt40ulc26DAL72GYxpdShUC72BBsGCJXd6UK5nfNt
vze+Y+2hKciDBuPw/Kji7YufQ+YfUezYosZ9dGumnCKIZwyNFYPLoWn9qRfxlR6XsbmodfjXyiTv
amhLvjbWHKfUbzdd24qt5HGDoWT58gQitvdl1H4yO5tpOj0vZQCZCA5Og2rpnqZxJx34THBPei8J
Efj/T3XJOnwUeHyfCrpEOTF8fB5K/83Fst0/3JicVHLgI+7O5bM41ccdd4fjsNm0vW4881u+Hgbx
fxPLzAwY10gjooAtQGbyZ/G2KRxEDf1enr8fH8gzetsk+STNoAKL3ggutTQ54sKLuDdS+DA9Nvj8
Vdntof53rMuohx4Ev3s8RAnW3WEFTsLXVHsTny0fzjeXFEpvfC9wa1Ytm+1k/rnVc112EI/6aTN7
MxA5ctQuW7FF7k5lLwFtChxOblmrGmmWoLDEXu4hCp95JYK7AZbedNvS+cO0k8VHIRq/e7r7q2Gu
bzCZXSSeUORONb9sLN9sOu9vGRl2VsLrYRPWz29jdUl22lIBeHNq8YmFp7tYftNPndjRwuFOl0NC
3r3e15QRRDood5dSM9Q/STV+R5MxYHY4/g/Ha71nF3F4pmaFLosmuPmBsM6Dtg0UNTnJEbNh/DCp
JWRD0Eq8UVXNxNlJE5Lgd6tfCyl7hPTXQD9UzLqavRWmf5i6Ga1W/V8Ta3eQKUMPunqPj+pW/gAi
yFXkJdWD5X1eyNIZruJ/HGO2PIPnOeSW1JdbgyvKUE2noMRlqmvKwjpT827wolQSIGTqoDk2j8VR
LLV7bk1qlBlYzzX/AWEKDX3oCVF7WTP+rxIo19CAccBvTp5uW3c+LdEnVa0ESQ34RgGSxiivev3X
y227wS2yh7Ubwhs7+yHyOVeFsmb9d0nXFsOJaBG1x2j9rpdPsK+067DCRSQix+rkuQwHXhP/JRbp
0QdM97HoC9PNqhJx4BqTFocGBfXZSudRw0Tslhn91fbKK8K1omikLbqbV2llwbc2hNRU3Q+tx0m4
YqlMEOspTcn0caLP5X4CkVReTeqBPQGgacep+jg61CZyyZmMO2IGIfntlHvfg2ThJDgBO1sm8X0F
ASp7qZmG0eut/J8BTiWC5xtpFyYSCr0/64tOB7ZUC1zuIY1MiYGbPlf4gHz57no9HV3ExnMd+8bQ
I2H6kZSz/qlkJSgGPPizVZD/Gv7AflgrTlve+drpWw/Ngj0x04J6ovF4QLUBwPNUlTBro+P8c1Bg
ElSgHJc0agCkeOeSbX+R0hNCvel2XWxrdhOKq5GaxBYPq485oimcznKBcgUG0a80/2HW9evTdaVu
P4YnXMIwr7XXZeRdgTuGXwPqXDeGZcu4rBjTwtOtXuvKEjpzTKOTPUPY8UeTelmpY7OFkxwmv/gO
4j5YrptjLlE61PnZ8GHITJtHp4eBVPdxBVoI0Z0t5miz5TxGkJkXcOHVac55FY+/lmH8YpXJoSBP
S4CqMl9OJo1E4cNkSoBb8mZg4hd/LrC6TQFIHoAcBsPjBz8TTOxVPZJgSLsZH2lzLTNq0DZfTU0O
oCkhuISR5fAP5VjjG5DSKxa152xYu1JU3PisVn4UcvZFuCILpOrYJvtOwf6CiiCn63cIpbDX3Ccr
MC8MEX0+SGDJ+NsCXZQeqd1N5buKqk8NlHInj03sprJw2IHPV1dRvnJvivRQgrnW/jqrPiMuYZDy
hNnUbEyirfF3YEVuijV1vzt9KWoOuI/vXhRXK04VSYtn2vdVUXFKen91NWyxEf51Wu+Pq5VMG4aQ
h+Np24GrxeFdZs+qHajkEX5Ccs4o2u0OWEO/49dj1N3Z5jqXpXUHtXsSdMVpp+cO+BIE6GzYaDqo
ej2iXN7Q7nvhcrEP6QjkNiMq3JaL0U5UQVU5vV5PgFJ3QRPFDsQmhG7YF8EB53TFnroX1urACg8S
OhZBawNiQkFgsZ9Okh2pmcjdZ0wLMQkZs56K6B2cSC5q5CBvatZIi20xlOvYSUailAN8HesWjunP
RSo2O4tdpUA+RuNSTGmo8h5dNHYuP1ONrLevrbWRT953sr6F76IsEOawbre5948JEOhIF7FFcB5J
lNPK2mtkvYaqa5Fe1bUmC8rLu85VlcxLt8BcsHjGdGSWR7KAkL02Tt5/SE5vfKVXrxQk7QRm4T/O
DKOcDAiR02L9QEiLkjk2mqV2KemPHzhhA+gCVXow8xoqY9ZTVTmmmSJgxpOXCAVt0kdMu57BGORe
rDRMnkXP/WqXj+HeFA4StkAkIRYMdXOM7Wm5kXGg3s5DsEFmRQ5aLCJYkGqV+RDtH0vRaP6W4ZXz
2c21kHAI+yMxPy8aN++tPpR7e6MKZ6gRsOP8Wbp43Zes2uSLf5eI7Bo8wG2lHG6m6PyX3SmKZBH0
pve3URB/RfqUlQtmPKMIPmrz+ddYiZwiWpIRoVeIxLpEY2V5gofxFkkVV4U09AfRkH8yHwqx0cpO
1f0jcp8h615/Y+JTeUuD6XRbfTW55G78XpIX7BU1B9ZmZU7lm6d9lvHetJ6/0R2ArEzZAPBISZsx
wKdk2DSta8mbkMKZvYvxuGKi7/OfkCKrsmIyL/0b3gjsMEXbyYBqnk4DaEo3Z2x0az7+AtHuW4Om
0fPk15sqbwbo+r2TEiJ8YpN4UwbEw6MhExqRG3KlkJlhmbzTsvXD5LaZysBeSYXbVpFPlGVf3THU
rN+msIi61HZmx62w3T4kWkXbD+x6eWwVjHkEC+I/+1NOvgjr8+fAYiouiEhocYTL2h8ryyWmTqWP
hF7yqdLqFeA/5mTL+vpceyCtmUJK8dI31UqDdPjNNCcR37Kb5Qql6QNCC6KxTN9wy+E3fg2kNTSk
YVGQxnEcsiBsED28Yh/oKjSlLHFcV6czdFzATyVfPl17DlGEvk4NHOSR4ztGB2AusDqa5w5lhcxq
jkcmY2ge94x4/dwgF/lKqJFRV5EacoqDsewyPEB7NHhKKlECm2b7LwXXTAhkJVlZYFTC7nSARLIX
5yR8jXHhLYo+pmfR+bMqXoGN2xydGR2kq/MdzXrt+VZUhN1gZPG9amknvERQiwxvGqZrLBeumPcT
aT0QwUXlX0ylbvMn+kuAxkHxBs6IBSU4F0awfYBAd43ChzxGVmRPtTYpiD1V6vbX9OQXalKvI/1h
3VHR6k2Xunk8rufItZmPHXqL3a1clQ4pMsuM21k0ISqcJWhsaRHALrh5ejbY/hluULfY1lQP94Pa
ziEbw4UV1PUwldNw4+9HLV8gOB18zqC6F8czZW0fMIZUbHW38F+F0byPZkCQREacA1fpx3DrM+zI
Y2T155+EnrP21pwzZgKOtoZ4r5wOO5JKRUxADivigUQEvIzhAFou4jna44RXtw6rMrLLhGg8QOb+
zUN1YxDSTpKbGVn65wb0SEJ06ETFBSR+LYoQjHgaTiHpvBXBFIwVSfHuPWf+MppCdff2p0Q5ABBm
iMuuUIsJ9ufBalAG4eIZuza1O7M3fNK0CXTTqZLMwNfyiJkAgq7gKUGQ1Z01q219c+4GNmqb3lc3
h7L3Jx6ClWEelBTAsxWdmzZg9o6NoXiOZ6zdvS2B0tQYfaEwNRQUcIRpm38bSDJH7NmDdB5+pQRU
+9Gv48rbnD1xGhHtZoGabPm4PKKk7AV9U98Kuu1QAvF2dHmE9OSAjtHUJSgK/993iHelpUNfFUse
53mwTyiHl6LzEeAARNNoRXDFmPORqFgivanDo4bNsuXUVZ5asF/uJmL284x0xbM5XfYgECVJLAQ/
T1g6BzKCUpsf9NHZ+K+g5jo2gfQrkzAWSJCTI+0DY6WRSTrrc/LfNRBrbikjxF1PMvZnXAWuiHA2
fj2D17yMtB0ROULxq1h86KqJhBTCyXh+XRXZridhGInOHxEPnYvFmKw44FHFCNjha43+lmJj0WL1
Pvs/bmbysHK6J0ZZ+8+SnfMTpl0+dqnJIUhhnwFOpMNiszRsLfngAhrDfq5v2JujxbWfE3uuEsbm
WaLy9VNRn20Mdeu2T2WM4SzfssJqhjEWbcWU600Q59yOqK6+LI950gU4qNAT5iVmloXf6isYptJU
0WcyqpwznNdPPtz0PbXYoi7ck//FRDi87q94ynhcj3T9Gj0DPHnDph7Cd4pXq543tRBYJko1SfrV
47cqadENkhaJdU/gxjdQg/dX35YktG4UwDC6HCxvAfFSeHvGAyJdo0uRGqZiecyR660c2IHRVK5C
HRMd4Sw91Yan7FABLofJilJoGFpeINjYgqRB+YYedXDjrqOm3Y/TxeGFwpKA+Mntb1jyrlVQPdRf
QFX/ZjFnmNUP1iKSUm/KPbHEKu2S0hqGZEll/YRVPJ505Zu0jyoCrAmxBldQXEMAzHhzgGTJU0BY
IsUOAuW33MyAb7FLXqlNSxv/TkLs10wQZG49jcafJK/j0vlJjIH9YdevywfNClv03Y1HHxD+ofV+
61RIaTMyC8pzIT/7Ko5zUgRKomyI7yeWqD+ITzQZc2stXgCriD8hgoCvN6kgquCDgRVnUxfRuEg6
umbI4BI8Pt/0CaQQZGcuWrHQHON8a3apXut4RbCbMhmnjVII5m9hpWuiBK6Eoh2vfwuZ6ba6mKwr
RjfXq6ys6mZGnkuOO3NIRlN6HMvm/f8eZGMhENAOp3U09Jl1yIuYnqwwpCmAjBVnuUJQf9nnYObO
kTkwPdhkGXn1nXmFqrAS8gnaDRTMHSeOyP3FqUHT1910g5JCKmmTOdTM2Ubb+WUNCtbZUtfmUmly
H8+S0wOgzOhJskKV/Qa+yKKI5tVBPP8QZ4bipKFHCdp6DonzLmV+PlHJTVzWtsFKEXVAxKYQMzTE
j50FcGc1uQ==
`protect end_protected
