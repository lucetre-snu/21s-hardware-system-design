`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KMVw0FCOv34cWOupKA05LIFbQSQzhdC7cNx6tCC7Npkh6sezaILAhlbFmH18n8IdW398pPD6Glkh
nmMHOn6obA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
r2Vofo4ESYu6AQRP7OJMqj48QN1X+bTn4JEjmARwD+qhEKSRQmyGOUq1t8l0qg8qo/ZIs5VwKYwK
blMPD6vM/uEwnk5Wez0Hq/jPY0aEpB1pCERAX2X6smsXJzU2JpDb8Bv4jaiPQ9/mgDegydcxJcW4
WBwS5KXFO7Gsz3oKPK0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pAbtnX8wMTjyj7ktuU7kB3OsG4J3geGiLG/iiwFlNsW8S9qlZpamsi0d4sQtTqmPOjyAT23RYI03
3eJflbWyfGtfT0plGK6bngtMyTN/jf3W4syLadA6h7j9E8mOIobqiQmTamY9g0KJUU+ANrgjfOeN
szhoWM9qDRgcJaJU+Cx+nAY3VB4tTyv43oIrirLgR86OBanyXXakWvhEt54DbM0vCZ60t/V6QWMM
5AfcUu990jo+nQDtAof4C+iUq0lq5HXoPve30kHeLheDubNTRgn2Av6hPjPsQ5Qz0j2WAarM6KDn
7cHfTFTSgsr/E7X2uEKIN/4lJWHSxKUq7PDxUw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rPYRq8HUEihuLW+Cu/YM2rG8TnDS0/Gq3OuS7DyesuYUbl7NRmqXiLHKzc9+77PQjmWHaU9ZJY3w
N6YcIOiMSkWEQLpbLg/pbpfex+DdzHHsSFs08kLH0Aeoi6wEMuwmutXxMSWf8pv2siWUaPA+NGwt
ziAvFi/n69rNrniM8mNc01TDuU6TvFPBierNczf7TfHf/MJ0sVVYEoNF80pmcX5wvnwy8yXBKI0h
aARNqp8ky5v7QanJDB0j6CtBvpVG6YZ2Cm249wygZ8h9+3OgBMbaZZew8UY3M34veYOSjAxxnJQw
/3/KId/WU24TWBYnFoEwhShGNnpuhsluwktCvA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H+vRkXrzIAXQKMevF01F0iWGRI6js2UlE0nDAE6dXjzlLvq3M3TgTAh1S5uwJFclzk5LaWErpkdd
bbGl6vqhScAbxp8N6yS+iKPZmIQgQybWc2aK6E5OT0qBcrXeLI9rd8c/FZH1E3d1/n4Ejgqjikka
Zri/Blr7vecUvt9ENOfmv8I2IwEibXrh+G+e6zXmAsiml/ciKeDtM4i+Ep7eUoVnlGB/uOC8buAq
eddIDAHqIu49VqNwin/vaacuHNEK0yjtupoIsxB8Fq4F8Wxk1tYNf80IQzD3C54Iz+D1ZmCe9IHQ
FU9XI2HrbdiAqeZMEgaa1bJs210sN9JTZGjtFw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j2xQg2iDFbFFI7+dDRrAxN59y4jd3S1Zvtd25yqSjv9nr/Fw2RraTH8/F2fUIIHYeeg2Wby5LkJ2
CgWtYUuRfFFrqGhr7jf8OGrKjgf2FYM2Xn6Ltu9TuJNNkSLA2uR1ibWyQm3uIN98tYI9tyOskioh
MJOMCB7MiE3RwcNOta0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XpqrVh5QI3WGWXCuXjnC9FYqu4ZL7+4Kk3kZlGgM/OdNMMdHTEE+gPHVGUx3Rt2e3mpY35HZ2V9r
iPS63FtPGbct+LA3iXsM8a26Sz1cR3DkQE/0Y7FY6mH9bqFXfJtntPHOz5eKls4LZH/lsg+59CjB
+WIVFVBGt455y8OplHxSSGYHCaWt0qT8zehnOZIx8jz3rxqduAMXu00jSfT3adACc+zTodb96KUD
xqOE3iNnyc0nU2JtLHvtKOuVLitKfLKEzKarbNEZ6kLp3bHG4da6dXCzxwe1GJ+OnfQYqkgJSU/b
hUOKvViAdP+Zre00Dm6xQdH/XIUwmpbDM9wlFw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
DaJbtb+J18eGMiCThqv115oFSAWp+tlQTsY/yiVYGbJd8YqLGZfqabJ8scpFeSC0Z0mcmDOWtmQV
6hMVY6nWFXsWkdPYRsLiz0wBRhpGJ3odEt5HaJrTmFg6isHQqk9SYiEkhRzBnuLmU5UnchMMOQR8
S3uQ0VfEL/2nuI8tp539Ws2I6y52vadcIg1OOq4l7LyBBpMxU7HBYM+EFAsk/XVMIlX8EymSrqDy
dwWVMtnmpaDVN1Lr9FGCzlwLmg8DZjybq4oxlZbOvZhK+FxJxHkiayjQ4+YJEI6jW5qK9B+9W3T+
7QmtppFlAf65jK1AF0LLaLg/QJyqZpmBFHGqx5lKVCtOq5OovScSw2Db21xcZ7J+7Iy1QwJ1359f
YsrsAAYNcdLWk0kB947Yqc8Dwb1kibkD3Xaesa30UKXZUCzO3NFdjDaRu/EYONqo1DSLj2/Fb/bI
fr4CZSTm3ynmEbV/bimdqgziq8XoQ+4ZvBjvaSeNcdmU/k1tbeLN6Vze7yDO92G2i33V8zGZtppb
KqCqSbmoR1KGIfYt6PpJ8RS8zkTFoPC/Jm11d3T3+96DRE5pbul51fJGiRD1hxb4n/8VzT3vizzm
/c42GO132PZSD3DLqqbSon+u+s9KV85t8d0+Nu9Z6nM6nripKg738KdP5K3RR5oAtkVb+ZHGYzu8
ogApTL/4WdPedwF7Iw4OAn6gZ1Gd1xyH/UJw7hjrkBCOFLJQha8I+BHRuX0+GqtDsNQFqmPUGVMN
Wb7zjPFnQZFTt9Tk2xRG3KDZwRuMqPdmctG9uu1KzgahQWMeA0aDcgnH1Pu+fIKnaBUt/PMqwGqk
vcdXS6Pqhg/oFNGbe/2RC63hfvuQtW+zxhmYAY73nEybMBYDcMNPv84vtlyXnSOhanSFNDcE99dC
8IcYQZTv9Sn4/qhyrDidKDiWhJgSB1suR3Q0IFzjSNdUh2nMfKmKETVPTFXhBwbMizH3KhjICdzV
7KtyzUXA5yHal7GsrV++Nx9fHtNvemzDMSIVLkiXckIC7YDlw3AZI+GYkSnGLhmXC8lKhDPg+QLY
nLfpru0bMnObG3wyYK8LlnlwqAl+wf/s5BJt6xIchC+laMCcth78A+iw9diHEosqEwRCEPn5iuS2
XLccwL+8TDjVZT5JNwhPAoikFtqqoWLeyeeOBY/bD+b3SSKUD2aS5M04mAf7l5lHKMCw6lR48aSR
iuSwL+M8dOyF3NiAH6+V+ZQ43tZHIeh8zL1KFYSHfTD+w20U9rahnNcTNFj9kRFXJ/CWEFuOv5fg
Dh3xZD0QK9DRz61YbLAe2oksqcZMHDRIrDyNW1QJCl7VijJie2D5SHKmf8L5pMImzXMKZyFKuT3f
IvDEmclS0kskC2I6Rdsb2c3UCazCR4q3uL3gEKmSSXGby5ZZ7R+jr19n6Pr2a0G9iAfVNhSwU3cd
RThWYx79f73kpMRWr/hn4E4xxtja2BXGWlX5CMlbatPyohwXwdH3CJFWvNjRgQMoSPXREDKzQhnt
0ohrC4S4KggiXrfefbl7nYADWvdxvRA2Ge2iImCgmiQbnYre2bwpU5mIOLb21sf+7O31pxsYA9B7
tHj94dApciV5ZLw1LNpK4NxJnR/0Mu7WRfH3oyexjPsCqUX4Z0BVdqNmThcU7hbCY5CTCNieac8D
4Noh8p9DVNj4/TyPEl7tlUq1YlZmLBSQ3oSQBvglMM/nFQ2rwEJjg+ONXCA2xaQg2eOfvo9Y6SKP
8UIa7jw0WcvCdwNTRl+3mMLiP4qExkypJVsp7wsw0C6ciUl1vhqePemxnN4VGLhh79n/zJU+IR0g
ipz5sj1x+8cwHCznFImMdAxzNk4pzMCaRwCeLkkoypoDY4smIEf2JLN8bMNlTGOd36tVlo+ZTwI7
xMcaJ/TozPidYuGpbVcTSw2mmNvWDsH2S40fth+5mUxrN2B/OeeqyxsLNXo1vNlNcZD+StuW4mGN
QvU5HptGjh282TMlqLs44YuR7hMMvmcaF1PUjJKV22Hu+hT/fhy9hOOZLoyyTTghLWt7GzYK/XFR
PXba6WNL4PMnJWU2DwVcuuObV8SPh1mq7p+BbHWPSbQDi376MEOW1Usy7jN209aZnsAIJlyQou+8
wPUWX4+GT+9JEjRMx84JoujhVH672P7t8IEeRYGQn/tdsBjF+vkSH94CE81e2M+8QcG3p6dALfBm
OqnXDI+NkrflL0YDc2SAyjMd7qYHT/hsz1utJ4Lne5y/P4yCj2/HJdw78POHORP7+Jn6UofVzCJM
Lsur4AeJitEYSThnveVIxlne90lAuRSFYN51xiPmWNZbomz0QM4ovlXUckqzbygJTpaCpOZbrEu1
MG5imBYrkUlLHg99ZZZmcjs2m91OEu+mU6u7DB8a1C0GfwjDWxLrGXUDQi4pAmKkOK8LVNDM+YO7
pfILn6Vq3xBvMZSekclp3GH31FsJL2Yb0HpbY8lvmfJDdSRGqqMHnaPuegAVdpnmmyHkpmbvzb7E
fvIaQq6iQrBnWmyF0NpVCVhue6nNiZE5aC2orDAuvY8PELpLo6WMXjC3yIx+cZTOig0gK8WkWX6a
MbSAarIXQ/JhKUPs7vq46NboPzhmq+x/A9L007+QhdsI5hMOXzgdEmNlhPKGNBoxI88H15/kBtlo
/zibXwpkF/tgwsGMjHD4py3G7HBdH/TSq9K06Z4KjalzLsxJaZbfYKHV7GrlW7LuMhGvg7tHOnxs
wqkL2VuFetJI2fR3r8o4SxIFUflc9aS9J74O+pFJ4r32Ph+ax0iDQP8oFq/ovKmIbP1ZJmrGOL+P
g+78CkFPm4HQzWo1aris413ZJ1ZyvKfDxoMtG+R+8zjyDJ5qkepeqyQo9ZR6zprH3BdWRXooXJwq
RWlM1I3uZYyBpnIFU2d6DQ5RiI53MZU0l7hHEiJLfkkIPwuM/mlzdk3yH5ZCH3sBgyiixNZ5PyUR
hkDl3akDWBlDVt5txrpuOkXzl34y9B+LNhkIKaBIy3dP8GlY+3qfyZH/IS1k3u0cf2EXo8G0hlsN
cOeKUo4gyFN8bOivJg9mViVxDQ20vQRQUzrqmMVJEAuuOD5mtiL/npqaE/rsSz9pgv9dp+Eh6iPo
f8TZ+08GS4HEqLavd5IJrwXnSDEeV8diyo/ofWbFgjpv9m7opksf7cdVAqSADN3WJPUBlf0VEVSm
2pgykYaRvnQ2j2LOekDX2PoP+eSzP2fu6BeMjv3NSUpJfPNbiTbBfMtf+eIiPSwqNgD8QSpGhLwe
O87FG+r6BEfairkTs0/wmRF9iQM/uYToClVkPgcHrNYIYjkJWwVUxWBKFQGVXa45bx44NkHtBO3g
aYl2xp0o1SkE8+EL1anpJuHWjZjGfGmXiemXUrnAl7vcyNC4VnFYowTDvX3NU1ISmoWSss+9tpXL
Xtq57BvtxY0T6E0q/3r0yPM1Exh9qmSZ0OWDK7M41Zt7arHI9SrMJduQGMQVWkhidUP1tlGFdWBB
xQdhceNE59GKazRVJuxZ4Bh/3TkkFnoN50jYnMiZmZfmfhc3phMnBUnmXnd3xPRz4sJAX39hi+4R
PRjzv8xDZEURpFgXpTdP5YqyLu+3Umh2uzEl87bX6nd2Yf9/mMw81iCjcus1U3+ZL6rgiabOF4kS
xcnbpVaiUvS+x9i9V47vNy/8PkAFqTK1CvmIYt0HmC714+DA9iSXV4fHHTionaqTnt3sRHl4rU+z
YYUw3TqFi4j32x1luwhUl//XHLhqW524IZPlhob1w2kmqR3h4oyYjB1toNrA4PawlbFFhDB6IfLi
5fV+7uHHpj3G10nxpKyQ5AF8vmCD/bnHZwa1nU8mDs9MEVjZ6t7hciAi208rBmCgTxoI5D/tQR/q
0H7uUSbMUSNwLyg87A1r0z8ftONK4BPhQB15qJa4Ii17gAq7TanNGfApT/pBU39rW+2vxc1CuESc
sUhOLFGIhOsIm6uaACbWpRvm90f7hvHC/zPjrfZaYzNAK/eCUoKOcw4LQ9X4sWBMY4HIvyNflIjC
zahEPzHUHUkw5v80wSE9i6JIVuJX5dDKc470dE23+fMKQzuzAvFLV2df2/SSabON8lGJYR8mMofC
OKV+mWKD32EF5WSTtbCHfSAjmmZT7AkQ9nX/qctMvrix+H3qjDNs/todsw2YEH569u3QXXsNACnn
lBUnZjZMKXaaoFfyCDLtrfaaS7teVnUpioHYyv7ZUGHlj0P45be1lY9Ij4q3N31DKF8JQdWU6YgJ
vZdwcwj5e2h2qT3dawrOwIWNfXkwE6RtsbF0ef0inah7rUUJwJHdELWg2OsZYDeDEseuojhtyaRg
Pj5BbqX+epwqVZuYSN3w0Zco3TMtKzzJfwVOy7Ou9rwNakbs7p1xeDbQsl5iEIiiDmnQola1IB+d
vxiKEVQ/oB5oUl/RIzKA14nQq3IKRA8gz7qRliXRbv9zYiaSBXDaDE1238ZeGiMsdauKxGslTgO3
FeeAYGFsKkFwyVPEf/hlgiJJU4MMpLOq291Z8d7Js9arADvR6VauBEKwEDs1KWRn96Uoef6Uzbwu
sQyJg3lMmHcAs+T6qWMqITdWj3Qk2TUJjk9wCAaih2h06HlnKkDFxC6AvMPKzPcPnS5UKFxiv7KM
VfDvmUODV47kiBxVNYKnVJp7C3RS4cjURUVn5poxTI5BEFr6cfDrR8/GY05btK5K75zxJxSx/A4b
nLeowNCsn15Igii/cokncnZSC4O5i8wjjFZF6bRpa999PahMiACKG/n5PdFYtR0W3uFlbDdMYtV2
yYo7FHlz8qYnJSURMJVaPlCOD9+L/GUkvUYtwAr1FV7Tp4YrhJfwRnSru4ej8eu8HOZbS3UnwJ9C
Umnrk4GdO2+essVgtquFKQN2Wrzs/QsLPFWHpjG6HubK7xwPzmf7GTkhJkCJzjhZzT10LX2cK4KI
7HrlAINsvEZUaLewKaB64V4wd+zGadhNUqGNjYbhy1XteDRORBDmyOkSvBGdt3TAv68/mHtQLbjh
C4f4sZV4YgIyH4mhsNfR0rOm85ACO9QS5308LhWpCEEA5rDtowPDScgrVMGDyVdM9+M/kPie8Nef
TdwT2BeBC/CiNuV5gK4mmgI1GEJVQk3LhCnIJnOwiRdqTDLDAiX40qAPIvBNWzr/rA6Okw9SLKtr
d4l+zGg/NIJFpPfZuLkde8lXKSXvsRuVzmeI3y64KOPCNLdnnWA2tgZAdnJnod+nr2G1elqHg1Cd
6C55yWnVYfQQyTs7y1/TUCikXfUSMz6o/wmfdH4Vf5ng1ah3lFg3ySG4djuZq5Cz2ckil4jvKfCC
XmE0wsvLcQvs5X9U9Pd+gWN1RUpPqwWR1GU5JAdn5Jk5amS98I5NbToBZBoHxXl72cTvD5Bcia67
7U9ODF3LIoZ7GpVqYajnz50JkrUcFaPN6UJ7J3r/W2E6THmSmnf1FAnI8tYTtxMVn++++y+pXsiZ
YINy2vNFz0Euo9toa1H6r5eFIiFgPcfWRil28QYFF7m1hac9aR3ObYYNzgBFbHJGHeOR27GF0DD1
+dlluKTnDv0XBo+VIkGCwy5EGYe00u77oUtsq7158QXmsSWl40gbAmudFgLdX9rStxXQ/p0PJ+02
pBOov6GNFqxTo+qi1Jp/cljlFkVDPeMqzthaYNSqGskz1gdnLPh1Xzof0uX6onjY7+VgwGGwkf1+
xqiXCMiwVk4/1igvDOqgSKkXot3M5qYKuY5lSG5NHD9OQSfRq2yyz4eMdv65RA3j47IiFIdr2fne
w9wP3iyZvaQPBrWTleWB4RtVgfvESZI2FTa4B5iMup9gJCSpJiyvX7wKOORhpm+IiC+Fvm45Z8PO
gos0CDi/+lkRHDfro0Em9uwuwyQmAPNX4TmHKlqNTLPQ6E08bSmzNYknORZO8vO26kvaASRFaptQ
OH0URzs0C+gLhh22rijT4E5BFJXG64R5+INzQDmF7rgZAZLAN4yl5kzP4l0Iz6a1ZNGBZ3Ia1lzA
3kqy7RvAPETMbiynsf8Hwb3NduxeSMn6jsjNWglC/0RxfWnEj9E3GwrBtMZD7ucDqtEemVKs7E2a
siyOzjNT5zVf8j980hZdcWGXiMZlQUK0EI4TLD3w67tdBDk+SbFJgFVRab6VoFqM557zj7ZK1n8N
CVRZTmHCYMLc50iVI7VYBdAm4tNlkjHe/PbD+knemthDx6xwBUQRX2YEk6IKzCiUPpPhPUzYCPJ5
9EbbigRo4skb9LX6aM7UTWNA1Wh/RQCWN5dRuswcBChUxh2xye+/FR9OotIYd0MmxnGjpAUDaiHk
zZTOOka4uif9KBc0OIhnE6vFthCjOv/vLmXTnGwSgAgs7S8w0wUMOqzeN4Cdrxzq0kLBaVRFukdk
Dk6uIrq+UhaMGcjBGILwRjmYspo4R826xUlJB/ioXCxcaFoCVJJD5KsAL8jK6GBSiAqxCsm8iBCL
VvLd4d5HTZggfEF5X6DR1cYZenedKoJHZOHk9Zb1hOyDFG9J2aQQepUpT+nMXKuPyGEhv6fkjTDq
n3mM5UBfPKOQWjfoYKREYGTD99KMd1EBY4NmYyAxM8HC3IPtRR0L1NiDr3skc4HSd0hxXrgaoytB
k1GHb7bLKFP6JdIRS+f7gC3lD7UcEScovaNtSvBq2OqrhDDa0HaQxzhRMVZ6bbSSEW5+P4/xrngH
ZE2PPpLi7kn/7fvkPvBKYoWBpMrF7s7f7q09Q+1XoJAuRHJy+p4f8EQhISI/26ybTMSEYC0KShOw
X3YuOc6TQ8WrwFgVJsgZI9KdmdO1ZeNt5ovmafHFK6n9nBcPNLv1mk4TiPrgl0xCXR61EtWGa3PT
QTUL16z8pIIywEM9sQp/KnWOPtgTU0UM9+6KH40iOVL1wzMvfwVYjEdx5wz8BXX4/9KAA4+oIPDC
fvH/uvapwrqvCdyDkf3cCHUBxPiV4jStElqOevDPJAlH0J14zjNQKDPuDOFW3rC2EftfUIVf1DUN
MT1tj7z1qAii408rpKYk+LPR4A1bt/L9YJbMCqVxxSAGoG4VgJvU3PznXE+AdWLEvfUyxIklK6hC
g9o0dn0rue8gdiLWctryjhrESMLnetp+jrlQxbUZYadWbBbZBKHskeuCs6lh+ngwavlejIaig51i
9VKKsM/naLErsW15EPRIwXDTRJYsI+44fsQNk9TwtinDEuxruk+sOor9gEcEzJ+hTd3A4bJv48GQ
XbVthXMZruw2j8zRJCqLr/GNcLgDAREMdvSdpip+5nVSz2/5eZ+GGzonPw+JIPq9FouKVXaL+C8g
oKQfVp5cXAMMHrN/ycqEPHR6yg0Iik/7WSn8SOOQYVbkrLbD7HdxtamUuioNDP4rpDlAsSIWq7Pt
W2Mni47wPOsE06qkyAOI9dXj7JxK4O8BHZRM1J95Lg2VjTAopl32KjqL9E4Oub7/XlCL4TTjtNEE
4qqSnjVv7n3wOOVuSoIzIlXZU3DwjaW1wGzhmOC3DaTDGsD0PGlhbyuJGtF8r9zaS6MH6L5x+Q7A
uU983ZE4ZQOLH5fCCsDMRaB9emk3Y+1aS5HgRiSZh9y4R1+avVHgOhEh9WlBXKlifbqKJS0YboQf
CkohtNsCjNOL52CxBqPIr8uXiXp0qEePbI1vTUSuc8FWc37JRo3j3gAt/upMU4qdq/CPjMedSkG8
BsfmcDRL+oFfwBeec5P6yfurl4h3F5jkEj8QFDdxH+biDwxmKHunhmiDyfFGB6Yn9HG4+EMQtiVK
huYvlBHeJJpgheCxhy3xFhcBUPRlsyloaIe/vofdqWSOGqbUwTacZ9u2FF0jFi3bkKQ4mP5pHru7
kbrgEAr6RiSm7wIDpaz04TBdDbqmNrgaJ90/hGgKUkNd2Wz/CsrgIjrCfuMt7WcQf7YXP1FHYjTN
rgnjjYI0zxOVppV6E4bBIiYp+6vNzV/im/LJHWcxjK7LjJa8fMDe8X/U2FuKsB/TdoVAtacgE0Dw
pIF4PMlHZVhUKob9YS5N6Bg76MpHzaKiJKu2niTXe34tX5CLO7NPAvfyvLQzj+9lngVv5p3TTc1w
jcYx8XUXzvrDS/tYQZBEO3fA6+Qh4uoXFFoIdZ1B4pnobfmRW4FH+v1+xyLPV97BqsmHd4h6j//r
Ho2eGKASGUgK3xB7L3uOVRwLIVQJawP/FzC0x92UwMycZkzVsFs7JUu20SVpRwUPNHEq12r7b1hG
UkY5k3EyyZ0ehNncAC7ORhfaJt5UvHgxjCQ6JgmLVYcg3OHdBIrghFtTJFoFjXXlL39A0sDV+++f
VR6EjSxEl66TO6gvMXoNRU93ZnsBk+//8ktQVWNPSMfeiJQMBahjo3+wWCYAI5/ALLBEdfebkckl
ZIIcGE3EV/Su8SK+N6yu6Lxg78dhEaSETF3NheP/4S45J1IR5ZMxFvifWLoMceJw2ogS41n2FE/u
kTI6Ha2mc1mSd3c4vkLPDWxrE0buv8ikI6tZW/hmq18y3Ols6c1zKaMzGD3JwBe1PiIt0mAc4Ci6
RDBlTSZM/WQmYH8nzZZJ0cDrUSDKVYJAFSPw/s/8nDgCvAx8Bly4stEGLsvgwUjAdbOs+pC0iATA
7KqetlmaMOfaHbJSb2peGO+vatIxXI/yTMB/Xdx4Il3RF0GIuDSvzdgcc2Lg6vQrrdg8m8kkH376
bEFozxsh/UU8WB7qWG1eWA/I9fUNWb7L/RHastk3A2zav0hnQyl+TjIziob1QAoRErYyeERMZyJc
0hI401ms9kS/rSE7dndAF4Glnzy3CqHM4fN0wF24+G8+owD0AaMBfc9JgUOFKSorUf6NAhR1Efzy
RitXuh5W83Q32ugBil10gxwvNC8IoTBb3UmrN3mDO0abh/F+I3+0YfIYdjJ89fP2plLddB2XhSPz
rcMa9OEhDhgZd0SFA9gfitnmcbL8MHZw/8TYMRrHp6cuY/+3FW4mbV03rGD73C+g9T1cue87AzYF
RDbRaVywzyvRT7ReKYPc7T13GyRU/C6ax4NVwU+aX4Vx1G8BFHbWOuv6ZjCxzZaVWI/Vk1lu/B5N
nE5yS94cq6la0m5waEZhkxouKcgRGWBzKVT8c9UVKsjmJJ4he+lIsN+908XgN2iYrVCj2JNJYPSe
kpDq9p/l/CW8WI7IiQklWuhDBWVX2/LQuFgdGF68pqQ4KiyikydN3PGQHqElhtKG2aYJc67OB4Ne
WftzJ/CaTZF585NMO8ZRWbdhnD3E6CxG8esB+ueP8GLf+mbBFy3VGjnUqROvTMl3GriT8nsTdjP1
Uv19ZyTje2ON59/tyBRyBmXHZgFsEVnq1jG1FuKLPXWKGMsSQ/07TlWi5fSpZH8Xgfhsp75Io0SG
GFciXY6GcmazYc4Xi31Ze/Qc5WsrKugpfe3uRp5g7qz5r6Kd2vMcXRVVmgJJLjlRU+MdB0B8DWR2
yXdABmF8Z5H960l/jHFfJUDM4X+zYXbaeg8uomeFp9MbCJiJh73djjRKJrCdbV6dTjBIoQFb72H7
b+c5VJe8knofJT+G0zO1WBhsKTYjO7f8M2E5Qn92VLNf26dAVivgBZt8Oo5yBaAsnLhO8k6SjH1f
39x2EKf2GFvX37MkKfx9HG/h36movZdOqNRVjuX/f5wLXyYf8JFcCnRorxCbzlxLhSnmje5i0HZc
cVCqknxHMuHd8qIgeAXJkKX6ea6KJPui/FoGD6VVS65s6KqrwMrVjrbYG2m+YONCdtHC3wwhCIOo
13ZXAWTIyl1TxKMTUBZEqeNzY6ryLR1RoeJAl8xwZiJer79UxCrnzNIJ9PY222jUHT4lgagKA1pg
LnHFILFLTLDvJVdHL5HU8VTDjLVCDy1ZX+54cbTOcwXQIalB8mjrlQR9mrQxHQhq4KEH3g3yBzFd
d95YAR4dLd/Wuh0yxcKYIAiRIXJdJWdXvNZ/X5bYVgpS31knz+dT3NMXEnVe4MUIC//bpaY49QFc
T16DhXfZeFUmr6NNySTCkILXE/Gt+8VJyDbAH1d21RWu++YpjGpKzdw5pBcL0g/b7+QecdHjKjc5
icC8kctjY5Bha7mJNwFGygXe0TNIk8PWbQPVfViLvN+rTbc/T4iJv6lDAGjkb5jjuBkmQNjX3nzG
ISfR2FO7t4s/zvy0ieUrqGZ9yP3vE9libkF4wv3x2cJYOeSa/QOeHKm/tIRD3WXuxxFHkJ0wOj/O
GkGVIWmrEzqDlNZ3+nkRRFKFSEYpBhj9Ac09SodKTVm+94etKALQEq61TFbWeFk0Nt2579U0etIV
v3VjjtymW4YZcewfimMB+BlAro3rBXbfpq3bxObqndpx+4N5knQwQLDWMUU202+s0+U/VbviYcP7
UQpy5PAwq0s0/U3yAni23pAn8npfiocqjH7avRZE9QdbeDZI2h8SWazdzUuPLt04pIiuERQeChzO
+BeWeyKFMUsl8qpTRCfZT9jc9lRTS1XSqmxKVWvpM56ppXU1Kl9qh52DeKPLZCIFM7lHmQrzj20w
EdYoG/kWfBrgDFA8RiaMKcxqLO+gd6engalQf5ZPH6gGX+0grq1p4Ba3S1dgTsuHZD4neZJ6JEOJ
guYbnJUvmyfTNsTKjG+xfIeLqt1CCrcfbw0pS2qvbW+imZASzmh1005Zf68fn6dVrguDa8HN82gJ
xNyJuGml14F+N83DQmYjAqMBl81UuUb1bf4ROt0kL9H+8RlsdKaV9cbE5Pm2r1Ihbo3Jo23fzeSl
A0YvpIKQn//a0n1iZ/KiA4zdXsH1mWAVEViGgwTzpP/WLYUqtrKtF5XGzcJoyU25YruErQZP3YKm
j7iISLv7fp5Itnvk7LwUUpQ/Ag1DLQtd1GFIMIU3UPO1li4JG2EvLwvc+LNXS+fKlcCbrscg2BSC
OEBs0TrdoWUZggqFcwOUChU+mwuJtH580OIO/8j96cu8XluQtEp4gHCDJR8Q/TIfVmiTlLyc0Vk+
MhsBBRpPsA1B+cmjV+KxAqoJFCKnatt/exA2ggjMVmGvf3prs8IkJ8PduFomAPKnyV0HLC8DUF4h
B/ISlqS83erRkevjSj9DlKORxQrQ1vsLUglWl5On07BNl5RTGBMyJO4a1I4bepoFTflTXbwfVGzT
lfvFe/uXzpT5EBsgC0lU0Bdc09UGar8bTQovzVAIa7VmSxokc5Y2QH+x9op7DXpx9XBf+B7xoTZy
JP71+2d75CbFTlh3lwfp9CK19AZW5DsjMdSDPOUq52OPeTq9w+4mx7NrYIAA6c66r5np97Qn706T
NLtDdlP/WXuX8ptXw0zC+M/gle/3a0UF53JyOA45/TwMzXV8TFQ+k5UpisfUsPdLrjw8CUOvgVfO
h+HWJnLHGPNu+hXUCXgMd4Wjd8nojqbNtu+4KR8p9JkhrqrWSG9iv448TY7oPEw8cTw9FJlzYtar
IuXXy5eXPFiPDuPrvbO8A+oZqrvI4kTnM6WwY8YesRtBeVUyM2R7UCUJKGJUpka1G31o1hJjCAU2
iqexr8udP/U+n72S3DaG2odQkQphsPFEPX02rvFWj4dKqDvjrKr4NLVkQwza3heLYWD02kjiiDKV
7ryaTk05QyjEJZRmSRf4ja4gjYZYsGzblNS/qCo6sIti2O07RBQGXpL3vuV54fAydH/0XBmUkkEC
Tvwqp09pviyT2FlPeIBtwn/QT3a0zYEdjAEPyHExbfHRJtuEB6zCwJ2eZOUJO+bwvPuGSDSWRBsu
oII5tantl/zWblCj0wDIiR0ohaoNVrddhmmFeo01y+rdBPSArQEslOr6GWab7ArcTf3RNVuZf4SE
zSytqVX4NkN4OLpLQi58TW0ntZXMcQshTcJhg8GX8cpYjfkgjqQXEYmUSriM9EN/4yMME9cfIlQF
4M06dgelAMT/THkcdlwxLWjSDDo4e5/zy0wr33KZ1/o6C1Up0T82h09aHjduC0sNUWs4lZzo0E/0
9fb0/yjwkadA8uCG4+XthZVY5xDWDvp++eJiwJEYKTg1vEBXXHaG4F15NVWh2qL5X1VYCkbjb6jR
7ItakQMZwLY9WWndB7NO6ezSe/h0iGitDYHPpPE0d2WTAq848mudrKbBH6ce663K+gui4c8yvJut
wIWnXabzUfpDxg5xKe0tbtBkV6nPY5b8+ADUM2ybiQT+tQ2Qj0tHooLmNkebfiwHW+1yf8mJoZSq
zwDTLsSTneNdMkfnIyUYfqmotXhqf2I9wVH9BZh14brNHcWn393oqdg1nvqke+T2gTIRy4E1BCcB
l0dDEr2xYixtpjjCreXwLeZkvCh2Bcd1bJyzAagCEtWHxM2bKKKTvtfaA2fvIwuc1TKzHaE6FRlR
LV3Ga5gen6RcmaQ3FkzYoENwMBB45KkezwNDY6QLcwClsTKM9tSN0HM1WGQjnNCZ8OxNOUkDKbcm
PywLrKmMskDrkFL64KmlINF8V0tTc2X+jvarCIBYA9k+PBHptLbvp4Qba6dFOCi9RocHUTCevPMC
UttCJoEvt7mO7rKuFsAOmyc5eZoUDKwEaR07mongCrjTkpY9fI7ui4LXbVcdLdQe/PtDMl3tI9u0
ZyqJT1mhSu1jt3TXZNMiUAj0kFd2ozpZ+UHAAfNMmfBMuA+EwyQ8fSDnS13ztIx7+AczHk6SeayH
/3IB2brPl9rGA05YgucerBi//+oX2rznnMrrcq6y8F4141oA3Gkp2C7J8k4f9RkaWLmRH/fiWACL
X/TkuzuFgAEK/zlxtjYwva7RnReDHjrZ2AWOqSwX5vK1tqzumaDqTauUrlwZbucCpAp6mVIis733
TZ7GkAqsyCxtvRIgj/BZg83nT3CrfvtBLnwmKkDRjsTkJ8yF93X6Scnzh7kKqLXo3+ZeqoxEEV5d
h1ZE7i2lsC3uyyRJcmFuyd4OypgzzOUuTJB3IxPCwiNRAaAMdc/mv0hzFogQsrl9O2sUOAGoknYR
xOJpsaD9RHp0OrJ4lMhvSUsEkvtvelu5DadQPdCsp0RMIVpHvDClRxtJo4/l5DcHa4N9Rg3zY2NO
f80/GfVlqo1I/8/a9piJMur9ZaFXyS8qpz5PIy5TK27GLdlE6mG/q2jXjCEML2R2A6KvRHsfK2J8
rKHp5gjyiGMS+saKa61uYzxqIz+XfvBng77yeQnXemE1BPcAlaQQvC1jU0H1umpAwwxvyqEQQedm
pI3TFZyJAuZRQkBVXFd9mKiExlZR6Q/Vd1sj616oCul5ZAvXh88xvbTsR28mCSgMdphvXPh8uIbs
yMlTbHpsFL+aUv2+jbEBGd0S5Ot8WqmZIFtAi47IAXBtqCDAmr+juvRMmxVZBgcWAeHFxr4Bi8RP
6/PtzTl8hJKoMstvSyqv4QOpnqgBr0JSbyipNPm5kJJhJG8ROAx15UWa/4GyMfZWHTRAqjZimEDQ
6i6PAEORIMH8NKDRXsMfiVwUZZ4pYYRg7hkuOIV/l0FGZb7MJCIXBp8TH78DrEW88vk5TWf0lcBm
7xFQVOFKXV9CnXSVQ3viT/lw5BHKSXk4grdnKTdYXMfn2gdrjv23fLPWdW/LXvciPDSDNUiJAa2E
GNJXwNIpvqtKvpO//BzdSpubyowAVg/AcYYrzWfMxDClvboMsSA0rM9P01Ze7C8JLMMH5d+P/WVG
sZkHWaDJ/Irdb2jMI7+CX0kbd2sab46GIFYpP11EgS35CFG37e6a3aIZYIBMVPAWLwv5D86ILN53
x/Ria1zdFOwGtG00g1htJ+mjWyAKC5AxXwLw924id1wSoDg4jFW8ZH448qhWVD0Vf8iYT+32KYgj
sqxSCvIbAV8hfS6QRj5IZVLB+Usi/GFPz9wDeTN3Z1Pi5rrD/rHat3mv9j8xpmCEFzDzVImVacMN
6L3hUHfgUcLJZtk57zYPc+MN3Jvu7FuK3PFYSfYjA5cuHepc+nl9OYluDbULDP/Vciuv55Sb4H8F
6uF/agGGXne0Ao2KsfZqrRaE9ABmVRrMPOjKOv8vgpCAj5s3YX5jMjN/u3FKtM3TJejceaRsgUmn
M1tdr/sbParCxos5UZIYdXQQnh+RwNBwePJJ2tfRp/tYageYfQZdeBapcXxqibBggNO1DLIgF79g
0fewm9pYezDrgdc762il27siQ6uSiHpbTYi0UKLv1KD27VF8FSVthTeuwCenGxjdIhPd0bxYMq2D
k18DcCBAwl7Eq73sFVaCcVyezv1Tebz0dkbekuplO+oqVJuaXJqmzfqrpOLoLoghjEs41KGEwhv4
IN6da8Sk2RQ3RVJkig0ess3jG7oAVwoDLoW/xyI2G2Gxm2HuZQRYzWlm7Sa7PsRyoRTZpxfwWEkQ
9ZcuFCg3OWabJkTK6Ti1yiMUMoZD9uosBPYBqvWy5icILZ0+w17+wQVEByFmMPBmlppF+Nc4wwhh
6mL661J1SfFX90ybhtZRMtUr8obQbUgO9ux8BJfZ2NjX/9AAHB09lYn77e3ZGUqCgrUvHXSB328J
p0ZS81/6xLjuyFqPQs7oKEL+/T9pA+dZODk5cwO+k05x8B8ajUDYpCkTDLdtKP48COpN5/z4fEv3
uJcB96bUwcdvotJLXAMOK3ULRAGG9c+stS/6HcpoqeH4+5ebMwi4gQ5YcVGThWEyfNl7ztX0COW2
I8qzurAFtpzE9wbmHLCNMK+VRU3ViXwv/PFZYUlC3dpHk9SpjGZaIsqdgMYrIRgnkupferkBz5zO
IDCPCB/9d1JHC6LpjXzyaATfy4QgEEgfDmCdrUGCYVpDiYpmxxL4+6xOzorq7nw69tsrA2Af7OFn
dbyzRTyM3nlgaUQQ79y9mrPCp9GRLGl2XraRZtz5pW0IfML+NR95BXJoVQmL7f4Pcoq1aCDKNJCM
gsVjoXn9mvnHPRPleUMRZrYc9FuQjuXubkw4qrQQ4QaANqM/EGnM/pu3skgtpwOBvJyVSs+S22Lc
V4Z8OkCyQm5DfmlpZfDu920+wrGgkPoVlE4Mtv2xyS6czRoXm+Ejd7WaFV37IDGrxKrxOqxs6shx
J4QUFWxVaFZN5qEKJn9gHkXXiIREHafFY4L526yB2NWoCZ4qhpT8SAXZCeye+z6goZ5VZLSguLzW
tcdV24Dgc+drMNuGBlRdQ6Ox1C14H7JtH3jdLVBkSmBp8wuvwVngcwmS598V9Rp7Z76R6JECTc3F
6XMgFTv03+MuIiZ3x/G6dO9mkrykeVkILbpg2q7GfJGPebRfZYQTSrO63UbDYIuf1wxSCW6B0EU8
an+86tgg6ajuYxpzzcNdzhRHdFSTrjNBA3Q9MgciefGmpC9h4Q+ipH81rpSfwVx5tjpv2b+BjXUo
sZNDk0uSrNKf9z9T7/DJ24PGv2jq1P2Tu8mLZYSc+MCGa1av1fFXLLqxfn0jjfB6nNCgEWU1T/qz
c84uUUyuhVyX9QnY9VbKblWy5rfE2UqszCkMfAMgpy0RPncLN1ZrgKdDojAQoVVhGCxBRvDcyTld
Rq3VOwaLNc6L5w96fegqc+90XUzdW3fYoHRAt463bFNq0B1gYDj0ovWGmQ9BwyqQzK5TXloSATKa
c8gPdfvHBhf7Jfbg85ZuDOo8dqXwYiUQSakNhaacDt0hoMVjWW/g2JQ3mgnFKMSw5pqjqwsHh1lQ
nxigp27CYBeeQy8JUH4UKZqeb9+GRe8XvLQzdE5vcgwGRgiwZiAiIy4tT1gJfeTzfEbLSXBuqoLA
S78DbVU5GciGrE9c9uxMe0Lmi9H6OD6ezvZPBy0uYw97Z5c0xBPQumshBg/v1beFfUHM+ISRJuXQ
WQAKzvIZ2xGpe7ykz+hD6AQ2mZy097O3MwxFihuThTDeyqAurWFYYN2yfI604U7BsvM8E/rqROgF
23htPI3sXVALSwNWeZWZDaj8FMEoMkJLLD2s3t6mQvVxkZOdU1Qzi014hT5LSMnKD+ktC/f+2AWO
zxkXp9Ii1fr0WBhRW/lca6OXiqfcuvKWQumS8M2B+buRGyYGqoQma6DiioccwhlsuSZyQ1HNrZUS
H5XH3ubKyQ4WA/PtDwOSibcAHN+D4a/rd9OXUVfZgqfgohneNmb9+lq7MQzSkL0oXt3Vkuwl1sWb
PnleWFVTqeGMDmqeemT4xyK+N+oZ9SBHND/A3fGS/tCB/ZtR0kuLTVkLTykX+WGUMyWUaX229PMy
aun0Y1BtmUR0YaFOX7n7sVfMScUgfcoRRAAOChYqz1M5KwghgRRLIDW0qDeO7tZiPHn7mlKXqAKm
HeFPoH2/LWPzoJKpvvFjXOQ1dJJOFP5gaB3mhYgvUoZD1A33AFifkbV2YRMa4/DAqotc2fm9KYkM
tWJzPKUjrHBLZSzOQ5V7QqlYGkZcW3hBX8Y/tx+fujQZEnPxJ1oW515mqz38xA84n7ix2saA7gOO
f/ASTWaQRIAe5WKEyGoN5uQHxJTNsWBA7nNv7lifYNI3BIWFVI0rBUm9/1+06Y9/rurpzsRaxw/z
sYWtQi4wg5lPZEM+FNpKK8ud236shOH+GnuPUGZNVFikl3I3VBxwNBL34opNZ9eaAslRU1UazBwv
K2Azsq55+ERamDg0mv0UYUDYa7L1ri6GFFwnHxm+yfnCPTerGOxJjdzILCtPm1nVDQ4CxYo+GqnN
yISGRXIT023qgTkJwKXyBmIrzpmKBqnFoYd6hFmlu8dDdD4juJBxDP7hr/WcMPSiBmHQbdSouGXz
B6pIAoBvj9W0vxa/tb2Y1UI/tnUFKWzUkFU5Kf4ewuZJ8xmFmFkkJYpVLo0W8J3OYc5mVr3HEgr8
C8KhbY76+8A9qEoXSYguxY0iO7KC/BYhKj74RfuuNQ3aXTlmXKsCACtxwT4fcqH6IIAxvE/2gMfh
YoJw2H3fvu4pBg6A2oLXt8KWUzlBHBZw0IyIOpspwfO7lpe/Hjr2tEfK5HvsWcJ0lDkwjwBo6ZjA
n4Y3v4u2ReMK9Dr0BrxObVxHzE++QMvDDMpOUUCagTLHoFouUlAFmVXETCrRDKB+tM8rAfx26a+Y
h2j5yKbDqEILnmy5C6MImu4Ol9Z/tNupw99ZpPWvnHrWWKRLqVv7PAryFaGLunp/iRSCGquqDuc8
zvpHXtcGufx68FKFvIn9yaM+7RhbM7bU6z4Uc3xszsGwk7tURFGurp/NjLjMWT0JFKM6GIQPYSuR
xrqICOdcihPJ+9yXVDwAutOHpUGyfkIVH5Dwv2X+G4jDW12FLaklV9lXwLPv+ZfpfoJ5TEEhuTk/
lPk53w9YTnHzSRT6jQKDCLshqSRExCnUlHLvnrflquCX9sATMGOJLPZJG3/kup2KW4ACM5R4DiQh
lOSiP7kVKR1R0L8ts6pVP1MKxxyrQPQobjNXYktF3lQPOu51Hro7qGsANN/VQ0ENH5T0eI2eV0Hy
3YbTQqKVLo3+mwGAS8U4enAptCwhQfKGDWdHVaVeMRVuxkD+isI8Strpx9JQhkszUBfrEWK3HOOU
j9VGUP4ynHK080v50+aaZCSfNPzabMdOr86x68CV/2/zV8ZRiDHd+/QnC9VKDxk0KzqzJJQE+uHH
AEeKKFgPpcMbELVvBvGny+6RHazuPJ4zVctZGA2eylwPgngq6IcoCQrHAaFrVD2+vVybef0AEImr
0XWtrA1RXzad0v3r+ESt9PMg3N6tKQVuqvvBARGMZsy6bOAJ7pxDan6ifORCBKrAaBOb04R8SGnT
7rNzW3byX+kwajKpeXMBV0GgZNsSLa9el/vmgXTAgItit1YxMaX9+d1ldVcRGdYVnKTecraWjgPY
a9gVUoLm/ZBUWzvDcGewb86ASpB59ehTP3yfovTvUUpQzlVl3jTPe7sTobhMjX+YJaGpBshg1oZ0
QHHaCtVkBjpvc/RUJOk6kMpihiyqwruualj1yBp+0AcjXy+SagnAKJAdN2PMio71mD7HlwYGtOGH
BHltuUWUIHzlpmadK48V4INkRGkKhbwXoJrXAnmll4Fmur20pNAFP2EC0iCA+tOdbzM9HFXRDLIE
DeJLh4hGO3biZVOSR49zSXvSVWNAhVOSMoFuOhuk5yR8sl2XM5FQ+QgvVEjLXZmHsVTHN4uDhyBw
XEZOEZtJ9LOehDLTetFiQzlz+lYk6w2hiRXNZZB/lxpb588VwUYdQkCnbz9zFcdQFWJuFwxDWoMp
rRu+BYsAaGFRGNPxHqLs5qBE28HI0PkOdRMHKEGsdFInq4ny7McCG+QDU3xQ2E4dJDEksN6H/3WT
G1TIlXuC4bBo+NdeBXHCZ2cAy+uhQGX1XLjQ1m5hYND2X+Ze66YT/ctYb6HzEA/stlBdRRDg+ALm
NAj8zq4JL4hHoX9M1cKFKBG3zp4eqsf+QZBaBdcagr7k8F3yFky4Ezpdd2hO/7Q8t4RpXrsGgqR5
+6zTDqLxsRSyL7vFBzMxpuA853u6kE7pYVWEto+lsiYkD75lqRyl/4Bxa13Ki0WzMCI9zbjsxQLD
ZidhjUXvTZYQgj/Yh/31h5NBhVAl/XBG5a/TdcY5Bip6x41oOxuH/kIiRISDSR9znbs0zdqHSOHv
OEP4lkWv9tQ9CaAPr4AX5TAD2jruGV8aE6gn1bW7yJEBA2Eeoc0EwofeBNOGGmdDq0u3gfsfTVAw
TJKfDZwQmCCtC0UzgapJTcWnidxuwqxcvMEeduhHLNNQ6cEyBWRzTyHTxfywi2aQYW9bJ7Gi3bbg
/JSUOvk9HZ4L4aqf+qkH+ez8NNDv2jfjmXArRRxZ0uVIotwr1+vSANCu18pO7JfDkhVOs/LipoQ5
ikltnqexy3cyr21xYw6hdqtRX5pC4iMvpuCqFREppDTQ/yP7AD43Rp2k/2uijXUHmwi5tov0b/SN
DkW8Fv82rW2vC9+WMcq/1EGs11SfkxnTuI9tgbierz/E6YTRn7EWbUNWH1m+ZEmsUMrL5g/byMRN
9yPwW0jCU/8HwZiYsjZ9H8XIJ7qlp6qPBFOH1VpEJ/R+ZiYPEss+gyyVMQ6R49kuZEjoZO0xZvxy
WRum0dUa+TG6SfsSQpgLA7HBXTLPXJ0NMpaL89Wp940bEjOpABQj4XkK5dC+94xCpOZMy86c4TCv
bu8hK9B/DGMqaXX2OYCUdWnMftg4sH63ZqNnnsHJOIDJSma0OR3pKdKnUYSKWxYjqEcHiOdXL+gV
Xxe94uPvehZT0TX4MkLJh7TzM32r9Wec0Z/ZD4DHlarKiJjRswmY6jhK4LP8XHsVZ9BRgQ8JyBQg
KpYGuHP47ffrhRxLbg3aNWJXiEP3wJ5Tfp1y2H7dRVJRA8T5GMHMz0JoXfHnXM47KKWbCj4CbOxc
2NS1Zu6lZ/4gY5Ix1tRulcHkzF1u8mrtbm2TnUBYhCNS6H2W1HeijXspG60PEmmy/lnQYGancGX1
IMu6OVfFQkTO80HAryv+cJu05rZHJrxiTX+Q6/JDDGobsv2DHEWcbaQNZYUaJoA8b8C0xEjg6ql+
Ice3uprQD3WK/JMhUkiXW8/sOHvzRuKgKm4MstcuRje4lohEWXEkbPzeFPWQ6eIFhfJufpnHZHgq
A2Ek1IVNFbkFJjQRm9Dk+Vjq/xps6/eNdz3r2Kdlxi6tN3TTcg2um5T9LcAk+QUFRnbNhBlkzxuB
5cnMpTSLmojBnUb6vb/zI+RujDvXFUGSM7g19TjcXpZOrOQ4CmWje849ak81QuH91TfII5H9Oq9+
lxUoH+PAiAe9LD/JHGTr42O9x17cRAWRx6UEKV7oXjz+GjtVCovTgg13E9sPcTa01jkFefGVTj+/
mPONhKAVe747f4jB6WKOgzqnLyX+/PrrN0GGigJlAA1htIeHZN7LFAdEU794HBf8O+AtcXPwm5He
qo25C40wmf/Wb61Ls+ji5njIxHus5jOqpg+DluGSEVSjoJltuWUzFrKsHl9AbfzJ6JzKzYr276M2
5u+QuwQ9WFqBXG/rtUJ+cQCCPc4gcz/Vs3G0q9+8EGWwS1/lpiXEFNljFS9o4Ni6xx8I4MVW9svc
DYRHERH3dA0MFRZzdboIVc4mHmwaGSdsO7uBMCQGCE+NE9oywM1RIvrmX3kFxMa1jWC5pHzpL6PK
q2wDGkJQ8Tjlw0pR7Q5MNKvfhh3SqA9vDMtFgu5NW9hvGO1ZAm1k20ouoZlZc1Re+a848V3qKjxo
0Qy8aDb3n8gOGsY+3rbSQiGuSOSVeVVDKV4Fcv7xx6JKUYDhGeT6lZCeieSzUsvuj0mlLYtwzYnk
vjnGUU4eNTHVJF5kANX1MpBUJZxEeXo1iLtov/Pw4BHFpk81L/lFgR81WaSyMNvxSbE2oZynbAqU
GZ6ybYUrtqkUvnAZ37/GedCsQFWdCOPifkt0ZqFyw+LhF/RnLgOz+VYdocfExYqzX2yCsRRlfDvE
IPG+TYUyx6t2JENB4qGHIRhXcIsQonPBwcUSaAm0F5m9oF8rN0LIo11dEpvhnY522lWcCvdyi5cY
A4eqq6y/xeFWB3Gl8vjZkrc7AqXUDHDWvqSkXkHyxF79vECYmuUqEKOZqljR35AEq3IUe8AHjjy3
laKMZWhEAh6il6vBq4A1imWQa+4bvOHlOfU9JJCw5GWsNPThtuzWflR14IvJLJD3SGQN65PrXpqh
Mpu6y51nAoNz/S30YTs+umn7XUlp8ma0vK0fPMfewzUbJHeQJ73G6BHQsdLCoTx/NXHgJ+lGDQQM
aQJ7bRoO4d/KRDpR2YsmM4YQO8b5oP9YXSefICKD9y3JqgurnysnA6v8UZfpZOtPzNzU7y5kIDg3
MqRZK+AldCUIXlwCyU6hEET2Z2s0eBLv4qxfhMwTwzlaNpNsqrSPg7eLdDPaxi0ojcGA0AerHdXR
Gf6oMA2llRKzsF3I0cW7O2G41ITWHRk0BJv8yvGaAsUzAK5BZd8MIvwMfGy4Jv2jmIjNQ1AGJdP5
0jbZvcUpG8sznSo0oJ09mVaysX6o2PDqrOcG4G+f3Qp5nRHZR08Dw7EOtmOqRQnlCbbJjK6ojqoG
LJfmxVH2a8A+fFx3g/wdVgZQmm7pxalzOJWUMDkgitSB481EKSV3iNW6pmyU97A3lxGSLc5hpQM2
HaNiTIgcej4bN6x6XTZS7KVVYWQtyNaCIJ+X0IB7HnjwP63LQjzYVCJLhEueSg5mj3aYOsC7T7nR
s0hauWhvcfkrk9vgDze+MrAo/XmVmBPaKZvcrZlFr3hUbfr29pFGpLp8e6cmdF0TKlu2N+uIxm4n
GmpTCnTOoYH7dYdGI1/Sc0Pjg7wVMlxXWYa+l69dtBNnudmsjh/FqquS/Nn1TDoVYzM1NXC7m9C2
H7NXm8sfezjp+sHEIs/TKseO2wgvaZYojkyHtPYMG2c22BrMM51ofIinbsSRB6rBEJnVtwWV3alN
hrlHtT2v54fC1FFwqgwG87OZpJv6wjckw/d5ts7/nRxEJvBLm2BzUblAJ5gzUW2CwGMz7vxlRj0L
dU/+91uuYsk8Q5ADFhfn6t3t21CUqAZQRF+GZ3s8+93hXm0VRkMfX364RDoQlNq9NNZ5WYJLs2CL
gi7XjaABDHmg3LVfobpM5UMiPp92J1nPrehsypt1FcZu/soZGD3ym27IiCc8TM2sDtqSIgI+7GMh
ggRi+4A1N9USYYBPzR9VvOePw0BhblWDOlSo0Ybs1NSlAYG9TtL/r2/nxQJo2enCDCjgenYCOHrJ
gOKEFsxHnZxwnbSgHXMRxQr3jE/CmgAv6NRc+aCeB9Dn8gTOttDU2aSajEasOWyizQP76eNviTAd
oDeo/Ae8sB7gt2Bez9owztwl58D5ebmCOfGI5cNTbsmJZf1l833Xe4vUYBXHG2w4Ueh5thbr4qp8
PnYbq7yPkVIRzSVBh5lxVw6Oja6ZotT5fy5/kkMMZ3ETJAB/l3dkAnbzVLwN6uruVI+rOnmV1SX3
tgXee4ttRQcX8o+InbwcM9z+53mRpp0vk9cgx7yqYV9JiGOEuQ/GcDzm2WyAF0O1rW7pbj2nek+3
fSFsuWU3zIZUv7O69AyvEmxyOqY7Xe6S8K9x2bLcHMWdrRY3frWIEE0WV7tjppuA2xeTwkjpL5lN
+39KwsLW6pqiw/d6iof0YzthakzN/LgrbG5iyYsKTJPqb3PHJ3CcEP4m9axui77Wss/j+u0UKgWr
zA03Dj2lL09x93eb7BKIrLeKbzhypI/GKmDJnKdFrXPMcE6elFS2T2VBqPVFp+QZhS0K5IhMGliE
2Wxwu2Rj413F9mdzdI2ijAfPT5ZcaAf1tXFBP67NtA+IbruFPcxMuKTpkiJnYaAfKjw5OwnHZEcc
kuWIcjn82tij5/pT3BYLNPK508jScWwWvf0Ea8UOCD312cmx3acBEeE4q8Bwb709GGLZihBA8rXo
6HCY6Wgln0otBckWA/RgXLmSX5Hx7VP4gfmFgO1v3U4OtWbPD4l6XyETdpn8BwY8pZfl+tNXuCYL
nwIPUBfCsRYoFmmY0qiQPd2Y1lDp83zxjVl1CUoX1UiQJw0DzthuscaE9pO8ACFsCptVsZZDKNsd
fD+qnwD8/py77SrSAYdPpaXveEFP5NwUj2BZXsa5Yv/r8Hy6AOuCsD4wOvPiAuC4+IAu/rr1WFQi
1Uzz/6JYD/uSX3IHkL3G2riNwUFowFgBGEyjVBDv2WeEwuCTL/4ejQENa2Qvy+OdXl9Cp4d4fr8K
BznRCL4/JF9EzzYXyIkmdhyEQpE9+q+qA5FiKhojuZ6tm82QdpgPUULT6ikxMyDhxAyPDI/wwyWg
LjfYvFRWlgQW2oH00NkSWkpYOxg2wx4n6WEvlU/iLyi9jJ8M9g2WPW0Dq07WzMp8sdeBpNct8WY8
KRSdaxgYlNoRXd+S6vbQmJ49AoNcjyidZjR9X5Oa0H30T/spT30Z6vEjMaMv7kUxlN8Eo1FjfTEm
nqt8+dJRz12oBqvNMnbMJB5zBa8UXytwJJ9PCuF/OFjG6rk/raabZ1h0XjgqhHOd58HyKs7WTMQj
eIqPKWPhyDP2qfYZHlrHJwJVI2Fp3Tih4+xKkncVR1Ng9TVD0Y/p/cI7Wo5H/wJSGZWn2iZyX+rA
Hjg/AZ9f7r7RbHmBLxyFsvHsBgMQ0tu54R40z/Fsus15P4+KnXrNB32Udyz7HEMzl4Fhch+c0Ik0
fetoIEM0TviRgttedXUAkzRLZfnjqL9m6Ujc5u584MAvQHErNU0AuBmh3SFG4x56/OIAo6dOehD6
zn5xURzS6a7dIlhg6HeFpo08TYvplA4H8Z+oUlWCayM3tdQss5dr3Ttb/ckIY3UgwNrCc5Hkv11W
sNCgn1IUhRGQuaV6aY7mzymNAfgL9BW4KC61Y7h9kne5Opq6YJg0rVKKsTi3flnDBtx7zRG2I+74
Hd65EtuRF4h1fFBw6oARkN6MjBgGG6djL6aNXn853ZxWQq8k9coYgmvEuja1befsAr6eYuNGjpAv
QZyaT09EA4hWna0ZojqONYpEnQLLK0bhWo7rhJ4LM4OefWstaLtqnKvdgYvIWUuZBiYCFhlW4aHc
tToF4eeDhemVK7ePfzoie2aZXoltilS44yWLC2C0OG/SiedTwZPYxF1CzYeUGbGS54zYoTupnV+6
/xCreDPDObJi9o2XtexraXJnW2qxElPZsHnP8WS+H9ttkEL5K8idXSp6YkKcAulKviDUTHHpt4wW
7mJjn6tmX1tOA9/vj4r7Z8rhZx/VrUfCyxNmOXAd8NwU+6VYX6MrUwF0foiCHFqYOt4UQJVWNsLS
F3RF/+Blv03gZZ6H7IN46OfJA6AaUHO2V5JUUW3MLuAynxvUK1tM7uocFv/jaZi+nm2x7nNAfA8k
s22Ww3qteyGCr/NME2FM8/l2AIcgh40UWVPvPF9uGIGJavyAziEPfHfA9f9NnSNL1krj4KZx5xfV
AN0lUVB/fcHCQU+oBCPxvZ3fGg90M+/2S2aMT7cH3ZJV15zrNF58tJHnS2yY3mccpRt1s65x0WJC
yOwknAln4Ox/ZYt61p0FuGxw8oqlTv589sDQKKD5SSNIXO6IQwmdkHjg6c5vSbhwbm8P4wYWoPKk
TPq7VBHbFSK6oXgSyDmHYPmArjDtHkQ+Higgi+t0N4+mOzapIHO08VFaWbv3DXC7GJoP3L+/JCpF
1qLXPnoXDhK0KAmX6sIP2Jlmtc3cLkDFueq8Y/CjxN+rh+3N0EgDCew1QVUYmLPnXGZXxV/nTdKB
JuDq5YyJmytFispx9rhaNH0327Otnw1IHe9uBrgpmNtKZkCbea5ZMPoFIj51I1GRLZJDKsLpACxp
Z91sUCJNyPrH11U8/Era+6h7DfpcfWnH6ka05zPngWPceNbyc5yjaxqfV3UAWjGadZNcToT31ADt
ugM0mtBjAd7yFrg69rRObwrhnFlyHzExUbAjv1UM40pgBu4V37V/BDKstB9of1jSrLZc6L1d7LgB
cL9sSjB8G1j4qJlhG7GOlKUqgW6Bo50/Mv1KLvlHnLmqO98eoj8OAFIESm9PmiVx7T8nIB+uPXop
LEeRIUu/06yypfFJ3UGKF4AwLJ/cfHlqKs9fXMuGtgLEislxDJR+a1sWkFRZ29snswxMBi6i1mbd
LJ5o3GlaKM7JBPmEjNop6yQFD0JKq6KVm4O9ru80veDJfId5CuHDtFej5fl7UiF7rVpnWVOYe/pn
+LFpjWfULdjYTF3thkENKxje6iJFYVL62InvpyMsI1v1Vlzx1SfbhUMUxTFlXIRaZxJ2+86GiqIP
BoroUAUr72KKUG2rCoQWPHCRy/ftDaRvz/GWcB+wuStIBDXYVygovSV3/LFOu6O62cZelM4ZmItU
hrTx5MGokw6jph2f/h6A+af54wV8FNzvbP6nweB4jTf/6Z6e3s7wG2MBuor6N37F44r4VwENmxBx
5Ki4w1Wp0oqtOzXv0r9sA9NU+iz5/U1c5qo605ngYPSp9waEyC8SrgJg9SwxE8PBaeun+o32W7Vz
TUM4cl4XIqNIbscJczXt3rlZo7uTkdWJC+6+1brM2FjUNMUP1YqGpgkAsww14YSd3nCI2qJgSgIk
Iz2lnh4K7JSRKqXueMLsDAx6OwvxKcijkH316LzwgORtbPYMDubPUexJIzKNu8+50k3RgZeYFWVN
+I22K7ovW0S453VcL36GAzPzuZrpigt+7xT8ax/b+09pKIW8HTljYLPH3J/TFsZ4/k3stPx6Dc/j
K+HN0v7IWuRzAfODyEVwkhQ4YVwnIzvqXyDxmaH1y0tMxrS/cZmLHLYohpbyAvgfg9eupQU7lHpK
WZBajq0FPfbqK8x6+oHfV1iYEYvn7UOXHolurFoawKysACTSzWVkYxP34kH2tussZ/nvysKNpJKf
4LOajD98yQ6+lHqMb82SkKY3yOsQeZvo1n+FTWR3Ny1ZhYI5TbW2EaXRDLcrESJRFydF9p6I+IXk
7uBFGLunOKTEXngfT+Otuz5NvJmuGnwtbvkp0t75rpgzRFiq3u1Do/xp7RuvWZj6A7SpyFdYPneV
lKSk5c4LhrS4gyjyyV5pOMKXGAz9QM8v/BuMp/hR3528rgpOWNrY9jH1GcL85D2aNnDWomQXUEPY
OKPC7bnGdryvHjxWjvhCCd8KAICsvSG5lvUPjlg617FJpMSwdyuw7bIB+8Lu4WV9LlEIqTPoQDPF
MBGfueWlYHuNK+TGjTTh5MpwDqzXFhNpk6LyR4V40JeL5X1zL8y+gF/iuyVan5cVwIXPPyuAOXTA
PXW5yHvz0urLkYgYAvbu7JstbfPkqhMEZw1M9jxnBWYesRKU92F0dDLGzOUAFcOhZXV22Lu+ir5f
EAsD+7WYxIA+iQk56QXTXeX2ktWpDY841RNFq+j9RXDnzi/VCJXoTiix3LKGoPGHeX5lsoJDTPkP
4PEJLxbSKQImPym1qcrGUjdmoLgk8SEdrXAhR8AJ4AVRhDtabXHBAkNTqlFHed364FeMr9BHs0KO
J/Jq63TLN6zveNpw4SOSXdu2fZg/ZHSYIjCmNdryHXwyf8qrO5sXV2ltZ0b3QPSzX9atCnzPgI8J
u5AzY/bVogZZRHhOGRFOPXhPEz9AyGuOaNQW6F/2RYZSgNxAqw7AqX72R6hv8x+Hd7NJ8CaStkrR
5nwQsxqmVEEbwvoffnHqUrX9xZBeFyQX2DhYHLp3A4WT44xv1cWLGNGsSwcBNNuhfUjvfSsnq6Ok
o3z9mYdHbDuG+LwPNo1wYa3De3H3JFaqKdzQqKP/cf7KVyhuggvoa2oArOKCHwrl1aTPeP1dgPEn
ZpeEx9nk+Lzpf0ssAEvv+u7Jh1YQr1lJZ34+TGUfQJIMo6qIndYljnYMtGbRB/yMAGkmilCIq4gC
AvNadaf6CZPvGPxTnBE0B5rkDzRFueuOBgGaFM3rxR+dtrc5yI76J17njC+phjeIliMT0hxJfU6H
qh3punVBh7aTLZgNAGqJOx69RC2VFp4HUavNnXt3eievj1tndGiYu6nLAI4v+xvJQsQFNXIOKIFh
NoFaLKfci+leFYTx+kR9Q5EQfTsThWnd1OHpTDRz1sAOT2HeWqwP38Nlxmxmkm3AMVH2H3pfn26X
b32QFvaoOPXVLzIXq1NFbSzQn3Wx/txgBPHr57aPmhENMmmzJzHfcTT6aL5hWhJ6SbK2nlSwpmHP
kPPAZTw0ey/kK0NSg6lwRtOjzxvv+cRTEkapiSri3WIJfBOl4vaUHphToq3DpwDJYx8Myh6tu2pD
xXkTyV28UCdTw685pLp6LqXV6v8ICVi8XjzWx9zG7D4P2/JRkCK4Y51HCoyoiSaeky4NSxf9xu+W
RKvJxaCBaGio3iLNkOv078elDcPQlpJQB/TKpCqumDTzgllNM0qtXBbMw19JZCoSM2om+zTK9gLZ
qGQTNyNisXatQtVeuWRAcB7t3hQCOdmRdpW/9Ag/iPryEq7kJPUoQff6SJ8jCo7XtHfqYsZrZVzE
IylNqpC9CECrSDkGh1QhFLcuAwLhnf33lvLL7hcq39PRTpFpX6N0uXYNMXRMROvd0cBfBEGwf4N2
22a0jy1o93Ya+mi2nJrT12TfQsNz0eSKF/VJVoNCkqbfWvAoNlvNpwXhhozJMP+UQApm2x+YO8eb
7KB9wQ4pclDF/9RhSxGh70te4REhO0vULk4xiAHCNcvY/xppJ5OP2+IPyIYVncd5xaEuFJnFhJ/4
LaO1u7HxMSqZG2CPtxVoK5dJdGHL1aTKXLoaeW47p7yqnNYYgCVUCvBT9jUDcjYj3YIC2thfCv+U
WoWTcp6HoBE+WbrfIkDrcap05zTajm0rTOP9oZOFOHd/B2nFPM/wTfGpGrskh9njVuGCreang9Ne
69lmxIw7Fdtg/23f1z1y2vzclreFpsktW8bBISs2jxmJ4FEOQSjB3/7kdHfR4H+EItghExT/V187
btnDO+c15+vx/J+BxzUm/wpvptak+HpuHKWjQHXe4u+bZU/Ii8gX31suo5yf76CVw5cCW5jlZpP4
aqhMoBN+H0FbA2s20cgl//pv5e0O/+fW3vC7KFvaw+/usA3Thi1aK+NLYvVeyFnkpEEaEmctftuE
Aqs1v587SUHeuYopXyB7lZVaG3YntXvNXUKlc73MxhiW50IBblvL5u7paLUoDNKidlR31K3vEkRj
SIZfo01Cftw5zc7fZ2OHGrErd/8AckVs5/buScE/Vr5wwHCYJyqfo8F+JMvg2Cof3dicYu7Zk9Pp
l1zOIHtLY6DNciYWENV1TndmNdsLq+Ij9nLhHnLWgEcGwTfXfGXRsbB1gZpHVdm3tqSkACgJLAqt
wWXDdK1x3h91DOGKSbK5I+eFcClsDg+QjxfhBqANG+G7sLHC4Y3WurXvCgWfURXNAWtOZmveiFfv
+RgNZxowc3vy9Hx4wSWKS0wwhY6A/Rs8LrU/KU2BiuPmQq/gPTcYJwVTDBVwO/A4hPIfTTUV+jkP
20/wlMEuBhmYKeM/HWid42DV0A4k0N3lVgKWaOkmdr99swXqoZl1+oGMuxwEb+WWA0GbzlGFqUvl
jKNBB1ClihzFrUA3DJAdfhd1DfM+nhsgmNfA20lBXM37BJGMHcKQrCVKQxunTHt+ZFdQmM/OoIV9
gzwOQ2Vwk4vFiTcMygJc1hk1EZxz2A0OwX51a+kWBTjVr6r+1K0hnCi1Sf8hrm46sql3ABZpyXkd
nt1DZColV7z6wlKJN74BmXk/hJfxTQoJuwwDmi7J2qlS/gNMZcOc33NYkKXgEvQCgdvkVfXtG0Cb
jqosEVr6oovTaUEKMaGWGyt+Gv82BBKT5XEQYf5fqb9jpY2P5hKxiAKO9MrSqL/y4GO4ZWlsir38
EUgTjmIQKD1zn5IepOwHsjcjysl2CET7WqZlXSpUsLDIutisb09sf8EuMKmgl++W460EzhW/tuFU
W5+Xf1uvEjMwLTHtYsgS3Izyrsf7Qj41O1h0GEvS0CLW52kWMfyzgCLFrY2LMAP3SNJM1JpZ0PVz
XwhJRcsm2wkfcivm/XgUYHuv0jcwM/JLxccaH7MnxWOpB2Lr2hBVgjqyET1lTAfuCQicClF+4kdZ
K/C78Ky6H8b6NqdDxaUJpheFHXGlwYkPRgP/rT5mqIew4dGErRWBjsgyoHYYFt1KCYilaStK5j5t
x6tRWl3XLx96zMK0SM+NAphXLxvlwPWQXPzBQATXt+65mNkyZ8yDUEPYpA6q+2QGnRji7roih+OM
SIGdVpkZP9tbbNeo6YiVA68gNbIVl7Vyg/MvP8g1E1yg3PAC+Iav3cQHVgerPb1f9Fm7nd56Lo0R
gJqNSUMxt14Pe3jq1Wp/wG+PhQ7U/Q6N5/CfQ16XtqS+FzSjXN+pxy3ksUdHFurmbv2Lmz5PGBgG
uH92//m2ONCBZX03LHL4QeeLM15jPUPEoNfNWUOL+0pW/t7Rwp/B1ST42NQUVre7K4HEvUzb30pA
sRSqtGEpGbSxb9X2yskkh+sFp7hmlp8WuuIkePjfD3zN60NkfLeiNyBz1kN4+SZ5t/Arqo/NSb4o
98m4FzX8d9wEvZytHtdZGkyI2MKQfC0Lkd5SREGbVVe9HwNTVk8mYjKuB3Zz3nc+TZePEey1xIfE
OxYidtlrIeHyPWGtLVmx4qrjMV8UfL48mMnPy+r50f52Q3nK5qVeQ7lVL+nQLNy3tgXSSo23BFyP
R3KxdT1NlsxMa1hfkMkbnIM9debW785v4Hxn4pmaA1hweTbRk2IGZa0ehuF4GlRwx59AWYkOLc//
fXZyyIaGZ/ryRGEwSpcmIlhkZuA7XzHGlHlnAg0/bUIKiAfZ7Wyz/jxxGHcrGmaDf3AYiyZAK7mp
o95RS9mkwEfKqgvv2mZT8y+zgYdPr5BEWG5Ew0b6DdMlD6v6BAyKra4DKSBgUS7mL0OboMGTFHjk
HZmSNbGiBIhBoMf6Mwxj9oW0QR++u4d+DMgWr5sfLhmCFZwn/Gm7DonoA2xmCxppQsIlwPrucwlC
gu5aJMMHq+xmd+mBn2Yjix0WlHaBn4PTMmKmkHOpR3giYAQj3Wuum0yTy52xWgPbeP7Skh3AGq7t
dOSXK63FpoahLsfzU2Y8QZgGK+6FRp954bmCkN2QBplA7mzhujDenthRC0/H+scM3FjNAVyQjBv1
cGRvihvCVqBE3HGTYbIQ3366H4ixKKbuU+WXyJDlf+rLXYMTWvwsUewC4m8wX6QZOSm5rytBz85O
ZKnR0kekkOslSlleqdFtK4OVsI+ne9ZKKPbUSP0s6RL/0SJYqraHf7J94Fh90nnN120qYL5IXDTD
nU8SEvruPQpOO8H+zgowvpqbgC4et6jF+p46XthMqqeoTeYlM6MHqkxj1upoCHeDOfg/eimxOHkU
1jS/4AKbitpEpubGPmgrAOJhRVLXuwyzBUqJRfNHuffxq6SxL/9CxdeXefimQkSUmnE5AM4kp4eK
YMpk09y1efvjnPSboMUgtzeMYJKg51uSy94Z+ZdgN2kqnyxNjn4RA0tjC5oOhTShvjZWsUBpKThM
inQMv6E31WYsbgpBVP5Ts86EXLATkdaZjVp9zamrdOrf4s+dxbkW0TQsld6MImJGrLPrIMDFRhaN
VNhrU0aHq8blw80KUhOdOUGuz5+GBFHHKwZC/k/+PItMdJ4NGFYms1GjWMW6mzO6lD0XVEARgvmY
mvYnlLrDAmxPWW1cJmfqhJV4m9q5i3MK7rskpeel0FYo9mfOmtfAxJveQK6VxTFDM/7svJLpDCGS
DvTFVrzY9n63h2hYutzaiNZgOL6+AFApxiiw2U9nHZI/MQ1nguzzBTHEGU5YrM+/u/itG8PqmwzJ
5eOj6iutBzX+Io2IGBcksBWiA4Bh99i/0CeL+T4VGIIASq0qc5eXxTJPLRhaxe0/5x5BPhNJjZxr
bOVOFMV7RximJ9/Ki5E+ak3zQO33RxGhTetvgAyCZRPFvMTfF+uOPNkcKWzbjwbGR3JVfO2wIbte
ghcxzJilmXQ7YfA/0t45wPX1Fro+Nrpoid77eoqqpeSdoAx5SL9cGcDNv1PNCfCBZD/SvIgxUyWe
/cZQn1s7tfO5LlZ+fbhDNurL2oOdmo4IGw0QChJNNH5GD6gcibW2ztIvG2o7khpS+oTpgKjq9GXW
6PsWrdKdWunn0UK1YsH04BefGMp3KCFE42GJI34arXDFeJTY0nQmUPSzzVcOyNnPM5zeJQSlSkg3
l+q0l2EFLzclxj1sZ7MbVmZlk3BCJl9cANpdq+pkz2OsXMcAhmvmpVUszUPQme99uKZSs4XNn8SA
Tx9qgSxU+mQHGgWwF//PBgS0IzvF6QUZWxiXuW7swjxJu3k9LHLfdEy9nREe94SLV6EMuhmR5yYI
Llc1Ix/At/pQbroLLbRizPzOfFWvu/uFk9jSfErRJoGFv8zib5vd0lT5ucNYn+hubH7r5cBW1OFZ
MByi+MUp+PXfTxsywZMrIW/KLTfI2VHqAuXWCb70cxadi/l+fzwABazMgNCaoIzfJNOaW7Db79Ng
0RAk9eAo0pIcWT65qFxmFnmeZO5HnRvKavdn2Gw7Ku4pgWPsMXL9ihPzT01HSdmsDGIYXUdr53hX
jA1PhwJb6H91amNnuDxpGwvTc9vmYqvfcTz5gfpewSAuaceGi8XrBdgzXqtQMKPJmDcu3Mfx9nME
cesFEN7NaPEqCPiwJCv58MLcPreS7y86gYdD6AlqOCDjD4ZSEP1bVKUtyLybB91tGtaY3mJiIX7j
utY+Yie+JFQRUOd6S06ugVZZO3PKFaltQxjhvkCkhcMkH0Q8eBMCp5VIYwsI4GiHUAxFeiTLDU/J
5H0XQMY7dvbgE5Z5U9Wi7qmkZjQzaVDBUPGQs+QcTkmdnMadHqDov2O6yBD3RlZzpHcYAFmM35z0
PGZdJpiOqhhf7whcvFHKrCAMA9JRN/pqJfa5th0M7KRdzly3sxbwgj/d0CD3AdTQmyhn+b797+0U
cK8j7K06ZlidZCbTJNuRwUoNVWZ+6v5zddnjXawNRh4+Uy7rQr1NQd/2nerOAZwpoGjru3mh1lLF
0mC1uRq0rJG3xvRRsLkTZQ5METBRjHH9fSejGO9aNhqsdkmNtDCQtpQpty0GkQ5t09YmqgInJJVm
1f1sUleuw8zawgheG78xGJ/TnmOlPuqYkljsLCNVMrOM9CpNQjODbfZXfWYFR6ne4Yr4hWFjH+NK
DFtarNGbpTOarIRRqGB2nuQEDFl0UScAlvhCIduF/35xd5yTxf7Gq7FbLU4agScg0X+LKzDs1cp0
U3WEj1UG4UFi5/Cieb5tPG7OvSocx3CO39X6xhn2VEiuFGUj5kglvRES7zFaJyWZdqd/cJjR2Cb0
3DczbnEMh6X/ySaLdFQWK3FIgI8DrmoAiDUPPj8xx1MAdh09GxERluoz+QC3FaOFISWuVO1OfBnt
EHRl7Z6LuNmxl2QbRX99eNoZqH5OlakuwnVYyL/NTFRv9Pcd/evufKHWmbY1j/wOfe3az+BeF4ln
/foe25wSuEaZm098LWTJFkvImwV+gOXEieehl5umoJAEh7kybB/SZi5LGhk+Pm7q7P8vKoRAISv6
sMVKcMMuu/w8pCMK+P+d5X+7O5ODBH62vK+9VCWORdbBLpcWbXQI//d++lRu+50mIcXKaeIvV788
KEUso1vO8S9SYmKDFaoSEKYPIrpIFarllHQDWd+naWkHrB4x0gWO3IUJwDGZRccFp76VUcrlB5yf
TpJKVPlAm2nXLx4SOj5OE0sugQtSC9Ck0xjV/UrtrpClUoRwIOgREGx6POQu267DcFS95jL9O++j
4Mp5q0w1onE/2HfMUZxTOKSVjE447ztdC/YsKOPrsh/4teFuEUJWKZBiPxsiklurHK/Sv8PW68BG
ZXVvnJN9TS+B2AErKWv3ccndahzRG+H1eH7a411520wweqoWu4gh25r3kIP8XMrp0Udi0SjuHsZf
FRYDFBPJW2xt6s+wDm7Ua2Wys6iiejxrQTb4KwCDD4Q/psUkGM0YtEc4ghTYZDZBPqy/ZiD8Q8qO
+qe9S/vG3ZOpSpkn/0cdcLvxjwRrK48fB5KyvH2kGHbT2ERxhqJVSx/UWxH7kCDiJBoisajvn3Wo
5Gj5jnpytKqrMTdjAWB3Ez3AKSugt3bow3pG6kbu7OkqoYvche1Ioi1iwzH2c/2wCjSouXUVI49V
CT23mEnr13yH13SIBx8BjTpO0CyJ+axiebJjpAY4PCzHrTuoXEvdL269FEBPAdygc2XCQM1nhZO8
GUvBQlKGX9impNgoKwk4aZnwOtEiVYXoGNX0dvc7UlGGnrpaAB8G1EwBJTzht1vVc3TI3YS2fuKY
TlRIqOVOknxqQQLB/sZf4BdtXbtisyhNvasgZ6WCGrrzi+l5T38iQIuFl7kCl6pGY96lfYJ6HPaU
XcJeLkbgGuTea4CRUWX4PWNMHWV7fE3rzBF3YOK9BDDh4G1uPt2ccnKQTZIr4vlSyQCfkTCGk6Ej
XCDV7oQPO8R+TqxbrgHkAzPQqxCwdboyC4+W5/rBVekonCPcsEYF+KQ/shp/tthzN2lPvSNKT/hi
SvLWAb78RyM9OV+LWr481f1X+e9yqBTtbcaJlFCNVls1d8967t0fQHnX4A6KM9znhAO4I5IJclUF
r3SlJRuSXYi8F6Iqvp+4p1aCUY8VKvtVwP9OuO4eXJoEjheOg6b3nHwlBNSn2deGzPCmFT9nZR/U
vcwW0SHDHJHBePIYqUyCe+ULPR1PUx+fHIKbknPjwIpLGQ2PTM2gr5N/ZdUI7QRHaaDUkd17UrGR
c/o6902TFkkLMfdO2BLwZZQmAAoMHHpcCGR+rcuWpPibpMTg/XHoQ32ig1p3fEUAwinOUtD3nCN4
nNo6L7QMHCcW+HSVf0A7/fPtOKkilIXAKOiMU0Eox826g3GLP2+mTKp/tcmWSbBIGE7KcQ086zbi
seR58KFYZXtPzFkgJdaCrJnTI5VOVb+VRRSavR7coxCXwOnXB8+qzgAGfBvaRTIg4NdGxg+OYcNV
SpyNFJQPgUJYfJi3SB6ag/9H7Sx5047BQIlmNR1gHbS6xmKtcXbU/EyfUhB1uTaMBeQPtbhdFG9H
wZz4LuksY0BOE+jR58k03MZCNDz4gLFrXCb4heAZdimpwCY8Og+tzM9KAQ/bZCjTMdgqfsBkaGjp
H0FOGZr8yUk1y0Yn+gtNK8GzBTne/jVdkryvuozC6YCj0cXX8JTfXcncFaeSxJC6GBx1XeOQNvhR
+UpJ3aPwNsl2Ulbgtb5Ry3hGnvi5Yq+fDoR0sNfEQXRKZQHOuPqg+NxR4mk43Ef15DcFfiNly4DJ
DhVrGPfjUGOy0RkVsuoq1uLMpswmAaJm7/510iF69rm6UaQQtXiwBMglWC1z/Ul1VEUKQqSZDBiy
7qgSf1NL5CzrRArm0EwnbRae9iTCE5nYqlgZnqpXCODDrfMZdrksvEahywUNrks7v8fVeGqpcCjl
YOw1H55CChNZvfRX4jzg/Pacorr4AgmOYZ7U6OcmkVWsm4nSmQtENF1wFJCoUFdCcamBvvyfrbuD
e4OJoyQJmEQ/0YefscZaatWZTpMWd2tDfh2EDApLzFe4dQNo2K8YFYedvuifx9kSl9Kaz+NIoUFc
m1VpJQk/rrZ+K66dHFX8+5K74WmUKvYmx3oEW4qxuRjGzBYa3GV7/gx6z4+fe/rJdi6ZAaw0HZpR
NXOi6QWzfOHWJAEf917uACqliPkTOoIfNiwjOh8McjoiLG1YhkuJvdktd4MQzWvzZ0ic3H/Y20Va
2GYQ7Xj33AmNFnOAqc9aq6XLJZy6k2GABPWOjGpodKfqLtqDPhFIhbdgMFgT+v5Q7oicWvPitrKi
OMrBO+0f/xnq2wJ6xCaYCdKQn1nBOJFrhP6sLgIlwD3mXGRv2sEszLC2u7nmxj0BiLsyGRvu0rDM
DbN68NIRnc+xIJNC+nAY79S2o9UnwwdwKDwvY5qCDyjGgqPSzQ4WlkeFrpJKXL5QXydP2FsrTIgB
L7QloQbCm6IhGmhHpKgYxY6pOECYCwfG7PEQPtDyio3MTU0wT10o/E/3liLDR96o0FTr1bJYDT78
tue1e/dwCOpO4nL4L3dWhvua6NbhjPdaexbNxfWrEWIubVhqDv9FuLQncbfBEbdE+7AR3G8qO1Iv
gsSwSXm4IYbZRK1eUETtRe+YbKkohZjj66vT06/fijI4QbS26ymZnbmXRJ9ikCnteS/FN0ky4z70
DkZ5VDVvdiOlHVP0FpFNIT+24VtLpp6LH7eKhDaWeLtvRGGsPAEVIokOV/+KKASAdM/ARqCd5ir1
gvI9XYHy2QPAu5Yih+Z2FwY2KSOVuwNhZ+OstG6BlrxIH97aJSJgLCNI/b9ZVdt6oDl6mxqm1x4H
EiDmki5csVfWV3JKERafGd2jDNRz6KaRP7QbnamLCCqEBc/4Qzc/1n+DV5Us69UFIE3a3kL14duA
pY70HwV6t9mg7nv92AQNg7EpKtCx4CrgxxOlOXMFSL4YvG0VNJSKomJ0pM2Ywp6d0jdMQFzKucvu
P8CvRmxVXZUKFdLKdp3oCTAHTrZUfAVq6aJnaaISSn8kZXfsRqi7q1OlJ+W1S23MCKKYx4rsFr79
FUn0ou43UqM1I72Hpo5wKrb3BQynoiUiqh9ZSPyWVGlExsqsSJ8h0wb1eId07bsjk4rz1uW+sO/s
tuY+Efw8AW61dDCMuPGgusDdelDt56cb1rjuqgPl3ZKY72TDQgOZP3dl8lIPJq4/yixEIEh1JBFt
xh9mnOxvo4clMj4A0lyVMW5pII3I8TT2rntLyVi5hyweMMjIHa5i8Oc+34IGH7D0rsjfDN872NEO
xMVF7pGwmThNeIoHAvjvRv6LNfHgFhVJzBuB2Hrrm8sfdEjvTdVdnejJndgGKJxGDxoWQ1iizzB/
NCAmO4WkV9Xl6NVGVfI4te8f/vy/qsLv5Bk4gpWWbLIFRey8fMJeTF2SUJ8ZN4/8HHd9XVkW9VQU
itMwMMu9SOUBAn0RPMteIXWwkS3wegwrhzUkNS+lM2646HysqowO20L8xxd0KYk/wopx3rYSZxF5
Wo28OarHjZomzKYlRfMD2xNMnUcaqtINqLN1gtSgLVlB6vbAAJ1xfJ3eTTtY/kUubtR1CL1g2Utz
3Eg875qKfe2dCr3zSdukD0eh1Y4BPXuECpGW1P4EfGVeVWNChCy1BwaVCnjnn11uchHdbwGYE45g
CNFkYE6FXaITVAHdvSNP2/SEDlc1HHEUgyhWFHrS3sJ8cDipTphFdiW62kEdHqOQCT6O7mTFibwI
QUhqwVPrzIkkIFg/OIFMlrFI6cPu0t3Zy9hm6wbyQCDxIXaElX5mgWaUTTT/DuFC7mXLJnRUsjSS
cpvmHUwDEr2S9J2xGgCtuxbarwjXye1n6/WMVEA46UXOg5MWqFnDHhwpstfhOC9MSEiIURAMPo6o
l7eoKWVHXpESeCMoYMEgEjd6p0RwGHd3WsbgIfTBtXmMTpdlFffSW10kYK0ElmsKghBXL78PWr7e
A4fGaQXA9vHEVA5t0VD5KBD6xDnsYI6KTWF13Ipit/Ba/HTEr+khIajwN7jgXT7wY5Ox1WjyhHB+
+QvCEpmSxURB+AD9pS1tVrPQnllZWKk9AX9o1f4GEcz6YVh5voaQQ5CluFqFiOLk6ZWSNnO9jCN0
JnID1vM15B5y7Lmg6EqqPZaqmrmXoZ5LSD2gFACqKvCLZ04a59bBtdkNZnmqvtF4HkWPGwLllokE
6d5gv8LPpTQlScEe/idBxY+GxYYkQqW35NvpYmxIqS/39P/GdTeKeWAa0yVvrDikOFyUqW55DF7/
qKTtQAMPiRbqxuuzoGK/apiq1wFNDSWU0skhxBNW3ar5nQdpTgtZJSgBw/rgCNRJYsQEisrswTxo
hhTNKXdMWPmcBSUTqVDgO1XZ9EIUDVWnWGGHF1YbQAxD62plyb0rYjWtb0W+W7o/gDww+SBMQOzg
CuRz3Rs1njKl2s8+AT/Gcgu4SL6TPL7E3zUOfUrQKB+KyXR7dpjqtwJ+REzg/Ac/OATnWPwNJuUU
G28pz5eWE0UVh0OQBkeWuNFaambtHeSwZDr865rN34oKVLAonYjUhADtgrteYTyAx/7JjIxxkVYk
lHtNK1glwpL6lI4tIDYiAnRd4vf4AX5/6Wn7betAIm8QEdYrT+aFN+BimanFwabbbcnZv1dP5DWF
+/4H2TinmY1yeSxSa5Uh97unGegGqUpt2P0B4pZ5GkEW7ftHrIEwygOCtNBjEhnUK6uTGReaHTsT
9HE8aVQ5xe20ZCn1Zy3kilncxm9bs5rW5Zhm23bt6wrA1cfubTbG7nVeU9Cwf8KtvGjPKlPSG5Tr
rzdKuLhMyv+ckKYjxCoMVtKbtf1Z19micVRkLwfPZuWSxoz7Rui3etS7eDSWXiT0nFjoxGy37dAI
vY87l7E+rPJDrzqahCXekn5uBElYqrziohLSUeaR9i3NPVQeem8LYZXxJqJi9ySYFpGk6N0tLZVL
Uj4/eT4kQn6XostEUn4lRxMFHi8ZpQ5vLIAJZNHVr3gu/jEPV0lzG03ZX9/2PPN0vyfqCg+J8Pt0
7AJUjrUZRZMS36WnfRspQguZ+CBNy813ZUiEzAZbYYkx3gsll54n086K9+01g/gVmQbxfAQMHWt+
z7cmDfPC1IXKVfGqndcfvF5yObU7FdHKZ2ddjbUfBUE3+SLlbvXVjiMr7ISL2MUaPFc9SEcUGVwg
QpFsq9JWPzlK3nr//iF8zupnuToy4VYtSN3zh/J3ZZfziHCqWFFvUG9BdyuyYmrzvadraLfIZqRV
EUY/RqlPdhDcB1uTgyaT40zfh5NZ00KSewBrIBfS7jQA6cosSbM9+GL4UH0+urkygYxnJZ0xjBgF
1H1GfpxmQXCnp+8I+strvE+i6IR9WaoYvVhh+c9p15DvwD7eMxES1pfXJb4lV25n2dOGNq5r1z/M
iWL2tsiUqy5ztJDy9JI2bOMYpTQH9okq9l3GZionxzQGXqV8Jg8DZsUS5Y1zg9FgJcyjD7iv9uuS
Sl4oJipYEyGpKzsPIbCwHDP+fUbOUHADfR7c0y+wX6f16PE9qr2WhvKjVgZbA8plQd/0EQRWiEMA
agoU31xqPqV2Bjoai8e/9Ei9tYsV18tm4A4MOYlEzJYWsWotE480d416ASStVaSOfILsokgak1Fo
ZVNhTGg4QZkKm0GWA4ziO2X6RPvPT30ewLnE1CxPmziAjw03O5pt2xazvz4SBI/r4vOHWL+lHrnR
2+jdUyVmKP1xGbT9M+8cA2I/n0WERTwVa3XQZCusHjbKsDpeLiuCZz9OuUnmwTefYklCNzdwFzVs
+yxuwSN3Kzs9Eml6Wo/zXY2ewQG0AzAJslnfsfh1vBD4BUwaQIaZeC1wiIlYkhovvy1RvjhWBDv+
853qeDS39UuH3JK+p8nhr/bHO6fiBj8pvxTcqTSLcw2ri9kPuEKcb9n6oQcBnMnTVPv3eeqDESsL
AGfSzxv5hgKWG0VGLFNZ9vFJCKnPTL/evamqQxT/pHpQ8jPNN6kqHsGWCnCk7+EC6LegeAqOMeDJ
rWdMjacRezEjQsFaHC7c6PeAWchNVofAzBQWQmPAY1HDiTMJ+6U7KESAiQc/PmfUujy8p0Ei3ozC
cEvbYa+Ik9Q2GnYG4WzDJ9ggdvP8ZyD0cYeQLzUPyfhElTz96dx6Mcts3Ochx0b+KnLS/gqRZMXv
ZQg3ryfW5fjrvYQN6xa9J13oEpsG+CK+5mdkmgZoD/fmfE45uTl977uZ41MFZ+c5HcnngYgsfMDW
D94yX5+n2o/sorn4t9SKsY0N0Q/lrBzyISjT9FGanWfh/hq8DP4hG7yjcHdJKSCJ+J6x0eTyMh8K
nwq0I2uzuC2ZcPT8dnT88ajwiiPJmBygMKe2ClW7dlIDrrCTRZF8zsqAdmNtDo4QEH3wHjfaH88S
0g0DUvPApQQgUrMi7n+KNL4upHDqmq1R/1FJj81IpT/YYVD0ln6MGpI9iUKdRxF98GnV5V7+QqG+
TdfRkh2zxyAdCrWgHVGrVFx7RtzpEMyfiNPuDPFHZ05LBOKXw3wn1p986y4AyVCLstfN0FvSEyAz
5/iF3nnobFq8YmfGEXVmbxFkMEdz5ijytaWGnGNBB4n35CqMy2GDU0KgRxXyfOWVBrcaOmGE8cuH
5qJeT59nyQJfOgEV8ln2TScx8/qvwq6o8bf2mnae/VOCOXiHkYZdiM/p4NP3jhIPFX24JGxK4a1U
JUxwQwx8/NXFRq9Iju20EN5+yDF/Fw8gS0n3dhcXt2uaToix+/yqDZW/n4Pr0b4wDeLmxVHw+/JQ
Y9wAQwY5M+x1Ai5sAu7KI9eh7Nj/W5kpyI6HsYkcrd0UJZgkyqH8SnXIl5DFrZZS+wqvmULTrxFi
hzWYZ9yKzGY3+fMfG6c+4cFrGwF6RZGj6meleLJuKgLTpDqO3VAsuGDgfTgs31VcV7b6Q+81Q4IE
H2YdBiT07MNMC7fRxGUYn1t3WLQAChjqjHclTLq373+lsOX9D2EnfsORNoHWbxSbaHceSZDJ6ips
xGn9/GUwYvomxXbx5HnuSwcEIIeYVFMAocPUOeV3uUyjNoBUKnrsKt8d3XEmEGdbKBlVg95m4Q1y
PSX5Z/+sNvmMVOSslDF0IvE8LbfYKHflpS/f3QKNVvfUd3f5M670JqcV9uYr1agU9g8vGrBrxhen
bFiFlyEyF3FMEL0ghf96kFVPXEFXR1pbO7/B8cxt3eknwaXUtAp6IopBame9zvkfl3n0dZu/hBAE
GXd+6q0aOk/4GnvHBnpAJII8VQPb2RLOMWINtq3yyrQvtZQKfzq1Ob8tQYWMWRLVfQtfOI7AtBCO
dPVcEhY0qPZpu9e/JjYiIk6PlvxAEs75+Vq0oItlDVB+7iBDL/zEuF4VNGHXleT/qCzXnqjkSEx6
LLViSu/3MxgHhsEZwqJx245BEg6FQlLsZJy4cQIKcdXCLevUA4d8jbSIijE6rF06fWgM/juz2YZQ
B/4q1uw3Y0Khve9E99kuDKYiV2qFwQEHX4WQx9FBK+ICxYRaVNhCTXVtMAs026mqjk053TavbRCh
xBGUbwYeBtIXx7w7Anh/WI3hqp9qaOcgAuCmPYtEsa0zVliuoxuEi2sD+CsyrduNBd95JVwjJ6Yw
LUpf6BOav5j+4eIdvRxyXFzLgF7KXLyxzgXFoOOPh2pqlbBiRStyQhP2XJIJjhqKdV+VgHbHboJV
fdvFSAj3027ayIV/QKf6P83uhfYfSW008AGqXAzoMFhAnffQt68jo6x2tL8D7qZIl9Hq4c7fCbf6
sslBQayzjTdXlFi08cHptPvrh0mw5YIYet7BfWjeRd+jG7NIEEK509HKenq5GHdvZkCTMlcm+Xss
aaJyX+UvU4lj39ovC21dCRmM1IQo83GP5lAnUKFYnVMsl7EcvkESEwwLmLg39fvC7yMXhgzhPGJ2
L0rQNa2Albyg7MsusyuoxQ5mxXM3QYvgiFtFAXnUStwLV3bRrm07rgNPsGCiIlmMv8LXFH4LeH88
WwHQPreIfbBjc6e02rAy2Pd3VYiigdQ0XTtADTCelYFErXAwk0AyunA12wD1xkzZ0kc6u34aNlx3
GUfz8JFkGLVZCnFi9eFGnNbU1CkZgLgVtaVCxiBiMwrMbZLcdAKjrgRxzfGUVWy/rbI6KOHPSclj
Y+1FzZJcC5SrfENYQBoyZmQxgNRqwBekDFN3oCvBjVb1tG7FZkQmG33MN8j/j8SzyVo6TBH5A5vA
Qn6DnXq6vvwcT9wk78+Q6uowVF2+t362g004jcbmH+pck79xUhQ6/sXJSewjg5+WJuKqNoOcZlMj
yZD6Cjds6W8tDuRJMv5weXp3wU36c9Ek8hIsbYKKVC7NrM/F5QTSsj69jA6HsUs5OuD5b3nShbb5
XdEr+tTjzt0s+2KTD44H6cUm6B+/2m5jkRebWtIVS4zgxipwDKcAd5KfxH3DtRTzjkU6FN30Ig39
cOKAyAOh6jsrFsjJ0378fyHnDNTbkBBl51zEZubNwjEiP1EEXLR4nyqUbuUYhIy6/xYgEKPrQeCO
0W/O73Kr5JJ6SzcCN7i4xAA2LAWK7x3kQ7rmsEtAazdNDyTiwXGDPW6PomsbFLgp7vpXAdt/J7XU
s8a0oXYa8Wp9x9dXFasgYUjbo5fPNKFMlRTXJUiEBMCiH9++Ojhc0XRvCllBMK/lXVK2CAseITzz
wxHHGZjIXHSGfwlYpRKp16IVSBJ1v90uu4pq1ueFoKw218dcdKctkg079JyH+sXKHzTd6jC3VrKE
bmemSYzQAIKBeITtw9uWDCQ9RSKIhzqQxPB5fzSynZTxUdpjpoKWOc9xIgDr8jeawkVSl1X2sMcJ
deKfyzau+aLCV9zDe1troKGf21s145AhMrfk2WBCGGaXFUiOw23s5fHg5FMfofZzgq3u23wxz56N
wNYF3hlQYGoXKc8AZxpT+c3je1MJJELtpJdCimMg9kzi4UaYuNWGyNIVmEkgyuCslVRS55FSqJAH
xotIDxhUB24gUYBx2erf0aYS3B14K20xOHBC0BDCucLvmvjoKOYn9ChD3//9PG9IVy8thWZSO9Bg
t369TaJk0ARIrJHiDsI7Ipu5Dp+vuuIeOiRc5zwKIspgHWJzCel7mFXZa7RJZkxPv//05gp06Pzx
Vy0sb+IudkYfrNgbQ4wp5vBrVgZC3cktJ0cd3ixWvSwkIo2hnNXvCWw+rAXkce0+MLK4170eye3r
cEZ1MtHHCNpFYENt+OD1a0UFCll/skv3L1PGoaGKoCnK61e3L3QwLZy0DvK3amNafxRnidHa1udp
Ajw93XLJ1EOx1lVKoSEICXmwa4LlOAxlJD95Z97q0E3MivSlK0iprVMFu0SD2JBcjqVI+VAD6NKF
EiDeOJJQiMYArpUFzVXH+sPuksezVDgaFZiFK5v20QZv25pSF3mxpS22qBXyNSdqozpksVhW8ywE
dlLEboskUp9coOFGaJQeiJNMuFA3EQABOVDyycdBB/niUPdxzPKDfYA+xQ0rSDTLKyvuMO/gz5Cs
K6M0hkjLbUkY4vp8CADZHoobzuIyVFPKdpzyYVOcdx+2rQSvUUsmHAXYrlk+8B00HBQ04mBzg8T8
qRDNP1ARW/lNz7AoQ5++s7ci+XRmoI3R/PztUBsihv0XDfA6PRZIcxrOYDQFq6BfbHBIJNEGAr0d
8QCzKpxhxA10ufItEmRBkswdTlQiylUZu54yXg59GzBNfzE/V15reDwacRKHzv3MpHKtBB0h2f1m
SiNvllS5C1pkYCjjb2YU2rp0rfJaTI363KBreYuXI7AUPSI0kdruVxQu9Luyirtq1aJWRQXJJA3C
b8KuwAOqvUg+WyZJI+8AOums9K6AdCfwFAx/KQtOzrR7Q+2OTmf0zZvX2l9Sy7TvP75LRcGo9F3g
1clv5XbBX8P2VEduFY25J5dK1pQ3rjioKY7jb7OutFoH2C9dVqEaBadDwMlhfz5ibEOkNsD+yv1r
IINZMtLmTyzXbcrjk45Qya1N45MKSWnaTkZ+JYLvkJvt59lecPQhiwLlEfrFkoRDR9ygTR4bus2i
xXSFCwcjo7WP0IwMjHEXNbRfxbLrvTXS3wVmIp3cZkhyKJdzSqbZJSH8MCcDc6vFZh6jvXp/88pa
jRNm2CaTva06DD+30efliTaYEGGgRCXHRmlWCNpnX1lrVUXrC390Q6xOTyAjz6ho/49Qqznns7KW
aE/zrlXWbmLhFF/oFLvMXL1hDDjf0EKn7BWm3IAdsjOYaA/5/qd0jJbCJdRz9FJO9OJVUNnYDVeh
CDjYrXAln3vwf7jr24vw60vzcjBCsf2ONDHnzem19zsEAZMcBaZTo966MNf40Oj1EBdTdn67jtLO
tH+O8M/0/AM5k6e+ZXZHmNk2NzjqLbn2rK82D1g0v8vUtvLrof6GzYmEqTdyS98G/KWeOP8Yf5fT
3lo+gBt68Ia4gZRa9QOAD/7tYEuQZB1LANkvxIO/dDhE66egyElOaCu0Tj4SBZaQiSyrrv7HCz2b
hWKI2n61NCCXyxcDE+zaO3LTtJiOf8dep44UE9lD45RhWAFf1zyjOmkdPVAgZ9MuNTFSHQ0aB+1c
PeIrzCG663ONDGE4Alui/iAUDEbQ28///4AATajLRXnZPGFw5WniPwG/kq7zGrdQgZlfIV2fgtFd
NEwSoJwoyB97NDO2NGjL7/srZmC1mreaUzJnvJYAiM/HfvlXvU61WpeRF7cx0qd6nqLV79g/Nuqp
T2FYn9KP30ZxNenO+ZxIW24ZdSAxRmENFhaZFfxRTFi0W43M99yfAmODd45gDjoqqH/w2SlrMIVE
U5lfhEprQI1vIeIeoE8kPBp2Fzfi4/3a4Wnf1hGQu+YMYbcxdTV6NePrOcoWvy2pImbKGOEn6F2U
sxDM0LLvITb8xsFGuApRa23nz9BoS2UedQEoBWWgw6E3572c/ptBzaoVGI+MRKzT4t6LreshERE7
GgvycLx8SCSjwLAqZdBLkicJY99aAGaL9mZd6HkDZlwfUNezJqF8BO55vWUaAZaK8OSl8eNGfL98
3OVkJcXxb+EPolxnT2eCKFMPVkoJTVEdq5htU57iVnfMDwmeC+q9pN/MszK1d498J/WWw/oipA+s
oZba/d4+7zfr3VfB+Wyz67z8jwzMnKZui2+sYL5VS4vp/4X0c3lrH2oo6dc+vpmXqDOVXhc4Q9xe
CjYE7v3KOf+kxfU+DveIhBoVQNhJ3IiDMy9q8Q7noS8+hF4BDDDsfJMiPupxs+IQhu+0I+LfKnk2
gOBwDnVTREnqu2JUDlTpderoIQ7sAymUTuprjyR9z2qXXP8VeTJkXc1+KWci5NMYBDEBkvDGcjtQ
tLuaRp15jxDTiiRtvVqSiqNMM8u5JYrbVwfdOZVitOsNmn7YNXSEyXu7j8VmFKFS8J5jEt+k3N0P
FlIV0Yk2n6OxGhN8Dyp0AXMOsbN5vVhYz8Zm0GHEVQ2u/7dmapJNLH+AZ62RH2ywucbUoC1iwDv/
4eO+LGqqo1SyaRXZEKMaxpJ2WjqYr3wFUQdcLsIhTu4yhylQpTzVJVrONXi9h2yURQ+GMxNuwcBn
4GM3QMPsne7uhSOXnXPuyOPWdm9/zoqUU8/CL43TjShZSUeNKEo5s6hZKx6XVpwHTaZ4ybXqcxxO
IHSyp4zrYf58b9N7uhFXXca8E3LaIe/WrLI/JWRT6C2LjwluAQLQzXCLsIqWEhwAo5wfpY+y0xhs
ZnzM5JNeddxAgj+XOBOiU0GaLWobSap+PSyNiVfMoGKvFS8Qrh6JHs4RfbKdidxqbRtCJQj8rEWZ
fw4HeN42uL8iqrY68DDSfGyWNa1SvhpJCTWD6PTZlEpPoRc+jGoV90QN/hmKsDnZRLyQyUObCwgI
ArfhLpcsHHf4OqCOH894t7Z3rJH1FBeG2OCgX3OoSKTk+INvD/BibQ4I6yZJ6sveihuH7/4jJxBt
kaL9HrTFQDodbNmKCF7eE4xuvlJyma2pe8sOycpeMA6HPlpGTKqLy3gTy/WMYEbcrS1BT7mHks9z
X6oi9/8/DgL2IDkAJM2RDmLvj/PVYnuTqxft7dkWrpL1p1OyUHiYzNvhWFsW1iQo/6O+6m2wt90C
ZMs3nGsh9ZLA1212r6rmrnZwcnAcRyYxWlRqMNHfVD2w50Jf+iFZ+T6QBl3JMXRtxvKpgagryz0t
s22uMCiD6J4/jnHzqJV2aSconlvujwGk/WBq72NaySrkLMU2Kadf1HD7neebjnD9kU8A/iBtYRIl
FG0aa9GHtGnXi+58dU7OiKU2Jo/vMSmIqdy82xfpIO/MuEH6u8GvHqxRdSUiNrAi5f8/uVKxK7qF
7eYJl1CQ8CF2RWejwyahdzs8Fl0+ew/wD/R4K5izSc+fvF0MnH5YeUlxgzwyNfEgNFY00Mdiz4/Q
RPTmN7P6hCgUIivVGFf+J3OxhTGzIBgsWmm4VguYJ5lHLuDBiWANGNkqImmG1j1MuLdc/xrR5wvc
D7RHy8ltIkddAbp5ExcqTqHiFuMJypCMtyPa6jP16cVoju9NOU6/XOVnqDGa2sMulLzV0j+SrcCT
ZhbvDZFpnfUWpZbLYomh4tarkoJdoIYIhAp375kCXZ+8iiR/ZD5DE8g6XA1n3cXa99Ms214j2J72
gC1Du6bGRsbRGvafkW/81HonuWVv3tp/cCIedXxO8No5tXIJ5Bxgv5wo0sUIiZT2oUPi3tc3sMnF
3tbPuOVzzBQB5lZ8nS2XaI8Xw/mBh/ckPOMLnbumI7TQWHedhqoQ08283e3E4n28WMjP9CZGAUGz
ukIex0RYXI6T/xNJA0r/e8WirJj7FSytPvmph5VCxphfnGm5BXCr/Tw+6F0d+qrzWjl8IrwgnQak
ianWoR1Q/OVCa5w2dd6OgDer98ZL0NVI5a6XI4nL1nLSuKRxOWazOdSpVrfLGFQwO5iS5GRUECAo
Hd6kQOk9hW8KfJTpKvr+5587NudqaOzyofAuLEWjCricq77LQqClfZT+wSHcz8fyt4wCdvJR0ZOM
r7EB8NFm/vFG+C9B8wh/6+Ag6FPFUpTL+dnDMe2OnuZ2gNf8upeYJdtszl/VoBH+jTidMHgbTh94
oDNeVEuOJ/UbMxL75iSEa2mEhvZdFb27HwMalAFn3vq/m9SUYCofNxhGFe4Sk4You2oPemjUJnhQ
t2bCsROZH8OVS2uRIdSzMRTLy680ik7gu7s87bY5H8gibaipK15Ag8B7ClDWegzhkgYS7OY/T//9
BKcjQNlqY4HnFopDkAUltk5goxLHFurlQurtnbooq6LrVBieplfGWc9hKPGfl7gqsYq6+yGs0pqb
33OeVDwj3budrpBihlIde+QQ3Ej/SzViqXG/0TZeqFv4u7mEsRdJZW2f8b3QLeM0ySzgp6BVHqvq
SqbWJL1pU4WljhrysQwo0jsBOcPvIe+hO63wySvzv7gKpf0OmQY1ORnqNSuDyMY7jB0QUF0zA75J
mzoYcKyiXAHomKZD/Z2OP834zwf1ypJx/bVbLfAlD2dahk56YfV30vn/Bpkkn2ZV0dboPrVRGS26
e963RDE+dsZE9b7YkI1TQ6CNsmZMofPjFrryNZOWQMIzG/zI7kXvZjbI7NUZRzUfHz4KYUdSafB7
Hk/k1Qp+upjtsoHq8IW1CFIrSHLGP0sr4GJH6Qo8bD051T0FR6diPQVFC2cW/pp1T5fXAgjwKNey
hBG4xCXLDnUdk4LCb/KmEwoWIBtbD03rXsMnsfrh93yDIRWzgwypbzzZVwcNvN43uD6zkfJ940Kr
kiYwnSqvb8tmkvim0MmCiJwGpfYra3C0DERqgf1wea2vBCQFQ58xAaW6yOZY5LQC+rsk8YG5C6gl
8/j4loLmQoxF0hmtBG/VpErXS+BxAnVPftQoyFvbq2tGksZKgL3dnzU/r1ugtxo+vidgGvc/9pzg
Uk0T95FVO82KUfPQ6qvCM9luEk+Zwx/jY6vMEYteXvwgEKEorR8zvMIg7aQHCTQzqREHqhZCiDF+
YYMhEMoiheREHm45baZSqFTFTcD75svfkZqyDhayHx7BVrxbRJ/wf5FNvnehoVaDqpcsuheUjgtY
k8I98KcXFql9I63tXs76sPrihYUqTUD5lMMPtl/rmSn+xHhj1nXIVvKFWHGopPIQqJ2kuKxwaltv
rODhMoqsBagBFxcoLRJqX8EkHYrf87KEeRiOoFGEZl9l2ChUOmFIRPkFT4e7asr+T7p1whrzw8Ns
BPZrgmAy7TvN2B/SjLped34jYJyeexn3T/AXAKbLHxOxvmGuuNpSdIfkuAAm2A6uoID6U+S+ksJe
4CwewTUYgUP9J4kdP8fNqtNj27ZdKDFumILnVxaNnceMQtv5CtBlP12jmqJVG9gBL5fI5NUcTH0m
+fqL6bTgx2tQJil44BCH/WGg60ty53xDh4/XVW1mWlo7KY+tJ1M+c3JUr0nxQHwUPFlEoqgA0Tx1
tHAuKUJiwgfDXe+Qe/Hs7xUys53S05czc4stHsoC9iyokbXyjfEfQRvdbfoRAVssNS0IqnOiJvM4
HpwAKf+teSFUXT6X/PAtIOoLnocNzXFllmzL93rJtwq9Jsjo6ixcxbHX/P6VtwKqDD+8sYQglTy6
1Aj2GBUCpaVQ0Wig63Jbm+eas7VOdPQvZYuZexhZxBUFlYYtPcpz+kCQKNSr8TNvRH5HBPCOLIbV
45hxrZ++MYyzVpIcSlGKRAFtOlN4mCXQ6VVyD4VWou9jrbyhnTuHbNICxAFBRg/8878WNYzSYkPg
7En/Y37v/JSVCvLB2VS06GPHvyt+qOZB9jXsmuRMz3XDp87st6alCRCgg85HtdJADyTxjGMCs/BY
z7LRbzowdsPmmY4Cwmoy4CkZtyiQU6nxOcsWLod9LoSAVKFM23zVZmSfp4+28WT8giEEZqehZmXs
mPLo9oYCBQHnPNgcs3lNRz5X9G+IXa6kWypHkRyzeweeSkPrbrHQiqxvTA/8XuMBZr7Vb+wkZoTp
TYd/Sz/iHi3gAyvAW4aNJ5PhtU1y5JTq644gPCC0qjLjlDC3xHfAYXeHIhyZB4klEsW79F+iyUWT
LDOu0aJk7OZfZihGP5p8FRdTdNiSBaqZ6p8x+KSv0bo7gPWV+Vfo3zJDYXXLk5lIjuxx4BjAAfn1
jTyh+wg81c5ombs2vjUfpRbfNKKfuBHR2LYVRV7cEKuLuTDFZCgvdrdYFk4g3Adk3F86XEnHrT0c
4AFsWzlrOcbZ+01akaawwBNJyXdj0zgS1UVWDSJz24UxgcpYF6D3u6BwkoJsjWHxmqoCi40ZiY66
1ptf8gZBL7iciJr6hJkJSVEPzufVM9wYsb/BYRHqy0vWk0RWaCPglOcPeLpTOLdRAhTK9FAU1ISB
J2qufSv1aKoyD4E0yfVkaa491ECkFO6zABGF+F/9c4t3gfOlj/wNU4B0/h5MkuXqI+GqB7vjkN6F
apBvNqnQO4Crs16skLYgHFp7Zzr2l0OwF2e0UzDz/JITZxzKg5oEZnAyEgIlEwb4eup5oIHSQPhm
UfdADgsW+iWAIhtwQbd2wTdbrp6mYYmIlopyKarlnA6oURGhLk8TgAbxH0hGdpt7kJtYRP7ioxQ5
rWt5kc9cc5I6yZcbRwn7G/kr2o3saQiqJiIffzAJx+fQXylVRZOadaF77/vmfqQdX6AcQGUdq8CY
ZqVy3vSSqyNJLkF/rkRZyulpnLsYix7/rX74fQemjmte0Tf/TZyAiV/A9WVH0kZAwAP2IWJapV0T
nbqzOTns48/fIZWopdtnEvhaX+5Q+UPL9JNlz3OGpE95uATEK/k9SH3HsjU+Dn4xHnLXoDH/O+9w
ZIEZzBlr5uDyBDfMhmTVj0VOgDWRxvIgtyE9fjsh8LQHqUhmn2EyXGsx64t30kyGtmZtcyz3Nk3P
43q9kFba3day2pOmIsP6OuwzpEPK6mSP6mQVW6o8YZzEb858cIg4baMaEwuu2sD8CgvVhziN1OPl
Cgb/vpJMaCK8VMCRcjNsviac2yTt7/cVzdTeQFPVqX1nvBaOfSPN1TYNanrFR98JD7h1R+GtT2wy
/mtlMv1UO2B/cpDGcsKMb/U/uD9ClUpLLRWAtykxsRqbstetoIBv6Vx/zFj9De7uXp9vWJsGRgz/
OxJdIndt+EarCiRi/X7Sy8t3SRnWLKoUYp3OKxqTf5dThXe64B+pc3ujtrWwhh3rd3SEmZxbWkqq
MHzPu3dNDIFu593PaKqNyWETwUU9yINkPMW9s7G2Gt90WUK0wla0oDnWZN10Fh5UNT/GvlLxpwg0
mVS8bpgY0nUdp49g81gdWJ3JkimtvnWg8UiHDA4XiEosbvlhKXW2BFdqKItK19joIB/3UwZDXz9d
Yo6oiP8bqsSnjlMJL+rFVI+v2FyJ8TguaWXJGnmtq9lmzUCYSmIwScK5s9SKGFBW4m/TDs+KYe7W
LyAvwZBXGScIK8sL/A0jPu5XPG8aS2uLPI/HzZ1bLvwU7fNm/L/wpm4LjIjJHu/oClYWZ/rJSXVk
nXFJhMWJLycNDv/ct/FnvVVbT8zOEKo4EhFYnmClyig8IlCu1Jy2nkULhC94UEoREVBqlNXaxZZK
DaGWLmV4ciuDIRrX7ZBDiDuYZjJkiGG44EiJOYX/XM8w7qKdwEUv377sSsl1RmCvg+QDeOmEViIi
kKtb3IWVSIb9Ge09YQgZ+ma48d4FireKtCOp/ylblxNmzu8wVE9jnpiF3xIBiKmf9jK3yv27PoQq
65kHxRUUBn5YM1510PYbAnA6PwoBIaoxuGRtqW9Ck9BX+YED2c16io8K9Gp9psWKHGBf9dceZipn
APYvkafVMrlJ5YLv+0l+fv/2GBILqs0nJ5OTxyqyzOkATUdovCGqZ6GZhvwuY7p/Acwg2O+t5gRG
N3xcG1PfNyfDeZzn0ok8vARnlqHyLZptFU65QVPbrtDjO72GqxJGy48ksKB3J7BbzMHIZeIS3rld
DmnaJNbPuzLid51URlyAtA43arbQP5QZ0ASyYDdwfYuq9lJBilQbzGEyGaX7z0hrQ74hYVS9Czk0
HRUssPUWC8nyId8Du9Fhg89NBw1yhP/JRyNdbL5giKhwNZp2IhAaUV9/tN10aTAk8lg3Ovp0XbIs
3MooEZ8u653AJvAAe4Hdl54oOs0mrOCU4Bk/QopyJIhbKKnA0pQud9ypHMkCYNMkUwX17X2POrZ4
ssT0IcmNYO43t/VtxKhZU77cZO8/FJtMkmTW6Jcc9TLDxXVVzdDHdJI3lyNnpE4eQeMRjansZblB
sD3lqpQK6zxGFJ5MAjRPu86IBiBtA6HyUeWU+TbCDSgsDbuOryC3iSROqdK7IvIGjuAYDiiiqTYN
RRFfwJ1yZgef79ggQCa93+X5k/Tv0pMcP6FLeUWtabBdsZToKxQ0IwqhJf/2bhU3SaSXLdtmm0bb
ABIuGS2qaAMOJPqsllAAdYxYusjUV48E4EhsAlrtW7ZMDd3kMPSdXVdLc1Zz5ZPJ2tuMmYHQaS4b
Y+nkOr5dVlWud0SojrJhzHwjPNftKOc/ijVm2ZT/wWjNdLvHhBGb7FchmglcOCrpSASF8isw3R9O
qdANWo1h5zbmGz8kwS3AOlZnTwonOYPZBw6uwrjNphiucfJ0/0ppEVvMsoHySTfd3dUyKUIUbCpT
SBLdxw1B7KlC6UKklqXpIMn05OYVjFuA8UJmXHLTqQjl6wTiib0HM5EEoxPYOZjIzPXuYw7L/BUM
iq3oStl61zL01wo8nkPCAW8FblAPOEB1ChwzYJ8Svu3yeDPg1UHUQN2BTe+8iEwdGWcXBwrkeO/L
mFxVGDv6JQaBQO+636gimSJZNbGxy10N10rRE+0Cw08005KInIsMPi4Vja2K5bBl1YRvpKFgzbQ7
tC++kveoc1Yb3AAQO0fCIxNZxuKVyMPVJ8BFfhAh4PO1HATMXFqSwA2lHpNLKSjhQDwwCgSf5//e
JFJQXH10lZ+MH/PK5JdgNh8DXeyf9KkFZxPaFKPgD916Bde5OzFBPGokbjZmqX3Qy9FSR0fpaRPD
BpfKF0suLTTAlr6FFe1fGnr1+2raBly8dubFMZoQ4ywf3pIjMRFCGZ/rPNHy8M7WylLzzIJUe011
KBDLpyjKPB1r3V/drQEjoJ99uBX7H3/5XgkOD6v1FymFcMpz/t8TAddxam2WBbHDXjkqbQ/3Lym7
zmP2A9YpHHLlgouECh7J/pcJKr3spNDw2ef4TK9XjdngJZLLK8wgjVN7fvTrtg4FaswoSokM0UdW
QXdQUnqpjWKXusEhrl0ve3luV/5/aCDvzFTTKzkHBODvr9YQiY7CY4GXUyCqz/eNT8bKFgjB+mTm
VtAv4B1YpVY1TyKwUJKp27zJhHLBB/yXWk3JSpgUHPvsMEZq/3cEyWNdaCnRdtfIWeS/FrNqPerb
dzS0ntsQuAAQ2XNcXuucoDUOFeXpLwkEgkwSL+0kQ02F88hEh+g+KzOXUU8LLWPxpDSp/Bu/7GKs
czrxQOKh7blrBQy7nlty27Ts2VuGXsDnXsy+0ckwymgZ0kxBcqmeqelpSrxQin59V9kINJIa5a7S
D7XMNNzVDlyVfI6TvXICKxXz2Nqrgm1LltAaO27h9c7k+pjJKUkl9HFjkWTv7L1tM4XbEIYtvrf/
VZFuAJdqudKyR2dFVWrbWyxqPkYi0ivrae9EgwS/5Yyj32nCpMfgcL6a3F8D/oJZd7bJI+8H/OeE
QdWF3lufu0EKs7bvPQDxsWypw50SSZlsFspGfQBv2AZiy0r5PE8nc54yw3gDFYdKDzLAi4LX8FYy
VsP1vP7ZoWwSIU7E8riJ5wIJrfgvYA+sssnH624Qg1eki9saj5ru3kPJp3CXnthJfg8QRO/26F0I
OKfg2x4a2a8lWVLUseobUewxvsPf5Kdg9LYrtRbmCNA9Oku3EFC2avJpj3cNzSuqX1E+dh+CZAKE
V5VZ8JCXZIqtPsRaBPymyOt+ogA2fGAKe1Bn3mDmr5FAbuPOs9sylkpc7xdG9Tr18aSMsPGUOkkZ
huk0s3IgyDTygK0Gx+kVpFWyiQNp7ygzIA9X2QCrGYgeKZbaLwcqSBBvyj0nFhyaqE3uMUO6Vpmb
xa4/WdjQJtQ1XHkyHDLqoKTlbkVA1ynocAre50XHkfRPsElIGPp77WstNNbsIGQd5aQBzJMkrlRG
t/PdYathGEbxkhJIplGHLwllzzSxtY6DVnJzkOA4ZFWbmcGpOsTTZBZyyNLR3hK6QuI4nVMwHys0
ix1uYH7KcZGK3uXMvYDiWYkCm+2zuJT2qrmRT7R7tSfqTeWB57Kn+0aJM6gob52X5iot36UAkHTE
m8pMmF/RgGIOdN2qEqFMHsjgr2dSq0J1QKMTOKpnx3YALmFtyuL8yUPfWXYHEOCd/VWiE/EbAf6x
U91CwxnckWJnmrBjACKXE6uQdTMPgavFJCe8RGmOWmGe6gIJf2xv6asa24YXYSXSRwx1uctW6ish
UOSQfz/4ctfTHBoeA3WMIjiEK/4Th+ExoKwvoeohdfTZf27gSFAYobTe0ga6antw9QhyUD0gqSm/
aYfsfXEDmQxIVzjRS3l6wZiJhqannaY5yuzCq9xr8CRnF/VTOtTx4DLzWR/d57EczQDw38jAjSTF
rZxcAPRSnKbSXF/iRX/O5XQvbEm6GJRSF6850vkLAXvfQhWsi1UIWIJvN7h9TpZhmb+5wL17Kq4P
zEiramosxhj/vR4q/r4ZcOuBfjB1WzYVO1V4XnELCK9/Z5mopsTJZH7i+MmuO5A4GpCS/m4IpIGb
J6uofMT7Nnwm759evBmkEobMYPref8SOo0YpfhVWSI4vrl8ZUsG0WanHia5BH2h/VpesGy5XKaKV
L7duthxoOibw1D6z7PEf1zT1mjDtgKYulwIsYn2NafUJYbOcWJdo/jTPVgFvGUVGY53dKDOD1wGZ
3Uj9uDazyNisFQAIqxvqk70jeQLguzpdGfBmf5h74QfF3WEHatQo4mceqV9+k9h1v6FBuuw7hWpx
SgOBqVmt6es51yqSgqovXP7oNKy4BWyq8pmxuLID+6L/eMC4/nmEltDP2vaq3szxOoyb2X7YGSRA
c43LD7BoG5izRujNwCLEd0kfSLdlt2yPifYZxeSzEuFZNrA4P5dQCfpygPfZWVhE37JtbJjCOmek
zsfHZZ2qUIu1WY7tAKsME/j2eW0kmjbvdBZ2bQhboQzTQp2baL7RftWCTD0pfA3DFsaqtyg4h6Ir
xVnH5FxGmWgNObvKUHdtjk66cMowophbAy1Q0kJHxAzFFePh/isLKn2F6xXaHz8IUrwyhwpVVWZQ
LhsP3OOCQzCwME9jmlPT4g0XDtRdyX+hZ4H1zT0oATM/2saTjBsNT9NitU85TYoTBCU6DqOaCZEF
9f3smVwYFfMUbvwjTi+i0u4rmSZo1OkOUrO08kcQo1JsOzYGhDL8CDyNrwa/nUVmr5JUuYGdMh2A
hWbwJd9LM60nQkT1oLO8Ecr9MHYox7sV5OenHfvblqOIrDdduECnvnIRXIEw6GVU7SM4uoWlgekj
oZqmeZfGuFHjI/Eu9diXiTdUJXDxggTFvrDNgnhvD1Ybq666g6uAE4t2WxT4wUiK9JXBCwtKvrqK
7q59R99tAYO3L/ks0wDIFpPSNerEbQl1WLf0CEcrWKDuNMbPd7UegX2BrxHAExghZKLfuWFro/Ql
m9i/CD9o8VG9UM48lucVaKN2kJBT4iF0EojjYUX10DxKkBtv0qytVwUFrDjx0eQcvpMl3UI7AmuF
jKwnJJ5bE6tPUFob8HxbttBYV5wsx4ZYQB/J4X9zf48XUKpsuvZFdkzZR/ItGIUuMxurXDbK+4RR
cBYnuLdIUuUAoif0MwhC3fWv1mmL7NKrQVMALDAF/ZfctDhAinW64K+AQ+sQf1qGhsTTZUWn7PuQ
5l40o5dBrnsW4UC7yxFAI4yMMR6jbw+/3O6Z3OtlOci5U8hTv7DaDPiQhYskPb0R0120AA3gzWSm
ZJbocK0QAjgxONbxZ4Emq7Od2PICoFZlyuBy2H2py017bJXeKPeLnYeScq+aacGrn/2LB2YYYl3s
7lXvXbd5eyQINjWANY4+B10n6XIZs2CzOjLkfIRd2snHtknftpYPB33NrPPOMJnq+uBn2TXAFy6s
b4dq/PwNgDpxvCw9JhUvKYNhTVnDS33YR5/k/377gMhioFQhYfH48Xh4YtWQvnO6Zy2Cd/FWvaoF
5TS7jM2Sr7qhmsmKVSwdJ+/dLMiolSdtHK0WqLohiflEMXYAM+EtwaYgO8FfJpkDxvpmTHczr5ct
J+lqdtJ/GaE/CNjM0eXd4mOe3mWxa9oEZ4QFSrRfqb2I2hji6SP91jjFJlLNmyUhh4zDIWhEYTI3
jUdpXBlBr97EnTef/op7E1BZUjYvQXU00aE6hnoEC4SDD0Ur98kjalMC/TV0TKuprrchR6deXohT
nn0vaeEBsac+cDJLcDuWQOmyfyaj/v9TD8yXwNBeJ0oOI8efFq766qufRVJ8JcYc7KSIFS9y5y05
Fo9ULcZfWGl1p0uL2z9M1wWpPKajUrlCZJkYyzN83DqakE2nrn2/5Xy0HWBCCtGS7w/eexfoEB9v
0AGDihWCugaNE7MgzMZwXGqFXsAD3gwENgVbvUlwh9ZDDZfYZh/5g1+vl3HzYjd1q6tHJFm/flyd
Cd+PORVPRC+ekuD9gP6B/OdE5dDErBkZZzejGPNkcjf59k86FjkTlY00o0cBEkS8JJptoMpbhG2O
a5I87j8MBCZ2GbZoy+u9+0yyNadpL/UsbSnxaa7F4Y8f4JBpSGzkmtTbQjhVtjHIDVkv6/d2jM66
zLf+iZ/2UZebkr6OAwRQFPPGcfm/sVlCHSVcjhgrnkQMYr4tY/h5CkpYcJF6XAuOQ+kP5UnLap88
6uRDP3m/rgQ78Ptb2QHJTXlOArB7dm1Z9PJUDgfqFL0VpgsaGKeb9KFg0/5PU7/YOInQ9xJS2Zh3
iNDkO3UkKjTqrgDCzbCckLyx6/Czgc5LRpQ6TeTOgZ74NDmuIt4uYg/X8dnTo2ZhwR8oCykY14ZI
Ubtp8mBfpJPnLjbTCWs1ut0FmXtBv4plAwJD1SocxQreoDEFMN3TqhC8t0GfiBgPKvcuzSncuHgY
OFgHmPeq0IjuzJoSonIDHX/4FiiuKB60Ta6g7zqbAUxghdIXrXNTl5GtKPHG8G/rIVCbwmGtbzNU
4KKLx2/8KqlB67ThmL7idjBSvHM7u/zXyD11pOql+WUieURMV5Tpl9+VpOIwjy+T2K0cvioQHOqa
tlbWzqgmEED1SdOyLsRjYXn6OsVe0bNY1Wu7Y86JupU3wIPZL6O800teAZ5rB6JjNn/Cvt7wm+lJ
0oC1nYpQBnDswwmLroP1F4NNey9WGHTpJkRzZnHPnuacNume3bYud+OLO8g+vRvXGvPl/R9tjYLP
9tOP7BQGU04/za+LxYVASlmuZXolcRJdW8hDWAnfYOjpP1hi791sUjON05eFUqXUDz0IakbpKsM5
6WnDC6vfnhIwUmX2OjMbKcSR3Mewxpc7lNpaEDxkgyzGezpyI6E+YH38OC0miTaQhS2XWjeKtk48
NgyW0QIC1OzLyJPkhLBOl3PlzNzhkttYSIm5sFeMuwixvhQPI+0XnVgOMKk8dVg+3ZECTJJxhq/O
7SBRTdbjPOwTL2DYx5pPAW/GtzTOiLEmJ8WtpFQpgLYLKBQ3KEDdPDgL6oyJ5KcNsu/yy4crvRPQ
XlQxkJTXvTrn06O2OCcABkJbJvXTPVhcJ2K/pAhqdILLCW6FMxR3FpDd/U6xhDV71m2haEASY6tR
IRrcRh+UV8GEbSZqJT3ZVow3Z00rwmAgpXxmXOzvloH/Y3kaxojpLpbrM6q+rMCk5Wn0VElXXPrj
c3PAeTXHe4X9HHtj1LPgInvu+AFSt60mlSwdZEx1ANvjKx89FdkTfauEGw2AqUazBx0kzo2XOLe2
PrS7+cIlBcjEFW30WzwlErPLiDVKLFen5jNMq4jumcp5s8XlLYe1WcMo0rSWbJhD7cfl0U/EjTx7
WWTnqdzeKSteIfKOyHNzXOvRcMS/gevpSqN0pmRQLPJGRFuWg9T6I67luZRRPxMHe3E7x9aWvpxH
3bgTyJ6EqOkX5RfXZqFkNZMOUhNdtfoKfgDMPVbzodb1BqntCyEeiKXyoTkK+rkpypn18c3XJPs1
GCp6bhjA4DD98ApevLYXOiS6HamPZpU16crJDnFoJJhhwv7Thu1a8qaHPUsYcyiVBkMR+zDngxtT
JMsdXao/8SGSp3fCJob2s/7adf2P49RlM0UUCb8LCQOwWf2PJhMecQhBjAGi6n/IEdfGkVQEXAd8
M+CeOcJ2+pzZ8JklTAV6yEwL8rXkuz4/dJuQQOoUerzOCVNC4yz04/AgzulRVEwPO5hJw+SFE4ee
qpdUAq/cwDhgQnEQPcWILH40MfxUW48muqSitrqtmBzyBZ5eoO8wxLkwrVAGJ9JAsP2odb/xOmPi
gp/sPiJZYAzS9hvft/Uce1gvVmeM+LxYFDgXZ3F7URfdZj9Iut+h063XR9//nE+moHkq8ovXvqu8
AWifcqG44NKl213e+ev1T1pkyav07135QAs7y4bcSqFEPNiHcYEyTxP8W0PDaucCLPGZNuc5E4z4
NS8X/zweobKV0gNRe6rW/4G4wRn33rQjiqiJQVR/3yaAAUgESsmGuYgRmjBd31YfC9iob4bYOk6J
w2dPETxp4FQsYhEfjhi24ddsNtmVBpdgC3rM8SqlezZUZxyGmVigx5lAyqk57iNbtbED/2C2bjbo
Li15Jsyoo4WduDhI0Qwql75sRiege+kK7ecSJjEXuHEB9nnlixf93iW8fC/B3c7tjoIJr9UL+OvC
5Lm6rp3n+Dh0NLJzKZugmCoiNDSw5nxTKgdgRM9UJCs3Rd5C5BXoIjTQjnFEe8/dz8cZUBDSE3O0
TahFAd7WHLCm97PWb9GmyZ7CoqQicX96gcSyd44Wtq6RmNQUSCcIdkCH6wgf5rjV2vgfPab4gzHX
Aq6+wZdjtgA0ynxls7POYKBS2HeBxxFOcyInsNcV9leJsMj7Yt4XU8zvDjNS5zrBs/zudryMvI1g
uNrcDL2pRP1UBuhthNJOFfAaMRzRwaAJRqpOnSiIxNevvCieev16f6iCLGv3HkWqFUqJeZ5s9FtR
m8d0KWfTxyHfWGi4pgWJY4T/kgeRonYh3leBctz/e1gJCJ2nHfG7hVcPSyRYubajgrUszCJy8iRZ
38huEA6Ge0weMAxrxzTUp0YLHeaBJu8Ia0nQhGti0VtQ1NKEG+TWkXLZjbxRbUVlwKIQALJAfiWv
JelbixdsYf6Ea1s7fz7uNVJpfaqI5vCKSPNOi+/mdL9bpc79XoZoQEPrz8cVDQnF/FVycEncGlyZ
s3diZiJVc7U0JtHY+5D3R7YVSLEx2RPFazQxUEda9UsQVLK6Cq9jS41tmsh5YEjaAVW4gT749Fpf
DWNukRxA/hYgz58JrUxLzu0MfRJ4TL28SCyog83naZbxRLScboGf0UXcx3AR96yGtuqX97W5AusQ
2Su8PTbw/qrPjHnC2DSEihYIQDld2O4+2mcCdAQvcRGRyeEEghnzcZ9dqgN8Hb6BTOWiyoQhN5fw
r7w1212VFkONpUMUBeD5wTRvWFlFieXNtKu6ydw4ZtjuPivQ2xe4D6mRa9gmZ7kElASuXKq0bFDV
Du8PQfjS7Ossqqmm3HdiZzJn+GrKypupYc2AUf1KsV+Ht9f9F7XzRs5pvDlbXt+xCbgN9sCI1c0k
IdBejCHgHIuW2MwsYDGeqDvd0kK42dnG5I9Zqgjry8jOfhz+JOjZLuThM8hmgCJ2TQahttIToUkX
gGU5mesvNzCKTkXWeJKF/5Dm6j+b7LMNX7FcKspGUUGBwDrtMZL9NBrA+BRxCA47IKdAWThCEBpF
7MEIWe4tkljbBdPkm0IKBAMTaKSySA4QIl74XvPCAVf+sqr6fVkMzxbULt28t8xP0IH5QvTDhrp6
UG2fO4mtJnc8DbCpNBA4GOJMzw1cI31RgB3rK/sVehYkmY9FthCnfLajM6ZsmW2F211lrYS5OveK
3DTLqraWl0V49v1AC2R+80IVMXy9FfL+pT6E6jQV65ySSbNtX+iEp0xEftT4Be5NsqTrRGO9KQ0u
26taPKyDUJVhXtdCBxW7gnAmPO75q/RCDInYTAEy47/GgtnfEx/twfcy9JJqWpXHyiWgKdvrNHKC
un4SIP/L5ONOeCHS+4ZVUAxdBb5ZqDIz0sUWVcMb4XewpQN5EG7sL/b3IgsoNvqaCl/UNSDWmDdS
0lULsL9P353WXTpzSeY7vR0BEhnL3hL3hboiPPj7PF/d03msCurgxb5M9lU/POdEMvbpCEsZcY8e
mYGmWcLlRLXLjoUp4ou6Zt93wvXJ26YBjswnA6ly5HVrx4jlwxS96Y9+e8HwjTccj0xmAJBaDxYz
6g9vpWDrYKJhiuEL4k8C1djULoi5phE1zOl+fi3mLWFxNkjWuYpcS0xeeKrFQ1zC6bTH7LIYYqDC
aViItTFbMjU5KvippRypy0+1KP7q1OaP3BhVZgCJ7gqCVM61k5DNe2o8pLKYoZygWpsEHsAzCfFn
owG8FOCCRrUZHNtOwC0hdbhj2Fq90OdvyW8hmKPk/asDl0T+84MkerJ7p/a4zqUL3U7HoR7WO1Sg
zaVAd58WzKt9GD7KvrytUj3T9xqLTLI1KJcjgptm8MEe4IEwYgSV+BQsfk+A6oPKkB8sBRm/ZH2V
kaVJIHf1tYXcULB7ZuVNQUdhxOS5UcaH0kcYXdByprtFZd4D5bDKgLBkMLk7bp5WxN3ZfpfeYU9f
Z7gvAWSeeidIfpIe5A2xnCMEW+SAjUD3mxm9zM8i8AdpjE6rtSYwHv40iuUtjjP4njSqKSBHmvZS
bt6wB177T+zC6EYt2635+N+9y3QuFJu1kXkl8ZR4TkIbRJGgFfCosmXhixbfceWWpqi8Tk766fsU
40JcwitTgX5JOhG4H7XZcx3Zl4YCsm/FXXVXkLn3/zGi/KRHNn91y5Gfvx6agt3ECAivmX0XtWQF
MOkyT1yJhndqGP54ijwEMtHk6WYVxh50f1kaghS8pDrYmlY9sM4KUxAvNr44lWYO6X+YU2f1zNGe
kf0J4brrdVMYayjxNpcRh+2LSTGJ0aBemJ1JrmjgKGNQOI7oACTscfU3sm74Ga7KwHxYIJtPTfKY
4tfr/YHwRIIx0LvlkbWUISAjiMR+4SsmYQEeTLLaUWTyJXuMeRpHxT73McLu05+K0QbNW17KG15l
1z29zCW+DvuOpBHQTnONFujbMu4keRu3VGbiOlU2PpnUtBS8w6T0qGmCNDcQrpxQFLF7/uWDrp3r
RwHaq2UnKigVJFBZ+AdSm7xKpMDjXeRsaYw6w9jYbdXAkNNebOnPwbaf02a894gcuHs+V3rKr0/4
KDHNogWC6S1sguJnV+Ox4hzb8VnGyt6OC7z5pwwi6hyQSYuA4Xh4ZKouV1m9IWnovskI715036+O
Lw73wHiiakp6dqUxjZvDg6J5c0QYiCcBud/7lF22hORe3PvFqF1nixY8pwfMeaacOsuebwra+Hsk
QqHwUPWjD4g7c4HHOXTYDU1o5PIzvA9ShL/V8FY4TIW+Ny5O99Q4ZymfGHOeT3jJ4OeD4m9PH7yp
Vle7ZNn6UbZp8TwzG65FwinXEhirldUL/9HW/BXeJf6Z6rkimx/RHCPcES4d2DewGXl2tm5MPFXh
S1k9OmO+UbM9+sBRLJsyA41xQ6nalmxTI+x3RfZFfCkr797vc5g7z5t0+0Mzr6oml2jrI7wW4uZx
nhzQm1Tyn9ld/OypVmZBs3ky02rf9j6UTxBm1Z+9UEMsi93j+iiMJ6vAi2xivgQagNgUogj15qyU
P7dycblo4ScD1/VmD/9SWW94FepSGSh5e8dd/8QlQgYu6A+jd1wChWGz31r16BhwevAbKho66DyB
0Hw69xfrSTu8AkCeVCQJJVwO/QpdtdwTDdBwLYqXU4ar0Rrm3R/TU0Udf+0qWlPNV5npD0dPQV5A
TGVSDews79sKewpLvnQi27BsGk+2DVI76Gq3UzSJ9wOjrv9+Qv2exGv+jxxv51B+Q+E6RtRdvxqJ
cLT9xNCf37xOKjkCE7QBnPfkrwY2Yq8+TIpSAiC3G4TYf21C1OTJdlp4J+KWPnCFuXYCXsY1rWFL
FWrauccGL1YMkLdj2BBmsuuMLv1e9qYUlvXABuSrGvl2nWYNZkHdNF6MQ2Yn4vjVx3jXl0wQYDDo
ccej9ctYaFVvo7Oux8S7xPiE1nSHzkqTyxZI2hnDQ5Ystk+bWpLAcBZH/cKCLIYnKACGaBc7A1HT
Dj1FAcHhCmW50arZIRmsjTClP42bAY9O/F0cQd3yhBMkY7ZhoQCPIvAa9c8pwJEIM/X+lAbG7bkC
v2MvM/NtLfDHHzJYD7PAn+KH1EMvKcMpTNjJieqO+gbZIw0v1JxoITBVK23OtN922wwGZjRcUbQ9
cvNZytpJ3UyG7GSg1+/e1vvMt9PfPJGszopqJozR6DueIfaJKZRvxm3nDLIy9AZDSJldM1WT5+dr
wWzIbSetgyVtH3uM9UF192z37oasBblM3dt+QHemc+ftcLeCFhra1Kp7YgQhbrGQKJqAezrgyuya
RxUoq2N78T8HsYdaR8EBDv3P5EgMG7To3cAqW9HU3C51t88uBAgksuS4XIgmkH+p46Mkg3pHiR8I
g4kFaNzCpU1EFDF6LKlNUDUa+MMKsbeMYHugAYyVwjU3HWJrxkeCU8q25V00RoCPiHYsrEyORTAy
P9IAuYCSTBJlIA/yyiWfJWv7U89OkaI/5RClgkp5/z8JCtuEdf/oHOkvszm0rj9XNaQ0FHVxMrCd
rSqjDr6UgWnyO644ML6CcsFKy0xDV65IL8iHX7e9/mzlwK2RFshIv79pchs5H0pb2ZI8FYoto0RA
FijC4lZrVJG1wQnR0Kik3+s9PBUijmEHkzaAuVFegBLknGTCjzjr90TP7kPDCduPw2U2Qr+xMUb7
JwlSwDWqna/eYfl+i2OXiQZXdzZVd5norLUx4rp0HyeW4Ld3EPujEWnhKYQkRFEYJsYNlYVyWI7O
L+Bng/ep+RhGfpEa1VZv7uxiuhNkzWFRp4uw+3pWxI2aK8j/l86AgLyckG/XcjUrWu5ufcc8fxus
dec98UwsHgPp03R1Hk3wXnsh4/JFjnn3UWDeFzCRM0M97qBghEpRX6F04+X7ZYDoQztRo70Y3DZq
JWPWGTLdE0fqnEqZgwrULDHUdlvxH+PFA3Y0Pf9V6oapaMn7PzVthXzH+tff8ZwjEl/rIREnZ8mt
WmvoQLQ48qBQQflwOG7ZhnNWxsFxoJKqguqPiwVmVC2aWAlhPHoS0r5dnrOXc551HqIWPJu+QGog
MAoEm9YHmA1JXg/bUC73ETyqoHDNMAE/UO/JvLGBzB49rmJm91OXnpEpTPNW35ZQ3uEOTP4p+vOY
/Hzv5QGINDbfHQ4Zqwce1XUPeK94GYCDaEQ8iDvug0+uqNroix6JNje0BVxGnZLN4YDtlPF8/l21
OtQ6vcDH5CVYidEc09eSdkQEekdfcrF6CS4CWYj/c84MkCIp0T4BtODgUwGyRpstlqqw0LQ4KtTW
MU6OKI2EMOaLKkOP/YamRZzNz1pzHtfqs+ooahOSmNj/0ZuyAYChuNdjlSCVfhe/5oBkm1sUmbO/
Xhb92i/gDHPA8pfbBpfvkQoigpV53UcpzMSsrtOWCCsVtWVGdYYZPuu95bpeYUwIqoMKj/kp9x3g
6SrD1Q1k1xHo+4ffCHLEkTFaoW0rzEVlrMySAgqz9UuyAHn5V+RyXCJEbNkH3yIvnOtIAVG/WpSl
6zQelVPeGv0ISdRf8uszH0HFynDGVBUmEijIjcYcq86R9POPyf2foOH690YWYvhW0mYO59qz4Ry2
RxnnEn5zgrZHqOHXzhBMJWZVI0HEKHHR2wxruwj/KkwD2ug4dW3dae0OI7jqzNSx6XSNgAApdea1
TjucbwLSnpMfDm9wvX1KPGsWkTOZ55izF38BhF7xN8v9beGZAQaSiq76eSWnrfMoZGYcnNv2UXyf
RoRKxQlxumWA4HKT1G/8JZptvXlqzmAQKzziFJ9+xPq/NRjskFy1aqIZwxBCOCbFEeZPBK8bvEfe
F9jt5A+oHESZmzZ5HvId1vB6CdsOamstpJgX7DzcFaQNA9tUkW0sJflSdNK60p06kxKmnGafWSpl
l5P9uxgLAM7CKQIk9o6WfLh7hmi6SIG/o7n1A+PmwSopxUy8s7wH1CB82or+/+E+eaMHoP+GHlzw
USpkNVFezSP5KKYHoZUeZA1FH7es9g9LOL6+RLWjB4A5ufD4ftw9Gy6sxD01pab3eMZ4Fpaprorz
oI+58FVZSv/vjPirfgI3do2MPRYLqzc0z4uxeaYtvTyJDCj6vAlktlV8C1UfxUbn8RoHLIxQWpMn
eHFQwM/O4fgLcahtgVUOQk5XCF/psLTTPFJ/aoe84TE+rsGhO/mXtd7vryANJxJ49QSz3vuwL2JB
zMMdtLn0xvvV9n2UkJZsP9eXeUHEaBop0ytzXBll04S7p0pseqgztzjE2ElnwQxVXWVcijhO22al
jbIP6zDjMj+wuuWj0h8/RbaHcU+szrVu+Po0ZCMo01vAq8cNOz0kDmo66xhvONGXTt59+has1hq6
FFqyOhYLtvVs+erTNkLBAcufBHu4q0eBaQ4svK+qFkUSJtv8fGlETU2twhOgwgo4T4E2C9Ngoozy
dstyfLoOzIkxAnWYfdptG/oz/FpHb0zRPDUUtb07UxVyvCs9VNH6IRigk5lMX1y2LVilzM7scIbR
ilYRQy2YT2muFb4F1HbLHZoDQ0VXM0ZkDPGwrLwuVuDKEy94xIsdG5DmbBrNwupte8t4TstHWJvE
x5ZHtn+0PVROTU3z+4cVsUQYZE0i9rsLYE0COuQzTvnoPxKCtdFm2b3iGgsYEs7hC7ah9HNPL8jD
6WmZdM3pzLS0LyAlbuzaiUaQvcfjtkvhKxm6Xx1CvKYrZQxKJh8xAC57rLJN4S2B1PNxxZNhFrm5
JUGV0HkC/4PJNl/JObUi/IDCkrFq3Eknu1RSz+m+T/ddsRx1UmdSBbPgpEL1E7CcRSkpobA7yn42
rvXkeYcjhDmTlGlrETXmW2FbdrtNpg7Ep7r7+UsZworQDB1AMUs/COnJrwjy5jbGTJWVq3iUXHR2
2pgd9kSugrpne3PgdkZbe8aYMb4QsynN1UUeIZLspyK3kARmo4Hympfw/ILEejhgZxp0psBMl5Ry
hsGEzR79ujQSR2Zh2NP3T1MFkVP4Xj7sgLA+GaomPDQOowfs1PGeuw0rZmyuY0d0GKnS7x3kPWjs
vR32mhWGQfetdt+WlmWz51ZCIx7MWmB6cUHrM7QQJGkzWAPmRGVHrx0iTyHYtHEcHQpbbn6ZNPni
FQY+Vb2Lns1EVtPRz2SHpWDO9Pn815tk5PnXKKgA7or3rJ8Hs2pxDulH/9v1F9c1f9imvHeGqB0V
7G7M2DstZrbR8o6iTDCb7sQG867pQGkxQzuDtd40JJSID3Kq7H/AY7tLuDJibGOnk4SLvuVI97wp
83PkkR8xPSSIKKlAs/RUxqYTPQbbalEMZ+g2ApnebxVODlUxuUm2nrXV7amzHtHOp6TZF6Tci/jo
sOaPQJn1l4exzMS9SMVFocTgR0X6DedhChBhddytEaoobLPkp2HDAbjJSBnZLjSVSzzpDZN+QEqq
DqP0yA4WECWAOLo79U4dk0KOriYvPcoCDogAvoDv/SNxQyCTd0D9ynh3MSdxkulAvz0aslWEWgUI
KzzYOLVe0g1I/1HLObW0tZTWg+dyK+J8HVD7cOMjP2AuJDCiIXGn/6V5VaGoATUtkY0SpDMArVEL
f5+zCWK4I/7zvbPwN7YmjHqIf0A+A9PsE4TUQ1LhX5yLo3emMVC9iJ424HQ6iDWKBUqjmY/ejBGW
eKN7kLQtJ3P7KiB0Y/xdluVvELZi6eYlBVIM6v/T4AYrRjCaVAmrs4zIl2xsLu+1i/YN5ppd5SzI
74Y+VgmMITIMW+sgb79kz8mrSnd9oWieIbba/82jIP3PQO78ZaSc5NIKjj5z0knH9cUKhVJ4UNJx
5SED6kqeu1DodBXH9tm/3W+HKJEFLe8AzboTSmcARkN+TyoGJnZYkfn3bJasnMX7PQonky63WfiY
LEeRNXq32N4//H3aC6OUMwJBJ22Fe7c4b91M7fPMQp2CU0zo5tyWZb0SSrNPEcg3vayDhoGFt2TA
Fj1j2giw+V/A9XNFBfsXmIgGIkthdRQhojAZnkUwvoXUodCmPpjoAN4Wve3VRpaA4kGvY6qmvd5s
XtGdBeXLVRXXbiwv8phMdkMWAVy4OHj/0sM8Ay49k0TZ2Jjavd+K8SaBFMbGqXybDTGq9yWAZmPz
NyMjBfOFGJ6+dprSLalOOIReDNzuKT8xTO3yEnCa2xplYUMahk1J1uDRD8VWWGnagOnM8Ev6VBSb
uHifJhOdGK7bPV+lLc2pwG0cxUOnP388TneIgGuFAUirZt8v4z3iKQWYNKX/sBwrQap5Vm7dCgmI
kD7x4iR6qhUEWtyL5gxKR+kMUMIGRfNazvpevJkhzNaGwfTKm/rx9BAJ+qVmetGcyaIuzOj2MbBm
nlmzfKPZ1x/wf8sK/h7/3feNpwf6g9xLaq5749wEg20V2QK4o63r/RENTZl1DBwC8TDqS5iPeDYG
mwSrwl7Z8+lOuI2VP3LfAiJ4LU7EfshrU801j20HVAAWE2KET4zW3+Q36ZgtzD+LSWRWSDUGSfkw
8svgcMphf2ECckq369o4ub4wuHf++++u3DE5ZjkOTjO5VrhEtoOmYvMTeM8uzJ9RW6TlkbsZYnWE
L6thTmXCZSKIHktuRyeLMTvpKrOm84IEsNg4UveFm6DQHr6Rvz1UVXWdjLfWTGFHKdkokk6XkZ1X
lBQ3uWlTSt0k5g4EgSrZBBJIJvtkymwa5OzeGffs4PKy+2vPTcMHYHz1u3F+DXaEwvoJ03eY/imA
TxpC/TleEpA7zBup8EMNkpo/V4aogYrEbmf7R77A4cYZqQJmlQJdUhT6pl5SZTCg1BW0WLTF1DQO
cdtglO7kyPL0xSVsRF8dmLZBV8tpbOuS7grGEjHoOtB0yKKa5ovm8hRhFLNZJD6/r39WIFFXb0Gy
3EmgdX+SOyBgs6BOMbGdrNroVf2Iqm9cWGgVk7E9M5S7FLmOwH8JDw5JJ7akoVv3tJlZPgv7dKtN
aSf2M6Xnx6gtlpXe3vV4ZWDBD6qmdchgx5DKcf1ZbHp71EYx0/U1mhTlZTBDiQY2UDANYqvl87qj
YJacD+SCIIGE1vHStgFfb5OZYe3ZUHq+u8C18lKvGxL+h45njMyiRAODPwHOA8V7OR+iR2mBL0uo
09/jmFtDQuyZlUbqVVZrSeaJqIXzcZpb1Ren8qZY2m1spZZANgeebqlIwRl0N0cHKfKAIZKXY9zN
9n0RLmipkKiv3pAcc7CUnx+/SLkyZkTjJ8B0ocy5TDXJzS7rWDk8grWbBlg9r7B+bRvS6BgJlomI
j+KxcRuOqONFMUYBZun/+kn2v8Qb5JzC6LQWci+geA8l+6X1pbm1aFl04H47j90rgRzGYiRCQUmK
J5QZgiXFZ4aRHHcxmWHpw/gDD48Xhe14p2HSgSvr4j4WILQs/J7dTQwWeyTxvungjjC8W4PLKpB7
fj/Cku9BfcXR9tGFQYjXOtKhnHsodLDh/Q0MlnRLTj97PNAVdsNPqov0755lmv4GdGtPcbIBYSgR
CjSnYZhGp0nV3gFgSQEWIm3E3AD2Ks0Z9p3ZUR07W2kcH67YGLD1qOV5L22nTsFLyDyFTADLmhWa
Lke9EnCX1FtogdkjHOyEqvhRvf12Z3jjxqNUvn6sltORXfXiUfsWg6bKx/l5DfJdwoAoCc16Djlp
yVXHz+vFz/P8YcjuTb7NgRRqvvdRJu56vEc2v+UMI/Z4TeuhadS08nwf+/a3xoJlcSu5+xy9iiXD
V68GMe1m7MxvjRLImqU7/RPbijcN5BaJWCY8lomnep32bQ2/RQ+50tWRgXjNW5g69ig+uFQwMZQg
eTgSY8gp18caJrfSJuCIpV6dtPaxjDWrv6qzuyNO70eUoCycChDGdwd5stmJZqMTyCWWwXDPWqrY
XXPacToGAMbyKHX2X6R8CycdT80otulV09PN3F+bTaDlcIEON8sRLbZk2fowIkNQsFbo+BaiQZaa
Khj2mM7NQRQ5Esab0+AuaOsOij+xaxP/F2eHgyi2rNe0TpMOovGnIaWW5Q1/soSNlskmrO+YvNTi
V7Kgs48zPgWrltQ/SOk/cZNt2d56ER3y4NyZI0udgzaTi8CotlTbcD4kDPAlKriQUqqmVDvgHLsF
riF+s3ZU2J6VRgzacv99v7K+MxdWMesO1YCeN9ICB5aNhGUdj7o0HRosEB4o12ILOuK5BL+eqe8z
WGYk5MxzyXypKSEdKzd2t5hc5aFXlqFZYoV7KZTid+VNtPnfRBBR2yPFJl3YT0vrGAdPyRuEEqIf
7IXMcjtilceeGl0JVxTT0mDknr2IhHQgMr7Ew2/tw1QTfKtkEWP3h58EXu5YpoaYPg21eDv8dXto
yEkiD7oavll4q7lkiCYO7eWE2u1lMFSf1SMemuBkrle+Pp4Su7BBj7iWR9WSWuczoZzwHCKUfalL
qeoAGT9u/ZnCSD/IezLUIY9AAtgBAxEWmFtYPRCvIHQSg0IYkI6922XfMtkAQbgCMk5b30BsD7Jf
Xcg0F/p5zduBmi7kkgbMFl9w3LO0k1imhrjm+SV+T09nJOu+NRewemID4q6TXnuzDRDwzEZIanh9
R3Ho9SV7yV4B8L0m3Eh226oFMsogHhGoEMVCC5llzWaQ+X3cgzm3KVTf7HPUoW0h5PnBR7nras9H
2qtMsW8vwdHE/WY7ZEatu+uYUs4IwPPaQpKfSotjWAsBn3qc27RQNUZu6Itauc5aibzy8QTdcfin
KJwTdHe9zSEVSHzjog5G62/QzKzO45h/iS/RQvmRcLwWLdmT8bVAi71/+Eq1gpIDvq+LUvtlGZJG
fptfNaLDMSYKJkJ2Vk+Mc4CN3W3hkWMWmeg1Z0ocbcuCqLnUgvHN0ODSRonDLjyqSkI4iXf0aUDq
n1LcmNUAn7FSxhq585teWB7vWlHlzflM4lPLyyJscdIYXY0fabM6exsT5dAe3mSyazTOJT/EyJGe
VctmDKIr8u8PPw+Z8oTAc9qFGTR/UmWSkt940JTdLW/7+qnDHuQkzDsPzX8HThZWu5QA/XG7zCVT
86p2fu8ewNnv6Thycu7T3aauXpwOBG8SIRjauzmVGm/QpUqSbVhnLFHtIXzUGoHVM/db5mjvSp4Q
MYsaqoQMa8T+zlEj803lzIqztP/ZVywTiZRn51Nur2Ed6lGnK44IzvD5t+34+JTI/5gYUUxjhyoz
5pfm5BH9cZ4Gu/eX4/JV2N0Guot+zFQAZSNZF+0MjCc752yd3YBpX7zE7ISqV9W5ZJ+8ViTtHYbf
ZV9TKSkmrd/qS2scv7/Mk51JXds9uf9Abb7SCA/KflfGkvn+0orVo2NIzdCewlYlyT3NDx6p9qmC
0+72HI+0z8dVCF0nsBXAhAG1HyqhIXW2Zzs1p0pgWwsFzrz7XCECfbw8YsCgea5ydgc0d/zu7VSY
46DI9LeYtKcZ5sZW380FHuhxQHW+YbbUNH3W8ZGTygJPf5ztVdJyvvhDYW9UHXOLLwdjcOT6kSSZ
gW4CT6qPqJXtMvd1rtar+L43x8wU3FNqPCzjQRFPIyRLe+VdRHY/fPk/tK5HK/SD1o0icae4pZkv
NrhCp7Si6BWWo1uxwT1jbFwNTWOAZtshZcato2z8c/S3+F09v74o1O7eFlXSAw8Bvg6JtnINvmob
iI+vq0cW/VPg6KdGAaAUD4eJrlPqxIt9YzZyYo+cgpfH0E2QgnErxpdghAyAS1QnHGL71sie4kgE
6eAXBq7k1xa3qM4c7SPwuof4BEPSL2wHGd1HIjF+hMEoqz9OCBn3f6Cwdr07MYb5RQqow3Ixlc3f
w7/UZ9izZqqzRJwB6HAzVKvlK7p766bKrB74txPedH31+fmJbRiR/Gn+EbAF04jphlDA+ukL0paw
j1NJ0XhFLSz2DJzbtENThmw6GU5OAYoR6r0pKjD9Wuwcz8PJSASV9qo3Tf/5RCcETx06c+gEIvn9
SBfmLSIWv6dUL+rSqaxJ/Zk+l6l6U1qXBWK6MhDr60KBt9qO6VXP1HOFzWnQK5C9Mj19GSb/oh5J
Q8Q4r6D9vGYOYGwV4yeGQkwp9tbuvfb890Olc2/CemfChOLElFseW4tSFq8/ehVzwG+4A9SnqPod
IOlEHWz7FBCYEMn/pEkmWiv43MrIsyibjdgw0nVlIgnS5OBQ30gLiOgzF3PkzMfdrTTqYyciF7DB
XBviBotKkt+zw4t3XWMofLSsy9IaqSOsXn6SsQxBB8croJxc/lEFJR71n2bqGZseY+xlS8a/87yl
6dD+7TDTV3g5CPxlrpS27IqrFygL53PTsW/nSBpMrbcqFAjnM9LSu2KDrMVoPiuj5JyRSeHQH1NZ
BBajFx6SuhX2Hz4MaH4oM38jomNPoEtKUSafaDtqvpZPFAD66W9IuuCQpQ//MomtogHoQCv8ZwiU
DRdqHQ9oXDQksenvcULC659nN1y22fmDptWsAM3lUq+9yHnJ9Fzv1WwqG3YV0U7z9P1T+nXT8ApY
kiEEr0pHrPqc/WFnJg/lKhXcpzBRQQUk8GQ43PdesUOpr0z6Feckl6P65k6JbhobVwx63l2LkjBQ
DRO1ibifeiKDM4MFRHg5XAzPMGHnYXpuR/xNR35F/fHQepfZ0P0E9CFi+mLM0xDCub/HRbjKmS7+
U955KB42zju8HOt3YcGxpD0wlPh+8OqXD3PP0djrxRYToTlKOyKLJPDgl9/2bmGSBw1eALKJTMW/
4JGU66j6dFedauhj1eGKJaFOCUAE+n3PSooHO3d4E8/cg6FfoI2+NLE5GxxoVA8zzw7iorMg4Y7a
7T1TKzoFlcPvXntvJ4f61460vmgyVjTkco91oJppOXprQybvMf3Ky8nLtfRqz9Sn+g6260oXwSpF
E3MPAWSjYZ18C2pCqzSq1uYLpqMuTgzyZQq7qP/2ytvDO+Nk1ClfmlVduI3CJ+JDwg1qDkQ/0djF
F7XSBU9dHtz5wFAJjO8ndX91dpmkKBiVB05rl6wU7IGQo2JgYOD+KCsQNEBq2ImZahEhS01JRXtC
L/cs/gFNjCI3uKpoZIAzbTCAr/OI28XJ3l80cESYnQtVUyFuT+T4oCnHJvrSft7SwLh7dXn3bzIO
gTS6sPwsw2tiHl3O/8tlkIMqaGVabhGtqp15/ogd77sCzOCRDf8jWH8KdCY8KHiAFFlIvIt/fAjA
fbkp+1juwlf9mWvUph9i/tO38QgU5W2miCwaOBRxWBBaSs4B1pyW3QQvAyBN5WqbKT1bZ3skieap
yhB+McN9mbM+eN8jeislmyzoMeIZua9rZoWM+1zeqGgb1QREXF9qc5I3liyWmRnR5GPhMVAuDujw
SYCjEC+isKAm7LpcdYnusgReaBTbsTUNK3d92/q7d25a6yKZUQYELRz7+gRy3kUiPsFYuoMDK5vY
WtsRyC0hGG0DrIPqDAqkP/NequgSEZ18f6TvJIQ2tuP3WQReHGgApEqDY1y1kSMy5M65FZjs+jjD
pCkqJNXhZCJn7dqNN02Go1X5jETIPt1qIuDt/gor3uAaYbnWNokEXjNGAcNxlFnZ6CaXBWQAWhTN
+VDMdDo6AJkQoI/hx/nV55mYwDpCzD6T73ZMcEOjUokNe3imsSCoNnhG8iNy/stqTjtjF5aWvb8U
fm9hb46g1TDlzC/KggpEosbhoOuJdX+sh9TVZi9I7FbCoxGL56UnRHCLiphHUwLGyl9iEngkFQdJ
vqtkPiRwx6q6qXwauQ4oFbffar++qWIcxJ+1w4mtK8xoWgADU2vWv268tkfW5pgh5igbKlDMzV5U
iKmRggwr4f/gM+dExxTq1vC9NVpkiwW0i/t+kEITH5mDP5mgZPh4+8ZWJ/ouJUhwOkMi0Zq5xEoP
zCyA+0MbvQ+1pkNEDKUv9mhcZT4GKeQcxmKvHwVG3X7RK1rQKuWG6eZskBqviVotcCNvjC03az0k
F+nEznkdkjYZpiiiWr63wZ5+o9B1d+x2oQKvPbnXTDTl84197yDVgJIFY+bt7kr5ry2QdzN6B+Ig
pspfDqrwv0oOWgdVsn98YZ5PQQl5a+ZPWQcZg/y8vnZsMsWcq9DmqjNms5F69itGqADjNlV9v4ei
eZv0aqFA3y37QBVxfbQuC6QjgYHfIVNQV7eYh27H49tD77mHWyRv/OlgVxsuCydXATnWLddX9j2e
e5DQYlcZSZFnVu+IqmzZDcbepHl7hQs2HNV9Da9GXBMOx/0YMZSxovdMlqN7YKDEbatdsVlpNWEg
DIeUkudSHh4ZUX4tY691QzSRh2L2jq/lkjnPQTeniBNGm+l9LHPk0a+WT5KBdKNs5iZ5A0dVZM5A
yyDmXcLX0vJsKW28fbuFncUWBTtqQI8YD2F9YMnlbXpoXjuub6SlKFjyl/M4DLQ3iL7NcOoJmsa5
e35UIVyyVLAimzMKU+Mzu2XvHob8XGArhHSQDeDK5ZPGuxjmuV0jGR3V8erueKQrZkrkPICz2sMj
Lvi80UDk7ymD2VHoW91NRaWrG4opXmd+yoiQW6pvCRNuKXOtkryKCKz7rAx/1PzlcpuXX/nIByBk
POokmJEolBOqDKiQNFEzVjhwdBpFrCNdEGyF/SBsRWtQmZ6A6HRPK2jL3Z3O9Ql8fpufuUwrI1da
6Y5BTgyDYe275EI8+ljokapiQVF2Ca2J0t+fKrnKR389yM/3rJ1eqeByh7SRQBNgZ67Aul8TqBv/
9NyNYc2MQUyQn8KPHF47mGLxiz3DcHOtWR1T4I201CeaPhOlvJAYLkIjxXlyOqyR+LuCYi+jvzKy
QkVAq1dnuu9z60UIwcEWP/gldklQ8SzXJmC0rLyQMrQQFpeGDoY6zCUrkbEDLbgf5a8C+Zztx7qt
clRBlQuJuYAa9y5nX1NR3nvLSkDgpszVGZq5Bj8/jze39ewwXPfvYKJaqnimq2luOLRQ0Q1hlXe2
FTUKizVTfBXRSgkuLkat4/6GT++sH74ERTb6iSNHjU45sX7VsP2E+jsvpp0QS2u82wBjzmYFE1SP
h6SRPlGpm2W17VCOyTxrEER2szW/apNTg96L4JyfEInKLEGdoJMKoWysdSW0d5OzS0XwbOheR0h3
/wxlUFRrFK9tVBkScHZD0V8yoXp/wlRR5JHifL65v0Vr/VB4eCF4vWTcEt7rp7NR89sKOLRf7+Rp
sVLog44JqvnufMjtWCPyET1g5ON9qM5n8HtF+7MENj4T7zWai6+K/lVWod5RH23eNxg4IMElkO5b
Q7AFcb3D7NhWTlZU4AVlVmwQPGL0OcOdwLIDK3UBkCICqHEpj0a0oEA/S5+dTPFBXuudsfk9/vT2
AycwI/2uD8upxWKC9vIgVf4GEfF7KG7LAc288d0FE9mLg0eoKvsxy3U2UBJ1BpaQPTJafdhTM8X+
c5nGUjN2VhuEP9mYi/djcD9HiWBKz53CTKW9UwVKnXLkYgJCTv3+zA3Nqt0TQc4Ke3ay3ICspLkM
N87wpiVol36CM+BTFU1XmYAhqBbPWVaYdUQvkp+B7yobIjy6zFAeiBeJtK3WUDIzdlvLZV4QfifG
byg0Gf80t4RNFPg5W+69gLC76kC8DFJ4sGfT1LIQzfay/mtljIZMlV+91/D/5T0FmozcKZX1e3Y8
am+2SEEb4v5AQz4X0i2IUvrVii9+VXu+p4irFIX1Eu6k+kg6uV+Z+C7i2BC8TvP9XN8ly0LrvjbE
r8B5jzde6u8ucqTH1WhJc4VfM9PkIodTLG5hgfcbDE/T3r0dMXR/H8s63t2d/jwG6nL9uz0Wi7rt
V2Mcai3+AvZgSHF4CfZiYP6tg1AlKwP3aklN/IWi9hAXRTh852iIWru8NKwJNVWkCsGNfzV3uvVx
MlHQvzeMH2JVba6xhqs4MX2UwAVZzj4Nx1dHw6EVM69mA+H7Cwfpvh79DnUNk8v38y2HXS/0D0Mp
ZRzzqaWJVYEM5KxzYxUWcm11dopGxNrn1N9KkuIqIBs9mCvMGIMHlEhDto2TLr7gFsEZZCLgyWu2
fOsPHebP8y6tbX7H/b6qFSZ4ACxU1UqVJJrpawat5AMx+2qiuBy5vOl6ppTiUBeuBWnxSr7SLZfX
IYOGuQXNsRtDsLiRGnijqo9rIG5AorO1CUaLPsc3pPJZ+mQ7pVYB/wY7P0kTvaudlLJvoG9+hnft
QAnD/yHN45Bb6XnvjBBwnFVpKzkYy1y1mRmgu0p7Q5zabz9zwHthLUjqGnDpE4cgCPL0hJJwE8BO
EZ4q8LE5YI8a99VLhrcNYDzVMKKwvVzy+6bLAJEveINgULL4NYoMPos6AU1i7AcyyQgdClxmhG72
2MOaEsvRvE757Woqe1Hi6o9i1SCM/qFgjh95f4jWz4J+DEdCNG57ZQtsgj9fXJmgDY6WYxFAfwXi
g1gak4MXNybJmCXESLMv8klxD3PyX/5Ym0kEGXwQBCcc2GOU0Lj3YD8A1eoXKEunBmdM3KbyjK/W
Q860l/U2a1AX2yFJ5p1wsqRBeU9IT23hUvTqg0gH2+ZEZGTJuyHssqkUaIMo4lFkXZ3/GamAW1vI
p8p+pAPnj7aztfK8c/NqydCt9XwcSud9tRB69g4F8eKT4+qeSrBgie4QotzyvElEBXOoYlCyvpVA
nRrOA8F3twOpbhbcwTuE6cSh0ona8th1QGXtMYJDv6ZUxmECUbdUjz2CqMBH5DOuQyAO39k8Ats1
C/pD3QimqhoFLOPXNgqXjfF3WLUFIKs/Vq08VBIadQheTaresbY4r01gXldurA4ww7dHZ98aKSnm
8Vud7TI1QtYMwlAPE7lR/17CSDj1KymmaSw3FmTVa0lNbWeOEC160GpdPI74imM0RkxF4nPZHueu
Qv9+mEDyhZChKHfnIgzze3bBE53bmUUq7FDNWOJXYQGyDeGgl/2cAS/kBuy4+Kp+H/stg35vifq7
Kz1MrXZjwWOsD3CW5CQt27mNOUb6DdKKWIX164WsEvtTEf5k/wRdiIZMYsMm5gxzQdY7Fo8OTE6k
kfeNP8MoGl4BiOb38HewJ3bdLYBXrJpmN8VioHLYvomCv4dcJtUN4p7VRTID4neIUwJstqLdeK24
n9DpyJuIqlxTPf7RzpbdTNfAk0UlBp9QFXg1vnpNfZPOP7pOhA9F2CN3y82SpNq3AQUFo1k0cCnP
CJvCA/t1Zu8R5tFPMwrypiwufHW+Q6aP/w7LuqO9TjrWwvFl9I8BOFc3SeXepwhOhDEDWyRRB7+k
jXfx54kFgmrMg/nu+JKmOI9wAr3bfFPDv/NnaqOYjrQfwmTPGSYLnhpHwDKCuIVHOUapI16cV/XQ
igyp0+nLqFf2ayJbhTfSTHDFH8iJRAMa/O5/ac3ND0JzVIcFxzLekBERNYVTY6SffA8TznLFFxyA
tmPucWIWnSD7HPRH0QnUbtO6ma+BxV3zHOhLtf18gZd37qiymPYHGMUqp5faJ25pBWLwYmcFO/cG
31uUK6nDz7wQYOYin2Jg0DD8TFBnvUZMkM2nl8yCa4oZnIeQYnfa/ot8j0vls+1UAwitWy/5VRNe
fKkQ+7EbNwQ56l9ys4ZGZUxdoIMOTNV2h6FPwCfnwugIp0/OfAQSbCq9dEB4I2WDv+pukqbSTpo6
I1ljiZVrVy3OKSBwjwmg2MYzounZs9KrtN5EG9aNwmPzKWxb3WKhj3LL/t9AuXYeGY5eUf1lVeJF
02i35X5jVh0r9mMaagMuccnVRezRSjskWLxqveRQ7arl1CmQfbmkPaBegQedAI/L36wwlbDENDBW
egjksKVluokEzM1kdHA2TvEcmzS2C55ECwDYiQOa7YMlDfAXgo8ZLHIJNmklwPUSjydLJ0PMf25M
xP7dld2C2+HU29mDKWlJH6rzWnCm/BgcTx7tIsnK7hxiRWHHMBBI/x3LqYN2iI1JsMh1Ne6suaIr
QmaThSnBleaxFtsgRsiaLDG2sp/06Y6sFK9IGAnzIWcRQH3OTiMBZNVJdoOf/1VpaKg1r+G74c06
t0dIYNoAr1WbJmwT5IUZSPCK9+h4T7+dUUCSMJzQ+/SueaC0y+BZCrvfOHGZJO9zEnaFlBFf8ITp
xffj3LoBUp0eb7AjCz4z5AC5j9vX72fEqO4lOzz1SvLBbWcv1uB1F9SqDTyuAHcrpIjGvxoBBt6E
gF/am9RkiQoxAqGAqKjwTolq4SzuBvD/MolfrP+Id3B4Pcp6K+sm8Nv3v2nzLx8LLLEp9xY7ctOs
LJyoKSUf6S2a8WkAcpCiG1L/27VJT1PIulXKp79H9MxRT2pSgFzzfyzWrnKCt3qKeVXb+QjUAN5t
0n5mmajXblkKXLw1xfdR8XHqc6Cd0lRB+paAKMF5UdmjuWrN2L0X5zv4QTc0fopwMsB4LtgRxRmV
buFWn5AM+n4YL9CSrB+qidri/8qzOqhRsV8Jr6brMpi2+pyPf/QGKWXa0uj+4tBUcthH8NHNRjt9
Cyv1cQSmPPtrpZA1TwHI3Yq6hnYM9BB50dGFIsEC4qrr3RXUxFSuBFOyxGSsteGZG25zqnkkfSfY
Q+QEj4fwYzSgQTy/h4RuBDf/E/GhX8vM9v/wukWSXwjWY1XcawDLhvPcD3AIiohnO7IccL5XaK7x
LJeKZaXFzjssNHWOQBhPL2W4lpx2BY3Q89+yMj/A4fv1Vk8fZ1JP6ELPbvZ9InlQLa7eUxSbDkTK
SHu+IrOwPb3nHGouVwHBeuYdFqG2RqCffd/eg8yb5vKqcwSLFawTU3ORaVTAOM3elZ94URqHXsZN
eeo6oBhBsaH1F/Jb3UWmoeyBdjHYVv9QISN7j52kNbyAs01JjOEYzHXF3l/KElKEDQH/U1ynmnpx
J5cey/NLb5Ctmw2bmJZ45eaOHb7XdyPOUv25vaZYoXDZAFvv9e9dJ45v6aJ78L8Z7vQyDdzydLYW
TkmDZy3InKAOUG9lGwC3mxF6VYxULXUIPFl/czm9ZjZYrsqdItOhvNTGceVDLg84PRAur0LRoxuT
hhvODmqwmKkxtOqiHap7io686xFB+bRGdSrULxslaYrrlGklsDVrkxcprkC6UijwbjsxbXdu/Wx4
Cs54CPFx7j1mE1aLBp7BFTYIlrnYD4UayrEzyH8WwPcT9m+uNW/8/ZLQ2gfQyGQUnnjRaHRN/Ewy
+/6EAxLV17qbBbafPZNAKMxd2YT714F6AgW4zgBMfQZWUEg5dRE6s+4HZVNVrlHxO8fyqGsyGto2
J/JlCYzyndu8tPSyUoBLnG4QWKmkCXrxS+QiVohtnlmPvqv56oJHN+z3Kop0/8dAroCw5T3ORJVC
+YsmMQa2vpfLSPA5e9C4vrL3WmR3ACvYTIq0CuNaERfhKhAjuagpXHAl3YO3Fg0MHZ2dAAKYdvZd
GNPEYa+s6Wah3QrS3swPT/Wvl8C2+l9CsC0Tfkha0vNKeInCPLpz3WLrrwxhmIf/QG7Qf5ynaTCJ
U46kNOdCWLSWDwms8CinfCwK15r9Ty6ohI7YAvrpgSRx9NSTN7moUTIO0NlHjoR3L6IGPNEsgW5i
tWqIiCip49OeKyTxSeQU5nAfT+gxoxi4ZRIe6FIPzmN4PAGq8E6SHyhIyX1KIrQG4RoJT5AbvT5I
BAFwrnkI43PY5v71fhVKn9MKcZTetI1ciNRHKycViQBghibv/ZleP92z7TXGf8I8vbD80GM/10KB
SCRfmYdfk5O/1sHBzgBLTKraYgm42UZ7Q2Xl74C36o2AbAJJXc6Qagx10AHH7GE+vpyPUmE09WZy
eDsKWtsKKo9h9y5w9vxqm1lZ9U92AHi0DZZY/K2Qa6GBM3UffCyV6yHu8De0to3vE0b6F13TLBLF
amFRZs4v9a56AlL27cYMT+SOH/V8uTldM+JD404NsCJb7czi2GYTaAdFJFIhK8F0S90abAKiPlAk
fJHcZET0f5ARC/oQLR20k0yVu2KpdRTAlD0lj4AjWVzCIjmKGcRQzaB/gec0O4QDliAbZlgQNOWn
EtJFlrXUwRCIFzLiipySAow/t6PXKbpyrbn8x9Cpw+A1OhtiQPTqc8rD0m45J393cbZrUAiDx6J5
OBwwG00yX1rLO/OGIAHcQngFri7YaCv+0UkKpibxaW9B+hrDwMUrd/Ogojz9o+qYGPgTPbijA4HX
DJCwVSSHmS+Nnu/F4As3Zy/l2tfWFgz6adV90UC7KVL8ArxnoXropuD8hQ89ibWIXBpejVhugKFH
NRna0KjQR/8bE8JEySJxrJAFQJLpYeT/fP+rmQp3QHmhEVKaCgjmzdPKkVO43w+6NEJgXtYoodh3
wAk21Ix3CMa6BP8uhn8TajVK2OEc9iAtF6n2/PyB8EKmflwLnoXWrcQpmSZcS3pOe3rNfSJ6QdQ0
vkBHvbsTYCpEqyLgjnGC84NwBjE93raH3+S9WPlRbttYqbzQLkGX/SmfHydpD//WvE+C593UQ8ME
UrC+fCVOVcKtbTAEFz7hKBfUQmkF4UtSqze0POY0uEZUBRwWgJkSAXVP9I30nkSoNWQ8Bx/9V+Aj
f3jaHWu5RP+i8DlP4h/y+J7oms+zUez54PqKMZTPr9pPbD5r/xLPFE5lhMqmFmcUklJlnNNFR6QR
9L5BZESR3bhFViUwlBR0SHGHcoiqP52/BNsIFFf/ao0G0PiKl0szINSXZj0WB3QqG1eKe0xjrX8x
R1t4tE2bQriThKBUlCDdy1ncOmGT+zpFpCQqv3tyBUeuxZDHaeg3jvOkN1wdPUWe6nbEWWF1hQLW
GBJ0bxyGv+7LEaYZmT1S1bxAc6DQLelvWPQVDck0/beBqESCT08FHuhnVX3KsKfGx0lo8hJks6T6
3sex2DQNyZiBY6P1nL7QEAuV1OW4vL8tvUZxWOPcxmpJD86eqEKiUz6XXlyWt4UHY1iNRANzEhNW
jUcx41sZz9iIp7uE6n9zDRFmDbHcC5PbyCpMOuij2XWp4vjnWmtfVEoY7kD/kt88gcPpNaUQtqn7
cUCpWKLt5uL3gZ/mMHKjoNCIcDRs6OX+PCQQ/nGydRZoijkZSS9r278JdYk7FaDhWKavNQuWMgRT
rG+FWBZrrnHwyHRJWHQIjavwO5wH3kpmFMOwkjv3jcN2udeUw50/Zjwn3WMb/DKzj8zmKlJzpRM2
6pKiznCzvS5h6/SwXII2gyl5Zr0agM6MhO1TXIaUea90/Lv4olEaSDIWSGAwU3chBpd1XE03S4Bx
5tIiiSq8XCalJH4LT2kuCxZTvTrYry8AN0mnJSevzx+eklSF2KuAAaJxcsZLVRzLQ6ElkNTKGtPS
k5OT2BOFt6mGfm1+bv/ZrGG2B2wClZ8g5P4a9/WHmbE6BYRJ+/HSxqnIiPskqfvGw06RttPIvlJi
cDzrWC7cinQHTv0k5Y+JtUOjjHM3hPWX9Krh1/NDC3PawcpZC5KkzlVeErgWibaumav+MiIK5xYT
wLioIjdFAs8GhyYqzyUqCmfBDIXBTcOxxCs3TVyoqcvSvp5VjCBdPFfOnJ0rgBxO7Rj6w51vRlAp
DXHg4dN34odiWS+2PV5vWPdrMemSb8na92Mvlcbmx7AJbsvTFaUD40uhYregV75ciwIeXaYAzpm6
BaVLFRP2G2UmDm7XLopjZ6Bm/Amn4d682zMdewvnJwxHMSiQbq8CJ8q1tPKwGeI9VXhHkw/3Nbig
30/sUXbC08QJrtTE/pdrOQxEyR0A21hb1RdVaVfwQyc5OC6NIa8mp6GQClONWZib8oaO0SxqyFua
diGPYlhfEvB+RpxLwTe18kxZpDjntEfxg2uD727w61NCn703GC+S4iBaSDuuHBjzOQyfbkxP43+F
7CjELktEXI4NBla0qrpFbZ6qvgwscx0mlG5OdR3zeBi7diUTBVcq/JjVRG2TLfdQoBCKy/S5uznz
dg/q15Pel27M41aFPbJxl9tvj1FyUIG9wrKJNx295lUC5SQxAtLH1sCeWuQdKhbGzSrGfOV5Ilgl
aMtbN1Hba2KdkmPIxxp4uVia7jJnOwRQ3pv+xGIS2v3GBw6qIkqMmp2a0w4XvaYq/ZqK0mDwptgZ
5L/3l4WhVxPAI2den5X+mNfwVImVQljRl5pFN5SEiF6+9gvzzbR1sAlqSyrHbl6xqw6zqGV/NVrs
O2oWb1JkdCtQBaVH97ZtX6i2WyaRXYzi4mZrG8ol87dHOfeTHXBxidj4ZFRk9FWFg8EDaXVVB7xR
KgMWPn+vEKHZlYoSX3Wm5rJGFzjx7LDcRvXQrPC/ijrjT7yNp4fXczSc9HFCSKz5QnkFhLXs0S+7
MG8SajxgvRdp6CJJtdK+LjqHN5Z47lHp1BWNbvHjUDr5An4NvXn13lpSdqR5ZNuaze3IW2lSiAsf
U6j0sXQE5ih1RZF869emH5GyJPIjax+sLYZAGTyrHrzFwUqecUZ+6nuUyTo/fDsB39LsZh0SZijJ
nKfwuWrbNS2TslfmxVW/W124Gy35eCq5HCSV21J4NbOCSzX+SRZTWBagrsfVmNn+Atf4YpIgSC1Y
k0vqMwLY6jKczepR633duE7cidPttBacmvaDP3X0GXJx2mNhXK/7Hin0XBQvTn442+q00lQiJSru
tWK5izPe3a3SjJoF5u48K6scAMxjE/Q+gd3ryyuTjARRi7KndvQc58OHYL8N2arHEOXYKKXvhyUq
YJdLekpNmRWHZgk8aGbFWHVMEcEu1zvX80iC0UdGyiG0JH1xz8ZgWLoHLo5imbbkOHQ6/6qbl1no
Y1dMjMCPbRtVCNqfFd/qrbW0sA2tOS7QB98h1h32c5XA8nPvGZ10c7/1LlO5F1frhpgbqCnWDQfF
csNfxRTPNu3BQhT07vyeSJUc9xSTQ44nGmruosb6MXcfA9syjonZlTirQ98XSfR3q+BXyyEzr1xR
UcNvOZr4YNI3wC863hAEHwIsKzUhOwCEoLyt8NPPzeRDi8XFKWy1gSu4X6ibUyNoMXa+5llGW5qR
QbxtBCnBhi0mX1FRjCFO6W8VZhw3RoI2RJqg3msryu46k2OuUFHOqE099vCJpFEAVSw9CgAV1ZYC
oEQZem/rL/JYKfEGIOL8cf6Ww7UyShRJ5HxIca7J+KqjFaot0UI0IjoQ2fCROTxMlpRfWi+xyAlT
/OHAnc6yp+BozYaKy5WvVQmt5koB0UYPBuQn3IUEWip0RQ+jK55nXW4OjGZgxzjr/C3RybpKX6vw
/YUYT4GDYJ7SjhaJklmjIvhq/eBxskxf8ruFv0N95yJkkfl6FIhXlvL+2pfIWCJcE6GZ+qpG17Uk
2YaJ3fyAYQbnecB+SPmZWerBs4pCVDNvc+IKwIN1vdCYTVAgglAd/t5zGBXyeb+LrgpHwxp7Jn+s
MjovxjbjMK3f074tFGcWOpptZxUkboIa0ItUxqgWnUDEU6aa+UbwPVc1lXeS6tHQLXSPKBXw4OsS
4JEWW+phEPNR5TvF+s2dncKaGkMCLqgo14c5rT/32W0W2/wYQGh98HITm/bgvw1mc5t32wO6nU2m
IPbO8dESCCqGwvf/KqN85EO4ekBfTyOULBs3Wo6vSaGhTWrfk34Bpcm0HzWVcOYBG8mgoORiDB3z
UpxQlXmetggq3t8IhzRBqgR8WhYCcsgT3X5GEV29UpUgtbLgcc2z9wtFJrUfHebC/aegs1noikFm
rMRCXCN+XG3QRZpgg5XJKhLKKxFssJqwNPPqseicH47o8cyrXFVnruJt3FQdZxr5LlVvpblZsiOM
/PmVX2MA2ljEiokhAXmrL3pyv7z1y5Do+KXukyuZx3PJQdBK+Wm4UDGYrhyTQcj5EedYkeH/ef/n
ZLMNbzf4pq42khBRF3jcEDcSfQh6vTTlYV1DImTJBSDho13qYhsphxYqqOvq582ZNN7aBWeNNeJj
olxCdx8jLMpXv6VwOFBktc2FULPU4CbKPGOIul9njzVWguik84lmLg+Oa3GUS4GfvyKyM8RQ3TuP
2jmRnYixTtg5z9lRSBrU5uFiRWoMPD9Cz3ORNR/qWMnozbRiUrBlOBBDvSn7kv0Ebu2K1s50Jxtn
mmvAAopIlRjfbGlCowNks1VYLgWD1OlYjrVk5BFwWX1L2rawnBl26S4oolEAolNdEPc+FS2oIgNB
41VzscCaU87FG5r3nXA1gMXsqHV8Vjrz3Ohjd8pDxYjbiCEMpMe6ZdLI9FefL4hwTPufamF3Ydts
JNeESjM/ODRxBdpQSKcLw0nJKgBEbKlLF2Phw+HLn7izlXyDb+oyEFb3Hd/mR+RRP1hQxnIVrlz3
v2htplbeIrGcNi8ug7R7nBS74BB7A0TJqV6jZw3CuWnGPQ3F9/TSFKB+0lQdDCHWQ6wBF+5D5Mki
MGmh+z72hh/h8rbm9x7q1oDiwF8iHAgFU7fLCQyuTJO9W5qwen48pfwjoxo+mAKGIGxWm+fM9OVh
0M393NJWDR8sAAh//mrA49Z04ExENs3hjUP14r0M4zUliBMke3Wz7mf9zPUnwu5Zqyonpj/3TgQy
yWU61nPPMz/4b4b6oKpBJSHPDmipjvLOZM4GdNEP4NLYYQSLBmtoElDYnBCNV06YVV8LpdAA/hzH
4fOqAwf9fZCDndH1Udo3Aj7d58e+aKWt/S42lxyioMyzMzApqkwfFf9kcMuIW/N5s6I7zbMiOPF/
su6eWpQ2Qexr8i/e0VRdzmr2w0TJ0jguL3uCb6auWbyQfcLmxP2UWtjY9uclNJMB8qaVWVOpMZny
BwLdDtoZdytfgGeh3nWb7U7RfSE9VXJrOQR0oFHeok1cOt79U3mc1Pjh8GSVv+7ZeseImv+X1/3U
n0U1HPnpvYwO4jqs1uK1lyAN+fJ35fFD1/i/khOtexlhRNiXvQt7f7HOntOc8BIZ3WCQGZ+sb8D5
A42M2MtDuo6izuq6k2UR8RmKxabua1V2luG9AGN2QGC0zVfsMVuViekdaH/T/r5ntbzY5YdPHaJa
useUyWHRy4XrEHhAj9DPFkh3Lk0xoYc/vbDcke5ReN0XjVdSk8FvQEp0aUDUKz/K65UgEzft/PkL
mlZ8OVz9xGh6OJv/EdNtqGb1k0snLwVsYwvyKosSWu41r6lCKnRmUq+UMX36nrxMpkjdLjCkJa7B
4wtFn+BIYg99UIUtxqHvfOZdzbMzuYcNpbNM/DVVRvegD5FOgmz86vO26Y7PQxcGN4aohbX4wYx4
rI/DmQGGD+ogFSPKKk39RDV5Cy2/gArmBGEuAng+x2RfNiVSVysSgyAMCFKl5HTRGiLUch7uC+nD
v595SFgdyqZ97lKQu639QffwB4fobURQra71ZxxgOe7rvhxEY1ccugrdtlSp28tpszYg0MEhjGLd
JrKchteulzzgYcCQ1bKcyhB/FmvLKzIZqsQuI8xt1jow0eo1fmtHMfJMZoBTbdPZyiJVJSTsceaL
NYqBR93Nwl+tkXC3H4zigCjIo5NAehZ73qr/Q2rSYlc1Pp5ewryN6Sb8eD0ufVxHZ7Y8dlQt2bGo
G6HNdcstLhflox+00SaP60AdZEkGk8ozRuycpcu4P7+Ngoz8ZVcBZmxttt6KhONUKL52+HeVKOvJ
lgcKrkMtOmK1aHA1k7VwgzboEgGkl27HAJZaL1aY2lLW0XZIWHjE9AtBZVF/3i9bAqocvvDDCmNF
5x7Gx11wET6NCLEloNBUiqVXP2Ogiia5NcnE0U1un1z59AUb2MYYuwlHouWMstaZsW/uyGLmayAc
818rHxNL07g6c3fMXaWq+EkUyWN8A1TtvMqvFd/QwWJXhTrPHWsATOiuWLAGQRwsUJraaWeeub/W
dlw6GlDqw/xKvLwB100KYcIpJt5m6pRpd/4+uTaa4jxmcVi0qtCyiTFSh3AC8zAoKfQx7GkYdISf
p/8cPwohtRMX6I2SorboW0h9tX3VuGKm7ehxU/yoROJbHXkNEYPwLDAUgm9A2dwrEuUlaMN+Fqm8
XTEDZDcTeBQUOQ3ZHaOfxjwR6BiFbZE10HVcHSGM48yuTg3uusBWOcj05VIyuLsFa6aOHSDZlcVw
v7wFyUOtYtLIkEsLssMA+rEqbD+h5ES7IEkFkfkZa9bt8ZbiTyzW6lMI+LtcsNugIkHI70zso5g3
NCSInogdahvoZmbLAtsyOFVngzkmGVpCDuYnkbzVyK/umcxMFy3NblhktrABXjlO4PKvuYqLDCXc
YiXhPDRa/q4hmn2FI7Hl6NOQ308r1d76tA3ryDzd/vTNs32B8tgdcHXBQH/OS1K9ObSHWXZlTsha
eNPtkPwJ+YUTzmqkavrnt4QfHZ0YkuXN4wI0kjHtIuxOShcMKKP0Jqx3Orq4oRlr7OLWJdlIjrYi
lhp3DGbMTb7C/a3QGvJDfAzOxAFuXu39UOWEqHYxU0jgpdzqFr0PISNU9Y6HZIyxxkW9N7sTuXN8
XFYeemOfaheAvePvFDoqCw36Ij6Jw9E9hCegULynxPxgtX5G6sq5lj396CYAmr6jINDIGMvKQD5v
9onhZZY6gi05WdDo2iDJdxwZTg5qHTb1ggBg0dRl3UmyTDMWhfR7XV4SzxpAKIBGX5c8X5qWdfb7
FdAxXVvCPHSTILvIRDaETUuwSs/OgjKHDHc7ohI+ulYT8B2nathoIIGGqEnD3kGhRD+BL045dKqa
p8sttKVkJ9r3VBas981KHaEDA5vwonLgZmMxeWQBggxS1nCJUVfPVB5vMBfC+4E91ymjN0rtB5t1
vu11VC+WUwqbaPMkCmMndKZSQ3hkxlNfmZCSYDwqy4380XzSgdagKdAlgGuAe2N2S6IubW5a5Ags
seXGdicJrIzU0nffs4SaPMGkMXSu/b06yH1UdfaOJnpAJsoYSWIQVrUJfURqNsBSHWDrI17pIw0g
It3a+6XVDm78GNylvh8XaarFZ0aQV0QxOzzwU5dp6KTNciZpqSCk2b3R2LrgFgEO9eRWEdI2Ny69
7qQjIZutAgvrVItIyRI5lDjPmc5Q5aKitXw2epr/icMm6MkcYMENtngydDWeB6JDBQnr+QpJKRds
VR2T2ZVEvn15IQVv2Z/HttJPy79b/VovWFjGmcvlHBLvAEjd6wcAFO0b31Wj0sabOzB2Fkx94vR2
93jduUXcoNbKy0ApCmpfEGUCdjezwVAXzfuxM1oOOqhVfd6xCB1c5VImYot/OYzpe19px8126RLZ
An9N5m9RkyeDkqSbbA5qXPHB75+g2598dmmTmyEpUtEMFINK6ylPkhQEMRpYFyBgP3/ZELGKI13X
EEYKlrjJr2thNelPxufPz7Z2ORCpScUhknNyxucPjmYKr5gJ+sMWBqYasJNeyYKIIeYw8qTQx4cO
+YNBxIoRd+xEvIyw6iAImpM9S0zBC94l2mzhPYupqkzo/aYK/T1Mf8NHyVp96EiYro4aN/2uwXPK
i6kzYDEmuFDP1RGZckeDYPV8NXF0yiqZqo76bBplX9/g5cJcXBX6QXns2BeCetuVUASruNYo8RAI
BulZVZt8qxOf9h/eQjIyWXa1GPL5sJJnsvZ6HsJow68bMicbBspEry3uEpHT2OlGq1kCLsTnm5Dj
+92a1nvXQLM3UDW+19uFq7fE2LAML4vnfhD/Nfi+mPRkzb6J3cXEiPfhG+ctHjDWhiscus6qHK9g
olf9JfXLwPPAFqFtRaDfIKJwk8kjoV741Azj/ss3KBdBJQfeEQQH1cKqZZ1366RDVJBcUj9iH64D
ojnhrRqHXH9p2wGVNpmsRGssG6G7/M89M1LmXSMatK6Ns2Yt43qAy3fmQ3Ucb8A0WP+gAEEKjM2m
/ZEe54ECQ5f+JuUpjGVR0aE0orC924sPYuUXJcMUXrDUW/JPvehfBmKlbDlDwEg6uASQ0o+LZrtY
Q2kMSmdDvB6RlV0OsJ4gLJuVIGs2olZG1eZO0Xv5led09aQ0iyYvEvFv9JsyABzbOQFn8j9bwcab
CeBDgU2/KjV0aVgWA0zRg+ClNvejMjYM6SbaxqImTUHwYQ/9d9WnwvRmwXM+kyyl7vIS0kafYLse
gEEg/B8J3vKajE+1SWDLqFhQQ2f5DJYQL1jHc/mx/EwhrKIH7PTENkUWU49leuDFvvp3FhhkXL5t
/RtOaJCD2G5lZMkcgSO/oKF/eaoA6jwGfSsOOwjYEvLQFx5O1wyxfqTaD9Qbo+kLdvyj728jg6kd
yGutnKDm216QbuOTdpNmictB8CJbCsAATH4vPZ6bCJg9/wsunm61h/fNHAFJRnFGcCM84b5iElRw
MOF3M1SawZrpHgpGDM2BDaXhcew3Rf4dznUal5p0g0q5PLLSWdlWxAwp00roK66oCiPCe+RK18Mf
43oY2DuYr5d4cOM0XrLxDoHHAASjJle9qIVqXKptYgbOm8pVul3EkdfmVFS9zAv0puS5U6S0mqRn
aYqd5hcW4ibaOaDbALtYEKm8h5dvnlovA5cODbkn/794nhCwRTM7tdWE11erb8BdUDNFiN3z/wsS
g7Drbb/tMrN4UMshiRtlg5xCq08on7AzyHqn7w7vvaCuiCzQ+dUW4OgHD5cqNtITEu6HwKuCJy1K
RFDxP6K5uQLUb4aI6Zrh0AymosJa5dCu89niwaxpVX2yuLhctefBzVgTjODzkDr/ptTA88yIWcp5
TmIZIaRguvwdpZjskTIolYsRLa7cf4+sgpJYXJbvFsjah7RJc6tCHFLwGw/ozKwHv00uyRAt73X+
pgGQoiBmHPIupCqKAWlx37ZAk3M5yKYeplkmxE+dKW5DcnmEVBEOZvgNB5lZ7kIA18nklFX1hfUi
fuEZCjnPvzY3+Qis7eaxyX2FfzfcR6kbG1mBlLIlFynJJaDbYPL9Dsd2SQ7iteTMBG3GvRqLEgWK
jn/U8JPUilPX5bqYH2zev6P2dm/ppXhTC7FuziTf0R4qrhLi6HdMrweT6jimTHsTPOLffiBQtpvO
UD2daLBgiXzJ4z7Y2qjmkwuEjTF+1dEvjIBDyS1NXs7SWMaz8pUXRspGwjwkmCjwCqrYDjvqyOG4
aDmhB+l3+h4sHLn9SK5F2dOKosBIPRXfuI9JNxXIQLnfEfY82idGudIR7ugRy94oz5howCmyrNjC
mktQH45CXqMaK2QdUyxmvMkh3EPLA6U10sNHANinva/an6AQmQYjMKyfHW0nDWlHqr0tzoOGsBv8
ChUBDYbuGuJl5k7Pu1EMos3D1cDO/DxR4XKOU2J/dlBfvbGLwWYpqNfA66BllQXvjKTmQGbkQlvZ
x1I+x6rMNa2ZPxB5UhYyU/3+1dalaWLwJa4bG2m7YtWZc9umcsRsBSpMHAF8LtaB/bD+1mTNnYe8
+qnLnR4waZ2yAXrlrUHytRk5kMctfmWYNmdb9STK6gc/n1wPQtjujAUW3pltEq8tzJSaaJVxH52i
oOc3qvBeTAsxTphUpmxzTzrIkejlhGU5oFRtCqd9pggXmQ6V6IqBnepL44Zs0zfgHHOuupdNFh0C
St+eZMvjbkhPjdcnBSsrLOG2oWROUL5tpUd6rDDaO2CULoIbadmJKKpIYd01SU/MrKavbk8R9PrQ
E3ilkSLlMR9nciPVo7hvMuKYZsYyWOqogzWtQWa593lFvWQHPxaB/BsDPHo3SCFziGxhvkN72u4O
McwnE2QlnqGNqcky+XvjIYvVmj7NzHSkJoqIfHqE5LTSo+w4k3h6i6jSxel+ItuRIMvjnCg9g9YT
tcCj96MvPC3+5zMlKEYp/5V9pSjAYyw+zykr1EaoDc9bWFK71x8w1jjc7Lol0LuK3MyKdZyluqeQ
5FqhgFf++tYl29YnOs5cprUp6XwWwGlbwJfYAL8SDZ+SkucVBlC/5QeSH1HPuKX608lg0/XRUt8g
n+cFl2mfsZYZN2QIjUUuvUlDYFu0xITA782zzTbVNcnaWOQVI0e/mQNOqFlGWT7G0mYZcTqM9NrM
2w1XuOzW7M+UemrnY9XKYx5jbQN9wsRZQq8mlu9p8yECnEb2iDclaZodHKzIYsS2qL8CpglK6z9b
x1NWmLmJwd8DZVAu+vXCnJYp6zBhMKb01BaqE40+h2kmUbcz1riLwj1g1wNEbq6GqfAE9yCaO1RR
9Fk5nTW9902NxDi1/BfzeNfYSzXuXpwlQUauE6F0w3UvcHsuj49R53v3WUYfuu3kVIFOlkyFjbLY
XY7uSftbIX/XR1KBDa6OBfj2nyJaF2kwijEZ8+Zo1M//S36ndndQDah7gTEZmjJGkuOnCuJlYUnx
tiGzk0H4pU9wq3GHHrVpUOYY/DAI0bSIca+pPM7CujJ1kn3MHNpFlOAWeiIv0lm0HxhobiiIMeo5
OOksWpA9K81YQKNiTvZUCq+PHYavnAzbnUH6viQwn8xlIoKz835cEZCnXVnwTAB4GsXmycKEMG0O
8iN8QRmc78uZYpySWxxBfuYF8qMRsrHXYV8laIyNGFWkX9Kf6FMbuxWAcgEsfj90FioB9mOZlJ4Y
g7g+pEutAPOcaHHA3LKOd0CNRLZ0fdy78BvZwvuIq9hEZ6i4gQg4sL7UIIBFwqUS3Ns1L0fjXbMg
wc7H90nqJhdf6vzd+CI4bEF41lABz9gNlvG99jyLond52k5ZdGfyQ01gBI8d8N2IkRPATHOSOrrL
KKJwbdmQhKEfJ/+oRWw2h0FJOLuKs4FhriFDgb8OtWS9lG61wrfzlt2INjaIIf5jKsUm3n2Uqt/r
tL+DXpZB9cxJsmNmMkKq2+ziIB3/k/eiT7ATuEGHHqhQ5PFLuw3ICBYzoe7Fmxm0KVZ7socCWcpi
FIYWJodKvFv+h6clO2zMUzT3FPsQ6mofkV1FR2sy+GU+L3APFQFiRbr5UuJFnem7XEgHHSEaQ482
4QiBo0UoNb2w83z9ZjiWTt72Rdnw5eEBUHlslaRmZu2wN79lle/0cWad1kfDFShT0duMTL5EjHZa
VM6ESncPqKX3tyQ4jYBlupbxbULiP8V24qWGOJYsHc89J3FwsF4hJQ/zmBvWBdobAGNtPgLILRfb
ZeXlg8by+qJtunLDTEhq/uH7JkQwjwtaB41J+drYBVN3UdGmWEGN/neRphgl0y80mPw/TI2q9lZq
9Y7uI4bmHWYq2rdVMi4RE0JdDxeEkzMoZCz48Q5sXriIdmQXN3ly0M3vOqyrs0UyG9xJTHLgbhFq
DCJ1/13Or8mCJecKDXcVnh1jt3DCcxeHA56CUeP3rUaZywpop00iFDeiKteZi25pbLnM9+T7rWAz
HvfRmyAdEK4fj9ZG0oW/DEfnBCmhPrt03FcJVBuOKk0iDTpeGA5NMyM2Mcjs6kXFvHxi6FaHDeAB
Rc6sEVYQKQTHfhsUxfnJceXGNkTY2NuUMxf+zctui/3iRq/SHgySkAAwuYR1wQtkWBnNAxRenJqD
wAZKrK75+pqAvtebgOEgy9giPfeBB+UZFd1zMcQrlMxf3M5DYMGbX9V+shm4GFRPeEaD7Rj54icC
WM8GqMfxM5iXaOSoz2vI+zLYWw4/K0aklc4h5EVYR8Qrz1k3GG1F+/sjDdITdAcMFJV28lYBxQbX
KipBB5cE42s5OZ5SykFn6mW8ziBeRmqMOew6XfLub9MNi+EVdCbDpeKUa27k752Gyc/ljkTMdGcI
8Th69pSYQOYqUKVMREjhkFrGQF8hVPz5SB9GJlPHCSABrXJLSs067LE3+Tw4UrWK5rU8s9CIAavn
HjDY2Yf3cUhFhKCjGKwYhVJWcaUFPAZ0MlN3Hdbyo4izkSMq/mIF+7voXE7kyaAoolHCe1y1DFHA
CBgXV8L6YfPYVvuLp3u5OWNW8WvaSPcbaOEDNf/Nl1wHWBoUuJlDwPYvN0JnYxbuzmcJ333yxvFx
CzXsYEpiH6reygEZJAUpF/Af5+1j/WJGk4dND2GoCM6Nzx4UtNQ2T+36D3rBv2jfZ3H+nS99jkkD
phm38AIxM2UC7hQLX6oCnb3m43IJutSZ31rT+TM3dRwXQlhVUBrj5/lSHdBPVWKok5NPyPnQ5UBA
SNhs94+uOiFGMWL59ru/K8GCxReHGXjLOaEk2w5lj7XAO7vvDgap0OhJPWcPshvdoAH2rY8RHshp
lndj/T0qgEGZIO0vepYyrXnAh/sUu0KSKl2BPruQLhDIrKkxoe2lMAtfFgxrwaDT5dsjsPMlVIrK
F8YPsL1KZhTMWXI52H5l7Kg7NKtWfIsUQHb8bfr77bxV619OlX+L3haXk+l3sqzZ0Irmsh4nFWXu
bxMG3xXnw6ZebExFvY5bSwBZZIO43b5+5FkBf+HZt8amXZZhWXmx4jgBjnuWKLfuKyQRKmI4fnC2
6jLlbN0sV5ei2t01qBdhcGn6iBEcgRoRduVVbpbv5sndoJfgO3D0IvKduP4EfNsXBTj2AuIRbk6N
hqI6E6VNanawKZtkvg/q0vI8bl5rgrBqjZWnT80hNHy09xkCVKtnAxdcu29f58mlYiJ7b28sjaTO
kVsP297PjHwbPZP1ZC+lKA/Xaz2zJUFzz9/BHGdBqT0bm2g2qbnoSTUGSTN0QdlB2q2bccKrMZ0N
ZlU0COGSUov/Qkh/7gWSj120EpDoPQww4oIYZRsSWV3cWTAXhIfvnFHTIuiHQpTd/QchyOxdliYy
h75dJPTb5i/kPcADqnGAZ/5h75szrSl6zJUCfkus8vR5JevUioFsZc2GuPhceWxjIRQKxVrF4IsR
U9J9Du2/Um+IEX8YsCvvZp/YNXO65BkXqJvzMvmtYJHa4ggFtNMSOgCNrhAUQm12Okl5XbA3m1Go
1N636JLzbsPF/JaGx1q/WmDtqdW6sULmg352p6xubPNO7/ggOdZArd26c2gbPzBOlBu/nyJDZhnn
z6VGAKn+JUf1X60P7Jdq8n1AL0gc6txfwz8lQvRzBX9mH3Eg5E8SKBnAj8Wt8zwxLY92OjYxsfI4
7IDIy8IoDKBgV5NuYKX5dbsPDkaKzXfGxCOJgip2UMkZhnH3rOP2Xc6TYtEp37kBk734SsSht1kB
86kXUl3zDV38uZe1VvCCw54ievt+H7diSVznepnh6jEcjkii1OFSeJBsSwcd7AifU+ZA/lORlpeG
v2owH4vuUuz1A5HdO8gBkw8XMYSefsG1L/LopDO2nZcKauOwGMrd6qJT5w/ikwPHutulRkpugIl6
HavDj4+YRGwpcuxdFdEOQ1H1JTJx6A3U0RcpJ9aebCwQYtyKJfmb/EIQim4QKkXN4svuT/h+N2Nr
wHd04tn0wQPVlAmHR1vmUC5if6VvuAMSRpNm1uRovpbL/wkx6m+X/i4KhScELXsD9EPZP9M8Rjnb
151Gr8luoCOtd7NIa2jmX8pSWCqBSJQUzM/4/hDoxrd+M/FO1rNAgojbZcvFo0RCCUkDpY3b1pVI
F5k90rER3Gvj7xPquj37h90czWheYj1qdi9XsY6d9qZv183euJQh2PopIaMrn9I+0pxfsvmFlxJt
QQq8057ksgp3lytCnRS0G9nebWUX4316jlCakbdhL6fxjulD1jLjc/7uCheMCg7twcvJkl1JyxKP
dwKeLSS3YQNaGRF+jMhHXeUysLPwMpNMch5g1R6hHG3LthCBJZSgxxHbf+zMgzJN2X4V8zUDopc0
ip5wZA+NfKO2Xrm1L+Q07mUWwZBqao8h/MZ+kx46qSvXmSud5MTPcL6AZwVt0ZBEdKfz6IdEO5Rf
YpYNqTeBobHtaYC+eHaNRLbKXZqAg5E7fuxG9n27OjqFUrMYe388kc6kG+13+0OqYru08IG5aVzs
MPdy0iDy1tnjz6Cgv+sL9IVaDMNIY6V8fnkHa5mOmc1h3hay6svvXTZGUmy0jBzT66uQ6W8Nfrty
Ekw6c2EdlTLDqVHtcBMg/7p05ZmqAPW7YE1s917WYLKMHRt2B6qwMWNb9naP1QZ0oMQvUtxXMmyR
5TamQrwpO+snGr4rQC6VkMEp2KxXWyUVLwyKlOJCJ4Ayxwe8bovW3KXHdOdppr4ew+AgUjdBsW9Q
bjHPjIihcSz+IVthXjFdz3VIBJYNt9b3GZWqM4FtAtzUKP+kXLnuPaA1R9eKDSzFVTViCv5t6B3h
mYz4B+ALOZ+Y+GKUd5p3Ich2m+nRsp/TEUbeA3Qj/oMX2gQw3bYM1FjUTyqngQuOSmcEI8p/AUQM
tGh2d42FzCpoTBjSrobDkkfFfYTKxP8qXEpXKnQn8EY2cnpj1tjSogbMIxVAM59pNg4fofhefh7e
XQqfACZZHJUHk3Ooo+YO+3gdx6xdhjG4Ko6GqMqiR1x1HsIil+q7PWyxHzgD9CRagkkvsnRRUkOt
E0Rmefdl66LK99dYwLpE8/HRcqFRaXmxxt22V8OMuhRbxk5FjeQgI+4My3nJVXx6A7trjXbt1CMx
h8ISnTm5XQ0R+z4OZiCWYK3TNYMq0WiRt+01H5YHny8I+S3I+vml+nIA61N3g6ESo10jMxD75F1l
IUbL11HsAxwtQ4LP9cFFIVMj3yCO+XpOOhWGK4n6+T/Dh3brfFZiz9lcuAv0BFMs6nzvyBleydOk
9AtQLOnYnQ1mlykqGvnkPL9qBZ8m1t8FccmpkQtRcxc6l8kGdRoTor2XwjNSrqQwLriuZNADk3gO
q4lS9yQFvKcwq4hvMFutQgas5E/wrZuB4C1toaR1CJwCzKcIXsFKP2ZEK5J+Q3m6rchBt8p0AnZP
cHMefch/tpO/09qmUb/icr9amXDkv9wbg0RnWM7B8LBblMFUOP16sNwUXX9ageGA6obmmd9y2DEb
n9dOV0d2uAjcwEeb64HghfXpDxMPu1IRCuuHevlHS/7u3dINpFzFv0NSYu1MMQaCuQH78sLZJ0RM
zDOu/ELKdzdxgjdVwMn/pdoalB5fSqZhpnpIi9IlLVTojEBuJ7bN/r1Hp6vFwEGUYOA3ERPnVHMf
d8ExuLAWirnYBc/a46ksrI4u2DlCU5A2M4GkyFbKaYh/cnLu1mnPazDY+BwycdBlcfcSFloRgn4J
PGi6LL4kDPDdswj3SwAvwS7iS1iivQvOXtRRZ6cpd9fwpcftwpJ4zxPawVXjdbpazD2s07PEcaIc
vAxbyVmX/AqGqIYn5JYuAnMeD67XqQe8ikde8cHERExVUC5aXAThgPO7PzzqC/av44VjQfhee/+7
+u/Cljidrlu1BtXWtvbY5zyv+WM9mJCY4dzzqCEWw5KNjtfDjtXlH9HeIlfKcNlqjBWaUKTjxmDK
KXxszY7HvcJRQUd/WPhuuTW+8Rr8ZWzhMu+p06eu/lvVRPgytx8X6Sd4RSmDyVUEAYwTZQIzCoGk
GYSMGzZIN5dwmc/uNMRXNXnBkpiNG0I7CreJXTCeCyoklGgndrtc0tVxwG/E/xwpXzXpGja68stL
D+PFPMF2tj9zu7VHBPn19KTAmhyLoQbTj/UlYTqxHdXzs1RC4UoTU37RrMLBHrNuLUn9IZ3DVV3G
SPvHF829FmOVbuE/5orRxSnm/jyz/KmC6rLu2q5EvEePFoV5tbWqZZxZZiBEyAfpSutsKn6EZtJm
e2XwMi1l9gIEql3YZ+e7k4L7mF8z+WJgnF3xK9l0FJgQJJFiGHXXy2NWDP41zK0bMfOItJL4TTS5
WSwb1WeSbbSZcxdaDsQRsyGab0yA4uHUP8LRhOG2R80A0ytznlP31YXG07IuDTPSBZqTrKJ4iJsO
187p1i3lfaNxlWodkKabA0OEtT1nSWyAYkpzU8YR4AvXVMW81Hygi5L059fZ29F60naKC+EZcLvc
5YHpl2KAu8//iMoM7gt0Z2Bcg4HgrjHJw/MDp4H13CPQlCYbwEr3vAkg8TBc0So7tSzrwyVOgf+i
lrwJavcd7vbQHdPXxIWVnvookE7Xe8EnuRtxAg6VOin5RZSzdSO/2KvE9UYUilmFPeXEQDwb05MP
EEPpdY+KJ59oyaY9cLanCTlEp6NZqlBR+EaxOKKUDKTPMNCEjh+3UFHeS7bWw6qMG+kwcPkcz3X+
8cyT1IuKvYiNWFvfIBvVg8QanXIFCh6z3hxMPLOgaHgIDp++gxy7D2msI016mrk0tRl6vD8tm6hZ
fZR1N3IcyyxNP9ka9hQFia8j5YzPzNCQZHNJkER9tjv8dJcu4gQDtOUPrgG2PZLWePJUVxzW+bSM
WeFdmrwE/kzFVY/JvmpbU/EPBlQaS+twbJe6PWXqdvkGc5pvewTM+EvxccJHgZeETsEBydrnKBq8
kwLIRaatqRl3ATXfyoTJOaCWFOY+tmJQ4VCz0DyVijcOh3hm8cvMPBPcug2xBoheDWlSShqWR3bt
lCjUeLfmtypV0sz6X1I5nqK/tkSZAgP+le9rdaBpYoN3LiF55qdHKq4NHiRzp5+kdfpmyqb0z3Kj
K79H4oxosvwmTBTddUNNpu0uNM2WdMc/YfYnvRVUp1HKWozR0ODktmm6D4TE8STJj6S4qg3VHqnV
Yf70OmCMgalE0dUHN5hVk2JPt/rPnLLn3cVcrxoDp8eATiBdA5CpkywJOPCzgXVkaENfd2EZm/st
gKFuA9PqKFK2GLGxu1ruuhcTt/e6QrKmr6RrkjnEmjBhzo71RGS8bghnZtjH8NvnQckcPU/gf3/4
Hh11Wh5iS+A7GymZjF1IqRE2KJEuj86AK7P50BF0YdV9qica1ZmYAfE6eA6k8Hi3NoS3OKCqHVBH
wsyKYygH66ZWJGLlSRm29irOidkIGbXsl+OvOMn2qYiBSwy507C7dcaOqFGivLcoZvbxJ9BSYygq
p+30mZiqg9kGBPx+B5Y1j1Fqkqcab+D3Uo3uG6OqtZvXIlFjbbTUuwgBT8RtJ7rU7DWBo4iy0unA
45Qa4R40Fh12OjsygVIGhkCc6FUoQj+0ExdM8PfPXS3qpJ9C3Aux/ZPiJq54mTVwAWfX90fGQ/H6
da6Ryy36aFLjaa8EzC6WPhpiCaa03ual1sTrNGyTJYObPWn1McR4AbTpzz/26aa74meYDalJjaxL
USy5wlgboJJOIHLd3v6Nr61Ds2xULna/eP6hmTJNElrhygsBPlzSic3P3hiic/0M7qOqAFN9jQ6g
yd+aUOYscHhOcv6Axd7EhsY/J+vbEioCbbGepeBgL7YNEQJfCz8JpadotxEtmfFbXaGohFzt+1Xt
ubOIKy5LfIpRCXw31fjgZmwhxxOiq+7uw6Hw7uQolqPkJmhj+qGANCf6QdyJC1swjFhf4wTCLj+Q
xrlE6a4iuIH2WfZrybFE3qVhKFpPsRSdAkyH33Ppmg5my0h8XtdvqeE0GjNDH/tBf7hLsoXkYLkI
5zXNPyBSz0Nwyuy3SA0VONH8YSy8m6iElim//Rdgd2yGC9/arToZpwCXfyhQ4FuPv6dBEzmReBmK
1kIHD8qyh0jiFR211VMewWbLnhBo7HJ6BNcBzfkSbrgTw9HCtuGhCeZC+9EmaHb3xjGPemombOzE
1o3TrmIQNo3YWRc+r0dYHhMYU5J3bgASokZTkh2zhX4nEXkGVGxU7IXOei594yMR/HceOawBzk3Y
XovrFn5oIreBP1+8ayx4i+diS4F/8k/xAjly10VhEmGUgpI63U5BxIN/eL7WPbPnzjTcIAwWsSyi
DXGuglBbT3CJTwlWcimVGRbkfDTlOYjqmLiKreLt3GxMC0XecLiy1plgT1vEvy+LIJ0pWtk3bjia
/+iWne8SlZpGHidvYItXdvHM+Cm6UKeF3G8hEIBbBHyvkbr0oIU55vCeS0c+8lzQBV1w38lIAkXz
1d/jobgiE2ZOeDhfdptsxeyfGd5OhOt6pxAJqjhqLC9Mier3ttflxhXiXyEGYg4CwKHPvhbxLNpB
kPJGXkkIXXz3/NN/WkqMX4X+vdP3f6a3pOuvhVCT5lzzXTaPvmeZijG00uM12H/Ef9qvYKZgK/w1
KXkFqabnYhkRU98qhJAFacfxSOjPqfQkdRzI5bPDHererZ84r2v+geI/FjItWjY2BcowjuEJq3ZP
GueBsWODEDBAxEYmSsua4OUiGdcDGXtJg965A9ImPFX3kJrQO5i5Vi73jGNcDwl1MS6dBc/JQ+xq
MZTXjxhzGgf1aczcG5MqtiqztxJm9RhisqWEcfMh8LuN2adDcZc1/CQxewKtdWhrRjao0wHT4MUy
eRwmv4QxPgUaWc5szGNT7s7CWGPlprjCmUxzZQPVQSiHBRt0eQgqJxTAj5wDzuiMRlQsC/T7WUvD
wVuHx93/k6DOxrEi5KXRdoJPnMiAi/V0EVkRcwJMizP0yM0g3LgLaeyStRBZa41BBBZqUb6z8Kut
c9ylmrVmAsWqlgBB56f8uP7SIC+d+mgcPRgJAiGEsrC2yL5CtsJR8qo/P4sdMmdZmzbmXzwmk1Xc
QvyI+f4Ee41ejYFxOMmX5N5HNEsTPEL34O6o8spBia65KrFdS5rSzscGLvSiB3Ry/HwWQ0/W/LlF
MGphR99ka06218qOeiWtpAKZRy0uPpF62gYD0j3QgtnDZDITK/QBtFgZppf0Pl4H6Zf4GvztzIA4
gl5Lxwgv7Vf4mnqTlwMljN+MV9X4uujI+jCO+dqSwx1wVU2L3cN8T8bqEa4bFYMCO9II3kHmRGO1
WSwdK22FRTzG6T23eH0toZQrcj0fGuPFJLCEEStIoDoO0TQvce0Ujdpclp29s80pPi86eM3pZJIK
oOJT8cxegiWsBrVU3Seq6aUu0xjKGpXYbchAdT8BBLWMuBaBS80HieCLtlfvWCpLeXyWonjjb4gK
cGRt8IUhK/UfLSbOCWZSQsOpcZch/8RZa7ZvzJ9nyGDQHBNa0zDKHaq4ZWm5CVUY0ls08ZPqxLKM
BGj93ucxEjYw0y7wmQtlVMSTXJkcRwv/gjYDgiQs4tJKPKd/ApKjhqXSO22SYHvnWHUHRlPz8bAt
ZarE60NF7eZNMRHry3YqywzEjP4X/+d2EK4pqSf1KrpI7LiBani6PNWSEzp8kgjzPeL0TkcSSF1r
I64vZyERD5KvxjU+IBiw1NiH4qtHiJC48x4E/MEfYdPpqLZX32vbWLUb/xJqc2IlJg8EjdU0uHhe
9O0Sl/C4c613oHSlLWDZDe5lVIWVty75ZkVc8PFPMwbAPO6FjgQQu8Tw7fOQXfnkGY96FH1qsIkT
LKcPtTYGa1rwcMphKNb6OyYsbCyan521Sbr3P0TFlaRA4X2xiw7Hq1YsR6gxW/ljLHZZMRVYXg1p
03ECopFgilrDuNPDe+P1MExQb1uovJ1R0Xi7avjhyAqktZuWblF5SBYKsxBwT0folcKdAJ8Gtvho
mb0Tx4VpxySjWSH1tEFRooDwJkep7IZdLB5FkRpX/fBWaFaMHHCLElrujmW1qhTCfXRJ0EqQL8Gq
b1Ww8qpDkicHy9Jgjz2f17igvhwI+bqamCT7AgBZ9iC1jcHpJ3BRnvrDbZebcFgN4jLdg2N6Y20P
TKpGzwk7TUHo6uDJBnz8EciCTpMa5Up0z/qK+W8H/iNxPsvE4EKdDr5xhsVm45d6l2YibMx2qgk9
+XZvwyVTcwifITPkxLKpubhQjHofCs82N1Ogtd7pm5EVGsoUVwafMimHGQw3EgnAxyvv5tc3VQM9
mOZSQbBa0D5GNVwykxFEHw9T4UT37GzQu/bwxx86txRFyZKr+2ZA055XMZADIdY7/cXc7hQWm98F
zyNJrDCG0ftHHBOcjkN9V5PBRcD4eWF57yLMKIaCHhMECx0xaUeM2LloB/7nwcm+LXHPCxwo9Axr
BECBDm6rh9EN3azkNrtxlj0QuFuA4oSBvFmPTlWI0hOjj2LK+miT4jaBnwaUgRXVVzWmsG+XqSfS
9MhuQfa3HZbiX35NI7LfuSGU6s8Y5xE9RFyRwA2n8k4pArhact/NUmWxJVGMDnRVhqrMmBzV5ao6
IQrUNaL36SK1hMq+ztmA4Ksw0zUZT/2/BJ8sVpiNBUCGUxrmxbWXdKBayEyyBSlxjq5Es1rb8d9S
MscDoy6+PGDGy9XjVLQv0G6LuOnmtuB5ihahqF1zG+0hRICoRtjqItNJB0azEjZ5+RZM9bX3cZwu
9J96hxp40Q2plx47r1zyKVDpr9mKjHH+vdHpr6uINChaOE9M9B/6vrv5jmwutV0fadkQROaWPrH2
sKpLH2HvcPqI0UrVFVm45bdgHaSBo6lkQZxG4r3fiponGWAqS1WHsXPwc2Rt5OOl1ns5ke1vAxoD
U0Z8yYj4C/9pAxoRF2T919Sw2bscvNOZUf1tLufgBhlQNf+9NxGOcdQumxaLvjDsGteASz/vewr+
A97rG6WDOR4m+xBFxLzqN49qgNG6e62Gu1nGIvB1iDhGtkTfk+tHiWTULcmp1P2yjF6LT3UUgSzh
PIJAnBHWkedmc7+xThQmHHAmO77rCD17SrHFEqmNbm9rnQ8aG0roiabrw31cZQD7LQB4AxIG8gDc
hnthUX1wwYdljpmaewx3VcqiWjA+NBgxSulDa5b7FA5paab307rz034RG48pirN5lrcbIZ7OfaZm
AJosJkGbrUZTNpnHKy17WgMFP9eQ7hj5D7c2oiUYgok0UASMeeeJ8Zj0w5/smAxKFQIUR33FSx7T
5dK4goOxqXHVEcuPcQZTalXynjSRtXjQ0P6q5DMbKzKILYJE9g2zJw8+iCq+pVSx/9y5YWDTjttt
tjEkQj3SDGxeaDZzFGhISvh89KtkmCTy2MkW+3lmh1uTZNxOgdsV/1BYO51y2YWaJdYp4+V7j5VC
FoKhzRO10fShh104YjlqujS9VKr28liNZF+qvLYrcxoCprnKq70joqymFaCcVygh8ZEHMkkUPDg7
rCHDWHw5jbNv43H7eAQvFGxUJsfMcUUj9a6fNm8NPaQxTS+qF4sibAeTfE6cmGxVEd4R4OSAeQOC
abozyYEU/HfgC70g7KvdCrOWwgLputqVD8X4DkmFFOiFaXZP1NVT2B4nJuINVLrSGXiqCv8R20wZ
Nj76dI6sylvekvbsY1TI+LXutkaYlyL8n79KLbQaDqG5iC/fzngQYXhKtubWCulhGxeKglkkU2hN
+/+aFOHtfHuWZzx7XXFnW2Y+GySeBa+qgIFNGoagEKDxCuOUn7CHv03Q2w8dhxm1M9GvsR8shC6o
F5soPk0tTo1jTtJUBds4CpC3FacXCdJGfbOtFCuVwNhWUVw8R5van1hyJ92FKSUqaVOY2ah7T0Xx
8IFd45Y95i7qlv77OMfS8HzwlP2ZpVdPOApqHK1GIfUIvmWn+S0ZZCpIcSirNVBwtIldvHV6CgO6
uPwxLTMOuL7oc4mBo9cDDykUZrvUCu25hxxaOv7NoAtUzScc69pLO1kWK/BHV36NoiGw9G8TUymQ
+E+KhqnLz/KgEPz5X4pLnUUsCae6E0rHSd+tJ+lQDzyF1UGIenZjvLI3JP440icUKnPsQN6Og4QI
yoh/eh2qHTdYtw33y+taJWFMRATBzCB2+YBHVjZUtPFtf3RJCZs0R0dGb+TVezYr+N2czX2Ad1mO
MBm+zWxgrHq9fIsFfA9XCaq5pp7Whqn6FfaPuMenhDnZfq1lxLcQcl3sfQxaUF3MYA+ENyW4PZir
tCr3ZUtBHvePVSfbgl9VFLWwU8C1lk+9vK60yTXHzriPSCJSSP+2XnfU/MV8srxykOY3ppQ6gU3u
tFUDuV4qxkbJt7rnZokU+eEm/oiUTFHpQoJayrDY0DxouiPkf6JH8POFvrGNnpAf4YVWEmbA9Erv
0EqcVspWLdbxvT2ru3Y8a/SlKu2HpXEqJ15iv1rVrDDfnY4sKcEUS6rp7UGWDt2QpTFWsoHLDicJ
iG7nAOYkbMEOBWF+W8GIng/oO3SnyOohbW9EJcBO/YdDIE01M+F5UX147u0erlnW9Qs5g9DvzoNy
++jZ5zgJweQR/rsQpwTZvkgTVh5qMGUwjk17BuunlI5LLwmKbhHs1phdLtdaGFBXDj4wDlyDwmYP
e5L37ModSGh8vLlJc2mc2ebbg7uNB/WwPxztuU2vLmduBSrkMzR3b5SZ6dxZnHTjxQSK3LTra3xS
okOiMb/Xb397ngUUMr6fTnZMgfDK2krH5dq4iLfKbfOBbvyF4yEjpYwJAl4GC1uThahwFGZZ54wC
PDrGM/Ow62XpgUV6l9KiIxe6+Sl0q3cnYsNjo4XIDvrJixdG05h/KNIw38pF68NI+rrZyaV2TV/z
QpQLg+CC+qoeYCUkbRpfLm6WKg+ISbuktmvRgvWbqIzy42lnETNGns1uI5aQ1O8f+0LPWJBu/cC7
WOCW6eQk8eIB2jOqHR/eGy6JHUzAz4hMFSEfYqwCIGT/EblO43NPVgEnS/CtZI8Pas9M9PbLoReq
w86/GN9A8Q6iPSCfO60ijjXqselsuDTwFly/CXDV1lyD6101tp7oa45cOpecbzFDClET08B1PJv6
zvnHnKDlcKzAzuUJVDIFhVH2058JQ1FvYnG8E9j3OZYMrxX0AL9Kb7PPvjPHTfpRhROkrq5wTLpQ
vXKjhU5W050fPUv5LgYDJLrsSBDH0rdRFvzIRAkLdWN0n1tbsvHvIVWKCtfykA2nujsXrHPhNxwJ
tQzAmqVoJ70/aWnOwpPWBmMqjn+kQpCb3A6xXJbVcV+dZ5/dPXtHSmTyYRiiFpg9yoGthkou2nRH
P0pUVHMJx07jv/DOULPbM/9ypzpOOoFQ3tbyCK1EUI0n9yzJcTbU2PiCzQrxF+1CfeTFIwVTIjll
N6FtjPIaPCZZ54kRhp1UxE/BkYoWnprl87uzztSZUty/Y/QGxbQJcxwkthq8XQ9K4C+rtPdRRdJ8
AT1hl80OYxrZUKx2I2jx+CBC0YRrZl34iTKEHNpDTVXc3VCUBRyqlBuJHzYIwwLxsXOJQS/fYVsC
728fOHhitr4Lq3Tvvka/CVk6kMoeE+aAGQbD9HlL9FxzYGRaXkCjwSNvLeQR0rA4h/is1tassmKZ
70QZ+vk4aBVwSlHOJgNCmcBKobq2JnM8H18RcicD+GoHltOjMN4HzbeUODrPbC1ACo1zGPyImqNl
UdB/ul4SScV3Y7O+n3dBKnxNCIAjYInGtn3MM3/lnDIl6EAhRoNxhCESL3QMFlPMdQROy1/YN9ka
ZQSC9NXEzYEBH5sd9u/eVUaMbpl7pIymfPkMhqiQfOqQ3rLpQ4yC/u6j/cdAjY0CroeMOWiGqdtV
OanYV0u7H9cosFvHxHLHFj2afVnZDDpcr/SfNWUUrPM29lAJNHyK4/rARg3xAHNWaTqVq8oBu2c8
IT+c2ry9aqrbUYHee1C1awuFD50VQjdC6+4YuWJWH4alVZow0d+Sj7WCc6xbMaaIKv7ZQUKJLTWQ
ikrSYyqw2fj5kruJQA3UB0w7TrDlcBSoRWCGDsscvoJ3QFRXzgcaq9K4LhLoxYcysF9Pw/sBMiO2
uHkDXtU8rkxosGHSY7La0C6h+vfScqyfzllfS2J/nOflnsUk5Ja5HuRsNYKTvlwOtbVyDCR5S/4n
UAoz+5a6kJELvdAzpWTD1YxfZCuXJZkgCyVhQi+71FPfNYL0ijDxhAo1LxSrrv70ezfPYbPnqBXl
/eQ/ce6+dvdYWJdeiV/xMwukdGn2SI0d77YtQEFCbjHeTzbyihp0n7d1cZW+cSeNcOFi9M7+rDaL
58LLRd0kv1eEiwZfFQETDQ5wg5/BUBefb93AqMTUtD2tellEMKp+dChbVzozqBq7he1YGfBq9Fsa
HAan4JM48onTAEQnVObJQjZ5/vIz+5t882AxlxVK1ogyulyV0XixuEmy/WqvKrkQH8kffvfAqjxh
3bwivFK2IxipE+VWWBFaDgIHzbOd7XvR72zwIEFqZ3+NcTfbdn50owWdPFq0CpCxtKSyrF2dJm+Z
t7u+RUBFQpaFy/O0u7BghMWhoUsys51MfyhdO0iZ8lYiDkRnj5xMYK4dnJ3OnG8sL3ZfvQykjsUf
CO6JvchmTEEtOYljyjy7B3SlAGCQXoWap17mUk9WFTW7HK/Z125VIf+cT72NZNEGcNdGbFDZba+Z
eRPhMm3z7johnjyKp7zcjTJ8KvChzSmbkaMFoKdA1Qk72CDgYu08in5OE6v6Cci+2Ea9+n0iIJla
AuOlVqJbxti9TEWNW4DOPUA+k/AVWLnw0mBvUhEWvQZv28Eo4Xjy4mKebjXJ/VEwYexuJp5UE6+u
QgJYGpPV0s/9ZbrZduiV62KsBHbajcfuPFmNY4SI+Vs47l4ij2+0L0Md9j9095OGqKEY7WRAS6Ch
CSfu1h6RwLyGXR0byOLGmfyzoJWJxmfRoA4rGSRvkOMgOwwTwjJblUUKOlMFnCZ2jA89mke3gHaC
TXq7jsVTqbG4Pk4Vd5Y6UTieTSdvzGZiUsksDxDWcW/TxHGIgwS1m73kwe8cMqRz9ECRsUzNUA7N
zn5p3A/sx/Ds7FHhNoQ7TTW8sgUFuSYRAFKL9mb/PXr93g8gGOknxrjjvCTIaOMCUnsHFS6rnHlS
jFgV6rPAOPLXYwfpE4UcyhOM6WMnhjO3jsQWyJksi0ZP1RZDVHEX2Iz4njuS0+I6T37ii91y5k/V
Bop1EsdqUG/X8rZf4qfEOujlLqGip7HVapJR9FdZKL81FodnDjRhSqVJSPeBnp1gwNNK94FZAtub
rfJj/LV0L52osPUNNPvIcP3G0H5Ee6mqw9769x+zxn6wO93PrrYtWYvxKYskcc0IEU0NCef4Ek+8
4mD55Oy9h+h0cDaEmvao7jls1/cB2NVaZ4WH2wzM7cZuOUVQERuwOli7y/yGF5jlBRXiCK9N3eTZ
GnORjASvN9d0pGNglz65QipvV0+GD2/HqcxzU7g0HyflTYYyQlzf/jjIAzg1ZiQaGa4eDDMYj6BH
LJIqoFIcHkSKLh/GMKZ4/GmwnCppEBNkCU8LqxHS3SFmpdSaynphjI1M5QB5oDyRh7TSEPZl4Y+Z
wnMexet/zUviLNMuA69+KrArWsPv1IKz4qGnR27oR6lG7yUVmwW8cWUjaAP0jBGZLA7zDDnE97ei
hJvUlikoTCSMgPttpElB4cekAHE5p7Vv8B/yY4zRgQ9SyQjM6w8GAQXRq+8G7W5Z6WFA8FgtZmVs
gS0ghgfaYpqy3yKKY0Lp01BUaYGxqNO0/qKvN1MYhqXwO5YaHpNOzOAFJW3aT05sp8L8lDMhUG4d
XlU8dEGEbwQoHf1a1SOX9SyJoIhWcnvtMDsxas/6VLXvKTH8v65MB/AIlehrRuCaUGch+C+LDQM9
iKy2KC1M8ii/LeY9TiPUdpd0srmF99Q1PwjrK6afwAr7lz4Or8iNsf/7MAOTRgx48Ht7Nx9RDlRy
sBhk/2OM3CNTSOFpsbFXLZy713yJXww/S2LsdlsUQLAgXR66u0WFzCZcMkjOiLVXEFvoEvrS6P6Y
mSyljVynOCS33O57msqhoRKjGyMJcNB+Wnc4hroHrZJmldI8UO7z/NZNFdSHUElHMuQANqx5wxO4
UgkdZnHdoEgltcCtcGkPnYfdn506lDrnCMGqmF3J57qoeRBrN6GBmY2odamQj6IVH8ZwfoTIeeCF
JSXGuhQ8pCa551D5kZoZ0epMlSxg58A6drhF/iT3AxW69ng7aVIalaEqtcqBTpLQf19xSEkmc+IG
YCGNnE3t82ldiIuM/1x3MB+ObEhhGbrTUoGo0ssMZ5jXt92ohQMdDBON32FL6Sj075wiI5tXtiyb
U++Kq4zXPkMZTBS/0DA993M4blf0LI7IQP3LmdG/BqfZIWv+YUqPWj9tIDyFwye5g7UPi5sCGWP6
Lrf8ZOp16OVPvKsIkpISlKZIUjao4sHIiZxtW2HPwuLqQK8N+GDdIgrUMMWhquyVa2w7DirKCEEz
64kJbFUH2nvsGzC/psKyVt6P4QbkrXyLN/su8KUpS0ERHaK96dVXvEvU8Sv3aXJZZiGmCDuDXHAA
5lBrGYnemGyU5jo5GQHQdGcEUQikn4Wx1sPrmPQ2VE8ZYvNgv7ZIiFuvPgMY1Utmk9wEGjznHL3a
0FwpHVADRQL9l+4hm1Vs0dqU9CWbK+SJfs9FM7Ml/r+Bj1KY2Gpq9XuELsCFu8Ac+aAwWTWp4Ml9
IWMhbQj/I8oG2Vpm4Q44wBVG8U3lo0w4B2eT8j1isSYNVPYaSJm5Hml8dIg28KrIVSMQVeLCbVKM
nTYBk5X7NwkmZhRnWkkg7k7irt5IIrF7QgGOZ1XnFYJwGCAeHcgPCO56x5HAcHHTgvxkURyv3iXS
3uxgovA8X+Qr4mGc38RnF9B+TAiHWcH4XxnchBoBF3ILKtAhmUbehQlLaspy0Q3TlDJxeXzDRABF
i/yS1QT9NtdLSRdQ8+ugs6BYCwLYEVIzFRHAXJvvBYlryBwFPri8ONBZZ7J88hyDOlFH1mYMRri/
XXFl2RNNH0bG+Vtsj+LXEp/HjYSCcK+NnSMR1g2jbyE2BtZpNxeTmyMoszwoGHHhNl1crFXkZTk8
wdAh7Rzr/EfU1/lS5T+e023Vgc8PR7uhaFG1/KdR26XAhL8yydMUf0kv0u6deH2aQJhOw/7ZL9XE
8WI+Uo4Em6ImwBcyIMcdnsHxVeG3R6Rp1/ME2N9HE7oYMyIE+FQSIQP4u8LMWfJzRPzRTb3/KMic
zSxQnlcyYrvy15FfsifxnEumSXV19DzoAuzByCkX61pNVQFCCRNfGlZjVFA6hNtgnJl7L+50wpoE
BJcFDPW9uGKoFV/kwP5a7KWjWai/YnN23kLdmFFm2rn3x5YFueASZyhg7g1laFdy9VmdqDC3qnpp
p84R4JlDbnctbJmmmC/IajgB9yXbfYE1RtMwE5kqinTQfyJirreDLVaDkRT6atrfrTdwn7IjTHRU
TzSA8AW8X4KjodOhHaGIMOqJPSTzSF/mOtSeAuRgoTlnae0kj2HbXuEmjnIq+PBCxMC2m/cCjaMc
dEAfrRlHEKAuFHwEBRoRGBUCSjo6jm/y6YIb3GTBnlpEqWvwtH4OQbRYuq94/+KuUBrjuW2eEBTA
0//oy5jSKbPQjsoGyYMPKmUfldg514cJS4py38/ue0ssbsTw1wzRCFsyq+GUxOfeRo3vzfQzAjBk
7bDUsDX7I99j1w24kf7ziMwkBmBrDlA66zr4k/B/nHRWrUGm3qMNrilRqt07s9Tl7h7A48AgdfQN
IisiFV6TLxGupvoyMh855vbqcANCs5oqkeUtRkWbQ1ns0iehl4Hd+cxvarJIksmEi/p1/+h4nvsc
DoM7VANGJwx7y8k0sW+uzoE+plUsZ3K8No+qHDotChd5I3dbwk7er0QZ/qM7SelNPYJ3UyP29cTl
InZdksZfXBXkXNi6KZik7fzi3cnfgGaMDtn+FyPx/muaeE9y/YqaobNirIB7+DDG7Q/Bfj0BvqFS
R4PhrvTuEbMmdMqCLv32c1U4C60DCSmaIx7SAV1xa+u5HUQrlCGHj2RpLW/Mj8XRwfhgJcG1plWt
xlGQXmrTfNv3b4lvkSSQgheYwPZ/c/xXMpklDWe240LKDAqlStU8p+skjO+Smmv4HHIbjYif2u39
EBoDKVFFDGz4vsw/n7GSwF//lWXWXwcnBmZ6TL8TbJGDdSaKefIxRuX9wE0ZDUEng5ReJQDQgUI/
1iAcQbwVZQRCYRUU8bn47gVOZnKJTGlbBk/KWjzYb/dqyBe23IPEoEflI6u/czMAf/cHYN7JQ8Ak
8lQkn+RAk5DuJtms2AIAGJSEDPMeYsL508pqIk5Po35Usb+uSyVgBLragbn/Fm/cPvuHg09pR8qE
OC2QGjM1UkZ1N0af+O3SfFnm0EVUIgL2jrhAOyJV29eL0xdycAvwub+UIKXMeIMvkwAqJIpGQrOu
hsBgpEi2xqMJHqjqRoeCb9s2jwMCD/RIswcpnNYOr9EBBqzsJY5yiG+4PGOUMyZQ8LI4EN7B/P+U
C3OBy++fD/GlGcVVbWnlA77C6UEups+LqryZ73Hy2XXyrb+t6Kz1RvqaAUCfGvlRX0XEMrC+CiYe
VrzSoCO2DQKr6HDuqdctPBxGTg52wLOjf7zwpPoru+1kpLRy7t7j3fCRL9kXBp1e/1gt6bVTCZim
XsZmne5vdzujoWbw4HrZHav5RYtUjLPHWFst7WQmjL8YbroFGqJ5elrYmFPkW5cHV42j7IdKYZBy
hB0YjLF0w1t8/RM3eYuLfR8u3CWk+KKUUbuAI0yU4X0eUCJtYPST81GoBYnTsxPC6+MixyIiSsyK
Zw3ECbgnjhRTc57GKIU2i0xdr7/sRrE0WjfAN3nleTxvbdWAhIg/EkPvFyuH0jcA8CGl7daQYqlh
k3Lrsi/DCkss1kkBf4KDMdlIFaXlne7vJQKb6oplqytm80xBHGveK3kO7C6a/qJaf0uzSIQ1is+H
k1bi9KAlu780hy2fKLQl1fxDI8dj9B2yoYLySeQBZT+KTANRrutRcuxtlqgjDmO+cuw2XRB0DcCh
M7bsZUH/HeS7XCPFilnPy0NiwVKbhljJFSubzXnGtFc6weFpMiF7JSniwImYb0K9OUZfLCxxzfAC
4P0+W73Swz9+00bpDtMP8GR1Hy/vvPbTYcQATvUEsZnW/NicodkA7ITDYlTShSSpqnWBdI7bjV9E
9bxWFdtBaG8Nn1gPqtZ3VeNnwmdm5LwSXwOYkFd4vjA9JpbLMKsZnEh+TCa4Rmbd8TsjT3IsTbKF
7kFw3HAZk9A/fqzjeM6Ql+/wYgyOT1toaIZBI02QDaPbsxJSFSrqco2epX/kpDz4cqzdiePMSrsV
lbEmGNS0gfeKZ2E0KjK8ockwiNDCBR7kGtZ7ZSOdCOmi1I4LN/NFt62iXaK+UXVon+Ygwk5XwSgl
RJyKtFZev+jKiC5Pb1ve7xrem9/j1wXSO9M5MQd9r803KFZ4vkHcrUCmzMJFjrwfmyJrlSkO6iKf
kjr+59uokwh1C5kTJWEjtSYFxBmbFIdFhc3SDvmcD1BrTaF620DIIZt1PfVUyD9GL40VDhqDh98o
W1J6Yg3oxme9VVI0+x97Hb2Q01knyPdY7fII46ZRgntGJOMcCJaAuBLDvf4T802KH5QvA2n8Yku0
JRs7a+1731MeNpui8mRFvu9iRhuwElc63Zk5va7AHk8HhTTC4GfygAse5afeasnlKUAz3TkAAH3N
gJOzRLfCb+3V/DGkYu2bqbRmELv8otYy9cYmOG+6bfnI4h1NYxlQ4e5qVUC5h3oucG84J9DKQ9Hf
wMQllZFa9Jgf7wSfVtZKQFgjcu3UXAObs49UaJb5FuA+TlY47MOcwkNlrYmaoitK2e9UNUoZya5D
caJ4dGZjYq+Rq0DFpizr8RU2fQT8qeRwIpISnfRr6ba/bRfgJT47MzN47s5KHvDablPaLo2/Ooag
Y33LHgombuzexRcp4vrM2NHlkS8LqMJJizxQ3PdoQ7UxRkmGoErEleBWqNS9V+4U9k3v5DdA43Fk
YvI7M8RdpSXdVl9fuM9e66XD2rVvMCj2felsLYz4qNQiSnHaTy8rG77jMpJXuyBRjaC7jwpiBG0C
mVJDOwKbU55otrWicjoKafOL9HmUMMHshQhXotk6izh/xfUDNiQveIYJtdB7ZUOV/kxcXK3aPdQW
U6d03j2Zm7GNYIi8WXkLIrPRrNg8F7iASZF7eIxhWQl4kvULa147yDuE8XOQDParszzdBzBVY2yF
4lljjdQuyo1l01XED0s89dtuWm3PP0BMdQjb6fQDc049cQFGg1Y58t6FsQOZpMC6Po5V58Y0TRbO
dPlctFt9wRkOTImcIxbIuZ/yBCfbvk0e4im6lDclA6qLehZSHMvrvbKHKIocm+pdQINzH9uGZWX8
ynXqF1ahieZauR+Lo2OwhbPIA1bwn/0HAl3pPGB/lHp41L1KJAridVPjfDdj6hf+ZZTLC6GPB1hf
OeuG8cGN0CRKYcpSTjPTaOo00flXc2g58qcLIEFv6klzgY7/clwB8ElaYgk8KYG5yy71/putjS0b
ST9FeCA9QtZHwOBQTfjUVbYMdhuP/RSUDMhc7I5dRMwE1Uo6dThpwy+NtQKKbNamHgT+vYKC3ERi
Kq/5Fmf1frKFt9ZnP4pCoxVaWgPz0Emmf9u0Gqmut91a6afi316oZZ4Gzvco5K1JfjeFGeUtCUtB
xNznKlMpF6Z1T5sf6fHvBBoy4X20XfkbILqNrZ+8zepEdphlAZYEcHo+EfBjJx2cmedVN48ncuNh
5w5jHFFv8VMhrUHUfTvfxN4jWcYuVIJeTipM066oZA9v3o8pdo+oaR4koBm9qxTJPXDnMRchHxWn
PghAsdKeyUf1SBvDumy86zrtPGok1xncJ0tITfDazxFVef89ap+XnJCS3GDIOLRoA04JWG8QPKGv
0g2UqIx5w9X8Z7SGElLTwRZcZ/NjO3rx0M9y75cn05fiajq20GDOkAumgq8Fl9krrtLUhe5dtKTT
JFI6vKbsZYjwELmFMNzuwgOifg8mXe+QtRq9nq62PtqT9pKJooxt8p/CNfHoHmztlAkxCamHYYGB
4obomSWfzsHLhvErzUMrKDmiKCpStWdDJ/nwlrOHPNkNBVxAUqTOPml1QT9bpAdzIuPVI9UqcJpD
6B5GgQ0ylaKdxGuhhObKUzWeW7bBCoHiu9WhpL6VxZaO8abnd32Hmn9WpkhnLgNoPEImp9a3ECw7
bZMJgYAHIxprca+y0bGc3blWcEeTBmr42ftdvyHxB7KV68WJc0V6PIbnkW0c6kg85V0EVpyWvIaG
oWgjsDIA3YshxOSpnvFqLyndIWKcie0LyWfXEZV0O4+BQCQdFNXbm0XdwyZYpeXJVPkVTisXIJcD
Ca8tD3vfKjyFYaNwuBIhEhxf5yje6sU0iAsO6zOO+KsuNFdvdFMpXJHi1AwJyrR9yd6sNRMajYmV
77EnbB3eYh8jaetLmhdS+7wPuBbfZz9s1YdLHbXZgKiXUJQvN+1vHsCAhGikSI/tKiv43FqCf+4K
ZZ8GZs+f1FlXRs9nHS2rPwz1nOZ7ffu5V4itbAspysHKKMNlNEn3cVJgtBMlK+IlQB8kfayZxdV2
cFwMGcz8JxclqfYQQo4u3t+CH2SpLJvSdE6w4lC9P7qKR2cgwq7Ie1RHEgHcsmsdwh8exWtAdcWs
DptNKpKmZvMe2bKXSb5AGqk3yiu/vjR3gMt5x3Xix2dVjWWdh4JjerTEqoVo+WkLT0rM60Anepoo
BhsVgtnnBLnYIEBBQPFcxupICjRnFkgYXlzPLT66JsC6bQ7UKT/uesg2zWPcmZTyAObf3dhL/iG+
KkldyWnT55je7dcM8U17RxS61TSGBgNyT69+7zPuaqRmpo/d7hhXy0qrCo+H0/CgJktBox64A46r
YmpIR/P1WomWG0dM47LG4R3SgFZgSz8VlKiHYl9rMn7uvg3iDstfvrPVOq6Ri3u0DvXt7bs/7gTe
dXEX6RsVwkRXCNu3nwMRL+NThbGg1eTVZolA503EAqM0VtptoytoGPoQkii0Evci5uBbqQ7EM8gF
9I+JGt8hQcuAnMVB6INaHiONrBuLwap+S4c+58Xk/4SWL59Xa/UivabHbMVPQU7+N6xaUcmRDn0z
p8lK41CgJ3OY0ace7qgKQouC7eeAYCnPA/NASZAdefTxxMChDtl9UMBlD8BI3mUjaqvV1riwQr+v
TpbBYJNpS3zvB9n6kvgDIHLYV2kRH+FfZ0xdsZMmA/pe/kXoFAbr8JkNDggQUElSyTbIzdEI3yhA
tkDf6YxDfDyL/yddb5ylFkbl1DIlUT/4kHZ/442qCFlkNeyw5DBFuyznYw0XAOrgeLCiY15Z2TpJ
cEPJiwUDEkcZxT+AFerSrwyydXUDzLTLBBLBXIou6TiQujR2pBkFikdBfS36CHlIySRBqeZQvQmD
9R+IpoUWbwzy1Qv33/Pq84Jqqs1TR226ktz9KKvlWgngBbNtL958POZquZt0o6SIcDH6lXLKDCx8
TASRdo0RfffzfjxkN+qAQsqECRUkDuoPeg8/2SBNtWbVOF3yzq6oZWYsqezmYUA2AHntQkf3zvnK
5MWA3cpm0nS8lmErMVUFE5epNttFW2VrF4s3ocNy0Bs0MRfan031Zx7K0XwgBZqM6iOwsKXeMBma
ef4xJUjRMna1oQ4icfXJww2eynvUrYQ6UL3ncBlw4+uKnwEKuptUMR4yQU//UQ/+Z/YCBv7Zr0xM
WXDO+/TuuehsFGyr6RsPz12NDMmQf8O+1VC2HEzTchulMrFVcux69QuDCmD/mYedQ3n2iY38lYtx
jT9bSNjhYP9mhKrLqs5kY5lRZpxICCCP02VJajHebtWFKTythRrwXDyNDqi3nQuEZinwCcEr++Z/
SgTOCPFnbskvx2UNKe2CoFRvZz/ru75V0kXhrQTZCw1tSo6hCgImamwN4WU7hOW72PTJZ6cWAHdm
wnigMODypU9lQDqkD7J7yLEgyEwq64I6+M7qODagXaSFiw5sEQa2TdNSMW4EVgL31EjvOEcy/8hD
WGft5mrwhQVOWEALebK2FCfnPmy27D5Dsh6OLZz1EjZfju4cc1tzyVTvhxEI+Ay/wl703p8WHP2O
MKHKT4848dEISknkUivZTT/bN6H4qL++hGlQSYbT49zj+EfZ4I7SIzb95RTrc0yRDZ9NQ1oE5zR2
r9746+sV/1BSV7ONbD7k2gDsWjQii6UdubVBuFW4M6UiBfHo/Dn1lz9Rmmd3kELh+wKH4MuB+ISv
ApSP0661b9Mk2Xm5oxQMP6Am5a2uaDaj4C6kb1Ky6leESKINAr3Z3mTQHZbw1C8LiQSVGi/KCk9t
Sq7CNRahSDCYX43EueG5/7XBsKg0nuKwzOV5O4IAtPBG2i1fL75aTOR7fhbqFOngtElA6AE0zKtL
OjesTJI9UhDTL49TKWj6bdpe3U2V/F+V/ay7XsDMooyZ3eY8jxIkDO47I5dVyBNLb0kZtbj28RGa
C/jsSwY3kJO3d4AcbSQzNzXi7CD8wsZQ4jLKwybx+R7XahglQa5JSfB+IqnfITMp+tiDRWfB+nhA
SNCrIuz3EGQt8HZWA9QyX5logm6yon+9fP7PNQ2hN3nog0jmWQm1ucnwht7iRcwWOaMP+ndB2ycK
OY30VPPj4wZvFRbNOo+dEXpdgtaDb4NYE9vmWZ689fWXaDvFskh+KCNieLnDfq/4tRgYDAw0NvIG
MXbktYRPcjqcsHeM4AIYnW0JQW+kAgRykxvzUXUQ80gExddnZM8YV61RUcT4FRowMzPE8uoBpt7m
PS0h7sTc3N6nDCs/1Lv4qApCmaZhLc8a8eREQTOQ4aFsVLWN96ULvxh7CI6p7b9xEuFQrHt+Om0Q
+h+huN0HI+fWriwCH/3837fF2txUXxBS9cOR3ISISatVJghswPloX9wQl3B48N0bM9NOz5hHdcm2
iydiRRkTKYaY+jl8nhLf2fer8qNSxIXOAQRoFctT/1B9X+b6t8iZp2/8m84XO3LGDdZEj5HAO9Cs
nVoxzHGU9DU/IyrrgLK2hCY3yXrSGGPxUQNrxgXrA2hQQhzRSGnXdT1EvNrK4itDVdHF4E4cH/KH
75pwRwo7biNrI4WWEaVaj8yqilHDb0RnB9yP3RFJejnRWjX5cUvDWGbUOskFAGdcowbRiMrhOdxr
pkf1bdmJbRIUfroa9ew2QkwwD4IichWQzyzDAXSvlpwHx7VbMSoWU1mbmFPhzIGG+ZQVVHhSjaOq
Sg5PcKLXS0aKEVEzfJxXDiOr/0ggWZAVNWbx7kiEcDOrOBptJOvtkw2H4osX7nLjncWSoJfUxbmb
5WOnMFW58wwBGlIvw8zENETrpnEalEkDlFKRqwbNLz9KyTOwOQugylMa4LotbJ/gIsSzlv7wyr9h
VVIZaMflTS6i4MFSXcxzXBCWb7HBBKUOJP9Og/RTHYw3JtvVdDCtXFQS7qSKMWDBJ60DVYL0xRLd
Jg+qxYl+jns0PXCnUWzZtIG2o82fMoDBdYwDz13Hdnhvf8jqZ3u0Ucvo4H1yO2FC0NiiC34Xz57/
6yd4JIHd+miwtRZ7N5mKEEDbZtGuE8QIJf8+6pMsVuhdFZTGma2N7ajn1dh30maVZ1HhjTtKUV75
4U+Yhhn+d/gGXK/PzKT8TBCXfx1G8bGNxy9d/V84QYziIduiBS0kgL0aTYXL/r5wnGAvo7Qpx3R7
REUg4U4dDOQswkPrTSEMW5kf4c5w9inguPdMZO/SJqB2Tpho5MDxlMHmotYB26pUd4YL5xobQmPi
3RDfC0G9H528ABqFNYdweeOj4firMP7QjvwS4aic0eSsSWkpDvH+mkSp3rZsf33ni84PHQDCmtpe
fWhR8p3SkbElYspTxlfcRUCnQMFLJfd53E5YiGgjWqzdKRBUSYFoP4Erql5hTxugmfzgas11TjoX
vD9S0Qawy1hnC2Mjgf4JmO8NuNTHYZX952Qw0zCEhhJvB8l2OadYyJNnepwPmlgtbaT3cBV042dz
iE1BxfFe4+XaTeiIXfMMCmPJO5yfOE9TPazJwOpDEgcUreGgbzK7UbD0U0lxC9AGPplmWcX677tm
3LZMj4pqzsZ6P7h0WHg7LOBElGNUOOFwd9FfLsueSOpul1kqU1j9mvFNTYZivfKm0m+2Oyn7d7Kr
B2Akro1dvHljUFY+PNKv6pt6oY2nfwullWPvmlpDfzoxAhylCzbWvck7RVZBKZJJ122lIuVskkqe
DT6e0wwO1Pi3B5rY+Il2E6bTg8tLtlTe/45kHgutzUMFDAd+nNFBmpvWd8+nfToOLFX5X8ggN2T+
BWqVCZuhqwCSJHEhl0FrEBOd2HofYku8WvFSc+OX0MjM1svrFT4+gLhoj0e4mXCx5QUMI13jItkZ
SRpqqLk+kSR2IhmxpQExNBf2eMI7BGUkHdLrHKkd6CcQS/ntlyrp17D/obQ5C1SwawlKOsyjYGrn
H29tLIrDEh1+UhrAZX6SnZypCUZ3Wv0Bf9C+xTHN6EilmvY5lmekJMNzNy7/kRhaNUJDJctx0Nbv
2ozVTCkZnJJs416qkr3PJRoQtRjA8yIDeoNvGU2GQDQku+2kSref2oGcEp4VjRCnFjNcfN3pHJap
5GBLlBluhzNI2Bdg21DGYphIjDJVIdIxzSRKC+acv9Dwu8On/2jHu+uJfLLH3Buukno42Pfl5PeD
xLC4d7qPth7jK5w/BPSKzrllsAESW6lMdqXDwZunSfajL+A11yxQcq6Vtne1kPI2yEO9iCpMwYvO
h0/Rn78yfhKywcg1/FDa+a0Bu1chggGYsjzgbBa0zA0HL4Bv1USE0sNz6uDYubBq1yZ6K8PkEng1
kcb9xj5l/cKa8nP4qzzlDGLdrTz15XdEaibOCLvVhPDcrca4vibaqk4FhltnFk5gk0OtQHM5+HEk
sltBHfPxCuP6Ljb+gfgzdBlFG3GqoVNJgypEcjdFaTQ/xSOLSK9CBuEz/Qq9hqbYMym/uxkuRf61
Bkl/Twt29pG6KDtmoy5XEcSSI2LPX3czf5lXagv6yFGSkp6sxFcPMRcmTBWbyKuiqGzlghl6C8H2
6GZ9r1E3OlQ8IGsr3xP+sPLggBnFE6on+aj6ZvigzMSh1+SuswssAKv1wK2VtLcGDP8Nl6YAB19g
iA3lFDTtGMHbbuyz26hI8eyEPcCqmTqzcCH6YS5Q5CyMnGjk0DDGix4Rcafp7W8wTVm/TZPml1b0
anlmqcBAqaq5GrhhqMX0qANHZc/yCYhgy0IFnYK3kcZzBh+ZUxILeslKv6QnNrQil6V7eIWZe4bK
7K9r5DKgc0Wg26aouBu/3Fuqx0utTPZnvLSobYAvmK3Dv80d6VkqFYvOZWW/miXWNHNZB9TaELVg
tes3Mb7cparhZcy2KJ730p2YHPl0U8qBbkGq/c0ZapAZD0AroSBtI50UthjLE+3HhwYx4XVqxpDw
pTpHdxPniYILODBOMJ9Oe9kgzxWNtcxwAcrOndvd1wzuOSDOz67NrMe7DvLi21z+zLAXa+N6a4H6
l3y8kU+4GYQUTTgx9maDYC2m/xbq873zIeyF31ND8n4Rykji7/ERAnLXZUTtFcciT7R3SPmSnv4t
H/Kk3nU0uIm2u+ZlQZxnB6RFofFSK0XG7kO3he2HIB0FKfyz9qheXpzyKfA+tchYS/vwk54kKc3K
lDpgOTPB2uyBk6QMm8LVZDCTKYBgvPDbnSvYrHBbdmNjdb0UCAyJIJDblGxcrtbQN0M51yrD9IQD
c90ukTnkCLDZx0Ax1XrAEoEMEVImddsVS+oXuBrVy/t3rAHceeKaFD1jOUFVb/v6WxgyWALJW8T7
R/A+qxz2F3mu9gNtLESnHsTGJ4mWhCllhXJM2ydoUjPDS64E4iyC37rf0yn5RK9MbjZNUi8JwxCx
AkyECFrbyeQYaB/mRoG9beqvn046KsR5yy8AIowy1YTeTeDhpGX9EIwjRw9O9hpNNAUTqPJOrg/M
I2CDrWTih8K+A7bcAX62mxrBnvNvfeSJwq9q7NIDjdLb7EYlzArIhFGKbTT9wGLVwidwrL74/PNz
TOFS3E9ZlmuE8CzKuPC9Mt3GUEwYGYd0t0CPxqEMkpLksFVQ9Pz94lNlgzPO0caarcWEMiwA40lo
ih7kS4K8NAcpbrDgQQ8flfXO9SdAXQvvyA4552khmtauvDmZ/i4NriBk9+ynIcyUOajeJt0pScDE
5sndXyI8aWWplYfuhJdFFjX7WS8dqnQjMW4+f6SF988jhoEd6tuZqY+Bh44necPStBOcHreS4gmB
kVB7eUwv1R2o7zSQkmo+cpdz9dqXrVEZLvq6qRI08LTw7jTSFD8ljJdHcDCyX3uTQpXAjPG/oWLe
jg3akNycTqZZe+8OeDG3Az+UWy0hJcZVBsRpfucOEEVR+olcc4txf6HhxYSkNLu7VyXvGJe5Q6SX
MLCC/B4TInofLgv4+IPuMUS+1vSLOslZoKY9OZlA/53FbH8yUlOhvFHVYWhGubZse4li/AyfG0jy
/YUfaBMbZV4Grv8DNDh8unzn7KauFqvrGxUjlrGL//4LNWKvJDW+bGJHzky9/AQeNrHF7RoeyEak
r103Tu9qOb5FbPdwhokboQxgDXQt1omgW2Ute71+nQEZ+FEj9Aj1gF+vlMXNS9l6U8QOcmxIzC1s
DivpuHHqNUhfRpMzEvcqqt+ekpRihMXEoxi+ZU7jI7sLuS6QzzIZjQYfw5FbViJx5kx3DgkYQ/p+
ABruRIgpovW70QAI8WGfdbDjvIw+NEhXV49rv4bfPgRf9qZAgMI2MNvWmfKQzkWUbNSTcTFYLHOe
xfLXpjarD8/jI5ruKFCVwzwZ/2sMhSk8EaED13ZzlTzWB2Lr8id1lKblbp+p36GxhQoingvMtEGD
a2WCmuHwSPNA3RsLcCXOuYmSJUpkc5iq9+qebUcHiz3kZXJzbaaCXgWxj7vJv5HuIUgeDz4Tne9Z
g0T32YW8o/jTLUJb7aceGFVeJVOfI3HH81ix0XddKd89Izy66pwsDYICKgL+czbyCl1RPHQ0B9tF
vzBOWNFrVedtzclhjcG1aWJUCQFTTiUVhfhVE0RYB2nsFD+YYDR8kDmF1fbG+Eq2vur25q03KEr2
13klL8ic/ZMgX2QteGy9RQNIe9ukz7yYq7/qI7O59YAaYYLHlAqO08fLVgfogJ3oupbD2bolr1Ku
fSBotfCZ6I2txmfzTVkr4To2aRCmO+nU4fF7t1hkaZV+oRj/gJjS1OM0Bg/smE1XCNtQzNscxh9z
MKMm+dhMXbKHpOpQM4Hp8jvg0zi6v4ooLwZOSKd333qYoqhmCmHoadmfTreBRqR4Jc7RNq0Q5oyV
QpOfao4ADJxaU3qM/RsuciMQ6KhRGuT1MIjWD53iZZqn+QwtRAOaxFpPEGqzQF992ey8tWz4FO82
Tt7XxgDiWMZJLQPmlwkoEa/CU7cobfmdAg5HyLrtgP4h2GjWB03Zbw6u1R2gQJ7vt4FvLAcjstif
pUYjZQrFgAh5DNUoZKrAtPdvGYSxtGUOrBzVg5cm1I319HgbOsCXGAOw/wRs84gfql/U/3+0Bo6q
FRiOjyiXC/uQp2H13XvMqrCxEegnSvTk6yl1N1AWUurx2s/QZOuz0g4hSt3ixS0PitaWostL5arx
MQz7Ja634WtLRgqsP6ry6B/SHwlDRX/W4bZpf0LR2V/lqoWvXWI8XChn3pC46SifS8VefAZkwN9t
mcGlVk0Vqz8HJpEu2z/KTd9nu2ndq8k9TNifXMkPLh6ITU/6JATxnWfbYer1VC7dwNaOMn+3arzP
LVLFKEPMRufTC+Nx5NOJhC0QOJfkPVp62elxNQnQcKl4HK6wVlBAIvPkG2x9GCDWsiGDs6bARNky
c+YhrG5tPiLR14thWkASfdr88C6hnvH9k75sRyY36910BsHBjbmg95J8qAKYRPRIZjQCqNQzXf6v
0WQlUE5c4IwPM/kf2xGCGeOwh9nLC4yDsebRWThGeMxhJqK1NJb62KHb+Huz3XJGJeIyAoX10fyz
9pW6ovXniCop0pKv12o+XdFjznVtKFjfT+CNmhmE0SdPr9HexxZt8vyZsW3Zj6GBDIUXKP7DsmY4
nJWSfAY6MaaQy8cSHZk9MZqPOnZsc+xKyG39xMupVLevqYEzBUoNBRgEAkDMitPswhmtdz393oZo
VIkQYOWM9/o6XEB/g2NsX33NrSEVIHRNvDECLBIwEx2u64wQu1kPECN/U/ysFnmjxX1QtI3xoLnU
kUvMJHaB56pfoSUMg3Q5GS4M4HlhEt+SphwXQew0NFdGJUufhZKj6iaOTOdCSelDfECvvZLmMM4q
S4qv0evdJc3NiDUuneYEB5Hf9XhBQNaTVcgeHGaHAvkmTYMACjPIit3g5LPd/PRsjwC5MSbAs2aW
cIVGdVGyVZf0QVuEY+k8FubbuKMHR2GK/XhNZNQPuMeYJsYaTfQWqVOKrdshR5JpRC/Z2jxM90D3
4Oz0k57o4Tyct8+s8EKvlai/xnfzex0awYzP6NmiO+Re/GiHqovYX+2zUm7QSU4ZCqGVF88V+Apa
sCVg17+lHVpld65NJBIQMuMqxHbknARmLIiyb1UJ5KmKey23+Lol3dTOuXsqpzOZ2YY4IUTlu3oj
WgwwKsrXMWkzJV1t8qNzii+vvPiX9yPxtTtlHs9zAYQqpGZfqrVqWIFe/kHPwIg8d/1iADJaGZGY
m3X0xOlBS9PMwtl3Cgoi1ryW3QHM8NWBGyQt8crF5cwEExKUX+F0MVkUu1ujI0gwlbqjTaqH29R2
mwFCXD1RHhqZvwWR+eX8zK+VTF0K6yrCnmrq6ukkBWykXz29zch0oCFUZa3d54az/1aEHuMKpKOY
5bvpA4M6ubpqHV9DL0cm2pXo/rWjobEnPZvkl4q0Xv9N0eZbyer1Y5Me20IjjgZP5SRaQgb8130o
QSNzo4nxlXpyREr8/WcM+gvpyfKrZ4sLn/Ho0Gi+2C1hM9S6OX8f3vqW9WLAAyuu8ij5vmGZGAHX
yUUXiWK0dp4wOuEZ4fEaKh5jbZXGvbVV5DI++OpwCCmUEORqPpK7zM1xyi8fs9T4NeZqPC94k6QO
ZBryPTH78AXHyHbfv0eK4yQzPGrtemG8Ss42GSUs+qJFgIP8PKejWYnafecshYvgBDedFQLzVDLp
E28m4lMJo74mcoAbLKG7guKdzG6xjwA31YYeJs213zPeGHuOd/ToSXO+Syzwws1oDRgLDE65+nPQ
o57USVkUQLH8o4t1P55rHHWmYOAMSOxMXA3rslOCuwenbYp9Z54FfpkNdKA30MU/rlPqVlnZVjZI
8YLqYto023VfWavGSQJtSKzWgPwCBaBwIr9v3wv62xZlBnsCW9feOY6QI0Ks09hNOAXHx+SuDh1O
J6ZQqTra9/wNcR9ZN4w3qYITEURmmtRv78DxYlZatgCPb664u/VPlztZdRven2Bycqf7TN4ugnZ6
Ed2ydQrGQ6UVFfe0+yanSHjqHxR3FlfZtiuBvtW+H3ZlMLP8VQaZpv2cCPgcw0CdNHNp2Zg1XxGJ
S2FhsACrxD/kGr3xXbwV8EBeZUudYyrkn6OqvoRNHfKAlfZRKyLkuOGr0AskCM+MYnntQKxQCEl0
iBt+4KHiRskaglgT2YClXdcciAOj2zwITBcB2uuWS0gDQs3ytMmYFinnCIDT/JgFPthlI8sMCuSX
2hCey3/TMrULyPQ0pL4KUo2HDOEPdPuv/p2S2S6E9mFk+VrlaBMXT9TGboYBaffsWdLHXQLiCWFw
gwnh/WqnGe6gbiOLxxQUDPIuCX3i7YkoNrbQ23mwsDiXZcCEySOZzbonziXKBlx6ZpuJK+0V1wjB
1z1rh8uEelDdAcm7uMast3kUFd0jP965uGzCohAksXXLLLLKVhKIicc0fObr0PBoTxWZREppC5qp
eum1UpKCEGIviynZ6Nz62qq2SBA94++Xw0ShXdQRTYRMYUQkWs059PyYnVb+R4qPQjNsxngrQojq
mr2pG+2HRT7Z8OMh4W2lnZxxC9+kgDhlvq+TD7vjFyZeAs66K+CnqDfNDBfQU3p5AqjjOYBzc5kd
xNBZSyJcQEtAa3QtEmlpXn0G4sLYrnvpwY5k6R1cBQ69No4CDuuluLoDpqYPSfSJoDr+Q6NVXrKO
+77BUZu8aRJ08wsP4Pw3FoQyVh1c7HAUQYSAr+cx8acEsfXpDR2vAPNQZ6skTKBbqZlwz2YcWhDA
pUr3m+mrgAc6bhs/0zbs4AbLMmI1WBlaUfnhsBU78ZyQbAFcJ1158CIWPOSuNSTOP4aQjJtMasGb
yFX35rlB5IMEO/RvqMuzx82csY4CLRi8Gq/Rn6c7U5Re++AonbrXrk/noulxHL/6RAFyRK5F7WtL
s0K+1S/bN8oRJ/VlX9WojEzOT2l8SVBxZHWIapY30YVtcPjM1tMTAxAzYk8EkBGwr7Z2jfac3Mh6
mB32SEK6abJ6t/yJmsSg1A4e6E3hMxTpGwWnCJj/S3PVqWFob0x/VGhx28mMQxX49ui+VtUNJoMC
jxBfkcm43u+Z6F3oH01EGMeHG5lEe10HLtwZUE9/6wwKZyNbSqxuljK4Gu4Vruj1AGmTUB4k54Yb
QzE5umNYjjLQvIzXMhEKNmmNHV/uiAABd3nojox+NR35VmpqMIT0Sd5BpQnHFL8Vh5jiiqVGIkcl
RG8nMmEdBO8WgSsAmOTUQEyk1vFi0jRaf8t29ZcUX3l9eEAH07SgDgh/PmFjclOmV3UqgZV62zSf
TZIxkQ6HwLdsGuXKVwr8TrINQd3b71TkR9sCpRLG+bzMFbJZXC11ylNV+5LJoViytMxR8n7NyaiH
2tSPVj9PiyMY/0Tyiwp9VlRFm9Kuhwa06JsetbVkG2NiFPmQ5uwzF/v7oCDYuarqGgtM3cOCRPaV
0w7uBuYSfBOLkNs28iN8clW2TQi5DA+aMry+Iqe89GTzGjvC38O8xsxd26TexKd/L0dnmszXQExS
XNGbzuO2kOIcFc/+B275G3+bOafc+w72vDI+Dr86AdeRvnRHukI1tkRA2t3zU9DCCRqq0bHYCsAN
cAC1f+ShdingHIX8W6VSmgK0P0i9zSOKFONDDYc9vJM8dnm730cJ9iwNDAbeU3W+XqLEnqvr4q54
jNUA7s6B9TBIBYOXybPOPcqcqvJyKn8bjrkQAsdIQ6Qtc5JYkfOjOB6nozEZf1d16IWGoDkujY3G
O2NbVAAr8NbFJDnWT4Lntm+1vq/1I7LMMr6cMvvYNne6bRO2DZd46WQf2PbP4+5Gk4xzELlRC0sA
pgLFL1XgXM+julCz5YzC8RTVvzE256BkzHARhybXNUKMrtTDAnYPEuJxwiobJTEeZytLL7bLq5JE
3EMNz84zB5N1ef7pbTiQCPloZ4eq3kGY/JTgpLkWRdsC8TCRK3Rkv/J37lAeIGVIk17QSyrH4CWq
IB3oc5h/cHNT5ZkKswO/dWfrpse8nGDtg8M8QQ8Wi2i5BJlxniJVE6Qv9s2sWXOr7bvr+l0IX44W
DWelKrjimBkPBhvULP/VwTo0dFqmZTnObrZfhN/5elNtUloxSKM3wWaquevODBBg+cogtgSk94Br
6TKXWwTf+Ptzo/Mrs5xQj9zCSRPevYfAgRN+oW9vRse0jyjkPoT2b4IxbeMdCNUMQ2gfI+bzgo0T
mmuljmNs0dpjWEpw8Otd1PGocFZSmNAVZtCSkYE23Jr0JEt1EAYYsp6yL8CtkamESHMCkVfdW2uF
NYx3BJOv7ipEFyJUv7aF2uFJYZ0KOF7KcWImiZFIu+m43KVxRek4SZ/Q6937C6bo1LW72usr1Nsy
jaGCTYTW/ynHoPao2NVR+gZat5ADrfxeVbTPJi8tHnVo7UkzJ8xV5w4OZBLVUMe9b7vSCoSaDxBd
iO3mpVBwqvDfSnRngHeyTqRQsLDm6QlRF5reZ6wYRI3jKhlM6FxYmwghQ8GQtqD/QgyvAS9G3Eue
6A3r58afn/j5OMpJnd/CA4p/rJFzH1XoDbMR4aKXoDmICEUPzL/UeKbkCUraWfGM2wM77O+08CQI
Vs11Z81yiudF0P9rUf5hsF3VSF3V/UFqLQgFGcNFtZ3B9hxv0BxX8MgZQXHrtd8cWOnHKzyx1B7N
Whkhv6G3Qk4L2RrrVzdxnYTv2t0iL0gy8w9TZkgH3i7iKCmwb5MRNZv2sV8sLVt9WHLQsQIuy98p
gz27PAXHonMlQe940lO3OpQVgqUHTLSz7JsOt4jKmGFbXj1XeUoLo+Nqe24fwGHXWd+7GvBgyxTF
0lzJhX3nq1a+rC/2mkCuvo4etn6UsMMHtK3lzq3qxSBX7/S5hBgb23BArV6nx/8txTYP6OmrlxRY
jE7u4FEWiNJubLHi61gpyCslHA58cBqk/+ahuGriPTKGFzandYecvdl313rrVWxKsO81KRgbvmwm
nxQwNDf+VhrplxKFRYNnYPxMhVePk67n1S707onNwuhjGd1yyzolFRs62qKdMQrrHUuDmElWyan3
C/jf5Mq+xQpH6hIsemnMwxyQjDWFmdo5O8W5Ziz6Xalsp6lxauGe3llG6UBkvk1A26AibKN1otpt
YMK4fhk6S5IW82tOGacArjf0/vp6b27atAojNv188SfeaB25gKDCzIG5wJI7Han5NrBRT1gPdaax
5jmDZGDxG0wkoPzLUZANFey3z3k0d0EUxNBZ6mwHRlJUVG6gx7fyW3Grwqj5S3+UXLF/QR/q3dFt
tuBww0r3ox8AdSAxAJfcosbSF36YK5rNaVcsZkul7fNjV1GNKJZobM2wX//Zaq40aL0pF+EGsLri
/ZpC98WsABHm/rwYfl+UMIzbZqBHp9rB/6yxLgSSEs+UCM3IaMjIZwsVHdU6ZXKZTBUoRR0OibbE
b3YY0IPwbyLWG2nPy17gKPsCYwQ63f235HU1Isy8dN4+nKti66wcoPouhppgLLelCMFl3AicKFCE
2ds2oLXKlNSdZtXsrmGklo9dvuD06IFS2qgEB9HlJau+zpTlV9jm/aI9W7t0lQZy+FfWWY/F00DV
CjZkBp+QnV1qSEs7xUOzQLy1rktBZmOzBrslXs0WdVrGngBFB8Wi4r0kIt3QfVjIeLNBrXjJMNd4
203RmxyIWatbC2BVxy5iniTJCY5j0gRat2IkoGjbQrrohsyeKEyou8tHtvJqvpCLpsfX4uJHuV7j
EJgIFTfsT7Dx2ar7EG76/kaKI5xr8Ipin9WRCIL+Z+ev0+iUBxPePHKufnGVyexPMT4N80ao0y1F
+u9/dGhW3iutgtJu3hK96w/wk9hjat3YYnvRbZgj4SL8WS67qzYyaZnKZ1pZx9vZzXX2nS1mkzjC
jfMs6zL7Y4oSGIcBrt8sBAeYnu7zM+YkbGkPw6yTyo0VZweu6Ra7L/5+YRCxiJImdypGjrUvbvQ9
WMbDkwcDAV5CqNN/iJ3ReRzLU8NgEG8ZgwQ7ZUx3TfbDMjDOHFSCQShmB6zXb2En0mqI70EKmk6t
umQzBazfLk31CyaZG9j5eTh3t+Tb/QQD69h/Tb7VUTLDvroplSjtz4ORdTO0alTyGo1czPuAys8b
QRH7P0yTkLuYaK161QYiGhgcFhIVRWWCuf9NQj2bywCDh1q4I3BYGWXkNpDLZYg+ESQZwT1izPTM
VxdHCU5uAWZjkKMH2zvcgHk8p5Sry/abnJgCxyyGJvPmRv6OlpKrlit8lnO8Q154dYX504UBfgRX
NENYC+L0XFW6m6XxC+9811WTFydcymIlUiP+yNo+4shXB3t3qAJ6ImivbvnIVGU3bNhOn3L4Fzt7
WlLEttptej3pIQuHnj75Dh4KsI2ZJLSIOhIrtKmh0kLXdhdHtNWj4pGIkGf/AQNsTXXL8ErIrFEM
zIk0opQ2NjMh5NE3y80XhNp7NeAGSgHTQgg31rzCJqJT3rdA0oVXCTT4u3oKD/YC/ui6hp+susEH
0/WLR4EsxorSrQNkoLjibTGkYBP6n497y7NceVKPqp76Fu7HM1MyG5yNvvTIKo22eeHidK+RYUIK
WeGDeMb1B/4oj8ZbHkrzvE7aKrwF06JpDQj0v2ApovZpz3bT4yuU5XCsxraCOWJGcb1C8/6a5Wbz
a/M4RqBfGVuz/iCUlASY7Wq7RKj/P/Csi90dhYfUQWCF5Lu0b7AT26u6s3/RgeMEKD8JMekLRMrM
AKK6+EIc511IlMRb/VtunxRJ0slc4yGNAPDk6oQYV/eebg/w2fUQ0/mydaijTBJteihj2TMGELZd
0psy2RzGOTkLse9/+k6yELL48km+Ic0D85iUW3tZfjuT6jviu1CumLVYB/JBH0XuyQ/nfLd9MoSA
Mkfh7CckZIisAxaumaRluescA0Ka4/BUMtHym7LwMcnLIsATAGf4OOAErFhDPKzt+3FODgZ+8+Xn
VxT/eHDilGxlTJqSfepQWdwnnR2ZrgiFkOBcDmMU4VKV5TX76lAvmk+X1TUx49KCZIHV4Pr4yqR9
+jF5DdCcD1MYqm4V2+HpylRRcXS1Hgvlw5nSOOYEvuOkpvbkgi1OpM1ohY2Dvp5JwtBAJIGnpBIv
nHG/lNx3gkRabGrGyJNqkg/nnF5+Aotz+6ZboqEq+AT9rIuDa2DpvEIDUhY0/E9pQNrKYVqQua+q
vHVRYiDOWKUNSi/82BT2BJlyIXA9aQdqGpuEONdquOo9fCU75/uRcVo8dlS/wsXn/SI1Rm4Y1eDs
nOXQ5enj7/M0CIOGISk8baMHjXH0j7uaKeuBXOTE6gMPBeg0ajtHW9JLtJppcbIEWDFImS6Mjj3p
W9hME47c47ltxlOqHg64Bm/s49NLf1nr466ncFtG5t7CBlp+4nfAGn8vr4VMhbMIl+7klOnNtn7R
ag/caUm/TtVQ9WZtA3HkWI6AhLg94L4n2TkESRLw9m8JDTdQ1UGqHTgbqpDzRCLXyT1HTJhBT9CD
ekYA0ylbytuC6L2Hh6sKDeGyU5fjMOSW0jX7R42tn7zO0O6iqqHADH3BybNXv8FM5uTydGkosY9H
8hwkGMgwViyq7nc9lmCaTJEAOwnJv9nWt144hSOvlgEvEE6AwnExV4Z47WIjNmHsabCCcPOfMGKH
2e9MrOIIVu8sayY7XygZOcvO1iYLKKSpZgAWbYN6lLDsQKCVP3baBOA4/hN+UW38ML5hRZvYnRfZ
NEo1HNFB3elgirutooaBpki26+vEUujhCLxNarz9TJpPdHSEecH0PIJaVypArtmWGYN2fYjZyjT5
DdObvTITPklZA7/kcmT8poaSnh5KOUfN5+OFVwulPmgibdd4vMl2CCeC+j1eOs8amm+55qIC0b2x
gG7uKtwMGS4fl21zaSyCFzxtxO31CgDavkgQgQub8banAyFPUHMbqcMz2dgw3EbRBgBr8+m8f3mN
dxQEBsQziX/XNf7h6CSpFDTB2XZ6SFTucGU3w121fBIjxW+5lRHzFhQ7ganLcld289RwHjVo6am7
8tHO/rzgFw/8o1GkePicPUprn+fB3C0P3ki1oo7sQtjwE9cJ/4MBr0hkZ3zr6p9hmwllrTZCQbYu
wOezMUlV2+JGQSKocNvDiSV74fUKw5GP4rTs9t+eKmlL80CUFO7ycR4P2S6MWK8W9aVqFJbOaoTC
l/w3Zom1Ue9uOdx8iwwSxDVAyY3MY6sdUz/J5kZYrRrN3vEJ0GESzlU2FOkGWM6TAr07Gk9wOjrw
ijcAGBkq7GZ0j/aLfHXaeRFYKMFpGJXb5kqffWzD55FozaDppJqm2/++G1XgMPFQl8PwzKt0BHJ9
4HJxUvZZTq0/3wI1l5ucfwjMYAoWnzwNh/O2NvuKzgUeJdLoVGMNWAoD/69GPPr7R8Kri5uSOQFS
RzZ6Eu/tZi6yfSuMT4Zx7fTrIqyCmUhHoT8hwNQTFGrfq9dUxlKH87MwHA9QSSKYb97gwPjZpBdY
aL7PRIyWmV+YlX2aroTrVakvBM4qGhWeB2LwRIWOPQ5x6DlrHIoMrhULY3u/PCrTKZvY2cl8hELN
Eo6VHvg83ZN8t8ggsaRBHLLgKDPusS6s08IAK2VccTmPHJ3A4nqpwWAJZNKRY5Vu98zLvIpDmQJP
wu4gJq8ita1zN+XSU9l8OQiCgZ5ExalFOMXqMKG/jxMvHz7Zmd7R6bAXipMh+HE+MKLaa+pCoBBA
d8E8/3Y8WmjbI8OrOCYHGGWvEYqpJxM4Nq9KWiFa/UiUskkAn1vKs6arg6s54VKKNFgSTtgEWvbE
cj07ap43z124Uepuk6E0suDLMDxSO9AfZnezEZIo1go5cz4CHD8try8mHCdBEeQtfBAuhtL9I1yu
RDU5ijNdfwTzDqOeZjkXWVqGiO/ZLANDEb0YRyDATvdRbyLEsfPJY1X5ahBx7JN287T2w+DJin3J
fVZg9C7clC+2Lpf/b74j/je2Ny1PAVNl13FSzgSQeRtwhY+qInPYvLN9Q65K2X3e7Af18bJJCY3k
pattX96yihAT9VymE+Swgpm7OpPswwvZ6DntEPpyUcypk2ZwMadMbwKnwxTwxOsjRCKcEf4xBGEw
qmxB9BNxQsTVX77k8mrfZGUL2WryumfKAcx7z2KyNLEIanv9W2ASnwHDklIxqKlxRDZpScO/rti2
3+HF0iiy9ikgLz2HzZlI6NfJrMPo3EHLP6bLnXw0C3M9He5Ta6aLVK7sTRlCNFk8bCigwHaK1Uj7
WvBf7ptYInyR0/ikG2o5zJbDNkBdxI2bxvYpaPLjBDYqHAB5wr9qU//pztbruKgtP9TrX746Vl0Z
lob8dcJIfrr46mMqUJmGM3laY1WzPlISUvZDAgBMPO5X/q2/3fr8zTgxn7KMkl7lX/42nYJmSwa2
bdnwfz9o32U38smGsPnipOwyIUe+Ns6Hi7L/Qusc52nVLmDN7V29pqB5H05ucKN3QLDOtyzm6E25
DVkPETVs+74AjUVM3AInTgH59g7UdqbqkH7n9iRJzY2EHnvXZaYvk9FSjaWJXirOXHfYSaRouyIY
fU3bntQUuIr3jeLCsMZJwvJPh6BQCj3mBDkXXui7h6lKLMsIPUOrXzyOiuVIDeosOQAJHtWDutWE
ZigF8/Tvfg4N0Reos2NplRvc084jenqkHfObiGE5OEusq5jfp2WjcjftEho/Ckc2IvDMYFv5EHRd
reVMyPh1euCBVYghYqiFaUQNitjvhcJBfAOns4hTdJUw4BYAjbunQxJUUANqXe678fKqApK4t23A
4a22p/PZaW4rEgoiSYgoc5prEUZYjQBF5QG7rqOFT4/Xo0f3FqmhjxUnbe/RD0CIFM9qnNsQ3RbK
d5WjssqzImbbkktT9WSNB0e6puK2/C1RXcjv7q8BHFw9M1Dziy/t/7qZ91ej6Q+B21YKGq3unVqD
ZmPjTEU8lAB78vR6TQPjrYn7mtV3hb+9rAA4rUFay+YmGFovRQd/wFYQMonacTud8Hlp/peHXOEr
AgpcYEaRwZ9g34Ahjax1UR9O0c2VZ4mmxs2Z8F2BrLF7t+LFbi6E0iyTRZEIAGic1EQ4KgQbEvh4
/9lfP/VTTSz+gU+vCQdkFL1aLUYyGoCQM4wPFQuGRpI1aU5VBI4CxhGPmzOOFcTmL9B9g1iUJtXu
zNGy/anuAA73uFVcXgVshzP/ex9/vD/d0q9ARK1B7QOWD+z/LD2OF9GffIpbrxZK7u4+wuKMm706
H0KX2DJ1R5ETSVOcr4exMS6mYbJmMP/tPZM+EBo6EdCK0YQlT5D+tTxK3D4Vp8OnKlPBTJDhKLie
mflVFz20ZOenBohBUNyR28FJeyML4HHoIQxRdRIcHO1N50b/emiAPdGu82JG3t3YeEAWNTKC1W1C
E1IpmRcOrJDGMc9oG64IboTjGSopYfY/kQiyjdOj7nXKWZUQRSdsvzb1amkF0k8DyBHl1yZL5OJ0
xBOJbYpg/RRhyrcGdHeMH2ZggmtDlIxP8hL87QOdSd6znYmpQlyMWTWsS+57IcV7Ey9NIAozEWED
jQ3Cs3n3koDfo++SQI/gZ0viUI5cNzFdti0ClpdKRZv0teKB9/yBRJewr0HKOt+eHYadj+wF/t7C
POa1T/v8jlMr1AgNwtmmgr5047OX8Q7q0md06DZXVuEPZr0jmPXP4CEF2S/NZys5u5jLOGn7B4sS
rteYaA480S61tt4MCFnbFmf310alhNxydHqTef0BcmvQ6IY0Qz/aGMtoZ0Kz9ECIH+zXbxcKq81s
GXgNmraFrTwUj2fZVjyUzOUps3UXP+jUF7ePzzsdxlVv8roxwZK+rQQhrW+Z6D7VPDRVo4F6197Q
3q55f9RIBNubnvdVH8Fcpms1KxsE05tJ8+9QHwsexe2V4VcICCgWH2922kfxkp6SXz1grQBanCTa
5cPq6eMlIhuyIKldVkLAUrI+0vpwt1dejXBe7DEt0QJJEy3J8Du9F2rDlJhLhCqK9sr6rUDDcVcV
U9k3fk6BVULzF76ikFDKF/tX0ePBSSuCXreybxE3iwHueXVJ5vwX79JplkWzqzmpdIWcI6ufY+ji
XXOKLMI48Avf1/ossSqKnQ1Mwiqvqkrcng3Jh/+chWMMOhQS/tWaMHcuphS5181Mol2kPs06JiLD
zT6EhuWvtm0ptCFaKAV/K9zw68VtJrUu94fBPB/bG+yY900gtTNRDgzW13WRW5Y2nImCzF0Pet2n
QUITl+93sLClnIeEXRX7LnHyGp2eEErgs8zLAfIXeP+pxgySbFjXuPXdTo0AFV6goop8OxadD7B3
RTu10qyaC1Bnjh0TFxbiCugSc0uFwO+9HhfbV3J5IS+0/qsYTtnw76gYnSLpfYyfmN1ey+lupmhu
qltu98rtTEtErPo6cZcaSVZEtC45ysNtp2+KLLKdrCF8Hnq/IDBJA02s6NDopINMHq0f8tCvvstb
WpYCH8c/IqMkJBHWJ6exTfKvB9Jrk81tYuXZjgLK8CGTA3Oshm7qt/zTblEF8taQq96n7f91sANE
mFxcNnYoeCJ2nLfSZr2q8fK0XsNm9Q8AFBFr8Eau45pG9T1BwH1EXLhRHWGyibLQbXegZHbFuUiJ
6KNjgL3pKz42C+wmU/eLi2blWIfqSKQjfr0YjiN6pn1GbJVnsInca601i0D6shHitwUPnmpxt0X4
Pr1N93KbaekWd1IqJdraSAiyeU5AqzXrO9MrapErTka5SvaRIZxM79/Zbuf6dupFQ9xBJusYcyOM
Tb2Uv7vc1mABz9ZnvG8Z8282xolXbSh8SlQyvrNNMZM4uTVS7t04ZWAfjbKYS/prKnWjHCLmGrBq
jXipOQDvnNpfy6eZAy8Sup56aaFvxJKMtdO1AjnjiX0+zVuU1LhJyi6YzZlRw+ROP8mlHbAPavkX
mkUFcSeSZLUTvrx4CQ35WPyT7uN73Dq4weCZ8b+Q2AoZZYI8jXc+UAHSSBihq7GOJM6dHnfyrr9c
Z7h/fw4gsJ2sqeX6Ey8HLTDBC7l+o+KUKTNBZghfjhj2AWaGcuV8Cc/ys3NHe5rkxi2D459OaRCq
AHMJiLMTAcND8y/pagb0Hw995nxBHjD+BDnoHgSDwhcCv/fnF1yQ3SezJX/Qzp67y4YCDm8oLwnj
8/7Etq7ZRYnWQ0GbUZHAJi7ARCq90tXfijPTCSeGOltb7uCSuYCru1T/sPnQ7ys9CmZDkpmmt0/+
q6UqqPIN6LkUtSJc0Sdsw/BbcSDUxl5kqqgWugFvoXhd75ETMnWlCDyNDsCIT9ZiOeYX9+Di8fRQ
324g4GTcSDJdoQQL16EUBMFpylj35M9a2meLJtopxh9jtKD3Bty16SHV0wnG+ecEsqk+T2Tsj7tj
tyERENiXUKFUFlIqyylS1ee867A/nNc3RkeHs4CprtiFq7QYEajCCETGqwpN90bHy82Xpq9foaK3
pF/MQSwCRzTkX24RH/ym8D1kwYemmDKzDg0/ge6EYozfPDWPsaKvurJ/g9Mzuu9kX/qDxm8AMJSk
Jlj7QuMfi5crsblOiKHdwmlt+F+Ae4dYWgn51He+HbioPQSWZ06CE1xTu54leylGwmUwj7Fl/tCh
BJvDJljGxwTr0yWVa500A9OcBEdIx9TW60i9fmPm9m+srCTlVfO2OOE1wVrQOn06U3otwraCFqpG
xK5bBe536E8GKZSlJVSziuNxezI9cNe/THcdEBgoEVfsvS1B/+t8/fL70PH+bVU/V8930rAolcHT
aM5kcGrnRV2LqNpHsCTlXoQeo8ibKzxrZNw0jsYkTH3Rdj9JdbIZyA/K/Fg26d2NeVJ5iOTnw8jL
bjfbSOeyLdN4nS39OvRYbthv7FTdZiGbe8TvMSZCT8sGyzYEtf2WMm1RdWVEAeMhUFoAWERoIzTW
omSZn1mulBcBlU9YvsUwF4WmNoTuxWfq7SzhHSTEFzk7KwrrlKBIVB3Z8X/UYhK3YP74dW6EKLBP
iITtmhxWyOVB4Js8wOcoI+2dtAt5Hyd09U+WGFwhugiijGTphz1vTk+4kjn5QTCuO5OcvEbAlo2C
6TWrS4aE0EWFViB0U+R3Y883yB8ZP+7EfvqiQn9XeF4Vg4ugpIqX+ztumt9vGdpxbYws4wSQMbGU
tHcBWCnKimW6x12dx+8Y+45ER4eS8sGiGkB151Tt6YsDpjJVX7s0RTpuGxuX+RXVAurLtizO/NX8
xDtxvvjp70vC7qtZnXdIh5vARYQfKKEIxghB0NRRw8AgS0CbeyqIUUgTs0dLM9vZtpW4UPca96iP
OrLVzGF8eZgw4Chw6Jywgmbo/zbDeFNnh7QR5ETzaKALPnqJkqgvVhGebO07alYPglT8/BeFjMls
U+R/4ghQiLXVeIR3tyOgJ03YVle9w70hsrLn21Lk181z4QbhzuiqIT3FkKR8U+FVHLzkKVpji6BO
1anfusu5wK3hrx7cGdKI7iorTEe53XebV0oe34BA/nbyz/YLHch7yx+Zc2CsV7ry1DoLPtQXtspR
5fMlLm5dD5SFIVXp5Bgf+4ry5EMD5un2YhRwRU2APwrv0BPDPc/JOSd6r1saO0rWFJV6qpnkTy/q
Fl9CkNxVI5LhcIT9wfrR7/d+f31m8rQbgNnr83sZ67bHZtXBxxKwVAWhB3PC53St+aPTPMxwFlzj
GEuE4WgJjasU9QxaqXU9o9WOcZ0JKvf7lfHf+fUUaUOZfRNUXp3EwZUE9HM0KQQoS9kAYKFApm7x
xRjgeh10AmG7ug1r2LISThJsqGXz8yhOjN1L+5J9b+BLpgTYyrudeJhNs9JFfQgF91tzZ0Z3/CBD
hKVjlDQLT7qw/y6Gvz+YNVbJvcSOdxn9X+GtHFfnwI8vyFqvA2/k1J7cV1FLI0r2Ptj6DQNNnpHZ
gk6iGHfrkgcXHkTmMitLRkr4QODuhI+I4S4hzaY0HxkrliHjrxWPnfa/Src7yI8AW82spbpEG1dd
0pr/HgUKk8O4EtHman0SFE48Zxdq/ssFixSLzE1qBw6VQhRzhySxSwyDlu6heLvdLyPZM8TLxt0C
lx4Do1qgJVWOHsm9Pl73Y0sXcP4CHpgO4Fn7UHMclFsMdBna0Bie0KDvoAqBG90dKwKFUqSb4dGW
bModDPRwJmhhUpp91+8sSmJD6v7EJJ8x31jg2v88S/e5qmoiMfGjpyNB4VIM2JGfAp7lhhsaQXmK
RPJ22IRI4QQPJD85dIZsS4WGsbGW20OGgLLKjXhm1hGMKShGCPQTjA4mft3PwcFflCfhDhngWzkO
BFsC3qgxs9SsK4XH95+9lxYV4AIrOq8ccA4Ws/pIe35CAnkxFKumdoVrEuTsUvYoOunDqu74EO63
FpyGH6t6QAHRg3M4f5r/a0jZQQn6koNEBKmTnqlscXPv7MOb94x9mCE/4otmKkqXlYnI8A7VA05/
29NZHEuZRxlxoQQYFhAFuplzJkTntsvmQtB9CbcBKxMkX6nlBJc/HxQrnoCUHb6MZ03dgsXz+1gy
a+x4LSktOQrJiUfyboKhlE9maazKIE6+3iHWLUGevScXCZDKC1PgaLj8yOT5EmPia1LcfRtZld2T
oiibJVfTtEbyVkY71qLq3gXp0eN4tVGIsSwN6YVDBxPGJFHRbdX413gpkq65yBwWYswTpbiUDAta
G1R46vHnqLN/x1AXKXsk33vikyPSyKIIzek6XCALS/eWNW2BySJth4LY83Yp8Xi5irBYuSjKJCoe
y5ICy5VteNzqwJu2kCqEYhf6ZfVDVVymbCWo809Z8KC+GLjWe01Dr7LAqagwdm2J6GhPb2HSBie9
ZdmVPp0wlqtNoUCJE5jDmBX6QvYYwK/6E9ebQrP9A8tMIrx3MK+O2NIWJacmjDPjP5WJcQ9qemov
j1rZ0xeko6NBScuhRgkYy+WPF5+7wQB4C1jjOoRWTlfDM2ZdR44zeaV8E9iV9Gj0o7xyJYrZS2b3
tYUUqs/i+41a15qp4mmGWkbSV4m7pMceZzCxCI9ea+Q7Il634r8Y2KmB95kTpWwVtE/8Ez+4a5qb
289xgpWhUH0HCdEFctrVoLfC7wXnEf3GyJfRKNtTmZfDO9kK2sfADlwtS0GV4r0jycyvjO5Ijhkw
Ozbf+rNVWgDkJl24kPmMaswIFkOiibk8m/K5vf6pHDrcqampn/I1V7K2iZh7WhWIUFK71FlgLP6L
RisuZRAvNiuycutKJcW7yi7/EEcK2V62y0Ymk3bwhDLhXyEqbJs60/+Ym/fR4eDgRCSE7GqrI0D8
Fs0IeF6W9a279Uwp9RVQF4aTQxXtGV2ZQlKPFYtWNv+p+tA160XpRG9TAKcX7nd2mjuc1dG1AvVu
8o1SGDHYRbyiGpkV3Vuj61lXDsg8Hx66HS/AkMj8g/jJIM9ShavURuHeoDHDAKbB8kvBZ+FXk1vt
mTc/XS4PoRbsoNc0ra+O21IHnQLtPgAS8Nq+ovX5/KlygxkW4Iqg4JCOrsauSknVsv8acc88/f4t
JHd28FtGqEsaMSoZs+dIWk2UVrmgB8mzGZXxO0NGKxVOSfmAZ6KlctfoRYhvmOyC58SzoAUGue7x
daeqwqRMN0ZDGFLsfLam0SWeox0y1LDRCoHBqV+KjQohhuZofBhbcDbXmsZi3OERWQtpYAGV0XS/
O+thuqVxZnne1+WMhclgW7x8e0AczM0VclgmOHiqfsi0h4GNWXr3j82Q38GQYLcmN+BJrmeIb2P0
uYdWJvyW8AenoVm4DB4k/eIdTMKOMCN7Jhm5YC0vT6vj+MQStnfH3g5qgx6ciMerKWy4gX6+QyEu
9xytOtYRpgMdlwpLkGqCr7vCRCtn5EPVU5DOsZyK/+PFQMkeo8OS3T9T3udkjWQSHJbeemULFm9O
BJxq1rmrUKQk8r8VyfScquwA7dZVV1KDYxCwnyY0VAjVW4KxA1ffMatXFXpCyzQxdaQqeD0T5emK
BGio0AdZE9AckNjklT3xhnANEsdtQAKUwayKP1F+unnO/WNpARi7EcEuZOBOvln5Bnujlxh60E02
rlNAYtcgrzMcuSzmhL8by23RZ6D50MrO3KsEmA9pPb5S7vNgLcWocKyBd6IFztGLvTcNDzmQr42Z
s1vixIhX/bz4ZM67hUP7fxVREkAMaQXzN7ota18Ys6v899o+uSvPRp9iLMIdd/48oIpOO4LZlDPQ
ay4GLYmAEeSRDOQQZlmVK1GzkjT2wM1FJuMFzW1iNtP44Aojz/k29R1TPXviLQb37Qe8wwyKld23
G/vw9OUDJsYGd/CNb6VmT8e++FcgxbUkDdwIQTGmykeAMuiHFcopOoRKQG8OMjjMitqHj1ZDRF9v
uxs1sKRsYE/SWKmtE5g0S+MidCxS4ZPYbE5kZB3ZyliZl8vc5zSEYYu8aigNDQu6lvHPG47sAYo4
NadCbpDetvlGdY0vsK7iGo/K6aWm86dyAsApVsyJ9biBb6S5Dv55w031XqyrFPOclVowOLN5WmMc
DJyunfjvgcH6Je3Dt0hQhPtmUbXQGkH7bq+eyZLzPu6Ola3VGPZ29XdnhOwkCXEhDujdW+/FlySK
hpMp125qzDHx9k7vhKk20Nu5wISmof/VY/qGp2zGDnGS3oS+p8zYom/8Y+OOVFXXy+2LtKucBT4g
vZJHmXV9gIBv/MMzbMaJ/BA586XLVKPgE40HgK4/05LIW7MZBfq4ptT8AS5VBgXb2pEiYT6MqMDF
ePg9GCggzzB3jV87NVJ505AFoGr9lPQpSHDvbQjWQlFXxj3ObC5hVCDZkahCGaS1F3mDAB8sVjsv
dTJrHr+4vqaPGfbbf7Pfg0IAu9CQR7iDzln2XDEjgU0Teoy/Wt0RCIYuGwAEJhYvh5WEL4gK1oDH
6bWHC2MgRDgJU4kBUHG3eUKT2XpN4oPr9c3NqQ912jOz91bQFn1pCQNYVEBPACJgwl2Ta6PnCcbW
Mjt79CO9iwMmrcfwDMrzVkPsilqnUUXfRUex/TBMNS3V/4fMADjENpujA6FZOsdyrj3r9quzKIRE
Hta2QvA/mhr5QqUrlgx9pojVHVlenhddVS0eCxgozoZWCHEsCht/SOOiT6ELPYdIJ3cK9Plbs6WJ
DJizim5mZXaA8zy+7gLupYmrviyC0gCknoBLetFXuKZDYLvvKcUmCJnTsuX5Q0I2QJdWEehWNPq1
fcek28+65EsR5xf2JeeyfC01GoFAh8Vgv2dXNw4mNKKr9Og2HivyMMJkWqWduuQeM30g65cKxGWr
jYx+I6zLia6aUACrP6F28Zd1tHjtGzQivsjBdgRON5mmHHsokL4c1la772cK6WgufgoExt0xNWux
6HvZPmoJgA40x75EPMCFXG+rbqa1NXcCJ3djazoUrTBvX5OJW6QkXd1oEXVRgDWMZL0vRZXYfjtk
G8D4O1phWP1B+YvnG5IpAbnR0wUToHyrcG5YGNGPrdGWLqMW9hI2+moRA1CE3wb2X4bm/oEyQPhI
dC2KWFDtVLGrlHa1GOIPAk3Hxsc5EFol/Qe1ZiaFKuPlXNc3xqR6m3Fjfc3QxhCMLBy9ufj1wKOa
HJKj7T7i95wydM7oe0+9RWyu8o/tiK518TmtsiGyJHI7t2erxwdWm6Y/b51XQXc25kMJKitLBu5z
NxU/XAG2L6x3G1FyYQ+LOhf4vWqd76ADhuetbiNHSHLyFclgpa+xuvmubdXfm83VGGhvOpoPbUWV
8Db9hf1UeUPR1SCZGiWhOmTSXkZf6C5D+B9sqKQsKluVlONX57EBmiSdskM71Tnf0oCcHzrtaENU
3r81F1M6MNMQy/OI6ecx5J7wPXIPFO0nj77QlxGu9CWNji87D36HnpCvCcwatq1uyMPO8MMrT7Ov
N7/LXT3wrX8MJbLlYwA/Aq//Z4bYtncsVIQexcXQ6/Uv2Teed6OKE9V82OeG+VCNkLbYAMdP9oeg
UwxUPe5k4WgkEfF+WkX/ReGz7dEh3rfNbaQy5xvq8BEBLevpuWZkyjToMJeFU6X/F9OrCTFRxQuB
33xdjR8DZReNfXJIbrjkNncN336jLcB3rO434oT6hC/8ifL0riNuqwlJ9BZFsMmPbS93rZYuNwem
beKRgXENkK1jUInI11OIZ2Pfxlda9LHV1NZrEWUqD9K5JeoYqTqKWO98p5t+isWVz2o/6vPJ7Um+
F9i6mGDL9t8h//6HnfWtBAVnA8XILCkNW+id3S9XMIREzHWkmXNNzpnxonPRBC4gLDlqaQw8j36T
H+srJ51kfRdF1GnYyKILysD++aaHOmrpkjRdpG3KK+tY/YDv8CvSsCoAYv32jYBeg2DNZYG6xuyH
gP8rqR7HALlbhQLjQxoqHZmg2Z5IDazUwSiKfbSVfi0d57WOQy5aF7Yi69hK0vOXxb4LVp7aaIcS
V45YW4XNDVphGU3JpbeWLIJ7OCjk624JAyJ+Oj3VC9U/OZzSfTU060wNMG3Ji1hsYXwgiaAjcudJ
MjhlvYJaehriJ+HC30p9dgum3xMZdHN+MKDucdfMQuAvZszBB5r/pAOho9HkFyZabavqqimGsX9G
GWvbXivhqGkOEboTp6dQhobaUVoy9avsts5U+SY6g/0cGuedUh2SX2FlAfgLGr7ab+BQswBji1qm
A41kyYrvmQQOpQd8hDIE7lFB3wvR4sRPkcV9kOxIWJ5K+FwQbWfFx/BP8hOGdkuDd0OA0MBDQ46O
fEi0lBUmZyI+kphA5ha2YgTLEl6c3v+W6gMfCXaY82iDkeKyOIXE0s47AF5LLdPgIgddDLYjdXyz
tAAIChRqzndnszS8ahVALPlGeqgKpAr1QTIJVkZ65qPy2zeYUVWRQphDKQ74VluLfsS7OoIUwxfb
gxeEVUWu0zT42dcp+szw7rw29NPmrWa8glLUCQVJAUeOM8UuVG3IgUgS6MRoTPqQQ52pjpch0ifq
zrbVViD599SPlxLJ4Y3pRRCRILX20ETF3/WqOL7F2r4LB4kTjH0BIEm+IN1NFURky0IVVSzTDV6b
5E/dV8SJU55cmy5cyomDLgT4z0EtuStklsQCSRdmX2WZ8bj9cdZPZcPWmqNFE6STGJo7WTdGPiDH
rOnzPFwLEYiy0cYN8/Y0ZA4yGDnO8MrZckFjGQZk/M1g6pRjYaG1IH7/mfLPa4DdadO6T1gJ0t1S
wtiRDF385RMosh2cp/hCrpTP0XTlIpEPCvsQACc5Jq4wYDGRXqDMWZLkcZAZJPdejQ2nD9nRnu6+
AgO5KfenRyh2PMzQqKP8/lEJVTlKA8MC55q9lxzsd5gGPNfT/ZG9q6uJVpACFowg6mk65yW8gnba
6dx612MVBWCsX6IECdAG4IHKPWeFYW6vDmOQst5pevc37OUMcp8gkekYfqeQtgT/5fdVyF7fn0cq
QlEqA03UMmuIi5rmw7emztD4iNyhTiQKAXOVOxW/rff2epn2MMe5CmevLRoUIB8R8A/78pn2CIgm
8f/IxQ+6MZt6UPyyNkvpv8iZFolyV19kmahgn08r8FJMbA4kIYbYw34LVo1fYtOt9ufy4cSvZoPk
D7+WRv78I4MAHbp18HmEL4HK+8oQgOzNwz+Wbd+DSXQcy+E3i32kYm8Lzc8YiiGpd8d8BNqLscVN
701erYWoOT0col7DzDlrqKI/BW35pm7by+Ewon/FoiZz6TWAYabxdangz1mFJQzO3c3v7kaOdXTc
gaes99zW4E7MAjaQFLtr++mwPflll0mrSGUy5wdq3SSnXRIXxEphs2DCn3fGSHxEP/fG8zcURhwD
ud15iNH7KpQPDpMa5D8jiriwBW2Oayjj95TAkQfmKF/YbWAnlBcmP/VlfnT+goZWGuyCVzjzc34R
maaV4gLqHHzl0Ygx3J31ta5fFzPj1I76vg4QwLBqkcxhzZVmlqwXaUjNgGpRP9vsBN3IGw6gYYAM
xAvTCYx3ekYmO881Pwm3PP0e6d8dJipsTG6xOJ1hkn1+nJZ6cc/soPmdP0kLbDcmOEta7Mc3bAcz
4LeQX81TgKqao6fZrOtJYoieMgOq2L2aGtDwYUvH8NV/Eqh4n0xB+rKuKLvlejixLYIRcqFHM5yS
6TqKFFYD1xP45aaP4+EIxAl16C0tDOQvw+5Z6AE+/U3TT3rA5IVsDXBSM4tINZbvdleiZhzYiFHQ
L+NP2SMOwK6nYxx7lRpFt6/XIH6epFRKrZ8hP1t5zT1gh5YrUT1Ee1+M9TLn1m2lpgwHcCrocav6
u4vJamr4lRTG12SDDawVkE/L1MRDUBAEHP0K5QjHr2bQQnyPliZ6+z5Kw8UdGLewQ2Mpg5fYQIAk
0mPW6T5qD/QAgKlFYpVmJ8oStcajEOtntPrlzZA+vAH76NhFw3caVh79+tz1/XaN1HcLWH5WzUvM
GJkbE/4cGceS4rWwsUyszoBilvxyAcjPC7CEoaMInGX3SjRkqI+60fGlB9AIQkvo5OizATn+OQ9+
gKlr5jlqVtBWC58YTWttEoyfknsLP6KOTWvXsvgOrC1MHwm8tyfkGBjaU60J35DrfRFw2nrQbit5
69kPK0zb6rTyV3TfrgDtuMa46iEP1oj06wTys1Xlq5ssp3DRnjTxXc/sxYPwhQcH9tqTK7o7o4L4
//FtypJ0Znk0g5NYjBuu7PB948wmcbbyjKvKKYTQ1e7ShjNcQEzIcvxNbriCJL4QyCe5n3TkZmrd
DpBibJH3W0knVms6/yN+s6CEfSYqKaLUNZe2Opg8zW3N8EOZ0IPp8IXC1HzHEoigfPWKXEg0rVa9
hcb/0qTLyJuo7LZoYHjm/e52tlO3Y9CSSukTGxUOtKH2rfeMMY3a6l9eCQ5kiugg7qsWckYLwRmy
urWkP6wWdSvFS5YFGB2fMuJYqPzgavd9bfHofUbqyQP6NgM8ALCnqcKXBimYQAe9QB6PS7C8N2q+
f+lu01ghIOFg3PMTmcNk9P09vxuikxFlNfAqp3wXQH+JVCFN4tZt0cVXfcDQcrKsRwPnB7frdJWB
ZnrlKe6/yntDRV8ZmZse95okGSykbI+4GyBe+QgxPxpzptrli9b9v8Z0Xi8KdKaWsMbOC5p4wg97
UD5D2WFCNbMGaCZHJCi8vLDG8ZcegbfAkhjpnN8epoQ40lqB38POSdf2hWteUoq/8dJ43O5XoCha
JTh24sKTwgxY2BGY4UjfLvnypblqIGY1Z3qS4AL+6ZG+MW0bRQrLvbOq4Hi93MjwbByyDS2StKrC
269XeXvBjn7ZpAsFG4C22SSyBUHZtq97dnSTBquwyJZCMnuuz54p95+4QZEXp5X8jlQD67b6DzZu
KZkyulaY+LBNcRrMeNnnM7m2zvJEcwL9pgUH6jJ2DTXmhQjKkSvLLzbNEQ/2VKL6KNRvED/jL64u
0lHKMyLBJT+2oYRQvwUi6SHqlZbkCNnHLnaNVlkPEw2nMH2Mm6vFVJOmibEeEQ1njr8JXPYkiMPX
5j0ABFprXiHxVFIlUouGM0iTzR44nunXP3zmutmcHUDgrSP7cCVQTtZTBvqotwuCU58dCN4Ug2Tj
wbkLfSiGVXUuwazPQBYgNs/2msh1xM02dyqkZwMmrMovrI0Rn3f0DPhxssN+qrY0eeqavKfF6/Np
1NBX7OnpYhMNxOT6gkeJ8jYoNlRGeDspFAeZfC6Gn6qlZDQrl/++j6qZpsZfQq9E9dZShb6er1LG
vTtL72A6GN0NKtIndYUq2cKwGWJ4ikzE3TuMKbLoznStP9BsxrKUN2HIR/FjL7ND6kJ+jQrPoIvm
HbmZNs+ZdStwYHdeWsiXFXE9xYqg6NFFQeG7VDNt7FX66xPaIYEHtLaURUDUfMV5AptY2nLQo4Zj
a4it9OpGKtA07EJxhnFOTQpu3jz0Y3JJajNJ7WLK8oGuL+qi0WaBMxVOlBv+PfwVVpj2S4f39Hw0
6DbQNTm8J7706wtNpi0WVJEjIS6v1/2V76xXxtL/0BXV/6Y5b459BSOE4On2V9ihYo6XsSwtg0vu
DtGGAhvKhzCmRNuLCczSPqURNbidDkj/FmPHe/ez7N61o/SDwNj8TO3PcD/ayqKzaHBGjYElgWiD
gsb0Trj2A+uoVHO7P3Ht+YZGRm9zw1l9jWi1rSxiLKdQSW/VtTm2hWFyi0OE94GopjJg28VCqKDf
8HZMkawQFntmu9L76HlWGLk88LbVfv/KrZjj8REY1duZ4gbZ2ZiyvWKA3ANF3Jyo4tHblCFOqJfM
i7/nJlBQcq3u+LWCUtg67jXlS/ieq4+yjGpiqrHB9O+pJ+/RncTCtLWZNFyhqIJ0Q88GM8+gSY8J
qqsM0EyCW/TMoPAtVfsutoQcg6qYfcUPIQrzsPSgDa1+Tpi6CCy+gyw1Xg3tE4lfLO+jMAGN+ltK
PSLHNZ63WJ+Q03u4Mr7+IKMeP+SHHOapnkcoJeWw3zFJbOCemVbjzzrZ2XajcEZ9FmUKHw1puPkN
xLlM+uP7jZbzB6+KbxIVRnRAEdWDHBo/7SjP5JOYQOJHeg1s7ej/l91y50rg3oy961WCPB98PB3o
lIYkGmkox+ql7TB1eP3vpkmPZtXNj22pVAyWEA2ZbJAStnAlA4S7V6ZG1/4MNwQLTwfkI/WEjE3N
pbm0kI3Sa82apwQDj8yWR1ZprUy3tfFsRDvOpojGiqKkiKp7MJXT3bWZWKV6aGQZNi/zRH0nDTxh
axJiQ4DdRcjVduhtotdhn1f48y7lHhfGcTiAHhk8svKSxJJB85/SXphIg4pTOHQ9I/2xRRIFq0d+
gxINkEaXoy2BVcc6ivUGfhTcEAwRtjCWVlwfxtHUHkcmoVwxDBQupdktR14obpwrEYyMkyHijAp7
cbo5bRyykKDG0n/QkiIu80BJkqKt0EQMstaWzvlXUYF/kBqDoCqqZJmoFJWFC5cWtDkRe+F2XT3o
WNcpK8b/CZQLoOXXSbkJ+XzAxn/+ORSFJpzdtlLCGzX7mI2th2JECLsNDN+Q5ut8A4zXQGp5myED
HKO1j93NrPzuImTwjb+yPae+14i5qJhbEkLueKdb/QmFKhIRxBOKGQ3+h6O/1sAx6f9wQG4Qz2q8
M6H4wrEfqcpQ6/pWIlDGrxyeZSWhJObmdskTJkIre78927GQkERRn+qMdeQKuUOSkmKDObKFkrl0
kEuieAjL1yXAOQaR1Ij2kt0cQSwCvtGLqUSlwLY0PkAKqivunL2KRJTh4+xb60QyiAE7E125DSLQ
/mjv+4ozwXSkk0tw4Ppg/F0eODOYAg2xy/eL3RBzOnWvkKfpsormfq+40/Q58DK4pMCRD9BVgI9g
Cv9yV7KV4vHpGZ8n673aJLBGr84F3//GquHi1AqfVoRhIKgtqnxF17y+SAaqGMgSRUB7GBfvrztV
i5EQSh8952rxiNLoI1vvLPB18Qj72DU2qF2QHxlNmfyoQhgp7eQ4E1QPBwdiIJVj0rT94IvnXMou
8hSTkoYzdzV3b0DLyJsMuzioiY4faPu6gHrVEPEiYxWGeXBAZpmrUSjLRrmExrDht9vs+aILIglH
pMfEVUlpA0WWrsO6IYgWFVJMXcM/ebzT5/jBNIKAYUA0q17P5sjeygU5bI8AE0F5j9MW6KUChv0/
in1G9Ea00Jk5GrFsJYhM+2HTwiKo2xmPG6vVUGCeFph6z93iY8tIaghLn+qcwJ7eOLUHpUqp67Pm
T6ykTVxtxtG/CXcE1ihvyEXCllHJ61GRobI184rcJPTw9fjjKNQ+N5rS0rFgeoNEueZX1cTCHgOj
xM1gUEVdNtckBcLmpsfxkU0VUlTmcl/arrFW9qPcAhIZOEZv/cgWBHh/1ys7PCIG58GILIBB+sSB
YPcGvLVgxXElxKBs+1SyzcKf6wa3bkIYLnAqxF5LhWnG+slvOyfkuCVwNsjMbQmu55jgTn9X5qC8
vWmkRCldvSWE9Etf9B8nObHExIFduBGR+5YE9FOqH6JhXZXTzvFYRTR8eTQHMpBXB8rll7lyV2+k
b0fPIeHLFwRaQtjkRmFDKUXyPlNQN4w535n8CK8Qz8vpWbC1bQEVihyXjQ2sLTZavriKuNBViyVs
uLS0t2EV4WicCY+T8Cai4nMUtFaOl3ljqoN4jT1Xeg5rHF/Ux6DE+vMzhJDx2g/1/R808CxYXw5s
yKWzLFVNjaMVzN30CsblivldoCVWbRhfYXO5rtTT3Ssu1XvYEET6I18vEk8rWSOPTNmG5i+JdNv7
c8Tk9GX/voCLDb0Hh/bL9GDECrSWGmfQOJNEZ5nQuNJJHwqHSIhXf5FofuMTIMAFVergUUGhvZzY
6LiOqSsbmaio6g2Ri3ROKPVU0pIrl9x8z9iIIiIGoZSHhRwvRvTNxotJMB9N/+j6dor1Ypk/KHiU
GoIWjTUBm8pDeJDrSCel51RjD0Y6VpEvxMq6xco1VXDi8RcV1CorCl2EBn7HOgqg2xxIXybxH58w
3seHGiUcsmnfcB0gvJ3fKoIbNsDHle7eXY/VbvlyddB7e9nAQj0YvjWeNh3cnYc7YaHt7VH+8Tes
7TD+XKiKDT/XV+9lhUFdLscCfuEbLvdoudTUF3+X/2ituoAdnUC0RvvMhNvy+Iun16EcRr2UzcbU
F077ETHpP/ne3tqYi0cXO3bNUBEXR1015e+SkZBHNHXhPCZU96dt0u2QD2W5Ka4NSAbyN7jx2/yc
uuffx8UeiubdVkUM99mDuW7ABZmyi6/eukS6F8mhr2fPXRPAp1TmKmhDVPGQh1u3Qs8xFT2lM1ZG
vksrxGXdnl18YrH4i/HuaBHHHekk2ld60g7Rr+lNnHcusoqyK+p+T83f2Y2bcZ+y3Dx4CCohXpH5
IjmKLEYb1G6ou1OtlUVKqGdRddvMBbtMnHsmbfWN4ksKFSw6IsyckJ9+E6eN5ZgiX7nPibmd7mv/
0MgurKHdGI41tTzpcGZoIvxpg9mYF3o4DVyDUktl+IbljMRLk+3ppQeYD2QlWXqAMbS5bpD7lTMe
27zp2YNd5gFDUEc/90VBw3UnbfgSSD3k62LDF6FF3GnBKT4mK2d2JV72JpBTQsCoaY5PqG2rjTUX
ySnsaKAOJNx87PD5+P/Q0kt82B3fbX79gaeFU+tAFh8sG5/YwXDgOwpwaKqP/85uxojGDXZ6v9kD
1t6QUt1JkNlmJWlDsr5SjEJTm712JnEWrIigPOBd/nUTSY8GwdOkphUDaPfZqe5H+DQed+iO+q1w
3KExhWEkMsJNymACGW2dQYFuCbqyjNnnPe2x94iPDei/0jhHmnwABwxSbIpdugn77Tjdu6rXg9dF
ky9I7UFSR3qW4GLtSNFEjCPsSgkPmC+uEFM5H3nmyoVOy0Lnkd6HarwkN+4QTKwBCnU7dIjFrZW+
ErNi4zDEtiLVOZuZcrPdIreZmwz58zc/MOOIm+1YOTyxh5bHzSNohfHimSPDl7uLH/ZPoRqaGJdn
wPLP/RRv+DezCZeA+Zu1kmQLSumoytpVo9eOc2Xy/SBPmVj0RqYyEgmSbNOdVKwnAR5m8nEIM00O
kBL09dezS0Gg1CpNyPPYbrZ0AH1vi+paF1iXTA823r/zf1unaPsuHPzM7Hk/6MEk5zmopRkO4Z77
51laFBr98b7eHXhfPy9yWH554G1dBZTVUJs9wIZo2P4UpJFrDoF9u6ghlmhsRVoB08rGi14qMdtU
VLnrL9bmq0o9jQ4m7Y7KKrNIfESxIX8c/JEJqI+UM+VvdCehHoPkyGeU5G+3WpB/NS96G3TSdndq
e+DRZtck8DpYoZvojZ/gNAvtTL3BwQyUg0fob8ZxT+2/06ODEh5cpDeaOxuKXzYx6SilzxBOdu1T
7wCMMGtS/ytwFW4j7HAU3XvfYZ+bTUsrGT/6jl3Lzguyue9/9rLRqmH68HfsZnQIxzT/3qTbvyKn
ZPjGDUCoBk2LGuMEkHQJ/EVFDPPc9u94kTFDnJFURtRLWuT9sWggXOuX4brbg7LKfWEXWtYeOevU
L3FVM7Xzzk3ccqxO9oV8Waw9VqXhRgaOGJ3D3/5M10gx5DAQDdyaZei9oQ8MjqsIgJD44UpOJJ1d
WWU22f4zYMVEgbRXyt5Ww0KH1H2+O0znZratURCrTQmnt2EoWwE+5H+WwDhwamyV8No5lRyCoDEO
vzmfta2JB4GODXKSBG63vgOITsNGxITbcFBP1IF+OmVPBDo5+k/+80YuJYg0bATF/VeSbCg/Yb5y
mtchNblEN/q+3SMRX0BqPZ7qMPsXp/hE3VRh1tq04FglzQOqp/v45iyFkSen/gMDiC0kWoQf018z
VSG4vdzg4kOA304IYG887BUvzA0gK8kZJupoSoHTCYT0tHg8rwingG3WA+FytjKK5FWYGy1J8iXj
wvMpa0vw+eO6Eys82PPxS3tPuF3X6/BViRfSCAADFpEgdl/mCBesdpJ07duGIK6F0//z/hfmJgad
zoU+4+0qiAMA4ruUqg6Wlhyyg5JIJOdj5awCRGcK/0gtBBaMdfXAn8E/4CJYbi99g8PZ4j0l5DHl
+5D2ab8vUGhozrGOgHZWS77rCBOYI4a891MOdy/fWY6HdpdCsF5k62RyVrTPlfooMsW6wo4BEoZI
AwHEvYa66loa2Ukc9ZD+/ZK96pLNXILNYrRpK1fi59GGXnXTkjvywGa+ce2fXlQvWMF9duYw1nVr
gsv6yjLy+3ARiTBhHzUBafnAkMEgN/r//yILQgyQfVwzsYYaBv/PvdJtrE9y/3RPBpZ4Avh7gOER
LJEodEsuQlxcqOrQx5m9cpYyehcD1nFfPLx9MGXWdb/7aW6hD6n2XUSoC0dPs90LfUcbCJtmmeZU
CHqPOGaIQnNWhjmsY70LycKVgCB1kyotznUysEIBIJG6hJbyRR/gn8yh247NB7/JsWO0Em5MzDD2
CZt32JLSfJV/6491xXu9roIeNEho1emky2uXb/m3lUjI3cvPl17Gm6C09Y6fnuY+l8RJ/JMTwufH
IFBHrjVUrJJ5tP57/AvSeLSkpPozdnCJAIQEPfEgjJ2JiL3EQegs9cPYuW0b7Z7Q657VD3KjLSy5
364hXxyiJjpyKozypp9LeaH9CPDVDzsv85cKt3zQQq9Q0Z3Hkc54DGQQKPEK6e5TI4JZj4zmNrDi
0TtDZUR9V0mcH5LZuIY4F1JxuO42mBbv/N/ofq6A/0v6f5NOitb2mWRWElwD3IqbiST+Ce5TggtK
Q4VahJl0UpE5ACQHP9QuGkJtWOELiKlJyxpgOo+28nRoGSK71zJ9Df/tZEbiWV0LHZvrIV8qyQSI
8omYEB5Lcaape0ve/lSJcjtjsU/rDDLRBcozwaqzh/XRGFHZ7VX3/u3Dhb5BNt+NZZV8MHh8dClh
vb7lxEkBkBP7Vgu2v0+djbA2BAkTSWDdKgDlWG6PvTW49OEj/s+aWJ3SFIFNPT5fTgt/W58PhbX8
4H4NGdxpWYnp1Y3vpRYf2z3sc35Xc19uHqb/kJSSg2SsJXxulowpuRt9Dvy7cHVqTPfFbAtM/2sR
ZjvutA9vkGCh1Pt19Us1UtqWgcl4+PozXwrgkKqU2QraIbsuYSouFpihkmRqUBUJi/QyGDveATVC
8iklSd3Q7bAh2L1WF9WDL4n2v2JsU2UTv73YYxfyZ9oXRrYfWOVLjL3bhxt9+ZL3dn/vG0bl9kWY
d+jFg9072t9N491WX0enV1zQtknj/EHGe32SPD1mttH4mylooRbAab3bu1SzgBRl3Jl2HVFYoGZI
qxLdEch+eZey9N9L63sqtg0LbpLuI888VejsnXZfDI2dfajEsrdpdCAO+zio4AQbCxRqVKk5AjCz
RDvjnCAnRZ1f6bbwAAUp3NaKA7DgpdJQzPOf2MnJVoerbKvMskXICTHEOoHKCyW3/4ttrc4cDx/T
W+L8Yl+3cVP7QRZvWFxjI9YFwRW27bKNxqzRuItit2cwpuaJVDEj5nuW16JEmI+iZlnP5Mjwk7Yv
VUZvd9VZskHXuuhZgc6JlzuF9zPnq1opd9q1XR+cO7SPgvq+RtJRXPEnH16RvW3E4NUlJzOkKBjI
wxpfw7vcF68H8h+G4qx7klSr/uBD8n+iiqFoNlkTlWHsIhQbjUgL0hlOynua6ybD5dv6TFz1wdIh
LJ/42OHDiEBWEEgcPFCtYMkN+uCIpyOIRvjztpyLA2Jk5nrJxz9Z97/ZjKcoZP9GwRVgfV2jsSCU
roGd/qKaKQeMO88Pf7dbK/ittBQ42DUvyuEjqW0d/VEKZiO9xlbe3U2CP3jpegYTkl8f+p+PwhLy
XBoj/lcI6K0Sl36gx+xJLbHUSsnY3cybE2PAMifpeKA8Re1kOyvOlnSym8BhRy15ldB6Xwf4/JsA
t0YXWGYTGMg6qzOfsbSGYPlnn4lW1ZPDJh6lNZowenRat2cOgtX87/Zu9xKidK7LAmjTSD+3O1+l
MVZ+EEARMJnLCb9AxBYQW4vECNtIBqpDlCnTMGJ4AIl/E5eCV8Hf+Rcy8C9hTuAGI/ydhUDDiZdT
rkU0mqapTrsIqlKWYIb2rL3jzpXfD+TR9xo0g8bjGxcYvgTy7utZgAv3IsyK829ZipvIFBeY58LI
AJRm1wBwJif3D9pdmyrliVqYgb3FVIcyoiBbayaJjY7Vnc+lzHh9CURiVQ81wUCAf8WBjR3CENGp
30LlJE5+/xFCuM0tK0Lcsvt8XYZBwe9CEkMFuA5tfLG27QHzaknMpbB9hwg/mto7I0XAwj3qKJTM
lQ4pmF5qcqanQULWUTQWSF2IpW0o/uytRsWUJaiUegn5u1hwOaOMtkPpmUNFbJ0n4K2zTBA3MVb/
gUVLYhuumeoogPGsvXtJvmiOEVtWpAAxASfJsqDtfAlyX1S6fLhU8QrZwTQIQWV2N143MCwdnYiD
8fgzftssP/ZMQfgCUNDkuUO2DRpuUQDsv/8T2KQd4nKyPiHq0Vbj515Zwl2qWh/6hTVxtSgU9W/X
XxWxkXTOQLbpP4lFiwNLi11gydfTT9XJks2guJfhnUD1weQpvb6D0qF5Nxj7zguoDNCr18snfyiN
N/rtBY6TOxSSUo2RoAkuBDXae486MeagEsCnrd626kJJYulX8gJWxncjQFPU+kdglnoLRhM1HqWk
zqErFFNY7P3OwnHTFPBnZ7P+GiCsfdpPVyLf23eTdTgDDrRElh4RroDs3PQs1UD0ZLrgY7hbt40c
MLzv+yIEfP9kYdr5RhT0xCOzZ7938B0AeeL4pzcB5M0wxNXhY2UNzBH+n9pMvg3x+c+07KfNjd4+
F7gv4vHY+QM+r5TV9dkkWFzwUnaeG+eyvQ9yA89Cj6rPnsNbQt6WoCmF0MKiNYvXQT42rvl8a3PN
2yqb0Qwzsf1PGFl5voQzzB77+QvlDNZSNkxYnC0aSW6aUK8GX3lOHLR5YK5UqX4k8pfV9ka7RL9t
EGDQBUjJ2QLdK9QxWjcN5xR3mRPeRsZj88qIqQAityzti48Cb+Lgb97grZS08q6Zk2f9CpfLa8D1
2wY+zu8O+MRysvZf9DYt9lj4riY+7PjvzBfv51Vwd5Ywi5cycyQkHRliT3bva/Ku2feAnZ+PwvIi
p610f/hGXoICzQ6irgrGN130DzETQvtRjGx/4GqJdsw+vxo7+c5w+hFyct/VLOgLEQCYWPjffZNF
7ewP5qtfgMyNtUaDduXr4qM53KXQxzabM8bJeTwhdViAnuiFIrgWEiUhhUs53cMhFH+dBSGgT7xC
Pu3A/baDn1PXQfzm1y4hIfuc2e49oyoPUlZRsy3ysrEpkIToHelTFzul4dvOpmj+NBq/jpfN94Hs
a2PYyrJBx11Rga31uwciSErdNHtnLTUdXNWqVIQthObIbYU1g5pO0Z9uWHDLi241WyL0b3LycMYR
xC681A+q/5IPVl4FFDwatCI1kDB9N85pAmzNDb6P4tNWS69awyqss23KXXGPnghCuS4anpUrckUl
Rc1hL50FguoMYciDAEQx33KoYiEQNUd4dtrV8bPLNzrqujSiV3/xd2rBKLjK0KHR5nCrZskS1aty
ryKg8vTtRpmwjTXnCfvgl2VgEF/4VcTVnKWmciZ8xyfMKLr/JQsyAnUfIimUv+ttQDQox/q0Wn1o
9Wg5d3OIlhSGhGO6b2TgD0Z+ZdfFzC6MIX/ZKMP62zyCXNfMtXQ/coBGgzEOX9Am0PQmyuIT8+3e
mygOkgyLDcFCEqBAbdgmpWa7hICVYqeo+x860wxPoYNuRrnbWy92KQqREr6ezlooC7wUbal91HE+
exOdyl5Bp3cmRRokm80BCYcqCEvweIW6SyZD4Qbqtm1rt8FyFhwyIhB1qLiLNteyekSZv4ObKrgY
vFZVAOoks8BX4xVCJUkJVom7OpIN8Uz+Pnd/1b8mYXj0+oszT/AWtnF+WhRr/iox7QdEnqfXA8Bh
xufWLaFegwEB/4DRDNfWVlGcV6QCP4bGL2/mH76LK0J/GrWpAAC7hVv5uoowFwcsPX3UptMu+ftV
zX+El8ClnGNZ/RO2yGANiaORYTllkcZg7vR87Nk+TVdEV+LSaPWx9Ov2VhqfoPhKsE3WdJWLRedP
vHnc9jTmyO5zDwPrKeVYFsYoTCZ6nLkcHaZUCtN1Lz76Z+xLf7MduCv2QNomQndBYOGwMXphaDs/
hyWRwHCyG4XD0HHks2E3iiyOLD7nRXKecR3JI/t1BDgDW18ZRk0tKOObkdNLUkdGPq9RkUjiHkgR
EH5pwRVAkL1jegVpGSSju3gd3AIVZZf/Rj0Xex0elVK7W4Jk/4FNPttTOKk8vilgZIC/brciQr2p
xrk6S/5rRDEe4MharkxBX1DCO0+FeNlROXmoUno8SDrg+brMJbEgq5JNrLAVMIGiG3uI1nH9pAeh
P1ZbXz+njQX9o3ATaihR1dJcYMdHOs0lKuAbKmgs4iQs2IoJm/sCwJgtH3OkN/yXveIaXEHKZSGQ
OyspN4uVu9xklAAMsL9No4zDbIAevmkjrD1jFDSlz5fvWwZnNe/4/5jvbIGgQ2JrVpXZykXzKIe6
4XAQn4pcjCc3Hn4FsWq2EaW8zypkdOIAeE7ZbjciSzl1ViuFVgr5OUsDX1/xrxI/qx6VfLxaja/W
xCaBg8AEsIUZLV7x3R6mOIWBaExbhR6XfEOpqSahr6WiJSFKC9JTY02Xr/4xEqqD5c60deEP7ZPQ
IjGklOWgk5voqYYMLvcbEBsDgkSkB5z7Nq1h/pMAWTYMBu1HL/i1HlWKEcXPZmpjt6IfbFO0f7y0
cJ0L4wvn/8gfAOTXdaCnVHTUiuhEElt8uaO5aB8L39ZLkuzU8HBa0DonKLd1Q0ldJigwmFzKFqe5
ZXhx73NOUqq65iqn4ICzEri4Wclo6fqhGjMij+fXLVbkqNTJX5kcMSYOKJwgzn2r7ey9w2X6xtQc
n/Je9pN2BPHaqawPxZnnm8WjgvqbnFkGq9qNj6tXMrREdTPejkKovyTK7aUNCu/y8gBrKxcpcN+Z
Je/FDNV1VF2Xl93uW/jviy8nEpzmYB0T3QHzldgc6q5zwV2h7J+0pPv73KtMe1a6Z5do8cFD/gY/
LxkSvwAMRyh1X4T7wuy/1I9cJZpPgs32hIfuBvM/1gKXZ2wbwq1qTb6ramnBLbd6P44brUmp31im
YUy1VIg9RcoVoC1zLs02zAFz87gqO43Zhh/4GJldY3ysNfhyL3uCH8UZOZx3UPScEjTZBdmLbhYh
ZlwOpgjZr5PkKYyzbdNbHeh+llMhStqTRs8g/VztM+l0wA/Bvq1tHp6bIquurFk8mW/Y8i+mIaF1
4nQE7QmOI+szhfh122wi59VXJPeo+YPRbWmPjMK3Ljn6ocbduOcLf/URx3eFZPYTMNFm6pk4UEQu
Wt9VkE0RTSfAAuWfpGxdP9+dpY2CZgjAEg+MEEe/j4+Fd5ZtQqFkJzPa2e+3F0QvR849M4CTEGdB
2+IrswAgavtvcMEZz1N/wGv1WtVniGXRuv+LtEx2WNnRCtxeJt8ErT0Z16kbBbm3CBabR8cc+IxG
FFPASV725i8apIb9rznSUuQCmk2O5nqNWNWXeH2wSLa9ApP4iwI2gDEfDd4UEWCDKbbm2m6hN0af
5VJhq6bXF9wHEBqGZ06tgW6yhSPPOVBu1ENTRSDBkSEJAIwoV3Z0SJK1DLl7rCUiYfJOz5Jl3uTp
FjNevbfL+bKvrqLBXtHKMdaWmaT2ZIKaqN4zVFQIBLYU+QefohNLiE1os2zEkVQOApqDcyTylVwn
MtV5moDaTFdu8975SfVRLEQJ2rNgFXN/ucO14iO2LwPpRU5jZ9oxDxtC4Bxu3E3HnsBJXCplHvwq
T1zENKiXcGqlHvyzXxGfzuSnu2OM1i43d955Q6eMrAtxBty5Y86v01crw+NtWv0qOhE0T7onGhfv
YCo2ZWVGjP4tCsQtnIhuG34HdegRuWcCJRJk1TkHvZ/5D5TF+0rprkzr02eiYlQRZNPWHx3ahFuE
4KkXFubsNm7c6Gudca8x0pzkcK7IaG3XhNpWUudiVQ+0KkLbnXARnxxE/oEY6ALhrSSDDewJ7GqY
QyqBjA+RJVMgQ5NPJq+WigHEpsVtf3xOFbnc8WAGRrLDrpOMLja/if9HxyYAWO4xC9PLL2Yp9SsW
nvnhHJXhmxGgLYZfyL4SIgwTDDJeUpNuGkf9OyxmatnxSkJJWlTpgbi+pfaq4OWsxXlblpscGCeo
CNWs4eMmxANZtbb+wkbEoBIA//8uacZQg9m0GSnsfGDlvhpOMGhmzLN9wyBrXKx6iF2nxWDBd8MJ
NUcrnAiuE+Bjuw54tI55dulS4FxtFEiK1vRxtbt1wXotx3Ei98aU1t9jSWbq+q6Va+nnsg2ScGTe
Ds7chafyqieBOYKxO5EyRl7+PnS/YLiZuW/7HvF0tWIK7i+AyY632CuATURzgtbTxKq45QRsovDk
dZpTWXgVqVnQA/2a36Iv7b6ajByYGmKG966stMf0cM5Kos1vTapV33fCM+S+0D+VmocUJp1Lorce
ComRZ0n3IKCKHCVuymupM6Kkej/szG3+He+xtjhoALNbL/16mTlHho37Fi+e0EuBCo2o6w5o2iMs
EJAnOZ/sx+2U1nkEeatcDDsQxL0Jdw/O7S2/4fRqUzlUqZRUz+9Jv2uLkNkzjyITmntMNjnX6d7L
AebS8/uK9D/sgHpya6vS71NFgadJRTrc3w0XUwnV/xaLY/FSfK95pmPfB6nCampizTX2pbHOP+ZP
H2wJf5TB+YOX5+Qe8qM2HbsXTDZghwg2djauyD0QUXaBDnKLzFFMWY6sGzB4lcAzaTIhwvMPHuA/
q0sxCznNauieie4+O9xNEGOAyxuKzHZEUOJrzVL8/vUVHRewexQ7GWftXgswMRJ0sO3nBM3PisRe
kEVA5M20zRZA9LswTZQVceiX3he6V4m8tZE3R2g7xuAb6U8ZPpMWt+mW1fl0+ZgO0FjRH6p5UYzm
Jf27nMTN5zzf2TqupXd39wJtFkT7aB1QIonTkZkGDH1vPnLUqrjsjD9vZRi1UhoPCV/jxEM0rJ1V
zqLmtWriy1md1I6urJEDK0VY51aRn9CNSLEnHSkfrbrInWULz4e/NG+id4y94VS/L0HJ+Tmsynu5
598vFZqMcarM9ZynjxS7LfTn1sy9dnpRi6SyFZSIYFyJ/m3tVmrX2MFPyg1bzZ/qV96lPVeqgpU5
avmggnmwbJHzG3DF8AeOdnQGCmss8SZysny2rzNkacfN2V5OiaHWYQuguEW+BDiDSnyGyOa9A/Pl
8O5akTPkNVsPQxnpjVeznwG5Q07CZl2I4BYpyvZukcMsN90FveLWscAKuKEKC0lA7XAdRm7gDacg
N9cI1vRJ6IxjaGLIFHWCbWx8Lh5EKbaAcO4N/qyQLBHCMOAzjkVPsT8iEBmqjxLL5KogAcy4P9wW
T8iVfxC4ov19IPr87ezyJPdMzkrpIGyBmGhLssxWmPPDkaonEouwpxu2Tf7rHxYgizrLyKU2961p
Bl8St0rdjn0oMGI3LFlJAFARkEeuuNXYeZcLic/45BqQ17ZXa3JSwiFCX8rjLZHqDodDH+rCqKX3
Ju84zBNIR3SJEW43iWXGYuKvCRL0hhTIwN7b38jaQ9qgD6Liza+jICt6+0CvHo3g0nWPHnIRJr/p
D+QTRic800q4f4Sp/n1aUVa8+5sPe/O8QS7xOxJv/fPMEhwooRuZZ/TPDhEz4mjzxVMQSDENO+KP
MeQYzCpa4DGrE8cfNvE1c43iQiwy0sBYi+JRXpgDGozx6URlU/PUfqVDYk4HRdQyOPSgEr+p59bS
RPWJVh8ZMWPQE0NAmAqlR75tDLfl6da0Z4b688jOCdCsWkYom/lXdkh2iZTyEeSk9VwbLdLx+8GP
Sa5tBxi8Ib+WW5NBPg5LrkEP3D6e93NtHtMz3y4ablErOuFyoL3s4Krb+fTAaDmRVrHbB9MyrLL1
M9BmyT+gJFtUy7EhgC5yBQxFo3We/DVGx8RbrxuleOMTY6TpTP65gelklxqjEXwP28lYVHHzvvsH
H5miZIf2UyOF4J5FAyFsO/crGZax4wG5zYTfRKCgBKfb4FNQdWSTZ2dmqtm3PXZhsOqbtZHN5pRr
LATzPAe9+gHWiZQj7S/RpEgBJ58MoxpxeUoe7ofCB6MUn9+11TsN5Oc07D2gfRyNzxVFR4LMCQNT
4VG8c5FtG/H+cd32K9nIu9u/ihvYChE+cKA0Mt7Rr+hUnqAKBLAtevRLqN4/Mz5c9/SDiW/cJgYe
Dw24sZGEEE93hWunZSjiJo8WVwa+Vm4Ed1EJDSHoNjplIRdmCzTZfXJXekPWoD9ggUXbxp+ZHpvs
rGzR8zlEcidCxHm9bgwW+nS8IG20VycAGpsyJKgvGP15BbRkl2O0M25v1f/G7PzTvIH0o4wRZI8G
oK5jRInExS7O9ILO9mKCnQRFHNIfcEQEArDocuufID339QvcR+5082SRDhkjDVPLLBKK9UsLlUtx
qBtXWh/OQqQxdHJp7TABP+Cuy+oiPAZArC1bqepjEEpzIKITbC/07nNf+vE8eQdn/xWfuqUuZqGT
jPOXLdTFROSD5ZIwZvTz+huB/FD6L/NFv83Ps+k1f+aa8/0Gy9vkqq5b13+qZLJf7S/3gkEdHs6r
RrtkqeSSKBsEFKdXbSOv4njlEi1eo/+2ZR3jUlbGbFPxCuxkahz9Il1WU+PtSlnmgHdPKNnXYhjj
3fOnvO302swMlsxLIUJCvp2c4iyJPXgEXOfo6I3jWA2apyPlekzSWT3XyIQ6gk3w4wZJGs2X4HSe
S235j+9em09GhXTUiMoklHpBAEqwbEIffwA/bmj788QGp33gBk7wQFr9QBVV0gf3On4dv5zN8XR0
wiOQPZ5X3rC/fHHxt71opNNJrVYJT6IwMW4oJ7ddGAsnETdVLNyzMRQJd4xkGRZ+8gXH2updFepN
2un+vaM4Ejj50T2VcT/LqUjEkvaI7/+nbbOXNLCPVB/C1i52wxCN5YK5WF8p0KnwqONshlsr7XQ9
SSs0ck7VswH39J6UqxNMOsVukNmjkt8Uqtj4SyfVBKYH/K+Ayk+FpTUodjBsZbA1tuii3WW3I3G/
DRq9fgbITPnEYa9fDeL9PeBMmB5XbMwHOZK7kOtLm7SPZhQOySjp/NoAK0ZZKLXplEtOhW60qAJy
FTbsy1s0GnK+pqSe080qlztofoSioMaH7XlaN/m3dklJnYFjJVMllM6jTl4if7aFryMlGArjAKE6
s0mV2kvbpUSbK6R4b4cMS6YcISLO6KC/VDP2i2hjH/hxKC0sVUZ33W7ccUcQWlZAbzFlAL4pOMyJ
i7F66p/YFy4eGmxG/N0Sjl3BL7bcP00C7Ir1IQkK+rqwZ3Oiell7mEAPNhncAXmJYwZewC8X60xI
/jkHaarGUaPSwp5M/lR1Oqyh32WBVQtuirRmgqPd9x5Ad2vA2MG2JMy/e+nQqEa0nmib+aWYXQns
oFSG7y3lcrbkykX7w6DUp5UWeBeZgXw5pKF05bFInPdwxsw/sZ5tUO3POInIj77ZSW4lKtqzzx6/
0l3mWoR5CrnsHuujduNs7/dslcn315Cw6vf+Hm+PoLvYVAzqH+s3gfvol/t/F0uT0/nTLmiESnur
7i+TtKWBAKuIW7/Iokoa4GBnx0dFgdqMHOGd4tY9KjCr6j3pY12V50uJ+WEilaXK9xOGlF6NR+1X
XHQgRC9z2wyt1OUr3jYYwL3xXyXcXv0UUwNeThGbeXx6butdjeWBHlT7QdeYj3fJbvG+wP4ggqfr
jOH3IQgWEeHNQILj5W5jPYbfPXMuVa/TG8gWjS69YdArgfypFXXzeRKWsPYNR9ryKNN4N+WtbcT8
3jiYdVYBQ07asNipgxgiL/oEwA4xiguJJgY+gHqS2PbnhsuQGWl+K1GbBXcLCsPwofbi6jBdp76F
XkBuawgeLYHIeGIuOpicjuoyycAQQDpRRwsm5MFhEBdlKqX5m7lVGkgxNzEMUnwmY0jKxFOlsIHI
xx+r6k3+cWPAgByitsekivhHQJqWMIEVVC99SbZuHCBRZi4c10GgKmBACunremKGO3Dw211VRtCN
tA9P8x9dy+NAvRjZdj/1Lj2+o+LkJ/n6A0u3eG8+YmdrF0oA87vrhJKvrAVD7KIBJNy5CeLGS9KQ
E+RLWtcwCFti1XsZdY3AvbCzxlD9v/v6JWzaCCAsL2tn0oQ686aMX62rIAIyCHyeoEarTOwYdzuw
Mt0+ieDpMyd8Fvfky1LB1NeoWogiNBXR0uUjSZS0+SvRkdR6srb6csvFPmNuGMOMf5W2d2n4vuKi
kPUGlsQ7AQfOOXFiuR1afPuFcW3eVbhMuJ/PogmBaONyULLTyNNBY1No9ml3tsUyX4gfU3DtUqrP
wALw20mzyKlyPoYMqlsCZ2tT1ueLVEenbD9OmQQa+foZoZeSPFdSk/a/TFIiiSlaMYmeKrzXkEpy
QwfyG4exEGAP5nOOxCB29E3xx9Ma2NqMgM74EwQLnRJg/3uLgTFki3QKWihBnqkF4k0yaAjmeO9r
HeNHegl/1tjN1MVVtdeRccfTSBjmCIx5lYapbm8UABD2nWujj4e6DhQ2F1+JQJxPF6wD/k/nEg4P
rS3b6Z9v4UPIaQtGmdIXSWjvzLSn3EPdZk+TNICte/ZHpU4j3Q3FN2XelhL2YqtYsFhPETNt35KC
BwM+/iTNloxWlSti7S5x+QELBtT6w7T9iaROkyhnhfXCaunWV+B/5liocQyOox+BdjngOxhg/bi+
3Y4UkFj7Tetm2kQEUiRQaZIZDi083Y1xIb4AajjWVX/b6naUe3jSpbzXgUDTqGQX3DEC4dXwK6Yq
cC/lPnsYdg3mae9n9A5wo1meFp/r7Q7R8D1Nn2e1O2hCfDXSdcwz9W3OBWVG7TM2Z4EpUgzjP3Cx
HXGzTN/bMOa9C4tFg8+zE9tcyJczqxA2GRdp04hZAla5caWVyKrGeXpzh6K17fxJvq1ERnH63Jbq
WE95JBEdrRfMTV9D28w3ExSRj5cG6ganGgZA1pXaPYU41wVBMtbyhvDl1mSC+4EPTdlnf0/AazUS
AzrKbhCBFZgyNpbw9PeO5y6GVOYkmYJNODnodAixDxpUPrOP1kfDZeasvP7obS9QufEFP9gGoX72
6/1JwyUfS6qasU3ZSeO143hdpBv7voRWS9E26T+mT3GIQNqVPX+x/5O0fhpp6QxbgkN06TK3c7Fj
YvDcFoxBlT2jljTBBTNoTxNi1D5xHms+o8IBKmU2tY/vZzWQuNO23Y0pR9LjfqJhkAFF1sYo2x3V
Sxv4GaFYqF4SZ3tSMg1m0MSt7+4aQMgb6SxRPWPWLQv8ggvVEiRyebM0UWmOw0GmTlTB6iB5otud
bGjVpuHysgGFENBE4i1J5DpF9HM1V6icH3lS9g4pNMKeN2AOqN8yEIXMckFKkbxS3JiZejXeSiDS
3oVI3qyWpVTCasT2DhxUMgYHdr828HdPjIrhNUT0AktHAxaMSVr2Pvv1HFwcwXRfRnNxTvppv5PF
1CGFBFIhKSedG9hadDP7avyU4aQm4V7Tpz5ZA/ATfwZhvYffMtSoEDuUocJdLzIfb85aYSzjTOI0
VD9C9yw5bOZxYOH9IRhxIcXvq2m2o4MFL4dK4y/ZzeSy3Y5YgT8vk9wE/wvk169r9aa8HwI0mGQU
vAm8tTrSZHqYY+RDrWg3QzArY9GG7KaYttrURnI4Hj9ESY8zrNwTYMceR4iDFanNQwRQWdDzGrqY
8rmQkJCoz2ZZZF/vGW72YU5PDiKEQxrSpPHWRnVjbI5SQI6H324a4e//NJ/tCr9kTwXIs+YNXYoa
+aMcHcxkmO4TNsPbBC+b0ZB7wauFjLUgV49ylBgNjXWGmwsc0jOsOaxrYcd3fLnR5nYLAbToKWxe
EWXgXd+9Znm7JgPGaB/e49zCFz/4Gm0tVsiffagIWZ4qXksQil+FyrbL7079fnZ+1M9Yv94+YojU
c1pVxK+nIDJUZRLqer3tEBbJ1WBLMgoS4NOlJjaGRyz7ofQsJZpld+XSuW5DY59J2j3MozaS994i
ieR6HjsuxCjnaYqrQqD6AAumOl82pwvlIgLH/nkSdVUoE1Rt6JHjRU9P0RCRVkDL/F5eLeuUfaHL
zNm0XxWVT2jKJO15kht4/G/Hppi3oId98kUu18KhwAtXmD3lOif5M4wjy/vvnlDjBGBsl7jc8pGW
jgYDNyBjspxC7uv2XtuDYM249I6QEkuLGFnin84lIyJM6xqnyTz2g7FWhIK55gw5UPWuvh/zPfXb
EBzzOMffn4OZazTz+tvGhX+BWflCojC2/otvSRQuSGxFtiTziR8x5jlDl/xzjE9KbBN01pW7E1en
XoBpnpexkh2fs5/l+Aq+3qIv7RnlHEwFwpXEnPmJItl5LVn59HruEs7W5AMaZ03Ys/9YqqATBqK2
oIbLC0JzFYqjiJ87l1mmitTG/n280EYFb/EmsVe0NHY9n14T3KFHXU5nUeytCvGoskrlP7SlVxln
giOUYqmMHIH6hhWzv912/d8tUrLWSPHEAFxEif9mTIxEjILlHYktjxQencH0qB28gjOQslDzcRzT
n/g4ECqm1yGyMYYKrMpT0/IN4p4gOpo5qr8YhPnjE7GaRoQT7w0JvwMP+JemAJVfHbBMwym7A8CO
btP9kfR6VRKmpAqDg+aYqD0Xaw901pTsgI1HHLEpWzDl5jPL2y9jHoU1uehBtewTOMZPHmeOcfUb
dheOSCG+EathHA8Qqy+OGogf3MN8xVSMidMzbdeSxZF9EMEycHKIVlDvt221lE4EWS8CXpsncPZd
0Dk4k0UwaoFookshm5JzzpuIr1MWSwLm79YMD5icZ5tojThbkwWijCxzmUIAmZBNkUWlBfwCuf15
BPVCipF1dxZaY1rj3gIpOdmiYvYDUjZPekvv0dLYevInJU/EJHeyjhwyFeXIFiUTF+XPauhAPyDp
RpSNkx/NSzwrn5AbrFrdpKhO+XEbytzjahR/XodKsUaQKpoqTrgsI5r42sH99DTTOgNALGRn005J
caJddUAxX1oo8GKINpVcXxxTjjtDEj1IWjlVwvoLU08jF9LVXt04YiSMGTMJx3MXs02u/0a/9gdj
g/Xqbpti8eL2SNPDzbJdZYxFGxXMGLFiEUurN3/PEaogh6hIhJxhicny4XZQdDxDyCtqivD3x/L7
Ssy4uF0dYeWMXJXwMmfwV66CVJF5m/P9P4hEfdTsVopeGC/OOVUBhlmaCz47HCyTTn4Q/d1GKeAU
pwp+SCts7/RF8zBJuUAZ7gqc5VDJjOXowjTABiv8Hl8iLkOZ3oN2ctk3idOpHUFbb4gJIljFNt4U
H/P19fj2U/s4HG+xnSF6DjO6kVD3h6btexmkTEAri5a7cjJ6BgNd0jtkNNTqYBpQmc0rfdDp3h9n
1BQv6f4KFXnNznh/JiFzq+uhDDexXBYu2RpJmuhiRvWqogdTqVQMWRT2h4k/djj+4spSjcYDZG3J
dYxGYS9aWqjEoi+0n2BxeKcdDHgjM9HNAoqWZLZLvJMPnPDCBYXrghaJubN7AGC4BTri2dYQQp5m
NLSXfbxbSn6VqfxUjohFGjEPk/0AoaWnDGqDbRmF+qtOINdZxBXyRZrPJmj3OCxHJMeJ6ikrjg/P
fjeGXhy4hU6XCApr4s+fwnyDY8QDyGXa/wLWgXByC2NpdI2TWEcZ37KIfGVEJc7xodC2atxfZ/Ua
29f5UuWf4CsxJh3ZTWN1kdL01Ps4FearzUEp5N53VN8iVJr1vvR9GnVS1Z2vakcNIj4VaDwWpSMF
fibCXq0E9fxeUQw7j2cfrwihq+ByawsxI3/2coFCjHsHmsQz9e4FUNqho1BxYs/ZVM8f7FQwLuAT
sxWzDhLa0gnEI/ChHFjUI1b8+ireIvzwQe9UlKh6nS4ZY2CJ+EWfpKR7rI08KMJb825NXZi2ziM4
nNT2rO6DGHW/6yrf2pUn42P22RVvJ3nmxSNj1q8P323lvLvK1SkWHoF87/TADmybkZcTkg70ySt2
HcBC1F1w8an+o9OEYTCWaKYRYqLkppaskbOQFcKhnHgteYKSacsic+xrnj2CcVDzcwZ2jQsHUAFE
puIJ2fZBFi4p3yMTxw05o2QPS5z+dibEKsLzIdBgudjGSxxvMwglJppw+ZX4e0zrzOSN6v8WvGY6
JH8DuSb1fCpCl6h+DQquKy9Cantfc/srNhbILmoR8ypLnYuOQAxV5AnPRPV0nFIlkFMO4M5ua0wo
QOslDFlONz3hF1CTt5xaIksOZcCM+C4lgNSbWNz0Z+bdXqLVKb6/K19aj9jqGVbf05xt4BDTEliU
73CxoA2+o80bjzOTxc9Jhvbs6ZJfkqSsUbzBWtPfmsYBUJZF0PLMj22e0MHlt2eoRBZszvXwiTfg
XlbT1eUlg4VBL/S+A0hk6+0injXPudBK23uPFrDT3PjHKLQL4pndfP5CPE10V7SoW7yrZLNuUmOi
qaBWOndYbYcycJhlLi4n2jm6DhtVLH2T7B9PPtJSdkkrfSal6Lid4Uv3Dh9XNsRBf11jOScIZOdJ
pjwYoI+TtJ9UnQRCx4SN3cKauPbkqeeiR8lOnWEFkdUnh7bSh5tg7oxsHADoaTfaWPTPmbIRMUQq
NtT+RPnTuOEUDz2a4VheCftgxF/xsXEubrwTAoizKqtVJmGrh9wwuO7POITy+4C6eNSm8CyXmuLI
XRJBeHttzYmCaEBtgr0CbcJT15QVYnt/NMivzBJHBjphUCNwqRLHNHUzDboVJfct11rP/Y7ZO7ss
nY/7gxjVKYTrFz8czKxXOrR8mVG6++bx6DuCcgtP1w1u/KOhxliKHHxNKZ8lrxl4p4LxCRpmeio5
VAI3vxu2YZY+15BgHHzrcMUUVNICvCy/yL+YAExDeeoxz6kD4m2apthlL9PyfR9lAjOQL594IWy7
pgnmq0rSP7vCYd1QFd+7rvYYLhdDbnbBhUW2EoiK2tqL6wXLPcHfU9CU1jTjEYa210tFr1Kdjtry
IXGudo6qbO0D6WOtwMY8R3FBUlFe+hiI1bVeqBYpHj/Ja6A/h3BjZI3zTWUdodiFg3x0xOqQ12Zf
gmlyfX4VbTWlfptEb7X6SeUAJXtNchCALVwofVYTVwtXlMVu2+TgM2Aymbzu8IQcPQQTeRmvEPv5
TQUJCyJqSUv+PL6CWYTCd1xYoIJp07jhE2B5GVRd/58wfv6+6w4pNYcewwuivBL2GT9OnUTFzTJg
cHu7V6mdu2hNbnwmwAez8yKNRcoIYFKngEN3LmU8CiPwtgs+hiFxXe1lexLuajV4RGRfHoBFBrFp
/hvQdPu53rJWAMCiemQ8KIzdnuGxmv9QLrzjJyPQOOHlfEPSOWuoTZpNQMXEYO5BQdSH2RQENRL6
yoDs9o1v5IO+ch4CaqDzV3HqsHrxf4bYhNQRTTzwFAwhhpk3CUsM+rUudgtpfFy5uq9/JcgBiaeo
p5ps61q30Y7Ec4yO5vIxgtHDKFTtPzhI1GfwUbuAqxQAm9nVwi3wFeJqBYM0Dm3gQhbQNmQh6/S1
yMWaGdmzMv6puWlzmNXqHzXVcJwWbenKIthOsYithIhswKvCrzbtlQlSNHKCCc9WR+n5RCSxEGVZ
JK6Hpdf/K/DwBxGqLiLoUPH81Vi8r/7lXWIWZpdyA1FwxU/H73b9EuqZ466eW5SI5pBrnboNBwdT
lA2tnktb7t4cgT7GEzOJsyBzEVGabq+rhOJH9OzLcEH0lEgjSLiv5IPCFQfW834rLgNPZkB533xH
4uSe9/M3oY31QTdWygbNle084qAbiT4h0q5lvGJGEpoxO8GdOh+Y0vXnVWju3En+Ni2N/9HQhUHR
ZeYD6UIMFWOnzQI6E0oSinyJuMDRjA4Tb0qk7JgvXF5xu4GyaoI8YY0ywPd2ulYGGSTKgDS5nc71
kLjOxrPnaCY1BVrlGcTaXQLEtCVH/EW7R52aBRo5T3ondpEspStHMzUIVz9isbAkNkVEOzpJttqL
2KYaC2/E3CGrSmx4NL7fztIOf9gcMEXfev/LyEc4m9f7FKNeCRFKm7hyC7faU/llG8m/LW4zXnSb
mNXJbMmvWAjJgjGpsyiqfOy6pLWg9LhzRinCr2mr3kkqe9hkvmVBllpYTcnnfzT73l+TPRFdP2FU
eibXhctVYKXuUXZvLlKlxGYWHbCU8Uv1k+y1NhdUEtbDPGhGHxNWclGkAd9LuKd9wcq6PoCmZ01O
cbERWgNBWC6c2T7yHYjBUL2EftPOJZCb3HBen/3npxe80+qhzVvJp5dzccpFMmMe2vXpcBkCbUU+
dXv2FnBeqPJ4AvPvMljb7gATX9biW1CiY6HXsQhN6Of9JPG+yttK4Y0gmX4TzWhZA6OCGmrknMQi
93kqUz7e1sdhE9gyQNa6M3EFCFijQo0/i5t0s3lFoD4BvV/Oi81gB4mCO76mIuE7DghkC2wHe3lR
OWOFTNA93lQ/AMbTOdbGJQ0+PzyWBA3xtxpgQgzaSdESTaPgJmPyzFkexyKvuzVnem09HN2hUEIY
qwyzzYvdGkxW18yLoW8cgcpjc9WZOGTumFJQxw/UeIuiJN4rRVbCtjxlAW02TR5JjdLs3Vtoi7no
aS7iShR3/iMYUGgfg+pihRWceDLJgdWyEQsQOMR6r0SBG3aj+mmbcHggqdnjlOAiouUIpIegRC0O
cA5Jp13uSA4cgAW+KGAei8EG8wHWA9jbTaJzkPbNcZ8lYtFSN0m8smq01bEpcHX1c3BXnwYW57mr
l3xfLabMTkRYt8uIlyWDIjtWchmWKf7KdHk7HxFACBRC3TQh/wFjbvl+BzVGlu95R4cdPkJE+xqa
Rv0beYGDKAxsUqssMORaKbhMix1WcEdLSzvbaNZ81rTjAkR823VtNWhq9pjCjhDQI+COHgLpTg3h
ljVyLcmtS9GDr2DLtHZ0z95rAUqjWvn9Uwewn9AioQfxz/QvYZMjTixqSapoGFZXTRweoddNdgZW
wzE3tzCxrytIKZuZhI6JMblciXLUD4eFbBau4bV5aaKn4v+xf3ILp6mrK+PD98iJVKU5UkdQSN98
Y+e4kh0VcC8aa7ZVkK+p26vuYfF01nZVzYoGwoUqsoPpjRAa3yJb71Nt+7U+m0aIl/7qt4ZeTK/u
HlBHYwTPg+rz+lP7ebeBXxIZZoD3E4BCyG0WxwWZqHb+rFh3nm05jKI5Ggg3zBF7fzrrxF6tGVsA
yo4U//Ddd4zDIs0/m2gmJH5ZFJlNFCumO6R7U5m7dtaePyOWqxd48FOVPjvx85fVzdTZJZ3bI55h
8dSmQEbbNLr5ClTJETzLKYZi+QcINDSgLLFQan/o4WOyfYpMgHBxaSGMtCWDRdw3TC0EKjlnSC5O
gZouITJ5LXG8jqQopf1P34CWF+mB6z5utsVru1DDrFm2zpyJ+H5eXBmifCd8UrIMaNdyN7L2gLVZ
esjoVG5FlSak1hDDB1GqcsA3hFd3ifiKNMJr1BgUZ6UxWfSsjYyBZSNT7zX+wqB23jlQ+rOFZtpg
46GzvZFzX9H07aX5R+Srbhc/gds3hgyzC2hiJM59OuOwgYbV9Cmm3xkhWxd2cOlsev+TFPOFW63T
E0DyMWEu2gXSIo+Q2LaFb454RW3vhFhu7wXMjCfnSHsfDdSJ7SlkpZZg0YNv9JgGXzK1nkZhAzJ0
O3WtECoLbU0WPNnRqQ9zZ2wchO9/DGsdIfNGB2pVULRpXJ2QtoSdd4g2En5/DaACvemfNaJk547/
pU4WRGiIyPOV4PihO2Z6ZUuX01wgibvqKAuCIzuanYANvO4yrlXoUAdh6f4VPEAgNEh7v+o0LydR
p89ouPyjOFg6tr/WD3+D7rNlXcuFV2ujICqdMTNClpH+I9EjYDO/Vfwnok3Thg58/v8E3TlgoJm3
Zfcht/R6Ax1wWgfSlS4ZO7t2h69NLF1ITeZ5M5q6EtiYEkuuiDQ2PoezkxvQ54Ya9x//o5W8rech
SJmiqA2DLIgnzq6mKmYI9EY3zrpJSXD/5dCoSfRV3EiYYvd/1XDHe3haAWV1cgTyz/f6N5T+IGsB
pPQQStXJQZrNJ7Ay9Pi6Whk//fbB2nzsQUtwqUhXqyHvKLRKwKBImXXUSLk7FUdl6Wts3FA34mVG
utCbLsP2tD6EzEJNxNs4vBMcVThHPZDekPB7eMiMhlNf12mPAeZbynhaVcGfzVULC8hoHb4nAPiQ
bpaGpBG5eQLtDkPR7jJ9gujLQYVdYIVhDiBp0vpmj9kvp2aPpoZtLRrRvyGprom5hF6u8fLS8mHr
QpkgkDZzmhIyxBg2/XHFYFlf3E/jTK9IDA0LKhRgO9sfIvqBX1V/FK37v7bVaf6oZsNdKQlA78cN
mAqCdxkblbbKsfUN7o39MUla8eHxTn/s0ytzRKbl4TlkTEHxNcFzLV94C0VlO/KnUt/ZSZR+cVDN
5XprjmNPdlu8C0++yv+b1o8FtOMvvFL0Y+E6Yg+x/FqRlyA6AUTw6peAsaW3XXvUGyXdArhn1yg8
wB65srR64LcRjtQjTzFm45hYO9P2YrkXLwhD4gydV1/46Dweqxr7FSrOghCnjj45qL8LxkjX6nR5
J7mJ/fFs/fGYOXlpNKRq03+j2OAeYz8wPCJQ4UsbsgdM4yM4mkqrtBVOQ5ZZmwN2osfbhwg0168w
e2kkqUggPVcCReAJKNwFBJ/1bMPjEYe9ZOkOlO9zRSdYRYNEPFCcODFCX9lZlaVO6/ccK2VFCM/g
kgy4f7Ogpy99qwxYE4Im8XsIvOmeR0jWAutO5LqNnPBS1MTHQwN5WYdjd3SzgOTzAC76JEXh1NQO
J/IjmWC/07MUQUFA0jr0GDJtpy3L9ZQhNzLfy4LAjsXtdzGyAe3aHvZvqrBaBVtwydcQa9N+uuXy
zKzzqlajyVUhwyFEUiXxS2N2rbkhlD6T7NXDuJnh+yi0OM+Y/ze+dSuL12Sc6jcQ5vb6MCUgqMR4
U+4CPvxZ97ELoEf9gbR9qpMadGIPKKoI/FDUINAeaIZCwULYPzq+PFbSgnK1W0ORQFdFO/Z16WFG
ObaDyQwwNB2Mqm/kIzLKyAweM5pJOfHr3ZfYB9WKOEerZY7rPVzDqDM5AGVg/nsuv4d/MVHfqb/c
qZ2+AIvUSTIJ1pe8ZZ1QHme808zBtX62pVXCxhSTRiUlKSJmkgfqVnDBhZ93QWvQKEUdCbPWv/K8
ngRCBFj8fLz74H29V21SteZHvnaEEtpUdFbw8WbS9SgF0LP5RrBsUrWRqxKnNeW8CA8f1h5gI4ww
LnA0eOgMuX4L/2U89QvOqltLlSXIC+lXU47iJO6R35wEV3mMbN4DfYKnOXa/73Nrr4IvcF3UQ/hM
IL882FgjjZqs1ssAk0wl14sx2xm5m0dIx4OIar0Tte9YjRHvJcNJcxS1hOmCKNMq4+n9ut7MGjAY
/I4OHjUVJLjEawcioxXJh/zUuqrqIHSCfs94Nwh/77+DNPsFEwNLBN54ObO+mS7gDQU8QuiNE1mA
ut5SHO/EzlaZHqfTt3LRNSOOCN4v8BLFT8q+rQQ7iXhSFmI9hjFiiXMe23KsBeLMOmKNswFoyhwE
Bo/5lVR9KUB3VsX8I4oFmra38IS7/YknBcqlPI8LaMb9eaVKdx8Xdu+ZoItAqw+e8u70o76uExSN
ZNnVOLAsKlaYk5wLHjxcgi7p29lL5Dzr5utfov5HAefompE6S6S+g7lEMitbLfaf4r4MF5zPDoAh
sgiHc0A/CcD7VPyPVyEK9J7w7u+qhLw+vlynUBrz4Y/ef5RYmepRqH8km6+qNw6G7yj+vspj5xSR
PAJOT92OHwr7/HGiUt83qaka8WG7EAtkV3+7UR46jOnhF7Ch6JsOGdYQEnYKIXYmMBIyc73wQwwI
LuIzXGWJOCuRI6KeYRwB/JvM/8wThqNtkLzZA3CEs4Ret7yP1iUy/Ob72tKFYyGW6205EL3368fR
gsFFmFDhc5ASgkKolo7Uo2U1NeQb45pHL+6oL9qWqZR3VFS71Nl/s5blh7FnI0gUefNsKaEYcwpk
/ODsEHidyBH7QQAe6X/gFRCCK/iFi0h58xrcWWEm+GNMt27S4gF5GUTe959WnFv73tEhZ9YOnidh
JhFpyMlcE+2Y1NdGaNUTIYVytaAPaR7Nx+cdd2kY3V09rK/xvc6zYDQy5U8XmpPktQP7FkqZu1Q2
Tyn1KGnHh1kXzwXcGZ1VdpmfJEbruSRifKhPK3DhTH48KREGw9XPIL9bL5Kki8QRBx0+idwnE0b9
CARjlB1Ckfem3/CT/O/67tCAZm7iuhiBElVo1DYDaVNbSJbLr2x7hVqBTULDjejnyO6MHwH4B05z
ymwmh9cQ5dAjpVxJpA9DxFpu1GFG6YWGUYugBxScIhbP2qQrDf0sS/m2HY7KCD2AfNs919shxFg2
STxlP/fL2LHkuU4EzNU4E9NL9qFc7aggcjxQTSkTSKwEXPpNAQrW7hZEwTXy7YHshfRN+hNGwzJu
UTAldg5TgXuSS7bNjAgGnLmsNaV21/KKjXVvAl2HlGo1r4Z8P+tfb/bGwyALVoS0rZ6ATKmzofGK
9OQ5PQ+mlScsgOVD9Zlo5jDsyCdvpQzXtQFDj9PMz4pTauGHA7zzFHoU2rKreRIStN2ceOnFsUws
oBHGpUmzKMUvNpzKm02s6GrtwkCZ72qZ7l4Q6SBCRJ8CJ1YsI7S4Onex3YcHbNgqo3QzD6zbmGAh
71EdbgVaD8X4voCvPCtCVTnaVmVSfG0DlbYQo/exsT1+IxJR0YvvE0jevoZje7Mlyjgzc25ULNsm
fOLvtGg8eig8gPI7m6rRn8wkdsq5aZ3ppdzuuLPgsh/6/nsaz91zM+nqCmVQePN7Dppnpfhiltvo
ndlVeFcr1ELkiyy5SXq5Zvr6jBKjB0Tznryeq6qXNHfOeLFBjE2dJ8kaKnuVklng6ue/O0ffDqgn
NyD1qN/2SHBIbrCoPD+NVfHVco+t614aobXii4F8Al1yHcreSm2wwL5r78qYplgdTcTSixxTJJ/T
fHgFOcBq/1LsS60KJwRNXSQpCbJXL22UiG3WC5VfAGGCIP6TRP0w+Oczfoz21NBWZiY6aF3T5ua1
DhWsntpw/PJcSqyIj/UMTm9Rf8OMeERgCNZPxo6Bh0PJoMI2BW98jdTZml6G0eRnRzgbwpYjB6ba
Dqrbn4vd0GAbEHN6XeSYBlxZ3VJZMF7fzJbxkym3yjHOAzZOTdiVqx9Ci6YBhabX2mHuNmNyHJkV
hoh2P96V3lcYUMaLtuoU01YGICSotU7jXa3ZyOd3I+gYQ7WUcYDDEjHNwajMQJxftPfCmA0Y8ouA
BqNQ5ji0VHdG+3K9uoHrsJCs5suzynxqmyZxGAIGaAVMr9yKQm/JYbkNin5UHOLIinmFfEjNcJ10
bcA54IntTB6Wrafo0NieCGwyScUFt6n0OZp6WPc5OyJm692YnnOiag9lAlKVWhsqU1hZtM8MeVVh
opAFnP0IXnVKvopECH34dGIIZLDUZSihSfwxIJF/o8SmDg6CBcfdTgcH6MfT7Gzm6puGoJoS2tcv
f1LfmLfwwAuv75/afdgWGKPlbJVWqdzNCfDPBGs6PIfUvDB1pr+8dodd4ggbdd7Rif9Qe3hzoMLp
jfWXnVFjw1zv9ahOGRjSk+uFLvNFMb9kWle6hQ2IeXKMh0MhLz+cuddWTZS93FnHzQgReheq7gKS
pg20eKanEhPyRx1ZwrkS1QnyHAYoFUG4C5pXLFuqUM+BcjBxifM9oKSO9Pv4TONiNbt5PB2/HvyA
qfHkupCPFp4IQ0Xf8UUkZ/4O/Y8AfHLnCxUvQ0QZbTljGjUf1j8EttVDASWB9XNaclkZFNenZTPx
IWr0IgiDWxOFVcRCakrTCBq2+OAOWxzkxJx9nqdRvw8ZUHB7WBzhr2JLYkkJyOujgle4dwmcqEpa
OQXAZPJqnVZ0APy00R9Iph1v+dKjztqTmHRADPD84NUxR6kcf7n77WywP6S2RnF13HZjsE3xs+MW
HkKWoV0WfX2glIVrjre0zECdRmUuXJoWLQUqHTzgUvdgWvzqCiuvyNxXW3cHicNkOmyaQVTjHJ8q
/y0WBYhVtvJZBCsOH/OoY6A5TyFyx8UD82mXeptsXbj6Sp6ptEk1tE/RfZ6bTtt0Dh21828BnQsh
bFNO8YykX8ZqDaw6ezr49q1KOJqmTsV2IIAb0oLkuzqeV00uX9i4p0dWT7PP7iDxHvpluGYoX7In
kKixQNc2b9GWlwO+jcnQISseNowGS6lvQXHRNyD1R957hz158wra87zzusAvwK0Ppd/Jbd0gGKpN
k5SKYn+ghlBt39GFU/pKkoWnR1A9TmUS5HdZv9mJ+P/9mR8pPiKAYNYkT5ClNXe6FzbBda1yAEmm
U48i9LAstr2b0XzNhNo8KC8wo6F80iqh6KjgX6Um2HYy8dmkZ10ufXRk8B4vfO1iLA93WVAEKaCk
IpsTK1Mp7O5aueobEM6Gk/sPv1LIMJI4OPLTxoat3ECOGTlgnrjeAkbWnYSS+J5wDt4vfSTBmXuC
LC0G036yqNo7K8+AGs/l9tRqdGskPvaoT9fc02H6EcMh8viUzB8agZQfVOrAizaKfRS2ipphRpoB
MGHD8iYpZorvLcPxTsPqHPhPdYdvhHjf2C73C5xrP0/bHCHkWj+YpdI5ta8e3+C3wvi7cRNK9dwo
jM/UFT2sQriHw24+M6L9SYQ82EOXVAXKb0wAAcTJYmwTtAcSJjpVfgBGOgzArTLDw5Ki8q3bi/Q7
QgiC7cXDEa8F3SZHwR1FPClY75XJ5AxHfDgiYDOpIrBj69a7Hu0uIXQpXiEzlnk3uY/Uh6G5mrlh
GMeY1ehtecJ9+k2mUX975AQqSFruUX82xYGvbxVmCFdDe5MOyN4NCcI7lfdrZBR2TUcabnELVoSS
td6MfxLlbsexu7MPPqKCqIh4BWl0TxW/yHpfhM+NFrhMYouZTzoZYoW+L4WXbwGChbkd3uCXsF8y
xt/tk7I8E91GX3u1otMglyEjaflyoSGqMkD/02D3h9em2/aDFPx9wjHfmrFKHn+wVSgi3XqfDdMq
WeEHfKAp0lI6W20kbkwN+mJidQTfaeeaEwnCcGgd7i8fCJu+pUf+cOWQEj0pYa09Z04hz2Up6h6I
2C/rkH+f4G2M3CMYZgATQ367y6/VmBwTY2gUK6E4uIpBfAHoOyE4mBJvxeJQR4hrKSJ3LGkYb7Je
D97EySFr/l/4KBncok9Y0PN3HqXrv2KiqitaoMI8EaLEzlXci+yWxqT1uYNTYbmG5rOyeTLzex3g
psmDm8ldFaEpuljbiGq4ie3DgeLIQmFtIBzLThC9QRwaib5WHrLXBZuI6qXhuaTK+r9E9QiYMfFr
2vNMiUWuhQiH6Fk1zk83UIpmD1TDeZrArlfChcyMJlHsLdNmFu0uBffC/B+Rxxr87JLnVr1iSV7U
vgPRCitUCGAqYvEGxldDssHzOe4LYWPPqc5AOr+6KjseOyygBETi7aTkbVTWBRS+KmHhOMKEbYg7
iGKc9d5vjJOtdShf0rUuoJIsn0pwOw6KHFFTvI1nvMuy1Vv7rDpP3ylS3P3QF6hZxL2Kn9VSdCro
g/+H53YhKVSpKT9UUVvgvYQEIjfLOufbPtf8hjoR8VQrDRyf8Ws1WELIduKOKXHyAaHb5WUmvGPW
iF1r6jIi5+98DNnt23+f2JkpEJ/Glv/hTCJ+US4wIZ9uq+Bw3PA9n8cUPhMF82kwjHPdFypeH5F4
QqJ1WrwGciS1pgQBlM2CRTb1oIZj3hvsB2ZSdb29b7CMxRz+laL//xLzQH3t4NamdfbpaGI8RVm/
SMAT8WUdM7auEO082pkLD9m9ZOTmCJfzKX2F7uoHLZli6ua3luTNLOIq5LgqZ8oxreLJ6cvZsAu+
yorT63FZTmKeTpuphbBUuo2JEIuncGtqGVvaXHKC8DMFcd2NUunejBMXZAEZqMj9/qIKVCllWOlP
bBg7yn8I9+gu6JBSPdDewWd9t/CZsnbIJNwSciC1CxEWWefmEcf8CwZvCJBOobZDeVkHqXReKdJM
8XrIKd+gQ+Kv9Qqg1ITYIJ5IAycxshb01K8HEGZyneGuKt35yXGhzoERZciijt2Jlu0m07myBwAp
h9gr8t910fUSWsU/BCTU4SrXfZAVzIR8fKs3HgNukEvqHYLUNS7WoY0hBX5pUDVxZhws2YnRlJn3
HZn5kMmLvdvIxlA5dyp4SkcXC+cRsxeHyZ1hxR7ESTUWWatLJJW7K3ES3EEWFlj0iyK4RuhDCwkG
eBpCnsEKhTxHqCR2lmHIEJFEAO63dzIMXZQfVg9XCxTPLKElZyzuf91aOOB9QpuR4um7f8JBdot3
KQ0ZE0/PvGE9mQU7Tx1TX9QNiO9zzHg9jfEeyDhCh2rp028q3rn9zc9KelxUjzGbj5NjQsRNRLlg
fFM/WN8LiryuiI/Q2J/5ra6padwj28wBA2xGrT+V5m3EdJkOv664823TTRBmZojX9FEWWgfHUhcE
WzNMfub7JtaPHEYmeQooT5NA3CUngBP4Yr4DGAw8flC7B5E/stpUbGPW4XQyrF6pjD/YNEEaD1Yq
aY5knVTSCQ1Ol1ERv9pSX8zTtVGqBUDtbjyXlgUCQtHfpHlakKozoM6vKJt8uK4DA+Dzy54cQXKE
OEVXcIoyUT2053GRGIW5orTgIX+dXZKniViZUK/UVi6kiE/SrD4dnGSaG71+6iiWp942WUYie0BX
e3gZ/oNKQ2jUVwlMniZHL5lnGtDna3ZKejK90OaPBjmFUSvAnMPPY/s9MSYzWjecCsXEMijNX52s
CoW45iESVcMY6uLVZtEpKQNmUEZd1cBBRS/6SbNxrTl05Si0IHBOqY4iwadW3WzvCMuZVx1Lr08n
yUm5rmZkFI+RaBpeKrFiBHHnAFxlRxrQ8/8ffAeaZ9H/g/G8A8r9sLPNprhGVihrWQ3Ww5IJ8c57
DAwJa3OvCW52OMBXKE09KQkzd2ZvBI6o1HqN4jwBwmrfwSnJ78g31pWJeJr4F25St1CmLFC35To/
Ty0KdBET08rt069LRxdd0W/RBnOlE1ujGdJe9vXxc6WryFJfgn1hpGSGcJonovZdp9etXx/imIz5
M+Grl8c2U/Z24C9pKz0SIDlgIDrFLjXnuLTcxgN6VUeanL7IcUPFa1QLxf9Ih/jPK4QXQGIW70qv
Ib/guSv1mzW6u7eRyRJFkMf3PuA8HMTmMt54dpOfF0j4rfPY1HBWRbDzYluQ7xurjyRHqdjR1GZE
DUOsKykct1tWmttt/BibEfO6Uueiu/gOak8t6ERI/pSj7X59gGpx6ldM+MiIPqvPtS4V5q8Hb1H6
NBDpLicfrJNg4jnp9nLZmkbbIi/NyZnCt1K5ScdX5lCPrmE4IKl+31+BwKUUYL8M6bgUslvvTONc
Tm4nqtUnpKrWpV+QtXMQvBvqt6GauFyxVpcrmx/EAQPONn/Me+GaZnEPEKiVLNZi89p/56DaqVl8
76foP5CdepXgO5Eb87w22HCEh5ewEVVoXUMTvN6EiaYdapFakRuYxKbyxb3o5/Di8U6tQc+4kIiM
P+EeK7tfqGIhfDljAD6uztgHW4ApAJfePGmRLCMWrML8wUriIIo5RMRdzPyGrl/sH51nu4ErENma
BdJI/nux10GkqeT6OAho7Rw8abZvMHLVoTl1ZTdJ+ttHrVmcYLYHCsdOUm0J+wlCmEOyZm1o34Dq
kqrlNWQfoHzRzFyL+2n5vz6mvHMMygZyzkTlPIfC8phzAPBfIPme5P2863KAtZx75+BZE5PzLGrk
z6+tlQ7nKB1yFHxJ9XmS41zpMLKQP/1zNgbSbGxT1RJlJqas1tbYRvE4DtYn3YblwnVDyDjBCM2d
qKjZils3fpjfAewPBcU+QF6+SflshQqPjhZN1LRLcvlajnr7PXutN64t45be+us+iplIT9OfAW8Q
dI3ddm109lGvxb7CO/kDVvT2pxAjbz//g1XKM0aZ8HylFT2Igb2qPSmqvKNJ3ly1QNyvVfry7MDj
z4YlLHmwcDhWy5ANUTbFFwU5vzUfXN35Achoz8qDh7F2YUIt41J0Xem+Un9q1tP8t83HlUryHSGP
qBJl3Tl+xlOWMycBIFf99PAJQg73KPbujU2agbszj9IAW2NlexXakWuwQWKIq6yD71EjDeZdDWGS
AwvRHU0tMCFSxOrzEZJk6/7TGJEZeZNPCUoe9eBRDrVPpMYUGD4iGZVa3vXTv7XFXxNv94HglyOe
rTaaP23vaNSBVS7Lqa3cjAohaBAgr89Lwk9dczoTOkkLvPpzvovmzhKN/4iLB7Y4XlzeomJ1TH+/
m+9XSKYXIhIFglc5UhQolBGh1A828GUp7C4c9jPkDaLPtCTE44CkFqSyIyfeZ6GNZWjgLfmDjPk2
TpurrFEVmjjwQbltkvg0G3ve0eCVUBxeXeKhCmLlatgOKZhfhMsSDid8mNMgYJq+uA3oNMxSCRFt
OPxNslcSvhQcPiEnsPqStoZ/hdGFKTfUzu2VlDwcBJVzuSRDyGg0uk60vsdTesXGH/FuXaQAbjqd
/QH2zP/EtFqNDLX24u6aJQhXT1ocTo9jst8iKMPQTqf8w6b84gcTlFNe609XDAsWl5lnDD88c9U+
GMjsGoLoYfgaNp5fck7LUsVQR4VVu1mcKKzE7uK8XEdA5+PBBcQhVMUXxV6Ccj8ovrbGQdbUzVcC
98IfC95LkZjRoRrGh/QJXI1ZoY18cUaQ7xZKh2d/CfHaC2JdMSsEdCounbqcAWNQOrtpEXznHzJd
v2/HeYihuO0xpajQGexqotqzhnYC9Pz4PIqZFZpS7/nMtFabS8ks5FmdxHpo3QHOONelVwscbtEc
rBItN87mUgPsv/u+EFRwHAr61g+zNCKzq/VPKjBH1CQ3kwCoWrQXjwDUmyxb4PhUYLkHkkosC9LF
mpX0S8qIC1AQV0eHAfR8u3W5ezxVEak3I9TT9INd4NQMGzbMeCvyRiJMhAv9OoNPYlXKpySdvefa
H56DWr0Qekok1KGy1rwRwbitvK3P3hszVxR0NThxI4ECXDYDXv+jh1bQwYcQoDDwIaiT5up5Ud/9
alTyw6gNwdorR87W/7DdkDzTal5xNEZ0GVNB7s7XoL1+i6pt1sr6wJulNnq3WmzMYvFbvAM/Vece
6vEO8zynX4XHsMwOJuTZxefDznCCubtrZCgzM3CxRL9M7MABq00HQY4/pR/OvNiCYGyU05wOFxaD
iYPfwuJcC21TYWSbUbMKQesSk8rdpB5vp2PDZyOWBk2PSMRIzkiU8XdOzZ1CXH3pMtk8uhllh/Z3
S47+pN6kX6GclCb1+vsH/eAtsM4CQj/qrYUxSlDqoWJ+jVuq58H84mk04FmyKr5fpASn554Z9ILk
VQpiRDwVRX83prSAQ00fJwXRcky0F56s44Ra5u0e64jnCK6KRyWQkraxuTJG3R4kkOLg/X6vAyHP
PxZTx/x9/FQTgjsGSYpkTbA//XtJsDplsv4f9zxAmsqG2sHpmcoIsWtyrc1jSvNfhKDd4ff3dMaH
jdlis3PGn1gaWGaKQL/G3MoaeUfi4Fu4rdkouL3vfvKW+FePvKeyfp8/ojXjm/ku1mJP7474bsn4
bHaBGs85QM3v3kELHCsZ+bVuHQ06NdXP670dk6vMTMxTcb9oQuLhP+jlcxfj5S5yOcmu9T+LntWQ
bWlL5/z78fakoaEgpVpO5kVsVldjpYudQJqJfffAJheyRVMP09dpA12G5g9QLDcqT2SQO3uW6mhe
W4M+2DU35puiu/bWRlnI3kdk7XIvUMYhpe7K7LdPfCqVIdA5bfgg9b7vk1aDjV7Z4WJOm05pvFbg
PVhrdDFjV8Ew7ZohPVNrzf0hSjkhstC+97NqGMD3JdrX97XBhWY81QfJ6qhpQqqziRXpb9k5CFI0
jhZBYL6dnSnJ4GpZCWnLOQb+PHfzDFB5t5e4/uZGUVhM4H+PBsHwTj4irdLsQM9WsjdocSSVvdwu
zvyNU2MM/4wwxU/cUTYFLBjgucKAui8+l7dcEshHjwRksqcu1/LONiYrsYM4UBgEXV6Ot5FKUjX5
XRpq5ymSnBp596APyabIP2UBw0NEaOu95zO82F2ULmnUpMD54E6JviER1VYs8iooqWRx50dOM8gT
DrGM6kSebA9eRwgHxcWoUXvG5eyHSEVuoE+hlAuRXBiRGQovj+Po1FyRTH2+gZ+Ku0JnYDN/Styc
yaw/wCYx2e1CGtnmfnAZScX5T3IDWqSMZ0M4FrKw/b1IBQuGzBQr8hR06JMMjavDTlkpyv1jJmDQ
87E7szwmI3e0eJQmvOEzUR9nKQrs0jhD/2N+vufCHVSeokpDNQfxqxP5gFwLaThqrJXpt7ati3HP
++pIuf+VlGC/853b/4QL4DzDPzVnafCYEHL2gSKdAlGcoqpRgHK+IVB5ibon9eBj6nB4ssTGtfvB
DJPJ44g36hKWq6EeP8fkJEYvjM8LZhf5PememkRd7pUJ6eiYsjYqlWIe+eGyXPv8D7s9sP7kUqpR
ULEFXeVX4eTPSJojWLpC1rqP/U/uqxWKw6brmzHR1enXHopk6bx9gxZEfWmt71fxSSt68Scnb0kr
PWY6Rkby3vfZlI+e02R07P5OjJXYPcfmiUbP0McMZTu84sic+U6E+FGzcszzo20teMJkolw80rth
np+JeKVBsyvxzc50zerOOpVwKrQpcGrtYUPXtF0PZ7IrxprKrrblQoPcjoFVkbO9ofQC2wQHJ+r3
6a9+/6r9FIPlj5ILX+eeeFBMPQnZ3gWMYne755+tICW5yjbInWGtLGCfhgcXUphYIlb4tiGFzPKB
Ti8JqI7y/cZq5Wh2pFCfDbjsgv8o0fkabk4rRmtHQ9cXIIYJfI8PDbiG71fJoDwKgDwsoLtx9UT1
aa+Zw8PXfNqnZHZJpvcVCUjbamSpROe7Wc6n8DbwBS+7ZagAqPefGKc4hm2ARGBXmq7Fevg5z4mB
JYLBm8olRjn6Mr7D6WpoIWIljOSXQoCJ56CAo0WZs1Vi0ZCgyusWpt6NLx6RLeA0h+Se9lrUntf7
eukj4TmEtJBeP7iA5522HFUthJqvZylWnwLEy7EOM+pvMc+M4YfpizcRJ/0C+1zCe9U4zQiimzGw
yU7YnKX7zDrsnzZlUe5/137gWjDatCWCLq1o1cZh+MxNC8CRQjVVyyc1ysF29gF1z2bDzj9Te3Vo
33Vzzk8vl8AcP+OtwFCvK49Bs23k610Nsd/gUga96y273Xgpuxw1LDC+17tsqg+XCUZB6OZOxuYh
RAFRez41wGqplGCNda754dg7XQ7Maamq9FoGwKJsvYi+ohRQKct7z4qrtGrIRpDyOOEjzu+dUREJ
mRpJuJZoeZO8eMcWxB4jRa0k2UAsgLPGUoFAA6lu8yaOaqqZHXx+TZodVMVY82FNcME2fO3MaMDd
c+3XTyF8d7wrriYzrNMCgVVz8MGBy8xX+LaiWTTYV6t/4MJzt3y1amu9pbJElvaDHMnqerSLMcly
4xa4nPDLJbhjedB11/6m0pfndm9HT99/HkgKL6JGMHxjp2IhoqFY7cCyJ6ffrSnGApz6OVuItJMy
AZByMHvmLTK9VNzJ3VDwPGg7ZWRMlZJdA5y4rJRMcmn2XnJ/7hRFJ2ej6y77aeu6rmXEM7Dve0M4
6b/ZNvPdXkuho8T2baFbx/5uvb/u+sny7TJXLmS5L09RuqJA717xUpN9w/JavtThJKABzRKbKUPu
otDOPOVEDcK5PPwtLmm+qPyA0eCpvKQ0ztUW1U9TLW9EydMz6KVDlZJ/99LWIWfEzPV9JcnIJtWt
wBqGO5SxThojldHitjJEjuWeo3dfSA2zA7i5z7P5OYQgHO/6PrLoDS+idVcQr3ohhTh0gAfG9SWt
G9pVBUobG2cjzCNcziMkpWe8McmJhu0g4qPFOIZoObpwAAum0VzItby0M+ruUlqfzIkootLiZeCm
OvFlS+rsQTraYbDk7s3vfBrGOicm6DZwfHDuroRPHtz4sq//GDqa/67BCoOcCfCIMJgYDw708Iok
+0GkMQek5mRyrmz/CuG12UXyRLrRjkmoUR5vU7bNAECFT8zgq9YPiRYainWwP/s+GX4dbQDNUXRo
ortxaGrBgt766qS/NS/BziE5k7W5Z8YuG4ROQ4o9VSYxip5+k/wuHpvedZbK1UQJwy4GF1P4QN/b
/HmLswAaNwr8NHzZXvnFwp3XFlj5pIlq0NPQCcv032L9eMhZl/QLRKkaPuPGCv3YtEIi6LlRoQio
/r18gMEdpZEp51UXWKgAkjXcuR+UnxwAxeJDGENz9FEdziYtlczCZnDPjLshgbaN+/Qucq73u4JE
mpjCGUlBR0K2TD0/mVKNZ9jv4TKJwLlqWyvLDjcBeeLEZ8A3uZ66SGRgfGT16XF+A5qYC07FD1hl
kC1nXXPQ0GvZI610Iq4XrTYTCgPTw8MB3RrMSpdYcXLzxF7cUUEBju/7EoCLxyxugtCr68MRFCpR
sO2dn9NzbMTFiybLKQS6ADiz+4pkMpG3KUIwxGCgGF5M+WlqqajzHNS7/zL1xluRDFhDU7Q9oGtu
gc2RV75/H3qx08qRxuBO7j+6WwyGkMC7oMnWhhmTF1D+TUmGtmCrgcU+hXu5/rCtoDreUxZDWOYp
2ZKHrdXlbIkkZsMqsOvvdsqnrWpk9HHCNRcVR5ZZkwsWWFi0l5g1tufBRwhYJGlE7GVKqZ7OUkxO
/J7Qj7kfqnK6FQpAI6lhBQWuKHAEWrN85KDohhAiFGv9ovmIjX4aEXasgaMTZjQztgzZT1Mq3zQa
lLTEFArWxoJxRtZLBAzXe5jA6zqKnOPCh2ZrkuYwuDR9Ul4AF+Unuv3HlFtccjvaAv1ytQEssGft
BjlJsm55Qx/QXZkuk5yIVcDVqHiJVkJwFzK3C1XADnzCEBxSTjg/WIpRo5LyTkkJfN6jwdyiLYk6
kkyc2l60SrOYSqodM+bXPC2xyIu8poc8kExIufJRj5EcNZYaLJzSaPm7or472cir1zxql0BLuN4I
ZwU2vnKkKWFx5boC4v3nleOCBDrTpH8wrxQGIxGAsoPvqOMYBMNb/EKx/J5EXbwjiV4k4dghtPB3
lXCSDs7NhScWe/xGbiVxF1gqTAPnUS0x9fi6oAt4mal0VY+ZwVOpkUhaxBYoqPPbNHgc5omdruML
+LTNrYUBIkV9o4fQQZFgcFafvXN1kY4ltaUcCBT09DGdJfUZDZuc4kTCbiUiOgEYK9ILqHDJvTsB
+oJtLZwjfH5LbkBGzg73q+Z3lX1hWNWtsekc5CKWRLw8qVmLoPEHvkVoZKg+HxgXnur2xRwbcgK8
oNAnzbCIzjzmzQuoirTPixr8KcsPopuS3XmQyXRBsYIWciYoZHyiFKpXFFPeZuq8cWK3UMTytFx3
L0zn4x4ARRBtknT4XD8c+mcyTakvD/TgrE00jY6YSjjdH0WVs0qxQofMLnpsfpUydjjEw/BCAhcU
m2SzbESVgACmRudynwBmVcdoAk2cjymS7M/cctVI4cgPvvxP+piuxAo/ROwbAVS/Koa1XkVfj6+q
cfcyYUUtWaj2ECghDhjyql1kFGkVxM//30+9ifEFeFpdNvsWbcdWcvKHy6zXfwsFUZqM3hytqwoE
DLOM4oKq65osJQSNLFMVIG6qhcHMowXp6OptjWX/+CHfNr9CXgXz4gPV80Cim2bsspAoVsShIHHE
vvV+yTx+l6s5tNtSGIhrLWcXQrEwbiMaVapEXVxLXq8VJLJrrbPtu5IMu4EAcPEpfKe9e4BEjDNb
NAzP+lU6osCnF/kN4W7GkK0NEz1B5+QhcrrIBKXZkH7CvgkXBAQqtYHxgfwz4LWCcsKljSz2T6yk
62ygeNKhMUaR/iLaS731E/YYnrEX6hzQE8DaPks2HuQ3ccGHfVidomPO3+LexEb1TcrbhuQMPXmC
tFvge3rJO6htLUAuEa/KwPztf7cTkh8Y6ZYCVjik5Tkkfr5VETErtEEUc7z/tK6LL4D4I9nntn0j
wdzWMHtYKM5RrlrfgblVUTii5hj/jVajk2tpYclmpV4uUshOosM/IpfPamZJUNORQb76wkOQ/gfN
DmhTcFs2oagBTiomZ6WB7YClUi81+MpeyykwOD7q25pae8eF6Lptd2UNoqZTC3iLkJXqd2amvj18
3O9+luOgrWRBLUod2Qtf8/0S5P1R7UNhYSl3x52zNgdtiYmz7ZG+4pIiqUBIHEGqHdd+aO7eJvOv
fh+h18m5xxhB677bFFvRAS1lHdFDqhzfSSCfQ693iQubDs+GfROGOOYhkEHlSPho9j8nvhuZ44Bn
+z9J4tamcL1CdwQpm949nCxFdkGXQRrdGVkzleVMknG2n4KUVwi5Gyq+BBs5jsEk9KAc1l+Y2miV
9pWPC9jGhnsQbINhLyd08gCjobMrpGSdpY2cIEcfSxduCcZxfQ0iqkSMUHw9WFb4HO4HKjwAMnfb
01yMmu8z6hY020cBWKFEZfD8b8bTfmue/ZMcfocHqEUvfohshQQXReuXYM/z65RbRvpYr7cwJ01q
5Ekt3IesKyse/QQMkh1wWYiEPKjWIavVra9t0PT41YVmelkxVxw2YAybZ/0kZIZPfvWPI8Pr4piZ
oYG3nPH+EbZy/jFjCgz7a/fHNyrCBzZ1yXSSU4Zpny+3l+DYxRq87qUbz370bT9yG9uxp7WqlIsn
Kh29Z4ezOIBHuPsHtZCoyDBp5WJULqe6YHuOjrVkAMkO8b2CGrQk2Tq4VuTRRWjrkUoiN7XAaklK
MShxVKPfrNEwey4cWr0wzpUwIHrxMvoN+mYgVULC4ZySFcG54b8S2PUIdGO/bEecQSAvUPNkK+Vn
2lBMuckZQkiSmkh/t9fp80zWr092Lj83H8L8Mp+iEqELsp5HcPKuC4rkl1mLglbUsSg7Ii/Dzjex
CNdpiHJoKo1mnZ53x9r8EmuWJsMzk/UNZDrZp0MICqg01VOK4VhX3iWuvmI6MRn/D0hr6tlHiZoC
UpFTc79RG9HMn5UX6FhIskC6ZFmGSPT95Uy1xgtefWYkqjqrSAGLJuCnbC5og5vKVVqphxs0VaWF
7/+dJheECLz5aASJ7iVot11/M9vm1BAVAFxspEh1gKilbPCcnfftIZLvZsDQUjanl5RnGFjpnNiA
qE+SD9U6YpHOYFsMm+lcianXAek2om/dPYAYqZ2Up6EmLIKOJTVxpuWrVfXjuywg40Q/AJJhMJh2
DYUZkAc/125e+qvfp+paQ/3BttmPH4lYEHZBZR+cJy5wQEJmAbI4m2l8NNgY2+qprDRdFM7rXbLY
tHY9ulEFo8lJyZim1Z/gQgHRv7pteJcNidhn069W14djFxt/ceAe/MQkU903cY71wK+nptT1qWrX
DiByaENqUw20dKyzH9eH6ESjvTkdIRN7Km+MKPJEojBzrKaKOtG2QGc28KS1kS26UaS9k4XwzRcs
tu1eg4EOzPUPc4trFvviTbFv18+RVhXfMqKubOd42E5SOh+1UKtfCHDgGlTW2stMgd4t/NvPrlOp
I2q5uCIONA17MWbVg5YOg5fbGztFfRJ2Bzf1GpiwPmrhw4Amwb08eEOpG0Rh/svsFsVAR1+yJcxJ
4qwmNN/6q4oE2gw5FdmuJ0Wg+K6C1oAl3oW3pAKXcxkvUcubjX0nKatcUBCliOsHa5yqlhUVNsUj
AxR/nohdotoXeOJ45lIIXhpiorMJQmTQ49pPwfIs8k3pR3pPD5N70MyOLdW+qAUsPo9sITqRcP5E
LLSxHHOtK0fonPXSMNPm4fVGve8b0mJt2/a4f0DV95bOgnwAPX+IA9XmcchLwO5zE14URz9dnFPq
QRm3hHVdEOnZYP+CR/cHNCu43h3QXWkOw6Ue8SNB0t7rPcXZ3bBYPPhwoVG+9lwqCK7xng6Fc7L4
0hjA4OlSA9X2FC5ryycQj0K2uan1qvu6eJEmf6GhRiOiFVzxYepYkJAd9AtmExevZMONBpZcar7l
7vI827V3g3H+7btG1GnMzp4EosRYzgM34Dv+pt1Z7EJqBVrFuHUEy27QT355X06BAQPIEgaPEJGc
/vF1xjqfysRcaDiwZaWC5JKnINFkWxXY2i14jOPIH7cNgDN0D6CN+AG4xZwzAmzSs+HeDxLpb5Yo
5tXT9CIq1Y/k9vmpzmdO9pYj3At07cJUUdgfsIC1vxHxC9NEuNcFVE6cVQA/bozq0Q5Of/xgUZbw
35fzg2KSue762iP0Rh8+xuJAB9FnRENQ8Ywcfuu6klvDcmg6ammZYkiFr2uD0W3v+zqdINEJiCcl
wbyzvnZPPQtmxqbFNAEHH0PWTT3RNvF9IYHLNcFpnco5daLr1mK3jzr5EB1kmulmrwlHh1VO33+5
kW9iuC80oVzlWBdrT+XwtDC2M/GXr12k2NzkZKUonN2BEWfODsvolB/XgvvtOksAdAdPkh2w9Zez
H9+xl/CHZoA23bYF7EiNqx9VwqbL2EEdP2Gn43hRX+ffuUtHuauJRMJtHICzzX18AJ0eIznGzgdf
spG58Gm0mDeDf9iQIPJeOQd6+gUIle+eOdMmRbZ367q8gDmObndVVLkfb2JqZ2q0BAmMz9RQ0yKj
GjPlH3zNuU0TV6sVJP0MmKHqFTToW2eT9fJpzHGY+2MlZsTKzhXvTfDETyl4LXFaaoEMKSV5ikAN
W037puv9qTaXjAE0WWKyd3XkrGDmpITZowCKMzMBu17fU+58Tn4Niz3mBYayV5sYYkzVc+w18ryl
lInYXVVB314cIfnnPw5pFz8SuUFWMawUg/GwfLZzumvF+S4mHuhIiAYmt6mGcYI8jnEVGusP1p0w
uShHXeaC0URX5fDYLS9Y7KlaEzEb8K065RyT37bLJB/PglasdFgQ6eJOJIvTcD+65J0s+qqDu1iq
UchcgsJyzBnaT8RY5UmynEmME+c5vC0CPdUqNFAIaLEVFIK2wSkRQSWZ9tSt4bS5jTqpjsRbm8Om
q9jWGYo0QBhq8VebLliMcDsnBhFWfCKh/jHhiPrjVB9kcLpwgpjMAqDTNndeYbv57oeaCxz+J3n4
Hgj3ssQ3esalkp11xdyT14u/UtFfHPOXBcNMD6kWs5D9NnQN0/I778awVHYX7FGeNIE3HIkJ8LBt
nPSAAa+dO4Ck6kyzrOupZV1dy+7DxLkZAEDSmee4/gKstLb0G7KqGk4sWQ1K6rr1xKFgiezgr3Ex
X8gDrQF1C3VMWaNBvxXPnFFysnmlOzDGObO6AoXfDWxFVRricDF5gNFj3XQaFWjVFuGDOdssRRmu
wQ+mB19lfIfrMR8SGCiLjv9duxFmAvDVc9ib5sEfnDHD94D8madclNm4G8gbrV9dWLXVmVZAHgtv
NZFt09XMtpmuGcjmKKhgqKju2TPCBX+naEiTFY+dIc4q1qyMtVv3e1G7DnTNaGGG3DqF7a7pBV/3
7pd/647Pf0orQEcYHYUH6Byr6W+qRkuHovsB6Ux07XU9U7bvxsTvfNdydfl/RimNkaNRGYw0154f
Q/28NwWfOs/drnwr30Pw058nA4WsBCOAW0wXl76n9HR1QJ7UwhCp0leq11erLk64+ejKhNBnEP6i
OfIjraI7xV1wp+TVRzLekXYBF/AkboKT+CzT1rorAC0VaJ2nb/rXUd/5zPbo4EZyZjmAjrDDSIvh
JjrV+g0FLAQ4WhJOK1XicUw5wyn76i6i3ROoACnOO4rjGPFeSSwEuMbNHHfcTD63GoCVe33RZXhb
mbuoiS0du/et/6eq63W+AcKSFcosxPPKdKVDH45cr+FXO5OKRYbuhv7utCUYD3TsgJPa2SEGQT8e
pBomOtDH0+2N9O0NyF5v/Bq+zLcfen60i2rC4jlYVNW0FBhcBinyKhjZHNKeZGM+d3x4Tyl1Hofi
MCBu+qTjzrboQ7njNYAA4fDB9qxWyjiygpOjBgZrZPdaZHdMtM/pZEUmn7DuYe1VTAnF8iRE2Mjy
Zr6yGWRpqf6i96T+fWDToZ8NGIvhMmoeAaMA92v4jx+ufekaMbO4Db44PrIS4XBKPVlFkS9diyah
YhuciAbypo9fQ4mNYNjtGQsVBdYFVajL5sFhWyU8qwn4y2CNJFT7RScGLwwmtoBFMTc1An37nFH1
2IBq7yPVaJKF0zPejVWxxuv/fo22KoS+/ufO+SrfRVglBr8E/9gHqLRSwkloVHQi5iLHIXSzLH06
7AEDxLARDQAhJ+yLyk5lBFGV3bWFURB9wppEiXZobSS+BuDkiQRNIZhCQQKrPe9X4frzXAao7sii
GClJd3Z73++sve6Sc7HYfTt/6RCz7myQOzIG+GBvmYAcL7JhH3f9ja4A9roRD5ORl/Dg2KiUv1OC
7Ht3tL2MawWnWjk7jHj1qxAXtOMCPBsd0Ee9Vp+chGDXaz0n7cvSniR5+GIkkCk612FmJKCuqRjl
/P6du5chN6kWc13ZQzQ/5mEC9iaNg3ng3xPsofVZFIvkMC8VLYLU5hXiH78uxwrlS8CPRrXAAdwO
+jhPkrgjCThPAgXiTJxUT02SbJEIJthXFChNXITAmETpqnWKaldP9aJR+ajr5UXE99M1aIvXnMVu
zHQ01lHXpC6HGSS4CxjHKWfbxy41sq/u4NsjF3cL0N3QftQNTDP/sbsKf4MyjBvxKR/pNU7YEDFv
03MIc+bH+hquLLBKylmgz6maVMcuwIBq6lPjihpyVaiKkJq1U4pcjnzC6kYt2/Facn9asoyrFeG2
V7ysNG+cZa9LzY59pe8Yg+zwbKrE79+jSzTN/e36kdmkndb23S6sjkIAeoGTI454gPnNc0lePM9n
VzKA1r089aunXaCT4vQwy3Fyrt5WZEXqrBR39IZVn9wOCtTaY3o0ExqvKMp5sU4r4RSuhzn5+Zwk
v/vSjSzlOyUlKfZHJMY8YEX0vCmlceHPivF0CGFIuHKOj2wdmhQmFZ+iB702I9SYxaruIwu9sXQK
Mjmgk8VXqC22C2YFgENRik4EKLXCA5HvLICCinmSJduC6i5G/ly8GMpI+gdEKpYbKn+2Z8YFmcnw
dwz1+Zq7cKjWKj8zn7w0PBNkq1yLoDzmVOlPEY9DsLbBI4vY+ug7qw3binXV07AnkWvZPFteigGA
izePqHs+jqIzuMuygWDsnZbGTgN4rrcTey+d8gBvbk/xghqkdxmrLg20TVtk76tcY48+/XsPc7NK
i53ErTV15+gtNfLA8Pq5RVLcrawXa85dnwVeQSQxCE+K3h02JEPvl7x8Bb+wepEiUqpXm3qetQin
2sWDWcx2c7lrDbU6umZmTNccxsP3kLmT+SRM1m86+yYPJlIOut6znlEW7iIHFHfTNJnwCjDrGe8M
hiBmRsM1Mmy/oHeA/zx+B7xG9aCF2yh4mRq1hWf8fwWkP6MJoFvTT5ofXG7POPakwRJqnZR+BY+D
n6kZ+b85+FNcomvWpXoqTdXFW5Ageeb/JRPFz16DMAxyXBxCt/7KpDqvcShUKtp+OLyvzX4bouvq
wCP1td+DxcONGP3sGSlhk46DCzEKGVYNGXTEMnp9okpGiSFS7boV5kkj7vO0ITaBIeSUgFaaoz0z
qh8hUpxY3RqI5pDcmY3zmJcbWTulW2Ek5A0igplJhvBAGFsM6O1gLw54R3AAzs3YwIiILmciAKMw
qgqpKV+WwtDkugttGZ0Cu91XbHHyTvE6oky2iB4wLsy8+SMzYt76IpCCvJN/D9ON6ejT2G8Bo120
DmsARLoOdzp1S5F773eiEeiDCrUfQbY1QFpHwZAKlavuiPW855N2lwpqhxFGZ8DgixlDJ63YKph9
1wu/jGHSHjWv4nZBPQpIVBOycdiAqJFewi/ca6GwAHDz9MzzYM4uIsDQ3QYY80RHtTnBBWxwmVI/
zHr0Qg8NdoCjyqoaF5csiEmgyG95p7sm2KMudQhncXDV0D8m5MicAmr9AL5+Sz3HaI1sJKKhC2vs
AYukUHJhfigl9BOxTaNJTZRoMgyAyOFUT4uSDdOYEHAdQ9oPFFJYyDopDAMKdUTGAapF7auCG0Vy
4+5uoHSv1qSLiE5iBaojUz9rhPwvKy5SeABcNsSjrzv0s6FbRGfc2i8gQ3ulI+XRqM6pI4hdtbYZ
prTRVHnGMrhNP72ft+6q7lC7MqnpK2rw+ZWKtvNdjfc4caZlTIExef/AhVJ1FQYW4AKjuzi6luaR
qqUUIH24jminpaWZySK9Jrw93eDJf06mbhIsTu4/8wWdnS3ai92ngtZoThRO3G7mO2zU9p+ztxNw
l5IzjnJ3HDDK6nv7PtgA0NSmb2AQY2yLda6KDL5yFjwvMqke4oOKPU1oR7zYbWbzUuguF7TqLgOn
vtzd66BLkDGX7pNvCa1thUk6PQQd1gLr1OHdcgZ+iePAeJewAp/rWiMjVFzIAW+zWFMbKGNpY8IN
lFm83Rh+a98+8KuvQeMV5rXw81bRyXWBXJei/WZcChLZ422VhwyMbuAcFsuTbwm9XKGd8nxIDzst
WhXW4RX4IMebyZw1UlZf/x8eLCKnQ5FONQupPds9jIuxEu/JltWha0C+I9OFbMH/vymFj4FxS1vl
3AxUzWO1TXzoVFXcgYh2MkgEVF+GAC30lskHvQww+8VZZHTxzzdOzaQr+TiqQXRuH+Uz8avoFWif
QIkl5+9NI72fZ/tvZzjNMo3+Ij0NNspAIbL6wv2F9oTpXi12Wi43yS0X/ahOj7OVYdRmIkWGtot2
QbE46QpbGMROuzSj2SupO1aTgES0yFkuZ/fxblVYg456eo2JakD/1Wz+N9K+7MlBTr9McXKM9LTJ
hiKG884eo7b1CC+qDy0nWVoFfQfx+uUGGSNkwrlQgd1tEeduZaudTjoqjqzaSczdiCgSLK9v7CUI
HKdTntQ+KyqEITMHOXOXQpbqw0pOBEoonE2BmM0Or+H9zEyVsZodInzEPSAiSYrRfKMTriVj5l/F
7qPJyuou5mndTAZflXz3zh0gGtR/STaWxYP//nxzj2/6Kd4va26ZtCeOW0Z1JH3RGCYjNjl9L84I
693tJlojqpcUt44P255a3DF3HBHQgJUtDu5frB8GmQ7oD2a25rhVpjRCDELl/dIfaTXB51HmyvYF
6lVKWEJEbCV0u+8mpfqZL+ARl+RRZk75utGoNtDbyXmI6BvhwehVft3d8bNMIxrAHAGlsLP5Q6dP
ByMGrjRLDFgar01hlmNPKV+IY2Be8gr2tGAGwC6Ex9M3LYvFdgT+3ATd4T2PBtoJUUs1OuiIynyS
/9hVC5qcoGdaoVBmSNO1L7wsH5oKX+sKPM8aeLOEB3kHCVv9uJYAkuZyXrQ0C1UdtOTPnt47u/Sg
llfSHEZLAUH+9/eZLJ8eZxIcsaqtA0Tm+CgKnfKQBNWnAE/tMHcXcvFYl8yItMkgytwYuKUV4g35
HI0JGkiXs6edo8mAmuRqCfOmYmaXBSXZLRvssNL+q8FLfRVOgU22MESiW0OrKTXu+0XpSiePsVWN
VbJlNEHuEPFhYw2Yu9fculT/QIbDkevW/N/notsf24NuQYhUTjJtWNr4u8mymmkNbB2HenTstWpc
p57YkOUbKsqQQ9jzDf1rjK6pD4A9VPI/ABqvmlI09wtEbQIdYLhBpMFGRAvUcmQ+suBwMhLWcHg7
ygAhJJqkUgavKlDbSBD3r8m/Hi9/F58crzIeMVf+vJI/cZpBMKpg+hDlk6ykcqA9kFweAr5aqTgI
SJ0fWbdt4jIKn5h13RQaAkP2HfRCbo/I7fZXdvKMyC3I4H1RI8wrEzbJqmvlDJ7r6BiiIeLSMyo5
74GUnw5mNxgfvHlrPO7Th/+nlcezb84qAhpFFAfZMdvACBZE3PrEYBkOiC7LPjpGqgJjWBZ7ZlQz
hgEK/ocUL5fYKD2XSqUQBTfTeWKDCMWcooE+SsOk0N+d/1qOvfFtA2/KUQxQ9aXPCL2n2ktSSFK3
DZRMoi/Gj8I/NSdDLq6h4OyBwXBVbGCJ4+xpuXs31wsEo5nVnBQ1v7qiU30iM7rLJCDVBvRguqI6
78lABQcGSNnWHfzxD/YGNOPW9sWXgDUSCZBtPg3CBQEb22KgqlAtWJUZO9xGydxgZrrfWEIl6orI
YjObjKFvJvuCuCKXRYoithKaH+tc4QGoTSJaDsrj69uwtF1Kp3003wuKKNeq2xvVp6C9z5IInU1X
oUC8jnghUU0KQ8aNM/s09aqKRcuq62cqUp4QtrkZ6scXzDetSba5pf5I9UVTvBCn3WB3Gky5NEmI
SGJec42F1Y02j00ay3qKl7YSwoOQ9tG7FF31aHhq3A0XCo67v9FLvQvK+dw/z3AEEzjOEmTyJZZI
0rOP43keTUQv3cughKiFxQZOIiIMl5HfVJAQ7017bFiN7VMWfYWRd8JxcCGsHv2fV6FPHIbFhBqI
PxGNU7Sccg82kl3Duu/t/C10mRbsVGUH2j0FxIHmi7GS2JqHfKKVGmCffq3CBae4BXjdIe1AlNHw
jDzq+tFPLEB6sePOW11ZNJ5VhkCoq4GGDupsHQEyaaizIjwrXW2op+CaSnl+oiCwAFhguvC7c/ci
PJi+DV4VLvI4wBpgwhG76zgMnrKLpi5z/qDcNJSgF2g/cwiTsB5fXBE39OPNKAJqkoo1IwU2MQ82
bktf1E8DFLUeo/d5bVJSCYz3l32XlotUxH385OIf5gR+NRxYy4NyYWqQXV9a8a3Voh8zJykBup2K
I4/k1U15PM3kOEJHQSCd98NkVvgl6adtaf/1y9QN1sTtE5DtUTRgXvv7mBjj4Rd24Fjqu0vQrkot
4EZ2KKgsqLdt8eynLLd/yZ23F1KI5LH7olOEuNmVnwJW/8sgCBqo7Knzk8p59+Mm/fdLFhL99vHG
enetPPeQdnGzOK1p3yD/a0uQyR0P+Xp+cfwR0yhG5uK7eYkv9yHYu40lTvH4fiSwpO9MST+K6rPR
baDTFrbjOYudY0Jrp2lLoQd1cadNR86cXQHIL8dwnmIwECyaKXFrRiHUB5TQAaR81F2iLygI1zbE
Vl8NG1LDNHmbnrmyIm0VPLoZB/xAZrDqZ8zbpfsTwx/mG8Qy2JRwRSSxlEGanAEjP0qnR9aJfczx
PqxNMNWbBq2D01Dohtdc6/jJ3ex/vvQLv/2ahBKfIJcFueF2PeawFNf9te/e5ah+UnI9+0Bfev3k
b2RHeq3dGxmImexj/or9+Xr+LoOuisi8+C+lrsWt1Vi3VyRyA6zcxX7gfo/g3QNBv6iXxY+cUHWK
SiRaaUvLj817XjjH/pZVKDNU8ezF92/sseYNCgbeAF/gb4E3Qsllv3zSfEUeRx0yHEbbOYayBeJt
0nPpRMd9av1QAihqDBqCl16v7cVMcGVZLUcnkJkXgpm/ns5ndlnWjyQvInl7dea+bJA0XpbqSGyV
FcP3htNoxI9ikH52ufCXdulDLApZoIwru9dw9i0TbKzbIRgYZzTj+SHCgfEYGn6IwWXhefO4yRr1
JX3fog8EdveWFyx3GGUpaYvaPfo230PwPoCVWBs5HJxJ/m6FzjrVpjbKALzkysus7vuxIgkNRMS1
3hmDDubMI6+lKsq3lMgcRAzq79e9UJ01kWpJ3LHsRvZBavGs9lFba+7thxBZPn+1aciostoSN+x8
CJNJnIa3zGxubDMh038EBkHl4iRvn3Qh5Kx81dK+TAvHbHQLWp59vU468y/mAD5A38JuKYq4seNl
IFudRLng3wsJzdkT4awAj2Y7RpsFbjml8Nt9RfXf+ed4lH5jdTpSIVY4fHZO1Hy5E4ZfImdmg04W
DGCsnNcwShi+zgJr/MUUD9HmlO5vgLfVvff6F2d2B0aeV2vIaoiS4lHacJ6iQ2Yc4qqdw5awf5Wu
FgabA3bcQ2OCQOMpFc7Bzhcbjd68ea7FUFvghaWXqlk+meFYhOD/WFKgvwQo9/35KQFg6T/R5Yk1
K9qrxUdg40eJD8/yIhxBdFOegV1K7dMdHTSvJi2TBFfWE4SSlwTjDH0+tyGegKlPizOKfrQSYXF8
82TRypKXlnkvWf7/yAAhvkrZWS7kHrCFARNbBdcnZOW92B1hRql8acZlwarLMo+UrOjrwb0lqNRn
yo50raeKCeGYsIx3iWAm6QqXR+Asg7oaEcrLd400gJ1rag4E9t5y+oLxo0v8pEThchylhRxc+O0o
cosh4GRQL2KQTmFiID1nGMi/PHCUrwq5xuHGD8wkohHzidX3H6KUwkDbPh+E/VYbndVA/L50bAHO
p7C8eBhomHvRbk4d2fA+TK21unqal/w1E+FVvzOc1Mb4CqbBNJpIiFMDPqUAs7KWxqsxYhtiDXyl
lUAIspVABStiXroJ6ZqGRSJ0N8sDwNbx5neU2EZNcHK41b5SBQfnAj0AMmaU7gQssPxFHM7QCd41
SGODBTj6sP28LjoixH8LzaW/z9R1Tv4d3iJIXOEaVx2Il/X7PTb2eEv5JGmNL3Tzh/G/UItG5LWg
a/w6J3VUSed/HePxEvm8IIf/eC9GZRhVO9LSwgq2BJQtZfaS3SNiJ5D0umYOL0VS7I1HmDDXmUTt
qroO/3hKW9BUtNf+v6Go5RLpk9IvCZBjzwNgxgEchNL4ZYXbGl/i4SEgtr9Fa38JZnqJmqwy1lXF
D97wepDmmowQJ5mIXOniZNIKlemxj3zSkRxmWebURM6LJ436e2PzlgDxDP7U1rxGPauCIaVJK0oH
btX4d4KoSeIz0qn2PYU49/hUuEktDJuEcTENERACZHtKX8UA3d5q+1fSih4xq2BTuYjgVO7ALiL6
RdyKHwbmmdvwPQNI8jQmSfOHcPKH1TZ3tgyYWSsiJf0wNcLwxBG1d4HSXOxYYv37AGvlT5yE2Hr2
x5vyXEnnTlxPm6x6dvBxC2q48u9VVNN48FECR1hfOcfxrBO5TA1fKgc+WWLxoYscJTH0PAO2s1ng
+1jemieqbpcfDyxRzLmzc7WN1VzKSkuZPoZrSTKlcr/rCHfxNI5mmBTRgMGZXwwVJw6FoxfcxX2A
LVFpPCDDOvy+hQT3ZlCB1apT47mkTOHB5z8DYlDDCoqonCLAPsLGz3rZxP3PwBAz8IWd7Gyj5abt
O26A/fnT5qYZFAqkMDMNihwk2BfehYvaSQlTeMnKQ0UGh/9HVvHaQuo2E4N8qlH96VD5FjAGs4sM
DtaQ9EK8qsNO/aHWOsqHflDeD4FOytjEsRva7eyVdVw4/UJrlN7B1rbsL6+LVIShDicu1tVUrPc8
qwhoFGysxacKF6LKnvRy4PqiZyMcAVG9gTWkQy1eqyKna0qyrAVqVXPFTkDcBj1itYq06d5gdyUi
UZhjN+2yz//wFEgYPZa6Hu4scV/8ifX9lAF/nZsZgz4bSUQIS/BNCqvsXAW0FTzgetV3ZTqolHtv
PqprJHGa+tBRYhGCqkE3kC2PMlO6/AwVlnvqt4FeimS7RKZpIhS9ViCcIHZoLl983JRFN6PmKCqz
Ie/syZqwH3hmOCOnMdOWcs6AeRPVMyc4Lim3KOUjXBxp0YSyOIUSvkaZkMNfa3FIh6xRtDIElp8T
4QKTiFCWEyD9XBriV5hvVoNbOD/UOjQHFcVpQLW46Q19rRQz4YLcj3zkd2ALOX81jqWmDJ5Nw5Af
2F1VekjfExTNcZ3+PadyS4fog3x8lcl10lY+V1H3XPGvkwbrOUB6hk2O62CISlORLH3KHs9PA6jA
0mk/R5yTjA8wA+J5nTC5I3IHiGFCLqacZNCMbsxrgpJO3RPXEAfyZQbxdGkOtdj+pYO7tkJZj6Fj
kkfJMUMJR/qNlEGeQ8dyWzl78kr/+hTVSUx1X3kYeGBluEI3gcyUjW+c/MJ2PRVclQ/iFcLPF+Wu
wnXrhB5117zRtE6m1B19zcVGsX7mQQkYffdhQQ3kfXBj9nKc/K3SR2MYtMze4WPHKdGmKiHrWd4q
XSBS2svukV48m4q48QX5ptS/50xgYNLvIAzHjH2JXsZRAdboh19P1yYer4EVoDqp5tlt6Ijkix7P
0gAt9Cbk5ul3ii6PT9bXx471qAB4mrNvPoxv8AQOik1Qmfu7hDZPpZO/3E+OAM5CmCt81DMWAIu4
ssKjaBP7gGwuvf0XTNi3gk0UGZH49D/wlkta6LANyTs9+TiDDdWTgh4ppCirLzs3xOg5e27htcez
GN2FMwVe5VTn/9fZ+jYKP2NPRN2BJ4VxdcpDYEclCFpNuKkpnGtRvGEaoB5pbmhK/L07qLAZC7lw
lVaemHymqSF+jQjn2VTQA7Z194fb6Qc+3iHjg7zqvbZuOZmrmyHHpIUCAak/twTfAqgLMX6uqDKN
LmRf5FfPr+QB7/3PXMh0ZGX1IZOouZlMFeca+kd+r+k2rkeJFB1D5auJautqqlPIZD3D0E653fBL
Psd0iMVVRvg52AtW1BspVBVe36x3sRZYNjzW6YYrpauAvjXOovvV10J/isJmjNAPbYBD3bqUXjQT
bBsCkJPb2xlTDG3DBWM0dLOGIRNugrRF7QsdND5lv0SW7/2DjEsWWDru0AoihPX2uG7B3VI36C1X
JgQ2KBOjZlMqK4IAWdQ36/tvHpxKabjRWyhoGk+pIAiEqVdWcRFMHbhPQMcoE8hnIIq7OOGmDz2l
6M69LEjf1CYV+oC8VAB9mwdGd0SmgNx6RLKZ42RmVd32zB36fXlGaE7LShX3G7tZNZnyzakYD9FW
dgsbOJfk0DiOxA+3umJgIISVhIez5XkcwCJTdje5qNmu3ZOTq2WDWd0ct49dK8oxhSaesUSCx5wF
UDmQuEXNimIiPKw5okqfyj2D6dtFntuVzMqu2AsY+OEM6W3l6LAAAC7M2JAhzwuyccA3IByMEm7j
S7HkhJ3JJoseuqYKyNQitGO+MHxw0ls+aT6kF6KqNFFS3OehlVS1P3ICRIUtWCUDH4eu8bH1oYhM
8pfoihuBxCoU91e6qMMreeZJuv9t27Zh3GoXHrm/kzleLQoabMIjCMwu3TeasQjaiUMDXsECEy92
J1ER+lZjvJwrNmPsKpyXgnibZGQLgbFRAiY1bisnt/rPqqW5cBS+JajJ0liTP6brsGqga/dIUmbw
u99FfPMItAbelbHnikJuPiJ/aA3Ci0LvOmu9kpFka5iPcGnor9DP9LWOslGXTgRbjr6JDVI0+7Eb
3q2b9Psy+Rv2xdrVXR9DeGo8dyCJHpefE0P6sq1i3nOtGjTZykoN61nlXIXhG69ZoKMGHpWZjLmt
R8eGrNkaRMP76+wY3XDGcbv8trxo782rZbSA9Hqlqgf53YIr9Fhn5gucFmwpQ2QUqzKGogoSp3Ik
VkBGfgRhm/f/cwmKLXv6ngkDbUcD8VU1BpgDTXBq5+nFE/YPlX9Dt2tvIsG68TLuxK+YiZXfpE/R
MzX9c8jdo/OG7p/nqUZuSmzTW2gZDACS6JiuMbVwo50tQ6mlk2D8LWxIp4a0vFLMpXhDHEsHnZHl
fD2hKGScPEcR0gvKLxWjYcd9kULzO1N/GERNhdjDjH/nmipXmQlrj0+00h3pGo70jzsuv1tr5/Wg
ZeGvcJ90eHco3xZY/9kcmOCXJZs4jkmTLQ1L6jE/Tqm+hQlL1iF6kqAk0dbvkm/gDk9tBYj4VVMu
ACRFQkBSv552xx/EHEn0sDs4WP05T2nTrNNt/Lgdq/+ZXTdlOEG4HTn7TLf9xy1T2BXPCfxeYnZq
4XUWzqDptpniA7HYop81axDsKcTjZpzNPhWqo0I4PjMlzP3IY/KIW86ZTHNXhsLhc4Om13AMrzpM
wGFvgiUsU4DJSAVvB0ucCMdiTBg7hpPJNrG/TU5/qiYs8k2Zu9iOGjEUIH3YK5CYHbHO3bpy3pqs
p2W1rIhpVPCN3Xw4x7fbJSmgLvHGBzv2AF9DEVV+NW6e0A2+dh9E1EPuQhVN+W/LqQM5tGuEkJXT
5RhrlOPwwmmg/FJsxXwAztAG/Q8OuH0aGwhswPFA3BS/JIiIShwnmFwSB2unqvvurfX+yUYay0Pd
cZI/p/rl2fWegWQxAqSLIldvEVSefr9jW+cOuqdxebZjAyS4FYEBhYlGQGvHS0gxiEolwsBOHuI1
fLhi7CElW+nTHWEQQ1ngHzGKRc2hvqnHN2VKMFb2FJXfINl9nDvY3B5SHploBaT9L0ErQC4oA6vY
JEXlBoZFeNTg+zAZSC5GPeD8EBZarSkFpy8e/163pmRWoL6TyDldFWeL1ZkcZLkcVgVI+im3sXi4
zHKUkh3vGjJoMMAYBHTy/O4GeLhV7uCNm79BI25fuhXnuHAwaRCGOwAUbbACoXcS0dyIq1cKAU0C
UZ2zumX54c55pGeMkSdw4cwHu8wcyR+Fj5kFia5OTP7E4S8Dm5Pgv3YFsTutgwq4Qo9rOTqZxBG2
1seIu05SA1E57jILr/PZc6cuIe6d38j91i+/0prhqoRPZMzBGCqPNj0o0Y2BUPl5w/izSL1odUnR
Mj4D64ekdvOdoI991EpGzBssKtM6hay1/TmedtgBdzhjJujwoE2/xmXLtSCRgkFEUJ4yNUt1oNeO
C61sU5YuoC8BWzStQv7XJIZ33bkXRDv6TZ0JU4PS6Se3R9Gr+jOkoHroswcJtK0YNMkA0QGIgMoY
TM9NWGcY7K4RsO26wEm+VY+Z780Ndf89GI4hp38fHP4SLdNr3E8eluschPXktpFoDBkyAW6E5pay
zcsJD1JO4AefNz8oDBrgWnvASQyJM2Zz3+VrAqzLQVKIQ0Dzdx/9v0TOAEnPUikeeBfqHGyMsSwL
IQrLtFmlyBG3eRCw1b52RlhOJUloyQyy1gDONt/OXYW0oxTgV58pucI8gc4FEI0dkSTc+Wwr8Fdm
rHRBtNzoX0eh6P68rqb3tmLM39NDLG1rj06vtOTakN6CTSr+qUe+qsNdDv/FhKvCcrDUrjICEcjV
CCSksKeCFPLvfg9D6+eEdHAHJ80/sxM8/X3ow/fRmENEM9EpN3kgzWeY+MSKpgCakutsUOJ3eWiT
faaerrCfA2ZAXl/x3mTR+QT+GckfkxLCUn9pEfbuzqpohZ9QF118qZQRPc8kGz539M+rBeO3NYIx
JHegblvh+CpBS7m0IrnDxvkwtviKFLXZ+GmrkYopEPho0Vj43teEykVXwCR3hitW6yD2fMCiFYtD
aXb5n87Z4Awz1Qg2C+Sf9hhdbUwqJNon6yTHKKyJyR1ItddZnpzwGsKv25qBxLNenUWQrPZJVzLn
Nkwak3oPc/5Uu/OBBiW6mnJAhhKH76ouva0UZRtJoRZHfdv7MfKQf7ovle0O6KJ5PiG4cvSkB1PL
sDmAGJ+CFxWeTRVHLCPQhZVAxTumJpDxDPEjzyPnrh/ANtsnnJjZ2PrbZ1szAsjwhekPH2SdEtPS
VL6FwEmVExtfGT+pR17Rd0j45ubHcxu+DmvcPpkSnT0w4lyzRzeQOgk3KTN8QMdk80WCmV9cMj7s
QilOPwqjD8JqInQf6uo6BirTiUXdzHYUHD/xrIAnOOJSqZ33y3Sp0CTA17OMr6K+npjXrU7Ugzqp
r9q06P2GPLzMAuUt7/X8ucb7+JRGnp3Mi83qNKt5lxIitlhJy2TMCG9X1Mvl6m/JICOMg5BkRrwT
8OTm646jeF4d7J4I5IDnUhwskm2x4o4bNdjYrwe51XzJ8I+GSVMkrNc03YKlkRq5uHnVQNVQiktU
bxn1qjo3yGx3VeWiOMeCqFwyPLgjehWm+HH/+ILClZrVdGemFia5YkLoYsAyvKxGrkqX7E9+Uh0+
6YEWhiXF2bmaRe4stHTf1ZdVgmu2Q9+fyM1eVJiam8WXi6ayRaCpAPWLn/N5xoEFOMGp8vJiEttH
CC57iygji+n8Lg9FXZXaBgJ6zxy33Rf4V8avZ97a6L3kL59ncO7w+Pm2DzdZjlvvcSHlHFLDmkTW
ngkViqbVoprGLOSYXYE5F9+6sCbSMAD+Ibm8hNM1p7q7djxNuzc2Zj6M4vH9FdJ1+6nP8E2lfEh4
aYhEAANww/QEywoC3UQQI+ura98T3jMgCYWE3ukgw4eVfnU4E08AHx7kELgN+uYbiFfK/tIvrR7K
PE6oC+0CJIXIGABdiWQsxyUXGCpAr+PqYrj5kmICyszu0MSCeYyEKuTmNlGtaj787NXglpQpYMkx
exhdm6Eck04msZ2Lwn3pc9Sk6PtBRlkh4ZpVDJjgDW+3nPiE87Ujmi0cGpARfkXSNRc32o414tPG
ctlYYlm/zLeVws91OjLdFloD0gisqykPAxDFTaidEI8VAxHWy8F2zeKl4Co9+VDxGBlZkTzZBIDn
ueu546GoFHerI+qmCyt52P5EqgttpeNsFbam8A5BmLIK7gwqk3O/ExO9kVLAoFiijjRsMg6KJYIg
U529hXlksDl+yKFg0byP64eH+SSPWKZXcrs06RGJ4pHs/pJiHhIr87jksSZ01UgqWSSa1IzciBbQ
Uc8THw4XWOqB0blOFV4LJUN29l8m43Qw8Y4mybLKkxY+fJLbMmrIacZCpcebO2ezHf0n0Hdrdm/H
g6rU6vT1h9n8PEwOsXgynw/GbixP+iCamRZwKf5ULAl7oixqYQGGgPrMGgqXZu7UeTqk/W00vP4w
ikF5FGMAqKy0nfbo4EaepDkLr4wJpR5XGBPjWMnmI03cG5xHMuOIbIpPdfL5LF9Y0r3WbzDzcbWZ
cvSixLlpCwLRcizBlCKSrwArNNSBvVpf+hnqFqxaosZtIEDMmUx/h1rTnvglx1ZjIGYht8uMYa2p
oy2yh23xo5tqZ+GC/EM0ALHafSLoumdOZ585G3KJIkeWrhiW3K3qSWoOKrblY5OvygfY9aB1ny/0
/gflb2SVVnSniRePHQKS5BZEwBeeDraQPLdsuDM5nZOWyn2GiFdy7uMwQxRYedD5E+vHDoKf0h4Q
bhaOx6SSjfw5KKal53r1jMeQNBGkekQbIhIpa0QrT/BRcH006xZ4zVv7WyK8ALUEl7CuxWdp3qS+
fGLWuh1Fc5dmMUl9wKtK5I7AHhA2VIEJHDedld08Olck11qaI8wwDLFR9X+AKEIKFG/dqcENtPly
SxDZ5rXdap7M4b7X6THMNz9V6AEwvFApvwdCs6b9uSOW/37idcX9CX2rLpYQDhQCVqoj9ZMv6hjR
FWwE23ASLyWfuRdZTpyUdVhfm4xuQRNBqPxPj7rXNAogyUt/pS+C9jU2Th4YqpTvuXws/1b7JEXi
VF/382MiqGCSbXT3CNs9okLbXEU3xypuTwno0Q3+3Fu/Fz8gDpo6CFfW2u1PIz6Sb1YWjMtbmBNS
yhZTVCAJbkmmzIHXrJTRhB2f3Lxie5BmynoeO4OxvXPcYOOPBAyo2XLsPNCkaA0VhFVNAcNp8Qw9
cQ9hOgy8ZsiQiU8pu5K+UDVxzFpQJcVdlsSx9DMAKO8qEVU8l5OYyPpVLAJUcgYqo1QQTHnb2+2+
GOl7NcqIsEvoH+mu/g81NRFiWR3g/j1OXe9R+QOTgdmiY4dqqbv2xI2b6dqrbP5Wdn/6XbraKNLC
8UAvCzUVeDI7xmw8y69QRP+NeotiJtBvnzYkB7X1iGNuLfLPuyct/+QDxHKLUN5IHTjoQPHmVlK9
V/lSN0zzBnsZxqG0Dn2Ns7P1rCDRnHs+Nb6bicX2x3NOhlpG19b9HWGCK/iGrpIs7o/xIYXhY12x
MQSAPgLYgqP21gIMHwXaEglRoP399/mG+zb+kfBWU6NKFaLVMtzPTbet81TIjMDTV1Ftq/JGFCO8
ZNznEtJbuCKkkw+G3iY/s/UE80q6/Adydj0DysLHUyCWpvlwif/lXzT2vogoJlIE5ItnigMjRlr5
BXRuCiSkAdnZ2SbycXouPln6vDHgXKRbGaGJjOyGNurs7hGDtJmStn3oRgCrJlgZoztEK/S+Puhs
UUCwSIL+gDsIbkUuFbKxFtg3eVPWanNs6ZIvxKUPaINzkqcF5PK8RrgQR1a5e5YucK6CrsX4oW4y
dndYAYmp6yYuFeApPLLLkDeXN9fZBhBqY7NntU4bh2lin99IHOAfudo9WBcNhwhnhOCtFH9LuZJ6
qIz22gJ9FcPbbrSxue8fQgxZIj/JZr+Q9MaFh/MHpvNTIezgzCIhxjsZ2b6B5oL/QoeqsKOiXtUq
kVRQtBacxy4tCADePmT68en2zvVEAP5yz+tjZR20j8yvPAlUXWGcNZB+Ttm2Mh7kKVGX7QXH8eB9
n5Su2z0js3mLnCD/fuzLiJGhsG6mB4I8kwlwzuvisVNq4jkZtumNgNdUKIOCEgSAdEwU0aWkIPB1
sGJGK3DfbRNLynlgu06SIVPcQN0iAmK+zhue60Xf5bt4HmFvuuHfD+v9UadZwaf2W/8k9gnVrCqe
C4tpH2liqmfiufJLHpU88kgQsz8XrTitYKq1i7KLPKSZwPuukQdY+jN2zsXI3ABgz7wlscwxWu7y
Y7EAm1YSXGEBk8EB7c4OgitPp9rLUxQuwRsFQ9pU5VTSolxq+/G4J1H4v1WY/DWseL44fYaPPuEQ
k2jJ+yeLlvQ1zzJLMquoJpnZOYqe9+Z85ENHRumo1PJYyjmhlZGcHyu1QMmPzhQiOVEqO9p0EqHw
kK6n3vQTrkbRvPRKaxEQeo9wDW5XRc6aE5uJp4fhylNSCW4dxRGR+1ZE7MPgG7qvlovRJZdItybu
/2x8rDplWG/zf4BZ/S6dYXpEj9lghosyW6KU+tc9y4uXDbKt9aGWDsF/HmuJKMiFB01ANcMk0JMg
hqTWvcUfPa/DefJ0EoRAhSTsL3bXYdfqh5CAN+p31wQyvXc6bXFVcfKoMNosPJwfZnAGEIOauTNR
OWd8rbXa7MPNyQr3/1lpacbeTXL4GVDasq7o44jDXun0EE5LH+cdpENxde6Z+H7PD5lxgMAjVZc8
c6P3U2XDapPm5DgkTP9erSGAPx4EP3ENIfE+ZxrKPdy7vw0hCoXsZS3xfE16tSqTNkcCyIC4pcKH
LxbqHWhsgeVG+x4+C1jf6hgAGY7KcxTJi+t9V9rAkOmMmqYlxC00EERmFeu9WLH0fD9qDMBkzxrP
Ss25Q2p/ueLI5Bkki27X3de/pPK+LaheHNTMt/xHetubJRSrbYWdEl6678zdE8camQYjquKAtys1
UtHPNrJJBmK4ORb1nibDMUAddzN9EpF3oAIDJhQ40Q67v6Gw4gbkKZIul7JIxWdYeqJn40fMpXiM
2/WsRwSa+z6W2DYDU/s/Z+sXj0Gncb7OYjiOaTeD94FKfgZtCbQSNcsqqhdD/M1g9dKHXlN1Y2gX
UM0WAlntPdPxEO8lfIi0qNO+iTq+bsJy6wzX6rbqOZzne5nmy+Wrr1unjB3lAA6qlt9W80Qz8sgH
MtfL8HmfItnYwdbhBKsPhQ2KkH58qtDZATXjk+xpOC2z0NN2S5PII05kceCkszwlkoMNLFFpaAKl
jL7I6nBEcNWIuV4N8vDUjhad7Yuk1msGEnv4m2psEZc4Vq0LnAcSSZ+TQA4wiJg9ICycVV43zghH
gRxnLT7h8ciumS/MZM5DSXJX4yAKOeHqVWNqzNIo0Wc0j7z5EVL8be3+69+8jxZR8iknLJDNQLAb
enmtGdQI06+iBBnh2nK7R9ycdjXxgJLAoA+sp6IScVDEy/p+K+gAZX5/yGZk47zyE0sVySHjEdOq
4Qc1yffEpulx8D0pK61mQyMyC5e8cCcxuSEYToo1XDMLq8uSzLZLO5K9w00oXYI+Fr62JHSNam9I
I7XzdAQTuns/NQg0HWtxSIbCuid3yDDWs4cYfLlibbvxuWrpdvFhQ7LdVmPOmGNxqvuSiB188D+r
B2JMdkAs+/Tq2faVws9whMYpdCEyEumIPZpkf7UBiFvcHhtBRgD3aCz31EqkP6hqVxAtla3/k9fj
TIVWo7+UqnvUO8CfG5wo4Rq0CW/1VPeuqc9NLTMylhBraC8pcOZh8WFF6X4E/ynoG1Zz05WuUgZS
MJSz9XOHP0Hpk+EDl3bHpa26O7ictd+Pu1x57I4bCT3djBBls5XIRv7XGeO8niX42vu5UmvhkoCU
hB8nrQYKid92tRIxGo7vUWoaDh4axxViBEYtEYO7ccAs3quU/dZVFOej0SYL6k/ZseiwNDcQFCNX
yagMtPxsv5uoyG6G/DH6vG23xkMFoV2N7VWHCYe8Hc0RAPXYHG4+qyXfaRS95dM/Y4C7EnzldEWv
NwZ6la93BipnFTBt25kcjm2o9i0yzNVYWmcvYXJdPb7kbVbTq31x8mTM7xLa2mihYItajiJbYPvI
VymaYtjy+otTcLJ1b7Aklbeh8ncQIIxiXxqvPVXbSv0khwSKDQXACIzNu5z1YHc89AKSSUh/4ddV
CIfITVFTeSKBLl+HKAo3bhqisbhqOZZ6zcGpqu5/BTp+Ko/cYoG3il2w52SiE2hizozIDypCbIzX
DTqpUZcNDmi5Hsn0l9Etob7g7/eZTLxPdWtfr2u8R/w/M1wcJ0lhHLS2E/nbJsyWpTWMQ15JMX1J
nxTIO1MCKjda5Yg2RDF8cWr/cIOd+u8RR1pFsOt5A/g7qM8HZS4oFYa+bYdvzxcf/kCFzYyLZPhM
lAKG4NNbzPJ8xiwPAL8PElEq4OxpQ9Zsxk0JfjC3jmaw+FJ8NkGdFDRmTTBtZAsUaPKPUqgfKAXz
oy63tXuiuiNqnJhmcS9M+UjUESab6o9YEja+GFDEZjV6CNrfb8jahmdwTJ+lVmdJQqlpX6TGj5cb
xFM/lpsf0t9HQQ0KzQ3z4A8M698+Jt+yixA9BuaWX7ZmvatUcS7lqxwUzx3gERbkOztwmxE8FI0+
ew7INTP0ue/83J5K48Ep/njTNR4JHEMyMQapwEiEd2yYp+z8i0zBbjeQrwht6W5VlWarfGxaljm3
kH5Q7fmCXCfZY+9U4GqZaZrtS1OleMGrSSUZg3flbz8g7JMO5m1bm0J8n5Y9yfEX/8Jvtap1pWzN
+TftVZUPBIuAhXaU6PSpSyZTd9+aZGUSOVbIkHjTXydcrYFU3dMuRx1rueQXiV9QhMJEAoBdAs92
DvOIpSdevhO/XKV0s7qFQXichH8fxBWWXEquyLl0G1RLz8FAJlph4oHc2qNWUGq1xSwfDGmHw7xl
j5tZjDHkw5Ov2mhqSUR+BIM+S6KmPFjzYw6D35Uqh+ewvmft1cjDf48/zld3ueHbhybZsNKXxZ+t
i29k7FPNhCHnWiCgJmRk6YzbOMMUmbiHxxvdstRh7brEsR7Mo2GgWYPFatzyNY4P+/TJ/fJZdmO1
g20BDNOnLTyV0GqAWVy321DJE6WdysVxB/z5WVavSfx3CeXnY6w/r/DMEoiRloDZ3VAcnaPFkqRL
y4oqVF0vZZ5yREz4u2DCWDLsv5BYvhzPyWoeqj05NMapK6JrOIArWzB6ycjEhDJRbQm3It4JIArr
HwgOoH55+ulnqynX3unpuI/8pceFn9wCAt9X7kO6L9bLJIWNVb9jHIw01uH8dYcFw2UtlwITngVw
qfrdnyDWkVMjdWmSVqDWSuJvF3lSw7l+UBopDGfVbhUm77kSsBo9tmj86k3JFCyceH0s/hSCDvtO
+AbEzb95jTrqa93UKpluHTPMvOm6QVwbMd1xupA+7dYrWA5B3rQf+TlnII9RC0SVbXGufOtyZ9od
+D6Fp/w7XniCjndUpcd8Cwx14PaRmJCQJgKkvLVUEzpQ1ONgk1w3Eon8LCHGkX0GpfQZtHQHbeUh
A/L/Q35OO8DHtAev62hNGVkA1I66azYMA2lcq6XO2aZ5bbdFC6w8wIXx5j6caVemDrFjlfL4aOgQ
5RZ2vAqzEJwyps2L04i1jLZZOJpAVquMtIG2A3O0C39epDJNTrNd8nZ1dBJrnrD4cB9MJ43C5bQk
8u6BD/gGaHW1SCW8bkX6jqVXUjQ5hXz+fCXeOvIbNjrNQ34lbPwoz6SGXxG81LsUcH6W/3w+MFK8
5C2QnZc7e3qzqPZXey1jV2m9kgtFOTY5k0grlSYD5LwUhV0bqCPkrfCKqql7Yfb8GDlVQz6IvNWj
4ltDjDSV39HNy0iyaymzDrb24WRix6M0WF5r1rc6LvXfePKhUOz+gdd7qg3E79XmBF4TRCS7PNyN
n26C8dHYXuLXS53o0TtcVo/tbIQgyPxUaDGI5oFSZzLk6u3bvHCJDh1EHNBGJ8BHV/Bfw2SX3Ti4
hjHFSvqCwOuE1Jmh5nin2AH7WuqKbNSALn5Ok1GRNgyLjYh/85qVNF4Yz+rK+xD4LzpyXMAjsVdC
wJWgWp7upx23FrW46iOQKyHONdCLxAeVCKvfSr/HF4l/S0GLoQkvCBjhRa6uKJeF3TR1DRWXgkA9
dIXRXNvmZJu/ZCAi5ohbXY4NE2ZdSV6NSPIyEzfG8Dd0qLXwx3jnNpSzlJZKSVreVv5jg1tkN82n
DsrfPf21gnOUzEm88SQKNKwiFaNquY03DfgITkBsRGtNp9bNWSDsQ0vZti4ktYQo+36eAzq7qKTq
NgELG4T5YX6ztbnS5P0dFCW7zPGFEgOrprUXlwYPgU6l2igWY+Z/9K9PwEKQQYrARmVG09OH+Dzh
4S30zs6PebhJH6xtPQhfkTLIUJreUl0OH4aWTrV2IoMnDQT0hJB5uzlFdTLJWHDXd8/rTU5mHjgt
FrGMZa3Pa2WjxHzwoPeu5zcv9yvK8JhkF+mrBsCFVQ1paBTuS1TlPgwna0pS9P9J2TlXKI7r7+AD
QXuZeVR6AaKh6mP4lvO/a+vk2sf/ySuTlWWFVFDJUkbU3E3Cox5S/p/YCxCdPQxRCbDsQi321WPC
IpIiiLK7lwp6dJgpV9fAhbWE5lVF2EJpShZxJFFvc6awrW3Q1bkUXyAMlgRotVsmny2WzZR05zT7
xOaoWOY1zkAbTM+NSLVYgPRpOzSoW+8H/IVWHFhNNPkX8rZeOQhBKokxI7gxuAAPTp0HG/kke2sd
XKSPA69YVt4auhScBPkLn1MvimoGYezLmZNzaLoSwBU8Us7o/JDD2q18ct1mMcw0C/yJ9spfvoLd
lwRC0deFG/IlJCxLvDaeFUQPTSz2q4pR9c+kkoO9pxyqI8fLJDsFhrdIq8ZtTUig+9YNSNnKsF0b
Ziakk2gd83oD2W5sMQShMr93sv1BsZfr7B+QE45xDe83l/i2HzLKWari4+HeEDejo6d33Gu5FwNa
5QfdsEpb16HG9gkdiG7ZAkRGtZMiNUPpsAy6SEBjbzWBeNMBMwdorLIEkfC3DtQQM6sR9/gQjJd7
TRE9WHpTvitX/eP/u5rGZ+fyc8mzVg61gmvtdCA3+ZUjq9v9RB2h/Xqab3zwe+oNH21aL8BX+Ef9
9MReshxYF1rmmVg/iUAu/pC8C4aGCO2TvdoA6N7JhNedWzgu48EUWFF4izHm+g0F4Ok6CEaYTUKx
yQ3m2h/ab9TZy3FlpFNRQkziYau58AwL028wcpKnjDKDyThnn6f0iljycezKV9MjPayOdZIw+oYD
eBVZnbouuZdKgKBhxwhME+MWBWCuiwTeiLFeBa7GMNg25p03Q3ukvTREsGbI3uKrhhJX5zQoEfPT
d/tRH6L877PkYAcZ67EqgYrcMWN85cPRinyVAJDG3y+JJjcxv24i7bUdzc3OByLLOkt0Bi9Ft1C2
bC4aJ9YWCbbW+Hj1NZrHq1NVuPtq/Y85gan2vvk9LX5YOp4SpfnRiYeYzCJZMiQo0/88IiZsV4I/
ayLI6Mn3P05rvq28C0Det5KADU7Fb6Wl2K0NwGMRPfTJAG2FcR2yEz2dOZnKnRqeQvFo9CuwVFyV
YLt7xYu4FcKV5LxYk/bdTM8Pmg2itWjH2imz1rxYxIJODH+vw/ykJl1FswPWsNkyPj0ULkGtwDpI
CflPR5GEYBQimEPNZlMhbCBnx/fjhjtD+keRU0aNSspdbCLyQRYmtYCWujLax7UBupCf4mjUyvIi
s+7FHP9NgXTFUzfwbHkZopbF+iunpdFMuMG7s/+N3IxMa+Y8xklTqtBkbi5tcRSFP0NHNql75/Or
8uF5IOGpINqalUeY/b2ljHVfU48fa7c4Z8SlUQ8Hf/nObtBZxWkx0UA2fWMbglLMwEronAkE3rmd
0zASgoI4e4wbPsAHCF8yWpHfWkLf9FGQdah/HtvznM64j8pvBro9GKAUuWd++A/n0i9eNw4uvNsW
7IzhfK8djbsrghvHyevdVqZ1meZFMwe3Ed2zYosEgdcRgJOJJBvO0LKGTRmf53H8i221S5AJkZ7Z
BEiV7l4bXQZlcwwVIfug5bRN9W+iZByhvMZ+H1HjV7M0usXBjwnE4nX//hRcnk4D05QchH/JyNBn
odT35DkYZ+IwvF+AOAfNt3uSBiBJ5pklK3PU1lTfVA+5thn43+dqLWawgPsEa8/Ho+vVP8HSa1kh
1F2w7r/PdCiRbngFIDfZ8q3E6DAxD6GeNTd3oZ7XHtTdUZf9bDK70fN8+VgnKJaZsV261ow1yrjK
5Jy44hp5X/OK5TMOKtJ43UedTY14clhD9I7YS322rBdZKR8bBySkVEtDa7sDieWf8dEL4F5MYuRN
SkYab30DnoD8pti5dq4oRpBBxQzFwn6xe8h+EaG8vgenF3xwx3odflwFJoU1w/pSL7W9Nl96AKyX
NM+HbFEwp0C+BInN9XMcG7hl6TReSjyLlI8ockViq4oJ1gGcX3fc+mNCxnyFxlvA852vqEggSOoQ
2KoohfIEK4hJDin/e3J2Qd/MbG4UmOaY2nyjyqvE6JBeyL7Koz1IQZMEzMLsBStxeSliHbOOZC2c
ayraWqo2GE+XtSkiCX7z8ZnNlOYetkuCe/bAsEAXBZVTh0oaziG6TQexbaZTSIazHkMhTvbZWegv
XVr29pczd6s2pSTBROt6iFBpukR8iBPyeKoo2xU1ig3f8yhJcFxCXQkyN/R/oBCNVgofCVWmI6qT
A2TLgXIQQsn4Y84WMV1ulRYMNFrLjzCGr6PKbOzJweucjcfFHZTXst9MmLaoTyMDZrhXjZNIH+tr
la41ALI6fWdSQgWlOZoBEbpy27DrQW24/vQvlzGme6UDX5o2KscRbQg3No+uCFYbou8orEht3hNj
GKu8Q4tZFJ53IbA7cRhCbV5e4KorjhfFlxVFSV6ndA8hh/D/pY40zl0Ta1Vvz8qsAE90Yz3XeFT8
2JC8/yu1wWaf20H1v1SGEiTs9wYKmjSuJfQSGF/shod1DnTVehaWqCreX+gZtrNKQezS5UrELDcD
g6W+qm3gcWIC968eMTL0lPqy/dJ2EZM+4EYEh2xrUe4vY/1cDpTGsaxum35ngKphFIxq1w6jwLyo
1TDoAtgLO+aImAWCMtEK6wC9XMzTEc5lPlZ8Ov1KEbKM0qaR9LbzN7RXrRcqQGKZh3c3tgz+yDv7
nuWrecCZ2x61E18gtwbMgq1OCJu5sCn0YZVaZuAWKJLnyddYqHeMkoqh/eINYqZ3tspkE0unPePr
XA3EnBnrlrMvywPruzAOEAzbAxthIGwYDjc6fvQ9wV+FV1PIuDH76I64ICp7oFkkYjVuim+m0QXE
rBPDtPvVD6owR+HPKzKDIJSMo8BKyAxJNzagqy5QrLUehfJ3280mS7QAtMMTG/8g/fMYicTzr0ok
tdeS5LgmaeV8p2ZdiVSFF/VtBnkUsvEUUdM5Yj2MTaEGYo+P6eoVc9oQLoV3xBRMA0VGTqBMtIfw
riXiy7Ti5SiKQCXGP/PT3DMuhlz3P0BkzMfhz+FKuz6ZUy62Sv6oGYgx7e+v0g3IVEG/GExknWZj
cQzfQUsek2BIzyStEu1e4brzaOKiapUfirHIjcxZUOO5mcYB71QyOwuHsYHdaVNveGgpAJ9Wniry
7PRNFxjUW4aEbGFrHDODVQ71oPWMmiwHG5QJXyAXQjWYF13Ja5VHOR6WmsNpyIfbiSGdIAf4r0O5
UOzp80DYJZcxCMmsSf9HofMW2RqJ7Evm2l0skVsGhF2sr1s6IXhPclaBVFenG8Za0/0Q8VY04/uk
GN0lJYMNPg0b+KS0pT99AuzhJEK5MPnH6lyO3108B6wW5ISF+wscBNzog2B6vibR1VSd5L0qHPdJ
VzZzofRDZkUhSWS7h4ZaKbm80+u/t2v4P6IksoY2HmOqiraond2NwsRf3q5EX01v+8KFqtpyxuN+
n0P/rPaDZalgnso6szO3HlP3dfKud6txHOpsZD/U4aGU60nXSZJYvI8aSwp/1uItveLtQO8ZPjvX
Y9hTy8BeaSzxY5LguESMSURgd/DRTpPwqVM3UD7Zl9fmZvgeBBRDIqoLizHFPb3xml81L2GMyQC6
7wk9k75cz6QvZAAIrCJwKB195kXX49dM1FsLngz3VNiC7R5sgQ5MMy8kdgIoJ9HCqlEBDI5CrKWY
qwaSKspEsxVYHRHd1EGT4kyOHchyVQmXkiIsjBR3gfyUIbB86cOvx6w2EOnpqGWO+BSoB7I9bQdF
dPQwaUDfQ20xExSBFe9e6JyVmRwKAhaoJvTIl5unisM6ThxbIGpSJH3qENyjUhTPiflqEKnv+JB0
slzrHRFFAgJPglDYItVct1mgGzxpSNbCjsAyV+3A1k9ghYZUu0aMJIrs+Co8Qj4y3KjQrOO7rFRm
eDbSUDYVbniU4y7S7/TmDo0BgXIubGc/Rfnl1n6EhlBPUeXovBwd2p25l7iVmfjv20M0s8mr4hGU
kZJBAIlevYbsyl3N+KLnRNVg6QtFJ3/HpTGwhF2Zg54+rhiDYsaJMM7VKr5+fxufMap8092Xwj99
o6xT9ZLjjdNA1qrq3TPcMc+Q5CAMR/IU43rEl9BDbdU02nvlDLeML++MbLzk+jeFeE6Q1El6syyr
bVzpeaqBXvueqHm/d7a1prN6McqGMRzZd17O/aGllTnut1mE/q+4lflh4bRJ03zXm+GVMNDH05us
n2btOFJDDekn9xTq4nghjNO21jHkw848/ywOfxVAdT0yn/p1w7dLzb26boPxElnpuxo82wnF2T+o
vE1HenE4xpQkDNYcbaqwWDxi9oeD4XaSFKphS0gmSVXm+lQyze+954Y+O4yTu56Du02l5Pk9Ag+i
RFsqqfIDZ/SUIBiUTGXkkpQxY9VnN2jfmbmhCYiXN0B79Jhs4ZYwd8I7SZhFdxehGouyZT0ljWZL
AMDj+MpYtqi8uHNp/r/49HcO/evecz7rV4M2AIbzbnLr0NFCtRFpo6/LyXTpdOFDuprBICza6/02
kWPGCBcEtPKaRnoD0dVtIuyaAGamYSiXq7qsB17UDr/CMRe4z8omlMXDuf1zkY9iFnfnW31PJni6
1H5NgpEtbrjJRArGqmZK38LOlh6H2ucna09rPvdjeIOOWvvP+egqKoaVH5HjZ2AdrMCIqs9O42XF
Q4WwWZ23hFIPwlgluuY5JbjpY2kuIKUUWfgJDsj0u0qmiD8RSwTSDP420tqvSpFtjmZGY7aAgwF9
C8sEW4LivmKlJ2flXJQ+vJXyuQYtIgCebopS7KLJg9fbWvrxt0mkW3auBR7pqbHJblYO30lyDyTv
u+gKAC5pbm0Ic8JsBh5k0/sGEn2c2yXcDdgYN/OVPbX8LUYacRID/JMoC7eoS3TQyPtOa8iRQgFd
iBKKlEoPPi+D0Z15KdFlLRtjJGIOaCKlegY5J3xknMccjfO/CS1LJ2Pj0mp6zdXpEeTnlrxjoytw
qrgb6f/5ifHuAtfsZVh+WirFoaf8booGOrGh1os9ak/sNtU3eCfR2wRKtqMB43cQ1F+G3zX+irzH
RA0J2m1Qhv7w9Xl6w+RcshvOJDPcWU+u5tieh8HSrFwkgTx7N8Kk0Eiq/J65W30wbbBy9N+hY7LB
fikQABYuaT8gREKQJVuKo+Keo4Jek3RRKpHPgwOUy4e1Gi4KGezuhP8tcScpU4dw52jhxSuahj9J
I/pW8a+3L8hy7DM+RcdxeJC9MgDzIN60+I2yxvPZJHDW5Qi+Th0N5yn0gKz/sp+1r5h7++zo6cWw
Z7K0bRmC/7QRsRpCws/xfME4pwgpEkrmABqSOXHp/ArnkbApPeSngnSki+vV/QDJwlW+e+SE0+o1
slBuLEFDVMm84WV4YlZcWJc6KLbpEqAQNIUmnavvqaMexuG6IONh6daz8Dzr4AZptNSErhTQmcGw
B0NEdv0Dqf3bGMiuepI1mZHrTKRXWJvuTS0gs4ewVDWaQHQ0JdMYED/Zrr7EoIP5Av1U3zORNgVl
IC8pNxuMmtHToiA/KTVQwYGntbeesKxxwCHs4KNQXxM9g2kfiUcM376Du7BF8EmowTeksKQ4Sw07
D5/fOSrSdCy5PZ50cl95u50uTWFyTBvq681A2Urpw55WbLXmmjNf4GnTGSxJwySFVXPyk/ooQH6m
WZX/3ybigP+obZgUlDjwxUxr9FxioWbJnnrst2gcvD8cPuOWglPbKdVfB4KFHzhAfCi/dUmzqAFX
N0O7LLrU2uwJYtSHNGFOmvCKoEMlQkCbLR32pRPHpAGEdF1ZVvZFsUO4PjoS+p026zbjQFe29Csz
Ld0oEtbQT9Xi5sJkAcun7xPxViaRpKYOJDwNxJlZQqcxvSypcibhwAymDcZye6W8+EI1DrjibVRI
FDZTzlXZYfvUw6DN/EPYu240HFAfXwz7fqcw22Ax/Mioj/zjLthQRvfGA/zuCm1gFGiWIr1H3B+t
Lh245L3Ih6o9VeBB99K8aKxnVRA4sD/W7Jc1zQNCgipCEJCIk9M7MBk7K/Yi8xgFJyuc67Q3UtZx
KxTpLVziMU8p05bTvbuKA1PAMPOhkDWfXwWktx/VWdvpyvYJ+fr9ej2q9MHQ9qN4tILnmdozqzhr
IsEjgEBEr1WIVu7OuZKApLDxrs/cUmyWiSVRbO0fT6E0CAuP7Y5OvhguR1Cj7TV+J2LFsTzJ1gmN
e8pz3/1998edbA0/suys4J0inhPqFBglDx/+fYygqJUljOGKr/NNiJo9WE4zHDOG6lMzVydtrwYl
nIWIKrZniU7Wb6GKqmDn2iRdZxEvwxeVBC+TEqMbmhzxs95XxvioANxUUJBst9ln8ctY2lFhaVDR
qDPanRbbfULADvt8/iSuSlH8ztRovf3HXbzo7/TfwKzLzUR9c6KMgLFMgho2F3MY6U239yK9EcgT
QRUsnXmcGg/n//Af8hjk4ubL2F5FKt2IBy+VoRog1pYqKGiB1jHwaKvTUhwKD+rwt1EhWeVnhrcw
9yFtmOV8v1mjVNlnNPpqEveOn8T13KvCU/+UJ2rHXyX5TGEz1bm0D3+/OnKUqr6V2c/IjCYWk8+L
E57OiE9OiFwUgJek0qR1uPy9P83RUMulQc4qYGBwnOzYxeIYupu3eHZqVy8sxAL3uANPhExONiVk
L8JtdN3SGbcuvYLunKPv38b+SeAnCuVIhvbU1mSIfJkZxmwThtJg0hvZvkw6TVpSeMHZxCGTP6MQ
H9ulvTkqO/48ID948RmwK6ZX0VDMlyxYRmLM4xkoXhDQsdi6Zi7PIsiEwTH0OEIyor8FGwZ2gNLt
0oqeBE+pV8n5pp4BpWWvzJvReCq5qq+w4jjhVHlRvr4/5rzMyKzsvdQn9f04SfcBFaOMw1LYhPvb
8xnXvXRuohJolq7kA97rKdkWI82awvUnQ11sgaKoUEzzUJA3Dv7pK/HXiyKQH4QzE67cMv8rWIIm
PofcnXd0zsjo61AKUycOTnUy9Z5B6C3tx5kwOKbeiulMy+NpNqDDxVXEVb6dUFjlXppW6atERziw
r3O9CtRuRa1rHHTyccK+YEEX8R7FHoxcStA+t/M9hh9xGQ5Dkb+LMOKo7lCYQan5mPJpZqhIvNxa
v7uSV2DEngPxTuGcKEaT3GX+i3KURZDwfEExR8++OXShIR9KHsh02Oyt+KISezRBmqrC32FX7Rt/
HWn5OoE7Fwmja2weRH95To3dnNHGDb2MUhf9wtbAT/dd7uu03GlE6dddxb1XboF0Facnk3y76ozV
RFAZbW8gV56Z2aXOnV+jdxYDVowUEY04esU3KFfJYFpwJtas1CmxtAi9VYAo21s3sRguhE73dnqv
qkYvfiGPC0MfjHZOuuvZowbUnRxMvlfQz1rDtICo1geGLlcx8V341C6eZWWTsWQANp+Qi37pK2i2
QcC/IDS7+ycSkw5K2aimyNX2W6C6w9SyeOVN4+ogMDiz243vzoYMO9Yd+hPGGuv0HWi+DdlfYC8s
/mq9u/QU+wHjw1P3beEYhL4GqmhCAnIdm4bV5i2vh+ky0cSREAMTggt0TlKdDMqYRBo8RUYhEGLb
a2lA/MYmyVIKl7aAx3YkaUdc4TKBQ7nzx6bjZEEkbCWqxeX9B/JRxjqh+2Av+QjYMdXkDBTsuFx0
/B1WrWH+IRiaJ2OCB8rCSrJsPFYFSEPhZEyLvvOyTtVy5XHnGCwyCyxRArbqN73n3EUPXCXd5DlH
y2fKKWqA+BWhhblWyg/A5qw8/3kUMINmortDn7YT7Byg5gDQmDECqn8uyo137Eh9eDn8+teI/Nbr
11vnFU4ucJVhkKByh+Pba8xhucr4rR52AXlJG7Z9HHJQJCr78HyqvLY6HUmuYW/TdVjDbPYKPIYY
7QA17FlLpYwkx9U1d7g0vYs89wkAIft0bGWbP8mWyw2uLyrQT7KnkfiGEgsSxZ9rcXRnMsfwN2bH
mQ/K9b9W/XLe7I+1n3PzhlGJqfcEFc9OAzlxsyF54IKHZVU4dihE3BvQnHCEo0hCetjhcvJ7gH6k
WSvjuc1Jyk81kdoz4PxIj827XZrMO7FKk2F1JG4SBnUFa/vejIS1zY0uFxOYDy+0Oyq/mFz+0d3X
HjqYyjn4+A8+G/ThF6er9anQ5SqWmrVoZg8YnUvI0RAfLp+SFLdNXFN3ZPoZUMu3RNPshpGkLBIk
RuQdmEzdRU0mLUJD9xWp67QSEqMADu9YV5Y7l/LS1DKOwioI5wbnwZGmNwUSk2x+afuvrDRVux8X
DO8AUPH0S6y1wTm8wi+HcqT9ryJ4+t6OHJqY5HpRTnU50xuzV7p9biUP5Jht17MXn7j4Yjud81/m
9o2GAEsWOP2KYgLiPmIJ2Xmk39BPQ0gc0f0Uyo/0PONM1IeP0etL736QVkPbO7cQgGbYNAfTSaJW
5VBmuvzzaUoVnclBjQahqf+1Xz2JBuEVpintGjdsK4Vi811Dkznc/knbvyEPnjIjSWz8AsHIZ9m+
iiGovwAH9+O6LaJivr4dJJh9gg4RwpJptCyJ4bam5QvJh6jzCsvTa2hqK62tkbnGi6DuchtuAc44
E7f6ISuq6F3K4pbPvC6nwngFpJ0hVnYhLqk5efGgfAEoKQ1BM+UNPDTIMO0tsC1bs8PBCzKRZ+2w
plqOaexUi4Ub9F6hod7dU8A4GZZRhS8M/BCInU8YBsaFHjgjsv4mmi5pr1SD2oqRX4JGwBgQECZA
R3l6JYik9gQH9LHL40cy6eRaTnY8eQODv++7EnJO6L738lxU0k7Nj7c0rgbDVZSIjWwIUEUFqIT/
nw5/Mpol7hGZQJtY8RibOk0+RuF68gGLo7ZkJ/uXCLjkbYQo8J1OcB66lSqxrmG5JiStBb0nlVsT
g7pDTNnv6KAubX0I6dATtb91JkzNnfa6Wftjl7O2b9GUFQWw+77PB1juCzgQCd5qz1T6Wkp/muak
RjNliwATTNuuLqHq5gNwTw/3WdJl7JUNolc2yyb/0SH1sHM4MXYSV9RcIbJVcENcOeMluQRiMh3c
/J8/uOy1QgBtQbFH0hmW6WfRmKFytfeaqc3OgFm2qFk5CtrAeCHnr1+PfkE1jbjjyYf2NtQ1u+3L
Awvnovr5EjT076dskc17wNOyIsQIMitfQNv4DoZ1Auccs+WcFG1anPXhignJsgqD++M6NJCsOdJC
Wbd+W87LjGBIfBH/phqngKHlFQ9lQps4UqcWTRmpJ4jJrI0FtL3/NHJOlBWRSPgqjhfA/3F3z9k6
v8U0lqm9AeiUCCBoFKL/pEdbaLJ/z0yoafSHMPSUfAVtrhOxDN6Tf+tul8C8RAj6JOgntMsguELo
FTYI6ww4XwQaTx0ksk9xEnhKZ6rU7toJ1S1i91pVpodf8eB/nM6bmG4Ur5y3WB7G3/0+KRsWIXe1
m6wfWewE1LVDZ1gvo5QuJHsQP2Ax1BOmMlnCCVmx5ODoHFCzq60fjvZWYnbbJ5YwPaE9Pab5Xq+k
CdtOne/LUpfYGO+QWuXY/hby4i3HUc8vG9ty0OhemR0zkZLMILE5g2SDj4Xv9fxtAr8jXQM82JtV
4omIIOorkB//B6Pt6xlBcFS0lNzR1oB6I4jtWGvJssaF7G36zPrABCw/aMXyVRQlYbvwx6XqqGr9
6csrMX58HGmAgWG2ngdJRHqSTO6qjh8fxeQoH9/Q9EagX/651Xdo/68q3xhzXX9rW1eTNobjHQ0H
4RmmSE2hMo4bH1b9VRcAo798bzVH6+x1FlrOE4ZAs7awwA+hIogJoJRk66unxMMJKUpJYbv18M/V
OXbX9chwN3g7TM/5z9jVMi+GxYS+3ll2WBgU6AcWoUl0IbaLvkaxm61z6v4AQzYD1yH5MYXUu7sw
/3VR4kU3dQfOJnu1Ue2G6h/LntPmL3buG4u1MeCmQwOb3m5g9sq1LYCOnDpDfYm6cGwZT4348PSP
AivxNPsMAUFmQcXacF58SeQS9YupJ2H0hxfHWpl+v1CKxj1Jrnv11MZCKb7rRXMz2NTm+drfyd/P
MBC7Q4BUMEDJSyagLu2g+HFyzH7Vt1KYXjarROERtIRkUSskIhszmkrMzFMo1uLRHflDWViKDR8T
Y8QQVczLMxKG+1yvVhkYmz8pHGOg0i8E6wuDymNqYym0HbcwrmKj22xJwXvC7sRZXkCyaPbtw7XO
N9s+gZSxWKnYoEe82+HwQ4KV6Eu1S+iZJ/Dp6s8uvWMuwH8C9EbDSaN2RWX2CgB8ETIlWoKZnqzs
+l7041hfsFeynaocKMQNYQjatULv2UvBMzjhSqgjQIoj1kcMWipRD52H98OihrGU+FWkb1QvJaLP
lnCc5OMM/qJthHlDcLOqWtcmxN6YAPtMZj919/ivFHpIZ2Gj93/UiWLgQYLELpIpn6EuWcJomFwV
CL05KGX+yql4sJpKxzi5JTVh5ungGjh+nb2yE1ch/QqnmSxP2FWMeA9JC2JOA9ysHrOAGgKYaD01
KbzSYtPjrFRmUWfRrxoR5+nu/zCVnKYDbx7MlHI1FzhiqPDMxhNlW8KGQZFc12OnmkzQvQ5GBs9g
mG0SyfPb0Fgr9/y7jpZ7BnwzjL0jn1plq4DBe9zBHyb1mgIULbRy+eyVv0vR2+4egEY/u/k0lqWn
kAOI74XN3lj6ow8avvfHCd7uFbQmgOPR0/Z2Zuia7tvi7pJOMg4H5fR01BmbsEXBlIK7dNYFi1d5
qRGo1KFCo9oIeOl1flbcbd1pQKpxg27or22A0G6dfD5oPQnoPY3WdiULwXs0yr8eUs34rI51A3FW
0IsWk59MDNtj/w5iNJCiHRS1y554CYo9NWUOQesQrVB4bdlqFeihdtZ2DJDuwaGuZUCqP4PxyAER
rUZNOQuTK3KcHOOVAEH8rMOHPOZ3H60cLjCYo41Tyo1dfnZLjNmHpANxYESVd0TNW2HTyNVwpApG
B9B6jKo8Iup81q/4g95EvG6ZXYrPKA6gOgs5VpOTX4iLytn2DZnOtah/VJvd7BYJN9tsSsgEm5FO
156NPDCuhJw62BLe/YIGLn7saHi8iVgpJpWszuPzrXciGN16QVsucheXCgnYN6rygTZuJPQ4aBQ4
dcdtl6EApxqxF88OxdHW07nEAFCs8zeIaM1of5VMtmMuAdsV+/YaWshXUtOilMBHHSEiRXRVt3QO
6S5l01D2UNNXuXH6Syq//x6fUqfqaaNNF02YgRZaS4OW6EKX9IPClt1ctSfR7tjbaSH5qJZtDWjG
Dr+oOAcG7qn3n+0+fdqat6Fn1sPYjZ+cktWCQamaG1CHD1nynMzPinBU8ko/2Kgr0wyHVt28PqOK
GvpxPyUr647K5dFUGoc3hMJs3+/rYRHoxlAvsoltfmtIZXdy1Td5mqV6DZ4RkKZYRPomHw1zdc80
y7TXVoA7nAgNfilivL9YTqxmhjpYhlbysRk+AoQEwtbvmMr+AyWqVquX2JDlHD4j/Th7Wl1jMRfG
06cCbaLEs7rdQfpWFdXP33iRv6ibRYww+P3Jc3oLGbDrmq+FqBRTVXgJDJgcMvQ6fADgSqcMy3G3
ma/FqCgiX5NE4TNdUupJ2/l0TgwlD8QtWwgqyBLLxFOBeL5FwkkMZ92qj15D9D5mj2tf4QK6ye8x
m3RAeRlVTr5WGX3LKQgH2ss5EeXGXK6XTipNeim2W3zCE8BoxieLN47Rg54CjwwyGuZOuLJiUzkV
LT+EzsStszUVaHjPH8VtEhLbL1RjVURuT8HFvcuAS2e97MEnTFdWdgN6xL+vnA5AMU6psbjgo+fr
wh5TYEfgDtpdFWCys8PhnB0KKl6o9top4Bnobio5SaNMykDGGF+PWV8LcInOMHAZVq4ey9sDvoWw
UrXcjm8pd/7CeQLd1s2UUrmfGNn3HFkWcc2Aggr1XGCjLJobH3COngWc/86bV4K7gFZAEcFcQzrH
h53Q8daBDgxgV8a/u2bob1FcdbBxdVEyPrKhcZXoaa0eySHirzSutsVp8MrZF/RFc0g7hV5oEI8A
kxR1gt8JY/eojjdcAPjsD8fMY0zdu248giP61q/tFCS+RI2ak6b2y00dOBGY58ZPxoO9zJRL5r0M
ZSdLdsLwYvVmWBR3mEuMRuTaU0LkIBHGsCbB2aB2dZCvX3qUDaYZMzoiUOGWzbNdk7CeR917E24a
sO0112lDA0WbDH3DRGCG7dplTpQgj/xrP0oUN3pF+1xrWFeB6MY4akM8WI7eVc0aDlnsjVxNDKnv
dkaf0lPnQJ7pamDG1Q3/Y2fBN9PdamAQp4ezRahovufSSC3Z1A0EMxwjIDOCpRpi6sOup9/vLWhk
2zzV+n9e2W2p8m8tFrFrYdBSF4snpgZoPZj0fk+8fHmiLfvSHuZBg/ye3deFg4PtLNrVwWj+HZFm
M/0ku3h4mpw2yHdRg/ISuAhPHFpy7uiIEplc/xrwZQNdi9S6vHTDB86mAF/MuvqakreExsWUi5Si
oH3/W5m8giWudk62TcV5PgUjzWHqhL5jk4Q7AWdXgmxNE+C8BopvtomaMqEUk+JGSfusIMwsSJie
eh36EXyoKdrZPfBSrQcfCBx4chpigRv049z6O5rS9oSmUVD8A0m2bjAgFWiISw9RRmLNRWat/RyP
wgSt58FTjmgeZNlpBc9kFYCoU0At7dW+lrGr2EjP/qzsCHXcxsGz+NUk1wxX3CVF4v8jz+O3H3qf
wVjUiyBUNH/q1Q4fNZcd9+QL5uTTxEIrGT8kDyg6OsGOzjzLvYp9SQL0tkxZQTFAnedFPGlTR9lQ
JEMfbjcO/Zem4qQhMRg0es9Al2XQWfr950drQ0pS2hO8uOp5VxfCGRhawgPgKT5SpEElgKvFg1aD
qReDVPlhpbjJRtFQQJm2j2yTY+nxtYcBievLfxAHo0WUG+hvoJlfK86wFdz83xglr3dHxrLM5stR
K+5QylGfLZf7Rg8irmikXBuWpps8bpBYmoCy6psFRddXQEL7lddrJ68sGI7BzEF9BnyDoi8gFI22
f/omoxX+Kfgz57nuAxeR3vKz0/tPifWtzlAEaorS+O7oiXKObZUL7D8lrQjyGWnGkTgJdK2Gmesd
2DGEUBuka0cCN/YkIHRV76VsZ5J/D6rdLU7XMG5JNbQhkQH0C7VaykH2zhaAN0duKAsqg1fZDXUa
MAkTF7jkgDhp+s8yWzw7h++TSsrquBRtAYYrZPlbIqHtx6sjm/dw9UeziDwWK1MlNAM4x7St+yW9
gRGXTAbexNT+PTPR2UKZBwHqCf5qhwPBw9Sw3kMPxE0RYyM49WFpppWIJV0eFG6LVgM6NWCTlUj4
j7k+nvnQjMdkpAliW5hwwOeBId6EFkaGpdmIJqvmV7taRdwT80g6TsdZz0Ur4PSLTCwjqLkEqMLt
L43r8gpyx46ce/iybfGm+T1+Q8d9COHrOvwGwR4fKKcFRqpOHyTH8mVo//KNjZcGO5Bqyot8ICll
MEhuf6FDnhfnFhUtnYuV0wNnUkwNXRr8kHoc6yrAjJwhwg+w4mZauHEsR5OdvrPuoE6j9PPyYsZT
j4P51yVs4v2EepQ/kIK99MKAxLKoAHOuCD0POVaFe1y+VWMlspPvshWn+bCF41lg2Yj6mXfwE7oG
jclr0mkDw+vwRlyaorOSpbXolCEkqhrSuo/OtSLBO6N9ZNAJ0BXZ7uCzr03eXkMlpN2MtacMuLni
qBduwm+9AdPZ5v7iPE0iZzLlBa1ep7QYl23ZptmMm9FyxSHb5TV5kkekzGamyGLuGmHKQMIc1gf/
hbGPJv6dMssLQQiu7IDYfqsQpeaxfRSfzgugClT3TOI40Fja7h2iWFzTjCXrogRiKnwNLDq5NT2c
AnBtr2Wlq7/nZPC/iI/yNSlB3Hv3q+2Z7ZKvz0i8NggMOlTXaAAdG9A4VLdUwAIltJ129SrR3eCp
sPftjPVYPiRBO6xX/uJQEyi/q+blxI2x3k9FNKwFzegmZTUiab/XmVucOZRoWmHg2axS7gRCwD+R
u/WvOTc5ISZbjd+d5Rmi1whwm6IbjaYAyclfrzU6nfeA3yFjWPPsEJrCO5SPZMmwv52hllUFix7g
e2wvBLNRlNugkR9zKMj0dtqZF4sMLM8w34CY9CvLXqzCcOO1yKmDHQqaMkIDKIOr6T2b5OrwJrZX
u4NIQgLN7GfzFQBReHfR07twdJsFhKqKmILaHJ5Qsp+DXA6WtmOctesGcLQ2W1YoUpTNSDfjFTxy
/HXJFyEPOJPzmtNdfOPtsj5tuP+8UAfgOgpod9pf750ptjTGcBUIgnp9dERd/0hv5QXHL8FwsM4Q
s1F/f3agx+Dg3IqUsDd0hMXiaRiumRJ8rM+Z21mhJCaQoOK6QGur723g3cZmV7037EDJ5VbRwK68
qjQ+zVB7vUM0lVF6CCjX3B7ACsQl72STglmkZPeJhAgwYZ6o0mBDzTMNTz0EBCEoutH+ja0gg6uu
mmfysJI+zVWIv01Feky8Piynrm8+E2muGV0pzAYOoOSFijbEwWk8lKKL6axPf8NWdsI/E1fLrzF+
gF3X5Q/6bjlhNDTBo2LxWGu3KvDlJyz/JyPg+MnnbQhLkCY/+3ZRz9nyQpEyl0T/5thwiQVV8Zcg
D/7S2/3vxKb2ruQC/ae8alNTimPOj+Fvmo3M757vIyD1HBl2IR9emtrbyO6ThyA5Htb2BqaMeqFY
B3AXvxfc0IoEvX+RUztld8024oncylJ26Dd38EeiDV3+weuTNOKdq+wyS/phXD2ihmbDgAHf1GG4
JR1tamI7osw7DIvbn4Olgp5vq/OdWGrdrOMa6VQ6IMMN0Py7BT5I6OFWoJT2+2UraLVyH4ewuk6T
kOP+Nc8ogXzVWSXMu67FuaShukLbF9dLktFfXB+E19PXNujBqpws1sU/DaeWxYtNHAbgvOGu0vD8
NxpHDz1mOZ4hRKXHdLMuaVdU9hLkWknSibV+tU0VfdQdbVrh01oRUbV08NUf12LGecYomx1BjTWa
C4Luceb8ts7DGcjQgUpbwcZhFH3j87PAqU/9RsGhry0PFn5Jk5GqL2oggl1ru0XETEPVulmj/rBE
GAfn1uHHJHRekeo97cjGE/Dn45c5Hk9cJ2LuhPM4o5MIUU3TDUcBboTNZ76zZBDaE1h8e6ruiT/m
VMLJeX4p5NfLWstx5Mqj8+gWpGqE42OuVryIZXiIy/tWqFQ3/214mKDisIgoAFg1o7KwM2133O3Z
I2aYaQPdB04S/y0TMYbq1eqa2SLtVAOMrEj5ByFxHRYgFlJhs3QedlgMsj2DFZ1/kTO5WrwJeVH3
1cFjmGShZab70rditSJQySCCGoMVoLlmjJOgWVXYAbrGd6+z0KQ6XKF4BAD76DfUQL/tOQAhJn5a
N0MBrMfl6q09pyhGvWhhn20I9gAZ+QrbaRqDrNO+N8CvZSvrylGISOG3CR9bw8z7/jm6nWoYrgcb
SQKC/my39zP/vMfCZKn/MmHJiWfHok7xNfXtAIvRij5XIxwsfEia9r1nZ/Ez9v1X6J6RDD8GVNQr
8jcAXDFbaeFdDuFpRI8CEJ2uqsgekMPaW6IGNkhnGlP1JicunyyGzZB5QsnEQD4FVBNnmAhtNk7I
4GVwS+YH2Gz/HxSWolMcp5LFZ2T0beiUJbOK3xv5D5aQs9NVd3mAn0stP9nY93iIhsr5qiC0R58f
x7Q21XHggxu5/BwD1ovUfF8URooML8X+ud9/G/xZbgF1mkHC2YRLJsKPA3tocvQYxEXVLpXOU1Hs
UdLc1/FWKx/nH+MW3KrmHao1ArhQFd1/12Sgz5AYMGP5i+DYEVVRjXwCd7j25e23XilrUens0D/i
+J/H7njuVtDS8K7puChpyj8EPkIww8klIobqkm3tC4YcKLAn8/KQtFRtdGmjxtkdRZ72RnmSkT3b
7GqiceoR1JM9Z+RvAA4+N93hOFXyK3k/qpb1nw448ha2cT1sxhtEStPK5/mwCMeTHh8G4c+DlE6H
HS1Ppew0jKtuGZNu7f3aSn4bgVlviDkxOWV8x3Xr8W0c33Sgh0e1dfUp/XPdbBX1Dvm6k4WEZTFx
31fP6Fz+15WRc5ne6kYenCe3YXxyMu/uZsFcJT5toKikACxJ6/+i9ja7ZvYkiGOehpaGv2wfk3Bb
NSjvRSR3iNflX0K9LvRCDte7Ryj9O9RE8qPK1okbUkOsKRv0BwsFLWs0oqvjwukAQ/0cmGv+QtBF
ATOL0MZMfu3bRn6SbTHf8NgbXCnAeUJTp+3Y+EdW8aZjDQotFu1hjkR2GuvXUI/qRsQ3a9E4pvcj
LxGwEsBWsM46LAzeM24xXC7yO28z1LmVA2MCMU/5P/lx4fgUxmm9riVPKVL+kemVc+A5clxcTDOD
/N5ctxvaLgU3JYqcAw2m33fBg4yAv4JwrjCIcz5Bw0R5BUqTW3fvfAq7/uHBsWYym2kqqlC6Qdf7
dWURKZzTvxvuDCMuFgI43BBrxEn3CpHnc52f97j1aSKtQ1rONslldrkEvt4wzUBrkrtjo4JaTNvf
0txPL4eYCRM3vgL/fEgZUNr4O7UpcRE4p712TI5z8iZ9OCLTsS404m6BdhBRHin0MO4YyHvVsh/Y
sM0S+cZYRhVVB64VlXLD1G+EuGlasRmOORKuxyxOEv5rALQw6KPwbrKSMW7oL2o8lfFXj5QVha5O
jpSsnz4a0iru1cjNq7WpxP8NGMaqxYad4FuptGlg4mVC2mBJQY9H40hMZxTb/66Lpjbsy0+LKR/Z
X8zTuqi34006HLUtqwyyiaaiSe4RAdZWKR1u+Vy0VG7b45ad2oTKY3k3N7ITZLYIARFo7rqj4fes
9K2l51GljNK/o70hYQ2nTlVlNiBucmHpoWmGy0NNUoljE/Ce01xDdAjUbi0c/qZ4K5wCPxiThwWh
9/IJbDuejzTYMwswZrjXHrJS41SOfJPHusXbt9BJrF5iUNxCMDxTxjpDKlpur4MWjQDjjYPopWE2
z0aJBI+LI8d1prycjejaRSv/2hRVHRdh8Qxq9ikra5YQ7yx/Oy4cdh5h81+o1qmErVa/72zUofAI
T8v6C+0ip66/wY4XuREh+LuHrR430zjAa8lRk+YUyXuiG2nxTKKNLtPIZiuJg5Wch51lHCv7LdrJ
OO6czkT35wvfXxKkYAuVsiWRVW5iFMYVSWe09iwgxIQuU4As9VjcE9qsSHREdwVenLFwNYHoQJZu
fEgsifZflI5rF5SBK3CBlZz3SBNwSE20AZzITC5T9etUW3yOAT2CLmnEJe0Io5w+Mnh8EEzZPy44
tQ85I6bUrMUD1ld/CwcTau4jCoDw9RNyYONiLt8ap+HX0/Y9Jc0nVRrthHbVOlC3Jm4mnemeWIJ6
DllId8ZDUU4LSr3IORcAdxvck+41w8goQSkJuUYjDU61vNuVfbE8dnaC1a51iinFM7zjS8WuA9hg
od8zfKERYzqvOeb1wG26JW0WjvWHyoKALLuamj5Gd6aHkhyZ1tfw06+u4BZmzztGqTr4RmJRq9UX
TeSKp+BhsBycuZgT+lhTg64lHcRhU5AAJSkCc+wpIxD7OSzNV0Dx/qLlzd5JrVpGXqxDpzCFofZZ
W+Se4euzdozt1AvyrlekdfmOHgNBDnQ9F1uZSVDn8LUK6fbwb0MNXxvl7BSK3jSp3b5NyZlSGZn5
zjDauM20XWW4A7WQyJqR7F/duwzMSVxeu3W2hBWiIu2pU7RzQb8OgvCXA0jDlcNAY7nagBRZ95I+
fdOhc51xsYDIsHkD6b+zYX0P2ibPTP9AdkHByAgEnfLN/BBAh1XJQpkR4rHjZg+Y5K/wn+cpwMhI
FpsdnhwGcpOdRkEFJduHPDGxQSmdY3oCQ0GYunD1Ij87aQNVkKVBIFPFNC54DaQOVpNZRTB8rDPy
FzU2wIuC0JBX4cTP+Y9e6bWAE5XoDDqhVf3FvMPRC3eCZKEpq2DUEpZFfr1Ux/iyCo2qnFG5RYnW
ud4gUeAk3+WvuJia0VWfXV/1WAx8+9tYz5/TI/X2YKDsdMF/tdNNIDG2GMjKqJzu/yoqalQV4WoA
Y66bPV60u3bUXUZvLALXqlV81rbvrzdhD8OBLo7vj1QhPJXbSBGu+ssxi/7rmQEw81jx3/f/+5W6
NVx6x/wwF43PDQJaqcSw/9i0oogVNVSa0hz1+hCT6aes5Jp57OrNZaAAkGflJHE8QsBg7Hm+LOEl
fyKzbKNnIv62UIZELAAKA4Y68Ms3BrAswWmA3l/y6w7CaXj665yeHakaU5TacwsECauyH+P+rf/Q
9QQgdcIDjTp6YReWKQhVta3alwcpREYXqbtteeWlNskItuKlXU6td2uiAvkEQE/OhKTTNQTzdF0R
ABPm1tuzBnocH26pakYMJHAk5CPRrlW5frkhxtbv+336IWRRiZlMf7mNoqbuUBY1EhkKEf6NfYhI
4sIXeq9PfoGcDUFkPfjmTsYyWKdj4U/PavIB26PC8+USCBdYaByKxWS0TjMmb5324vIgJMs4w+sG
SsR+FUwMAnEvzNatAenWKXt9I27xVTy8Lhf3JonzLaFUUNO/gCtvDgK/4NAm8aaLYwU/SnxLr+ws
Ylrmxq9KiRzEPv3n8ApTxPU53KNrWQHt4cTp6V/kwPM+JrOAwvvv0zo7GF6aXBnxoC0cSkYO2S2o
Y6+JlAOIoNe12yVuq6DCCy3ae3xxA8MlaJaqNr2LmbGOUb/jE36GoCLGoPNe+1J2Lsp0spKMmTns
GpSOyX809B4HpVT8plySTYgUwlkGCDw6ad3iHSEG6nFmnrt2qUwrKo2U3XGmzvfSg18f+oU3Mvww
SbZIQAabvR/zGHBEt0PZqhfEl4GJHD+B76NdklomCg9oudwE4XJzEO+HejGofQ3OgxIvPJIuI9jK
HirZtzuicOnPHIZ4silVC4sB0nmBOjdAiI7C2ecIt84gL998TCIwZi703kTNf/gzNcLaCYnfuER0
HCiT4QyKT6BnJVA1aXSD9Lx9DJvrnwSyifr/LWmgGSBk46u6LosB7qwJYJSt5jocn1vxAuaxUigo
l00kxOGuuZ5Fk5hZleOLPTXzUbNaN3OO9m1/tiN2n67VbnKEVQ/jr8Q8HnWBuyGPi4TRwBz6yMT9
U/datwZtH3qPIgmvPEOKBcu7kujoKZehkonPhm5Nbk3w2ejv4RLgsCQprSICe1InjADGvyHTDtum
6erBxwGR8Z+EgDVIv54feQcZKwTVaBd4JbLzRUnVE0+fXI39eaPM9SCvFvE5+SAeP2siF34SVgSf
rpA3g60yt+SVZ7Qb5eFcdkGhImz5eZc82SwEQvmj/AR1i7ULSpljojbGhJXiUeACvLLwgr9Ii7d8
wgtAQkJEuSqmwiRKjs7IQ7AaJbitDLUu3DO3PwQt8VX7+aRJg35qoagWX+FhrIjPL3UvSnpPvrW4
PfkBZb5pgDUCUkKYUXJ6fITa0bxTP2NK0pCQ+fwgqR03CCwjd2myL2bdWEDNKTw/18aG7cBiZa0a
BkFgQM1PVLYBYCFGHpdKjCsAmqsvsvQU6odKNw06nPMAHf15qmW2Rt2ZVXQTiVzZHPEJVpnYWKEI
jTojeQEbi2w7xvPg7i8GfoPe9DSjg0W+d2Ukrf4w+tsm0TKK+IhYKYN/TE8HQYNv49ih7kvLfiHD
TC5Ap2MFe9mYBDZY75i67tpHivBbtRCir0Huh06NND9USJsF5mxio/j4FYOufx9p42WRYifE013N
SGtB1JeXS8kgC9yKX3bRs14RIy6Bv5Q4lXW81jIvwPoWIDGVAFiH7s12wjicMF3yppScXuHlAqGP
00B3tYT+xGvjQw3ZFs1exNBdJForveFY3rzqPKdeujUqzuIrxE95+G7Nxv77QJ/SXFrlSZQlIscp
cJ4/ii5IvxvVB2DJRiux9cTeE299ZOqt0R7L3NQqTtTR5ARgIVgVN34yIijGyssWlMu9XJ46cOCI
P/zgd4kbufPYa1P63GDiCFIOnbo3MhO3w49VRRqYfhzIFJW9ylu02fjPqLu0UWbpTJ1yjxUtVDUz
sWlB3bVda8JqWZvjdM0xCIWxq17EBv6uuAENMGkyvTkQBU+xm8r/994tGnFyFGuWe3eOuZEnwREL
SBK/EPmgfWiU/DMgQyCJzQ5AnzGprRBjUXNR/FvBAAR2vs6UaZ5aqeBVgyWl2DFlB6/QCYi/da3B
a5QYGV56aVtfRIiPJo6tKDZ+CQM2BguRlSIONXvfCC4ESv58JtJNJjTnLpswYWCeelHcNJFZs1Gt
XzEhdeMm916CeHfTp/WWlfThlf/W2Bw7OcskzAjbaXxCZE0AYDr/2OH2WEXq7grmrjfkd0I18HXG
2JnBnHyTV5eVQRLKJzbLCVQSLi6wvaie3n2CEibDw6EniNdD3rJFbGGZsNGxsT6FysU+g8cgzF2y
aoHV9AYbjClrVhHaUw0Gf9ZHkaUqEEOO9dGNMM1UEWCSXKS6xMSyvoYWlEI+Ubvyz3J3R8SK/Zp/
UbInc+3PwBg12wH68MOIJ9SVK9kApGGqa6nAx3Ae7kKR076R6R21x9+Ri8Dl3GZxAjscCJm1i8we
Ag7H7WE5V6Aaw47RxjnEVUDdOWF6OGMhaFBAA5kUxAz2BNHl/YnMPbxV/7dRsgI+45V5/8rwjK3Y
MVMr2QdLfKSwBW8D93+OkncXBWQiz6jkNIpUewtYBiZw5FpFpKYTT+bNobm6Lxaa8ILM/bcaQVSa
c9jqiJTMd6Xy1LDNv3mr2YVqLXdvKtEmCT4mDzDtfno7uun9lEoDyvP+7jEdsF2eeObM2Kiqy+PC
FiaeyBYL9Pxwl8UlPPorKKyE3ceaPb94/2vGxojHY5gG93HjXtowMGvWQZgOPLA77HIdQulDQtSv
qiZyC9zB9Lwpz7sKgndUL0XEQwi5QPlllY8DxeVjVMdYHq7vMkXY0bMXrRrxzUgemoPj8ObLViHE
Ed6qd6lHz7bO1tbmCY176I/Pu80kSfDB+gaAQC9HQJYCjzX8R+E/l+xsX50je56NcTzF/PtqpK6y
/FsnKWuUqxKdlLkWN6fh+VJFPcZgbcGBF2Gqq/52af4oI1mtuUsQ144bvrGEK3qE4I7MVIALVs0R
oV0jpI16ekju9xHL9WKET5lYUcasZGu0eTqYCFIIpa9MvC5Cn3vk0Jb8sHhbPubL9Sn0IfbKFk1A
CJcsGKRYi0p9Xzo+CKvi/nJdjhhc3rZExL5fQosmb/edVqVwoJxnS2Hc35ZPVQMwWGTzAvbwpPD8
qFX5cZP0W5+intQyxFao4ODtni5V3E+ILUkOFzWKtACRbN+70lDqgcnEOpwHmeevcCjOdqIt7rlc
0P6I+5MqS3zlZc+o2F/NQg1YNFqIQHDR7hxbaEbMqw0mOaJfbOeNRDK7CI2AkX/1bjrCi5KBaG/M
Vr7ieQGHVvCM8b6I/IahFm2HT2l3GAYGMgNGUk3911zO9KeORP2vEEeQIpd8mtIUm2rWgy+t2QLQ
CIUmrVxaraFo/dZ250jieu8B/3bN8fpP+ca9z1SMiCi9DiGCb8eQhfyZJr+POGlpDq/YOBZDYNP/
rE4P/mDMz6X3mz4qYkNdGgnuOnW/reKwvfmJQYIYG+siU/nS+3fmGw+aMksK4Mwbdb2xiaVIhZp+
MNau7H2N+emQ4vk2E1lxCh4nH+hk+tEPZ+5sk1RpTg2EEoTSLzoSa4FulagBfISFtiIule/UUSwQ
whyQdLYaoDcaEEwXGNZaJj3P3dGgXrvF9ujcRCCNtHtq8KzOl1goon/BloKVdCtfsLQTYV4BL5eb
XzlRVHE2C36DziEpuxkPJXomjblkOQHv/MZ9cdW+xqGuBaiHYGA4GKpPcAcgwiRZCeCsk+FVDx+k
OklTch5YswagpPIGUnI+7SD/jahevH8LrHf1+wnB/rRJZ0SNovyxYA8ZsuM4X6s9P0gTMvJR6aJM
V0qljhqBwxUA+7bvi9IVsGxnCD0osNle7KBzfhsC42xZwl5aObbWRiKcqcD08EhZqigKKfhBVj0W
LmXT3l1Iyoz2tZ0gGp3XGSPwUYrLToegA2IDdkxKcjK68OXnLjdfeZe+Tspa50jaj5IcM1C8Xoih
AaM2HdvOfjWFQrE1ditRxFv12mT6RyIpfCltlwTGYz9uL/yA/QvQmX95hs0F9kaoL1tjCF+/v6n+
ivV5lpLx98rvfdiwyXBtL9vu6/CC9/Wcza26Vx3a0QnHo2eyLHnJ8cb8ef0wNWVfkGXYqQIKH3Fy
eqOHMlCnWCFLB5EP+0PTQ5kBPxCR5LSkbDiE1k1XQqh6uKm+5PUIGE6+bkJx+3XKD/2FyQyojLl4
6nZIFmxFud4z5VvMpsgFzAhmshN8VBf6r3a7hK+tgGVMkSgML3BONc3T78+nlxVn8bCDMQstsrrd
EUMbJFYTEAy2aBPGag5kd3sZh42OTzn7M6hMDIadcih7Obg+uE+4twZxByPkaaaaMgawP/clBmWc
Zr+yARGjQkhdaiU4P8x+GZPY8lTtFl4NqY3uckECmVd86BGQ0hWRlZ7G80O4eO7CUMW0rcwVJ1Ol
omWRAuRk5Fc2GFZzB3yMZRTWvg7uy4xuDbY4+64uAQRmeNSm+xaMeRdiywGFh3NoKnVdM90fgCN3
fbZV/fZ+Kx/3k8/0mPZbA37UhG2qykTPEJs2oivc2RO2fG2Ji1Zs7Z/V6IMf+exE5OzLc7x0KHjq
Ed/KxgZhz1meMr7Dhm8MYzX5b82BtF6oKMNbLyp0REG+JiJOamdIGV1QjsU5AcK54sW/rQzW8olF
FoHrC13SHUgu1g0NapF9bjBmrkl2XeO6zMuZM1KqV9o84HvzMi0pafLR+ax1Bk97G2NQYoItuSi0
/Gz+/yBcDa4J9Qq4UzqJtZnAs3zuif1kSqGEudvyXVklbwNgfj/y25w/g7qZCAjyNRwMEEs/Ia5E
RHOxE1NscqQhnMDdHHwxAp8JG1RKKf/nsS6xeVN5titrVHuAC+twnjG9zp5UPbPQXbtVDL7xrG2o
baAOW5AstUe+vm3KSZZ+a7QP2YapjJmaso+NIPIKDrjhZdr1ADtl1FzFNe6TcpSf8QQOc+V44yqe
D/5aBtGrflCdxPu4dzhkNVtIg3yUAToHGN+uu/KzlXd3+JslvS3JbJjTXDmOpn930zrjCEAf62Ws
kDkSKx5lup6QoAW3+MTlK4eex4qmKTMV1vZAQMNt4aZGGxgU9qMmqOmUi7Y7ncsJOrjZVcH/2fKv
TtKTmtD9MxOng35UahaXoPdU3/uRmaTWIcEV3yzWtAnS0j4zGi/BLAxq92X5cdjw+NFk9IO3hteE
4YmECeu9PAJV+jyW7qMLQfV0rVgNXos0FolJEcpnryqKnMvZJkRL2HoelZ1qSdAqNBJfCwX3Clp4
2+b6zWl44k6bpn6w3II1rzmXrLDMNIOVqyfLKwHCpxuTrSFi0NVk1XLjLOshnG3DooWeo8AVoCU6
YVjY/cn3fUmbvVePIPYx4AsDtb36HLVTbuPMRziMvZhFlsitNMvz+Ed8qKeJgr/F9KeWT2p3/7kr
GTMI6aNWxAIbu5EWs8GJitcKjRD+0WCdPsuNFVTcWxFTxZ+Eqwdg5pLbeATQLGb16D/8bFSlPMp5
Ewb3FVRj/AsPTv/2PAR8wpKFGXijsRkYOniB4E/S3j+F40NaDIhXboDDVvkXYFaQ2IdBYOLFXhks
hTJJ3WAOzLBlaowpw5AmWyOBlVLq6blm6rYF41V12I+CbGIolSVUSO9UQ4Z9ImmvBr0Yr6RZf4j5
yPMhySXGVvzXVCoza7iFEJRNW6mqZLUsOezpa+eEgIwyWR1h9tXuPOWHA2awHOZ9F/HG+koDwwUB
ZTxZ94+4Zy9zWLtC1JIyWiVB6Yi6cbvb8y3dB3dO2NoSnKUjx31+VkJHGA6rTymjax2mbpakIoXB
Jn5tlceDYUkFZIE7kB6ke3Jh9ITYUhDx3WPFrS0relsrRB5T9OWZ+N7pNwZWKbYWmC6MaPzTqB/Z
mdzxrFO8KWBFdAtBewOtEDzNm4yXrleTEBvTc9eYAAgnrlfYXP3AnwiKppjIMRHOQFlP3NKBDtnd
odo6NteV4/D08jYYsykxEiD8+pJAdIRvBDLe6BtqGNwO9aU0rEfUYpHpIsgl7HNZN5VQhUu+wQSz
fA65OKUw4DM0tyUj5vQ1klx9QyVPX90LB7W/WX/My7G0ugcFKuQDyKevlI0tJuIg9IFNHaIhqbex
6cKw8iy7bW9jxsPEGrE5/mbIqFemw120uyjYun9U8/TUkA3ro3luaP8GnY1B/DjZGDar3H4DQpIb
+fbnF1EX32fOn/7i91loXAy8LgMWbvuNWCHAZFyL/IJPhB/aQFbVHcqCQB+amQOlGof8ae7oYfuN
xMDqEHr0Bg3HnrPPZgmfbEnLKzSdOSgvvbqqiccsAvuDxWntjF7JYC4usJu2B0TeQhtoeipvN02A
NwyJ3BxWHaer0ZxjDi4YhpKWS86qKmHEI9DNaNJLm5N3/BOl9v7yIShKIXUXL7MnOIUWWPqjApdD
FuDwVwUeV9lE25I2rlgHBSduuWRJ8d3Plj3xEbjLfwIGYvVwknGWNm8ANFwYSKoFzDLmrERCKeMi
INnWyP03ma5ddR8Fms7h+qNsGiTAVbsECB8Btq9wmjv6i59KaXMP9rJxEc4TqGV210L5Ti8hBW7+
+OrVeTzT5IGaUt42Twjhcz6A06Rk2Dn5sAVxgdcLUTu34Vqj9g9sQ1OAoK1AUsuMllZ+35HEma6M
+C/iYGWMbOG/vSohSzR6sOQ5zxELE5TJ/49SBkFaQ1UBuuHP3pRHFhXGBkhK3BjBnkHyR+lD6gVd
Xjls7s7DWVsZ7RSrU2kf30jG3UpXhgmxeY0pyy6MjF90kNhnY5dA+fUTm95PvqVk1DPb5tQNIPsu
yVFuPQ/veYImDW68rId3xFz8AJBws13ucZ+HWFFgcMlpSjY+Lbos+LPLe97I73ujlFF55fLyo5p3
5u2EiNx3ZpKHcdZ+FYywJtDle+47o1sDoFEWEyJ3lO8YvtkrR1O7pch6yCkpDzwG8QzCSvB5nPiu
yP9CrZgYb4BpToss9wjzga7Dz5uc54gPwIrgQtxabZzapU5E9mhRqn7YzQkYt2bAq+ruIADCz/Es
bXjmCrY15QIPZwGLgSmi7Xj+VL0M0g8PfyIpdMkHiOEwWrjCMUJ0jHtEDcW7f+QL1WQaSGb+mHIu
jo6iv8bMtChmseWalbf0Un97UHhHvx7fDNZzeI31QpgfAXogP/DPmtVBhFAb0J3sjNaFiidmtbKX
X6ppSPJ/AbJC2S6MqRhsK6x39PZs7kguyBk8kspPpmJBvqohiwoQ7ZZiak+ldVUUnoJ7wbtmKGTu
gu6dj4xbKvb7Yc1ynjZHylk0TPua9DDksJIsHk40gUmubeL2vgBa+aorPAnCelP4KaPhDdyYI3cb
+b7+JIMk8hqmBLy4FughSAoegxDh8doO7Y/Pn7xaFDqc+qUeElmSqNAlB0eaHxLXLYFXri5Q3hoZ
WPSt8Uo3YNUPTnv0NqQkhvWj9kLVeVeYW/+u57GsxXBeC3XVtQGTtH70OxF8ZnwEj/mfkNwX0lvj
ON5f0eiFRjXx2/O6jh00Uu78qpZAqRoYXDTeGNemr99SLjVUmJHV0+1WEbgCrNoP2y12DxRtFqeT
RWzQR67n4+HwtsQs8CdGaXyXPWrn4P1zEiPC+VUqyn88vbH47rzrnYjS/Fc1/2YiPnBmE4u4pWJ7
xxvF4/nMaC2YdsxZhIU/SfWlxZpmaI4W488xausdy9dPiP1JoI/1bpM33Zc8qCVlwcEoUR2Kyk2e
YaGll+k0RLe8mfBbouyA1aDyP+QyLIR3Xa858M1y0hgYHcnp+GmbC1PP9ryH1WR0RYO14MQ2Fjot
PV8miKOC0IntNoKsxCljTojv6Pb4F4iJTbHe2+gCgfxQQaCzgD+WfhiTdB8TNw8tJRePffmnySRc
x+h9nJViBNlN2V19wRr93sa0TVeDszik5UpjssT7nL1wm14BC8OdWrSIval8d6CJgyBPUrgdQcJK
zJ3SUR2nDTVlSi/Wc0xBuKIHnTntJY+YEuqkra6N58GKGt1a0T/Aqt4aTtbylAsrKGwqV+O5oFW5
Qsn+iKLDQnZVfOlGtk1Hl93jkMzue1myHwMts4iAuTz98njSILbWfe3r+xA5hF/KsGeN6ZcrKN88
r1yBIAY/Jis9i6r8aXcbsXvRBOfWgYJRkE5ElQ9cr/6dbVsoaeyp5r43R4gibL1jh98NlEOWxXGH
tFAghZMGkgB3N/IeRZR1fw/basAxvl+rdXgPjnlml7MDKPp945dJxQwFSRLueBn9oBX+zeg1yn56
FzmplyUZ4d/VSgvoEjatFjW44IYw+mKzOtkp9u1/5E/Ae3IdyHHpj6fuOug08Xh8sNh8LzwbzJn+
FkNf2bDb4FcHmLWli5j1BnX82rXo4DNRRupIRaemv+Lr8qrSdCPQGrhg2i5EYIWtTPlK4AdB5d3N
uxt2wSd8UFY1+WI+ljx31H2BPULmiLOhSInJ/vhfFqw8geN2GPUTAW2uRo2lmAebnxw/0tntfeI2
bdjQnvAhNwya1NBcQdLwTu9hWBGo4tbAJhpCXCnzmoeJ9ZV+Swcwo6fkIscT/kyRFMa7zjDzQjZB
0ymUoLS9sI+BXvI/9puiN5aCVE2SP24XYo4IwlrHJMyYpSvRPW1B3ez2MQPijl9ctn5vP/XH2kSk
seo1p8mI/K2YibtEL5VQqD/miiPm5fZMb4+9eXtuMVVluVheF5GNrc6t7nZqmk/31+QokxM0nxis
Mh1cejXKOACML7HYb2IiW4orcbPhRcwS1iuMOuFwZXa4cyxSWiOI2+74l6Yrf79pLy09tz8il7H/
/D7kCY4ZI36SLx1F8UEAfBYBbnl+ARQjBMVVEy1f5i8U8skm7xXnrAeU0SfpqmR7bjitwMLQN3tc
lPu8SWF4pWrgK1teL1vMX5ahRlYvI20nXPBO5Bd+k94tspowwtG41fRB7YWhWUkIIY4igmCK4N3m
2w0+/Y9v4uEakSOSY3e3nU4odU3wLgXzS3wcOQtypc7xEHr2Bvz8p2tGg1Dw6k+gv4yKetj9r38l
3nj6u4aZ9mqLZa+Hd5LG7wji1649LvHnTttXC9U8JnIGdNabU6wIdLMfFrdeQ92s7j6Yod+ldrPv
PthB/xJhcZjkVYb2hDcajxc8DCT7ALS+f6d1k5RQJlbZj6muVWeWsKqS3wgVLD1G8fncdCkcbBU5
soV+9VMQFz5EqFxXR7Wzh8SZ3K+6UBRHUmGQZ6V+hlRNQqx1usRsJlrXE49Lvqtz0zt1VjtUtZ62
FCSgec2SirnlQAMsKTS25vMcH5+B1X8P0nQfNqoT5smjMVVX8T540AcyiWRUgwkYf4LnDjmwDx4W
DkPtx+94Ts/aNUcjZuGwhblUTg695s98a1ek60V65ZC+xBNSg8D+8M0uXJrChhOzZ7RDds4yfQ9u
9HqalhagipqrG86FEDZuPMFcIOII+GiotMthCfMXv1TnQgYwjW4o7g/2Y7q2gromYIdM4VmfLxF/
sD844yt0pa9/xSxAvZS+LrfpfspY9KyzxdnN+7Y9oiHYWyEkW2GGzXC+fHTKDS4M8qHa+Piw+NpD
Qi81vx7csGksszlwb7jDKlXqz8Z7L8iZjKTT746/+fi5/XNj2vegAMw9xQYchHO8Anmb7PZO5JXj
xpoLF3FSJMQsQItOh1J4vncg8oWSnaGkKUdH6rZwslToIezNXUPXxfW+C3jMAvUUr1LSFmDh7Dhl
W8CYELloWT9DVPQkJ1f/P2ZmDdVRWIj27WtKu2FrZe3yB4Tfsb+biSIPmlilDxfcrGpOQYyJ2bc/
aygpws8Ca8iuPZ/5k3kfE0cV+myXGmlGekaqBoW2FzmdhDRhWvVi/DkRtprpi+c2XzvGs8VT0KBz
DQNXAj8sXIW5vRy+fjXGXAaWHUqOUOGjTy1jG3ph1W9PhyiLWWEzhVWX7Y7HmEm42gMUZYpLz4TX
e4McICi2CzXJkbkuxTRJeJ4g1kUy7qZkuPodlNOAcS2cfDbc7Hr6PI6vwFlLXqdtjD3HlARAM59M
kazRB3f88IeuJypkr30KdydGZ/0FvaccjIJLLhM7MyF9tUQQnI9QQ/mhPhBQ62ad7Q2scIxYrkDL
L0ScRem+oT0F3cu3m6sYEJN0HVbq/Hl0i5wUfpZpw7+zksahtf5jXByWLw/ixuaDtF5ShgJ/78jG
lqf1NtKIr12SALUM0YjzBukMc8BZw+uXR963vJkZSWbZ1xp5QGr31y9hUKtOK9dgoYjLRUTuhvgN
zr7xeMfDRoM5jj3pc7lBGDFBZcEjbsD9tfKuiCdddy8dEGxI9ihFWnbgSHdzLQVa+U2Lpaj1vzwO
JZAHbxc5gD+leak3NhoYJ8VuHNbSEn7I6wDwhfrIALYDZrkv/tZzb21MFnDtS5zOTYH/jdIZiN2t
u3XPlPPwYAD2Tpvd6BjBto2Gwv6FRDA9e/uHvsyC+T3cGO137ZFnv8uK+DAIDIfX26dRdvLEcM65
6xvG4BOC0za308our30bPCxN/xQMTz7CyyWqUgqO9LXy9vlHVdIz6OG0Bwyyr/Lme3SrI+zCQZNS
wCafpmLF+fBSdcR17ZGSkzI4nhkgVWtTPuxV1Cf+Kcj8m0JgcsflAsdrQrYxZMyclrLLeA3oENOE
Kc0Dw5dH7UJkAznKLf+VFzo+ItpgePQmySdHrQp9ZEz1LsqdQPm8KrfBSr7r76H7+cx55B5PXwc1
6CEdMiW/xlJ9Q1NZdnwuZdrZl9qPslNQ8QlExxMWy6FQh+EXpfJ/+JmXWua4GrfUDvEIYDAOk95M
4HPr49lDa1X88n/qqKlOzh5oh6VTRtLdx0HNkXxN+8RmJHDwmR0QK0YY8mD+v4osY8+QK+uSKFUA
Iwv9Nbqq1kCNZZn7ba37Yn0Gwu/mjUidGD6BJZM8qv3df4VVNZX2ExUCXUaGilKGjz1o1wbLIlkw
NwUaJa/4I0uy+9mHgNKkZIQxBTSQYNBZYH73ZZvQN5fQf9Cuj5pNtFXLvETnLM20/kO6iMH11/QK
Vo+oDVvPiNDoN2NGiL75N4H8P8f4gbnMY5jUbYtWIithujKTn0hZJPITxrvLyRgZ7ynk8CbQ7bDh
I+lLfK2Q7HySzquhkzeXu8SdTwPAKTaN7ploPyZOw1QjENAzEgo6ZO7C5uo0Ci2KEIAJXg4ruNM3
GRsT/+SPlHo7v2RQAJu6aGD2GL3HY/Bwd/fHEHeyh3nsbaeJwTPQObQq8VZJk6mc2yxSSYJ2PeC0
agm49MzIVOf3R5dPi5z1RFwekvryz8ejH71owkUfTvT2kwszoe+t4RmzwFK2sSRkYHF/7KVncFTE
ZNUBH42j0AldnO6LM8twCo3V/idKORuQqJ9NKIl9tJCmmd5YNhwWD6+Hp/fxp7MXigKg7Bk9en2Y
QiFBmjzBotJrnirCd5DObNvgv/RMG7MM2cmi36QxF/Oeqzdk6a6oevrvc65mmW8FqF2n4JsSRRgR
Wbyxy4qPEaXFYMY5dORHxpcj2SpIGE6oPnFOcpgigf4AeG5sh3ZP2VOn7r/kYL1LsykJZYzMThv6
PbagK01nUTvEr1x08lJWBv53r3e58oV1/i+FfdGatNWNvMSWJGeAYPEzCswEbGPxJVpka7pR5vzh
BkAHs6Iai6MEdqw3pjqU0YiLIalDgmjYs6/eSAGhUROssHg/8kjbTAXfKNVVmLHHCC7MKT7OeaMQ
ve8rhYAwcU8S2D8QGImv5tooUJF4bMX27uXs2+SuocyrBNnOzXhCgrjgCHmQ6N9CCHFurcvZLO3S
S36bTTSDIx8DeADAewWD0H9+/24TxlS7ABul0Eau7BWt6TZvZi87wrNreGWL31V2m8KkjDLi5jxG
igFocTFErqXsyWOH2/yD22ApvY9YZJeABHBqtqDtKnAa/vWsFQ1wCbHGyydwQMj4MhBUgs1eHSY5
NVNn7WYo0USAMe6W1Nz8wd1sz4OkzzEEwHFnWj7tPQGvMhM+BHKAn+W5dXIBbm54pdP3Usu7Wu0j
eVWXUC0tbTq1v75eDIel/TsgihJmabbP5gBmT6b4tD6gmESGnuVPPWU090zwCgjUoTREKKfecUoE
BCNyXCzFGFsrI7lAgV7+rPlDmhfBdxVadzQD49qmPGkLjzFi4rqqQN0VEsG4xA/rz0BAtdr/Vz7N
gh52FWSzFcOXqm4a8F7sh8dkYettIsQHz7l8t3I0jKCGPBVDsd343rksa73gLvDnc0u/LF+tvvpr
L6cT7wkXUg+x8xu0WJf2OBxh113jUXRyGjG72t3mbg+ZDIvb9MCsrLDdG/eUwJyumoc6lTm/+Abl
4Of+ATko8HsEOJntudWI294wR/abRUR8JtO1L8qSpGRfvJIqO5yUc1oJZODIf5nwTBV2sIE/TqxR
kg/meoTGTbBhqtvxmptuCSt04yAT7AzoTXQqh7JkWAP/wlUTQgHVqMRnMpM9n3hdVBsgq+2gSgPH
kjUxSmQvf/zCRPtGcf4ZOVHcZG+q2PF4D+H8Ai8KWalitfi47CBc+b48AoVjKnNqJDvwpXQV/YC0
INdcETfV7febqJ4+hF6W2Ts3HhPcO3Rw8k9JeuitdWC8/2F+gLg3gusZw/0yOMCMG4RnOyD1Hj6p
StB0/AWoPWrotbbvVbzoFJNW+VJjJ2tHZUqHEPMwiVf0JqYtfic/mgj3hKa2ZeXIpPGMqD+EJulI
FXQDj1w/+9/PCD8lSwjHL5Zk/NkYylKrKOHJqFQgjMHK/jSfITQHoz/MvWvaBxN0XRTiVvpCGOBK
ER+/KsbVpQSaQFauiKZCP5qMozOm5v9Zn7CACAJj3s1sqaQ74B+sbOu2dH0Z1wuwiqk2WuaMoZwu
C0Aku5Q0IvaWeidBvaplXHIYsxV6n0pS9fUXKRkjfOTC7GxKnQvLzM2/0LH+vdOiR8CYJinHDV+c
EnS8mFRpmwPXRpBvrI9EDQL5nExMtEisTWz2h8l+lLKf5SQVHanbIL8s3iZOLnu3LT2aV0rceXWB
002xNPI+QLQjdY7frNffhIRJCaLxRuYfugWJVkDMpMWnG/+BXXwDMXUyvzXwNOiCTO1kkJJvPyHx
jjPDibWs7ylhm1Em5lE4KRrD5+sg+gVSHJQ/GL/YPdKazYEzx9iVuvo/p4iSqW8MmLq0xhFvhN/4
YIz1D9gpYZ9BUXd1EqFp8clYCKryPKrylXx1Hf4oV5NAFA7rdQgn3McRXKqY3rY2K71LsuktlLUI
Aim52C6hMSKo/9yYv6w6LizE9sW2oKIE/7xU7A7jqetunY0XUrk7VvCun0+TH3E9/n6TN+NBbBJz
1yEnpFVJowxAQyVylsSZw6++L8wkj4A9K5A/+ddZu0ZOWTmotzRdeIe+8ArbLmjyfRw9d5hpwpNk
+DqFV03fy2StbGxX/dyWbIxxi/GgZkGnO25f/DCmlpPtCRdUPZO4jAvkAuCQCu7H99nmMf5P3Gme
09u1LXKvuJrehEaGHsgS3VL92MF4subAkzP5BoOrSRv5Dn2EKsKnE8UqaG7v8nap359C/V5hl76B
3ZL/uC3qbaoDGPcOEyTwVHm6lOWnt3U8G6iI1M3YUEeDBr4CoaTTf4DQBk8s3NGHc8JGx7sUJGZt
Rva9TL08Q2UP5BZRpvrsnS4svJhUFq2MwXLJdsUF1Vddvk59W5F95m0+4PK96RFVNLGwalcPt1AE
Hv4tr/mo2+YPLgzoLkyyLuBrHSUTuv7/7p7md6Lb6OPthF2vis0o+eV5o5EXsC7YdJlYalI4V74P
tFOPcbM3dBx9atlZ/QF1H6TzO9hsJUcynrgnzYvXvPKPOhZe0xPf/Jp1I1WgY/MUXlX77KQZKmMs
98TdnRZ8DTssj9x880+/y84QmHVYXML4jh3PmGc2CfUn2W+MUl4gCvgZPEkIlQLg3fbgjTPr4KsS
fsajInQhvGlwrin+uf1pGdpInkS4NE4ZGZA7Uc1FZI0ByaaWoJUOWd8+2ksxN682ZtmNHwi3nm2u
mKCgKDxwpU3CWTNnIxS74MXqp6mHUzR5fsuKoKQk8nkKpXH2CmVXip9uUDa0fGZy4S3+QC42kf+I
GoqQ1mdQLLkcMwKmwme6CWIguvnIDxVJaq9s+Qy1dhieIOWZ/UCAVG5u4NUP6Qh9p8Y2+nH2pGKX
HTBEZsTzUh1V5l5dHKPVpCOPwW6ct+z7VWSXaEEOv9A0THiXRNRbT/HGXt+LI+AQ6laUbqzyDD8A
KCbC0P0GKGl2dWk64oSNP9mnqI7Uxmo+98fSTPBLmenO9uHaLQyWH29tJZciYLF6pycGC3nNWAIF
ZmdK8zK1LoDwy+4/JwdcojNVBWDTaPJN4mFIABYmqtE0UkEJzS2r0rHx5N7/3467Ig2mCqs7bPjk
ZHlwBjNBktqPdGwco80K/ebdU3aldmZITK36Pv/HMi8dmmpnZiiTsfT/pmjNSQE8irHsj0CA2LY2
ugb7f8qOUn5hwFs5RjFExuWyUFTGLPT/GKuOVNnpgLCP3EFV4enI2NdG7nxcZNKDSir7j3a+vfjI
rB/8tm0FfZ6i8SW0yYIfQVZm7GUctjDda4a/0zryRgek/E4/hSnqoJyasMpyTR6A8T1F3MpI2C9x
w+uXdcRV7bQgx1t0s+AEPQBmhGEPao2KhbHAXMc3SrY7gwamSlkNVySDaEz5ow+Aep1KL9EWGSMK
s92UIvUq1rwJzWYWv0tYlLWOityWXZmj9OxJvuU+aFfcyRBvlghBxKICMAQHaiEi7GyX3KwdOJPV
/lU6UOagTL1S/W0EFy0DL086wwGyma9dVzlZ6mJ7JlU5ZXK7vx42gUH91oYZ5pNCapCHQ60f0lXX
ioN5QhuOSA5WZMy8JL0LWR4Dhcyw7nMv4f3Vum9Duia8a/89cG3TqZMOTl1rhoF+pmltCuQNg8ud
UXflnNyKTZR+Db81/XQ9iFDrdgfLkoUOhgzZ0/+rPNETgmGIuFBXbjCUwCUWK64Uv7vHbvBkMaE1
tzor2w3Gv4oOxThWQxXl71wSuZ2dKP0766c8tIvDYlWjyBRGjrkQSs4LUGqTmsTLU71i55uTarzL
Y0meJh3f0zb7DPvNB7xU2Gd/KMpqeDxPdHlaqH1A09SIkvI/Tdo2InWX4U+NTd03JUOPbIoa+Wka
B74HplRBDvC8f/tesZfB/bM/dxV+qFFUyLniMUU9vIWhJMKhdmU7eTcKsWzTg9QksQ9ecImeDBxF
T1BdYkma5CIf5ce8K+7MuIhV0Byi77AbIabPPjGek/0fbz3ll4jVta9pDbMNpwCEURTVlX7MSnVf
xYGIT/PlLAEHWa8O95l2bGVRvrRnS0SF9QNpl69HnVJHW3Wb5JkXz0greLbEaCUaGwb3XoN4fFae
PnFYgDzVGEtOxmpsUhwygJOCxHrcNFO6UmiSU5Z9rDR4CpkDQJIrO5BXgY2vxocOEMZi7pGmz8/N
7pO/gUJbmcwomhGtsR/O0/nDOviTBLyo64kgqWLR9ApeS1oA4t7TSqK7JrhpOMEt4A/cOaH8WlH9
hBXBuVU37IyPl3ktsl2274eD3j3hOX/+o1hT2S8X0rVZtFI1si/GygIIA8/KVdOFzRJ1Nm+FV42R
FoRfikadZ6Sy7aj43PfYtGHBXGov3Dj1B734Q/X8z9kVpLENk8NwlfHDAN7Ufnmq3Oq0+BK71c4w
ZbszGO/VU4crYmJ80DDYvZOIc2TF4B3BVrHLK8084UMaJV0/AvWrqIp7oLJcOdHRssuNhOanhtN4
nCFbAvf6YwEu4r8bMOkqYzaGs+AnD5uYP6hRwQXU6wctuaNxsX17VdU6P39RP4ZqrsLsE371ldNw
h8NgL7E0laekzTcQGyUYi/H1Xaon6mkOixQgYYF302ZihKNgsqT4decXSjt3gXjiQNDRGHgQMcQY
xa1/V4X5/eNGdRFzuRpDEjWT0DMaueR/mVijwIshwyJB6BreS64lXdtRcm7qwcH4cdj0HKcTXYZY
6X9wddMDnZv7SfxtXNlW6JamuN5TcxpcfMcWy/iyzgeIvLFUtysoBkdOiqEFZ4iQwhJnxDf1HQNH
UyHVJC2hL6xYnlhqD9kuCgGgd//9QAFvVCqVZKzJNrU3hNS/I2dQ8Qe+/ngK+p0y1ZYHVOaQzXS8
xoMwiQhC5su+vSq1BxQEkFWSXCprTc/0BlxrLqMItwrCl3tzCFkHWXfpfJlC/qqIBWcUFMvMdXa5
KHcYPep8RYLSmdu22aLlMbqoybjvfEX0x90jbZjdpJKlAFdOM4IPhAcHorCHpGesQTglukRqi2wW
30GoKjitWaFFD3kuv9bN+UK5Dhc2OuGmabuQm0kytAfmSzygFA1raaEprCzyMGJwbiLq50rm295e
TFm8tO33j85RMNc779D0VsR27iZ8jsqJq083cZHggJJl4jlDonlfPIVgGoSlPE60t1Os8nfrm3sC
Yv2JlzQ+I9H6FaCmxWe/WsKB9xIJEgvYvns1S/BPA22UrSh/bmJVwpO709s9t4SGlwJhZkiet/20
qMRtVBIGiJMb/ACKzuxwQwphE5ll33wlhyZJxIt2Jc1IbaCE/8ZXHPlgc5+fi0Yk2Pn16VNnQIx1
CF3HHzjgUIVJxYokQ3Xhwv/Y1oVKqjZ/TcssbAEIr1QK+EjSoQotv4UZ7j/XJpLsaqg1YbdYLauH
sziTAMuI38Je/7iCXZmUrG0NAjb12X2iyUOZ0bOI7YZ68AgHjnfQjn3qMp4ouAvouoFsBPmLaV8R
tUcHDxu28M40rwGjIc3+n6ScYPeZxj2U/Se69JshH9ilANPuqepBnPG5E2e4k+DLhIF95A/eJKPN
83MV9wvA1j1BiYFxeT5mLVIjIQzOlnE1Iiw1EtSjgBzhxmRGru91Wv7xZb0CrMaJFr19O9r/zVKt
g0K4Nvsa3nt0SunXTvMqTHg1uQkBL2gV/t2IUqeQtsHIcOUEKBn2XKcsp2CPFfnIPqSD2jbI4Pa3
uDKd4oTDnjgmWiJE1b2j8fU9I9v5REv2HfewnVUNdBYRJi8QIdzBvgjGgiSqnUN2sc/uCItkSGMI
NIZntkUNndNgo3f/4SAtYiVwEewfXQ0kIwToiWsG/W9t21XFCmgu66Pzg77uE6x/cjhg5oUy5ADK
B2DAXo24NStfc1yOFcSOxL6TioDrohur52FgH3Kraz/oYn/JkiaXXM5ZVGafcITyRj0pboj3ckj6
pGhb7aBX5UvGk6yS0K4kgaUbcE2V0KJYkOJUZwkXmzcXprLiemXVgMOXhY7fAahUFgHHeTh3ZVO9
TdWDylwxb0OvSPHf7j5FgbK70JRKlC64hk570l+vaxG0O7Fk5akU5+nykOlhRQwWh8/P2FmH2JfN
fSIvtGo/EIAQDRZC5IyaDPQPbgrgmzQQjgXsaJUTfuAi8GUOJKqqyxjH9ZMADBjpUrBI0gDvP5rQ
4tifZdU+3RHiJZQFFhEeQmhCaWWIuHTVmq4Fjuh9hihQzqe/UNuJKUVjxPDcBHZthhjiTOQZhAs6
ehtwt9nrGeWDbdggAm96TWqvpD0l1Hggh1Ep1l/m+cW0sMPxVdNuG4dZ0iERDyXPfONkTrN54+GP
ePUxoQxTBlwEhqVy68I/WkkGestxPHGIrRnBlVufxwY3mCP1Y2fs4LUvD9azBOXmj7GHOgJrahnp
+/DfZbF/+82wkonwVEPEVVMIf2A8PcC07bcmzXQKRVjbUYcnXbTavAtlikUcsVXR9a8VCHDh0OMo
2ss8IVm7gxus+bPnOFliCjrYtmQ5zQb1lX/LrAISX0O/I/VR3zAQs/w1rQFwJhmgkUxNSu0gg/HV
VOwoNKptEI+YvtI54J2nub5URLYXTrZQqzyxHhow+DgLinAZ4emRjCbD7BP19YtZrEodgxNKBImy
Kq2XvgWRLeNvpIz4R+UkmG81xGzLDN/cyCOfkF33RQZev5t689oxJAfqK4OQj8gBwZwLNHBxZdXf
2+WDar4H68UK61v45nx+KfjkvwypoomwJcqWPLLB7/tLGZOx9gbPOHDnHJSkIv5N6BvlOpCK51c7
d4EfGAeQrj12KFes9UMxamw2n0BZMrkKjQkKkrAM7slwqgaVSbX7LNGgb2n6cBrI63ofy/Xe2bus
X+s+6jNcBd1viRaJYHKjfRJhV8Py1vZDOPe+6C58K2hovJxfccrpwwtKRkJmo1ZarsLMH6adbZ5s
GkwaSbhjOzoUTotkRggppll/8SPgemcIM2QJxAW/uFu9yqaBzwrcHLyLArxhNCJpYJl1lTjGN552
sGfDJuSuZsrfw8LP89agpGhLE6F9QjStUrUKzYhG96BnokwQJmCJWVmloot2FKXBRO9ypHTEBrS0
xVosK+w+NsRsIuZGgOfcplwjDkHhtHJM2I7ktHSHdJEdnNmW8G+PnHCK7EWBYZ9gzV7bw2VE4PVw
3RAOCDqcxMLA1LtT+CJL1FP9SXhFiVAEKmDszJFeh5Ch9KGegxynCHciSWULlIUwgFWUidSf9pN/
S9Rrgndvctg+a+C1GNfootf0RdFKORqnW78lZ7b390eIY7cMF3jJYAmqn0XpMo6lvxcw79cje+Jq
8j5JqLiE27BbKQ/jG1va007RThjWIb1IVIrWnYt4s1o/jz9F4RhmT2D6p0Vd8AWstbYfKJvrlTcu
IhGsANWj9dJMFaYCPvFKoBzlu4sW/mouJN6fX7/fyvMMDodD0sEeqVJbT7OcSnIBpiKXUvPu423A
3ixNTTgaAxA+i18x6L7vzQ4y7lAlpacNub45Hx/vbc2QYOILiMDiA1/RAsoFO1AQlbznfyHqT1HN
tc2qoc/MLobTBUs8bk8z4W3mt0yPnCAxaVi9xiMn6SfK0oa9rPWkmG9tEp/I0IGIlDooR/GpDM5L
2Czqvdlo+j1M+q+WoBkYTkBME1MGneCKGDaOoX1WO2KJjJsD8tE0m+KFYpCieNq8rTuOKnZNg1zP
M+QqNPKjYAQ84Dpy+sJ53uoPskrmuM4LjAHuGBULcZEEl2cpSengUhzSBki7A8GvkX9QdsjJzPUw
eLBHua5OXdUhSEzrBXDv5sZ25BpKsKPmWa4qphfnexcxA8zqxcGdAIrYOCFOQwB7rTrIRaGGH1o8
tOnKj9Pr1MtBsbwonwaPMEXFbt8wmoqAXZrxaSnBKJr7n9Y6TW1EVRj1aqfN73klxNyL/8kvJOa1
q0k1E4dADh/2Dcbb/ZADbQz1M0iQNyXCxWFEyz84JCtFhbiCZij0ciidKEEt4NaKvXBWYAbzK/Oo
j0H4iRRnhl4fbiXWiZ3uRSGttbEhONdn4psudVWKZZ+mGhRPWBSrFVzKh1ua9a6680G8iTXKgb5X
iwh73FbB3bJvuDMdRRNSvgpeyvzv5Is9P9dTqUz4wWO1JsGIOhFrrUEFPdXvYQ2+RzZ7xZKGTTTz
l1TyIgSaEHdDl0UNHyaEa8INHO9LulAj20HYs9BbbEdi5vn554lAyzZ7IyW77gB0FLCYr27YtPTs
Wodvvriddzp3a/tFexUVnUyr8DzisgMwnxcOLK4oNCOoxwat7GoKXczSXyYAAc2hdW8LcZBEzK6E
rTyb77CaiTJmiK0wv8XZx6KFsAxA21T9z4scEY87oE88M411K6cPIInR6128yMQ+msuAYs5t5Bwr
BSSw67Z60jW9S2y6T01lBpa9hrA/bWOsK5DwEHM/xijYmfn/b04jL1iH+mJZ8jc3bEpMiypldEvG
05OB2opDC9ma8SF9u/Pl10F7mGd20gjKMvzX/uRYytJA8yDSE30UkSmnliigPI6sCZXevXLP2021
HRnjDXb388cpvY9cd0YPAhvputRqIVKxDE29A+mBgNfEcuMa0nRB99aGCi15aiCqP+X6pK0JBueI
VpbGjPyuM6OgWRzlNLwFAEmFSNKV1vaiA51XQIy12Kz8CmPI53g1Z5QP+bdLTNZohblB5U6nXlOP
cU+tYl631VNR6L0dL7vQgSAoJNnI8MElY+4oYAGmKE20Y3hlh9PpVD+nfL9KAMuTkpiCXUDwoiTO
COxn5F7RQB7FIExgzheiIoD0HYEisPycWhXULFJmvPKEOp7rw3xKaNaWPGjy0X9+KW8uAM7c7v/m
N8FkCxv5CXXu91i78FSQ+YeymMujnY3sqpDM2UJtaw+pRSlJ2A28vo6ch89xkcdUupbXXEGrx012
QHLstnTb7eLqzlSW7UE+1x3m9vtfmhKYK5oucEp/ezJ3a8X4jaJL4mqn/C5iJ2DNdcT9tO18Wp4j
16FU2ukacfAvYKUpLm2aUjhJDj1WHA/XsyBeEKQSUC6S5abChjbVbtn/80lQEsyPLojBfAAMEMfN
YnHRF3vCMnCzdJoMlDOHkm5VwoqIf+mOAMX5l+tn6rxkvs3vG+w+sW8+Ok5+xU5E3rzfEdVri2Hu
i5UdcsSzegDJVTCMQwRzdc7xcHsZ+hFVclvmI7rBPiOOYu0/Yievg2qBx/wT1Ysy5V+7oX4u+rfp
DUILJcH9SxK5zAy1bTJQprf2O+FARiom8gzzdpg0qzrODeUtvvCzm/nw6Oige3gNPgiDOJfH/GQS
I/YWe32Zg8DCjk8CQiESPmCO1rZc5Ps0EOv/h3kk5VInw2BRKL1nCl3nsHwd+DNP5rZGj234KgCM
NVA+4d0NWax5TQZqJakoiX72s+leHxFjdQxBKYQNKLweXGokh5oR4zKR2ZiMYqBqy4Q9rL0qf9mb
aPVSqKYM3jjCTmVJnxPUmVBlCpgAiZX6Oj/1WjF3LjyyMfTYs1LSAq7S9jy+YyAux1VBNT1KxnB5
cKo4jri4GjC4HQwYcIGpuRBpka3PFLXbd+AyZjmD5gKtmLnpAHj+u9jSCBSARG/SP/mK7XXb06fL
ZIhZ6GAfBPgpHWcj1V/x8uwD7D/Wd38E7o0GPly3JeDLVtQRNDTJr5/y4Lr2pCkiUtlUf9LuuNtD
feoryO+92JfcexefOC0VYtj5HaaQKa/zHkUs9Y4NpF+sWwjGOFckVGzDo/h/12+/hoBVEdy9bc9B
irn7prxBSZVH46XZjtH6UVZK+97jV4a2LjAWurmLg3VoqJZguwOAInJ/UbwXHPiRKetpFja+RCWl
/3T3KCh3jWBsKvq+inpJGwzSvYLM8SxDt90DgmhJSadfpPdDkOPuaVW2mHiayyv1VPRCjbzB7Ddw
RAYBGwaq1oGnbZatEveUzzwKhxBJelool31z9xx2ZDHDAhlL3U8abPA6eSge88U3X1FRrynBuMNO
sYsIqiposmsKaulwKaKLsu5dFDLSTNN2wvZ22MZpAkTSiF+W7Vn65HJRakmN7X6V1GD0FGFuODIN
sjzvpwGtaDXJ2vunNhW3RsNwmdKJCBuKALhd6KxZFLUn9pP7MvYLDMpuHY6gsprRjs+1Yti1GSWh
RXtk07mdjeV1SUWE6hEn4F8c389iCM0RrkdnqlpE4uhRMv/w/5c/HyGK72WE6NumhJaNYfJhxMtL
sUamYvDUss0Dqj2dcxn0kq/jkHpUwqGUEFOy6V/7ZBfNBgfgfo3m4N5p7XCVPzuqA+hrAth8Cwjq
NCknF0PAw9w8uijZWTZibph/2Y5zBDbiq1rHqfZnjRhas8EcexZBGtbHwqN0I1mqrUf2Ffax4XCb
y1tU913F/GG35XYAPCxu11YaMAHjwCADW3JGznBdnGzxrVSniBQjhk2kAgRzcl4iLlKz/j+fPIxY
WOygA46MetXonpRjEJW7rfFzo5tELxP8c4aRcJhzzKtac45aABtaP76/FV6KnsEq8jThzu4eDIrc
iygLn+ktE5oqI1QNEbJT5/6fn9GhcR5lWI68FlF6p4xLctJP5IxwWpXAnlCRDUFxLVHpfD90cQC/
N1DKag0BSdYPQGGr1CXmWouAY+mBx3j9mWfZ79mMxAq5mKO7EExAk0n9anyTrMEfUOMTb6RcHNjt
rilI35kIFbri6LLs2hFUjDUeolaCXIi6tmsz8K/x470j3Fwi/L0Z798hhbdGBn+jmsbVHcN/SNb6
Q6egpFYvZgqJ/E/yOYfHzR9/Pi0uy5PLrKpa3lx0rdK4RJWiVeJzNMxLx+vUtDPR909NFQVnj3ml
Os4XTJtE+RxEltmcAc4ITrqMzjVECGCTAYgBdWdzmcgWKxf2vF+0NWfi2KXM8SQhM9++LoePH7Ds
YKlpxqPIpxiiO2VraDN7BFgQmBPdmQIr+cVhTKk19eEJ5UGG/PeeYZwUKZYSPW0cwdi1P0kfyviy
Usl2RvEHmD/kTHSHO/T8jtYK6fffhWKDFMqBLkixTVK9aLUQqFv6Dfkx245SgjBkuIYCEv4IQdLu
9lvvcqE8nwidgm+GSy7/0cw2tOVuc+YfgyuMwEhnEqCkQoev20Q6Q2QPd2SMkUrquQYnBRvjBctc
E52UiwRPOtrHOlJcNWnUGf9BACl68nqRKU8To+yCMh4/6x3f7uzgoFXT1mYfroCyWwRohESpc4ar
dqc4vcOvfCpngMcKDrffpsbT5edwT4h3PNl6CvcDM+icfA/dyMlbX1TbQY40mDTC98izlZOYDe8P
fWNEkeOMZOHtWNs6uymqYmLlmswXZ9zwGsYgwbNDNMIvP2SX1BxhSeFBgkqsRCrdB+IV50YJ5pEZ
ahzDkLERnd0nXb54GyXjQTla7y6TRxqYCHYeHD4Eoz4KoPppN8vN6hT5L8Zr4inK25mIFuBvyoHm
4z65vMaaAbDBRul4zy3x8AGuJ0hwvUF4KWD3B/YJImq/Z19ywzMi3VZEjucWTwrTl3hPNahYIBV1
htOrfxk4atcbj/AkBcl6ZYQKiF//s2adxSfJs//8FASmBhyC8RYUioXJk/hbT0BCDLvYPAiPmcD4
8AABAyxewTynNJuW5rQ9EqEP7bUL7TsdbHaopjztFUQWx1+xxpM5yv/F+uw0R7e8fawZzmIOmAoa
kQB6bIVNfFv3qOlXJKVL0mSOaKp+SVQlN87thi1fjc5O3O1WV7DtDZYRTtk3gNfK4RSWbJZS8zeE
XfRGbMv65XS9oSY/7V6gfDD/xzVDlbQYyV+s8TxZHDU9Dy4ntq71RLRyQ5GxP1tbTvSbVNpwUeZU
HvhfsoplOU96P+9ykvK0VKftfWsOIKEUEXxEXG308EySVVVpcNVS+KobLVjWvPUt9qlp3i+AYGZE
LaNBQtJGUOE+CbkEDAZAz97+ITxl/+Tf7YF5ZjtMpaxYbtHEl0Uno94Gd4skcK2gew/9Uyqiy4rp
VnsQ7UW2V5LLsZV7LqeEib07FmJ9wgJKvgRvS3Ki4s/7V5Ptf0ZZCkFsjZHeeo2sYD+PnheLKE8T
5nhUQ1KidYXYY8gUwi27cnndZLCvXC6wG8hKZlOBvcbi976uvHuh760NkFMb4SZ96JlDV2bZlk2P
uWCCUQGNAn/no2PJrAn7SZk9spiDiwJclSh/0sbaK8MDx8JyH55dFkdsG9NF7amXpGTxXwcScjAF
UV2HMX0p5oVaoKXfXBWvbPryBvmSrVrRcjuSChptRhw3HfETXnX53dLrocvEpkwDHivgWQsLEIJL
kYXA7ZtC8rOJBSSi819I9SwBe9DyMBPsQH2l5KlDAuLpJSf6vIPL4fv5GSe79FA08lTluDKbdpVR
cnw7ufvL46CsqJv7jpZkkp6d/WI6iXs5c2p5/r9DNoB2kZuU+/yQOthRuchpMmRcPFMmVZWuKwAe
6g6Ww+FinB4PgF2TWNsIGaiFcAvYF3KebWaANsoEsS4xqTULF7pGz9ej7Ed3vulqIzNlFhbjjIMf
HoD9eQPk/RHe33zRowN2k2Qcv9eI8A+Bl0uGnSLsyhF9yfbxxJP7Nqd/mg6Rk5KVwOIXx+WdOezM
97c9pt28WQhu7mamEHFvc2WNAdeMLlZWKywg3creg4+TujwqNMoETZXJPmockcn014PFbmAr4ZAK
WZQM2OYWFepO6PTfiYIbNz/RWCgsEgW2Xh3K5i+Vo+QrztFWidMMttOTP1miXu28SHm1L4H0jOT/
JlVmH1OE8AHSgf0rtt2PYDd+nD9nHhLrlfsNh+qvgTlZxl0ApOqIB22EVdHzzTeyOPo/Es05t5vV
5sJNgP/8eWfHY5y/mT0LNi6dYJFhXnH/IoleIeRSVwSJREDrb0G4C6/XB6X3ym+MUQVQ465qYjTK
tigo93SzA3tbgQ5Q0sVWIPK2PSGJ7MRzatrN/0a0tVMLGhM+N3MUHT8BiaAJltR2pbwBcbMKByZC
PjQkZoym3O7NnYnNKrAVyD5syIpLuyG6+Nb0zVnPxgb9MSzhpHo1m2SuDG3o+PL6m0zBbSGyrqTN
Z0aCVClTXXj4t7czR9nfW+E37nybeQnFPix92U12nEopBwdb6n/iOVdOZoaOo0tJXD/qxf92wcow
MLBrvREb2EVjFMU/QbTvuHKPo1msivZU2vO85pVRU1HVD/pKFcfF2Gt6d3+0uv4R1nfhUvJtlAAI
syhjltfPNOusSc2rqHUVkjYSJSAd2wGiqZY0mXAiCJj6C4+7WGjqQmORdarDkYh6WQjNdU0mvEeX
IXQfbSKyto2F71x77JMGfJMht7Qv7V1cbTyWM/obIZJY2x8VNCUP0qOwrKwTkV5vdAAaR8NjgZaR
iaWSZDfShwE49K36iKleL9xB9MuM47m+HSyheiRYnAoVQ6wNFyoEUZGLrNkJrGMNpCRmTgCA8P+L
AZqyIdc6qjPQeC+Tby4RN44PTmMv6VeCF/RSGLkg4cxdkbHgZDeC5kmjRoSdmDe0cA6iqY1PjKWS
45fhnJ9s2SZcH2tGGqv8ojCC46Si2qPTslyRSz0QB3scV2MwTab1t4jHduIuzgEF5oKyZ0zgb/uX
R/M+E4MWBmSxrzCapEt2RgiuzTepecTpGXJUSBeIF3bnvSgC99eKsqSlZAaTT+ahwL4GL225mQP7
pDY8UYRZas+RyGaik3mmhF5Zyce9rKOVMaS6ouzXGX3/npaV0xtEE6mz0c/O2oUAEX1uLBvBHkgs
Czs7kGKfBWP3y0qFGjpTs+q5OezCWs4HZLbkcZgjZjQPHB77Ntug4jUwZxAcpirWJLQ7DkpVjuSE
r6Jqq6qSyDu/q+gy9+2f1EMRc0ZfWHpAHiYKbpWPLKu6dZywOuZcavmLWdQTXSZO50+QTxyDT8b2
xgGZb0m47EF8u/mg3jbS91SHxWpPnPL2R1ogNeWrVxdTYiBMIOaBfCcR73nWVQlmUMX59eihmsLw
EyC/kg6qUM1YmQxYdsjdptawYuSiAUQH9/Eye5fVJ1atXf6Jfu736IgwWI+H34lc/B0ApCAkKrXy
8y9m9xaEJe086H1HzNFZM5Z1SsJ+MSdtigE+8FqUoiybWXVH13bQF3lfCpXi4816YQ04r2Yc6Pov
ly3jV8E1Dh5EDaIVf8aH98Ldiua0dnxw1DPwPOJ1y/poKbqQ9yFo/WuRsF6usDubPz4YrH0T45Lk
J9IYpj9ICO7EaHrHU5S4UYIJ5/YltSk0lH/UY0q+DW6tS4m2/B7fPp7BERrmJKXR2gKziCZrr/Qb
8zxC0SNUI7B57sHkhjteDqzd5oLuWFrsOoSxXp6B4V7cNomA42794ffBSz/6ycG1GTl5jOSh3Cqq
cafKasth0P14/fUPtilSuCdm9MhOAKv10HBKwEpmSkbpdCfCigbqmYuCR1qQ6bs9gRT7E5Ni1AeI
cFMIZyfIQUH4mUxhAMaiD0VGNBbBBd4l3l/1XgRt8iNpx26JTxMM4H5i4T2/bZGV2Qs9mx7rYqwx
uoOmqHq30E9pig3C3FYxBMGvLTuHlxeWGipTLvYgQKihkgLKOEz9Cy7RMfWDFj5dG0fLVdTeef22
MqaVxHjaN7flkni3060j/UN3yWI/NWjIhs+BJUWnqe3f97wmE0DuIvf0ETOJGfsUqZNjXcbegmxl
6XZn0lFp+aqtyDbhFaJGc9bcANtpK/bQMlrmKevxjUzX6NC8u/vwzI+leNCPJs6pQJUPuiHLhmk7
qAk6CrQXjzaS6dU8Q5Ae7UKckiGS1n5iPGrngWV6+ncLAdsqd7ZuIy48DbniwuRr5Y4DID78PpXa
8jq9y8WJFuakBggVEt14Sq6PONSnbrOK78rFQagXxPbY20WP90fyXL7JzygTY4/N6zADjAihuWnY
4/ntLdqBZ5ytdCZUZXNixkFF9pUEncXaD38Ej9rGT3+VgpV6U88nBJNNKU2nW9TRJkrOe3YSepjE
V/vVkO+Mql2GgpJ43OMquCEJidXj36UrB2MiMuMeIAWfgB23b1FEPaY2QqLp9Uf/eNmI/j9SPy63
JHDiF3FzdfoRzMALPTM7Bk+iM4FCR1BRlXOSE6s82EacevxRUQ5BHKzoqCqEXor1/MyiidMjB+qa
WnG6o8+NQ/J812a3rUaMHj1NxrTfSDsAHvJQQckGbGAIJ+eX79OGmaOKtsmBV6UrDfVTO2LAnSEO
VuOKigJKvcYmODNgDMS7bcjetfQhjIceOBqkUk98vctEboZ9albS8ZXT4s9n8bOgSAGbLlR2lJ0v
qnnrcuqjufg2ytZ9V0QP/CR0Stu3e9ix4TnpQG8mcRyuhafh8Er7srEfgMpfF4YWIMYgt2HNyYy4
oYOHp+AA20r24+lVvbHsygsXLraLnvw94TYlos1os4L3URHvkt+75nN1NxRW5MJzH6WMyuVsDWRS
fgXkPQYqIt7fGp8R/Oi6mhvLsJd9OxlQl2iDEIMeg0veM+pv8GKFjm+RkVobRGhFltFZIIdyHeiF
06M1OhqzSOwkxIYPfSaCC+r5pEldMZBzDPXRacUKl6f+lU1P8LvbHCQ+W+S1MIc8LBqGU/4Gc13D
fnrahKWYSIhJChqJrX0Xz2Y2TTBxDUsGmx0/n5jYT0YzlwpqFznXnTJEwlul4fRbi+1RjaoGNb6x
sMlQj/3KnFh86J1GcZkvHEA/pYoIKK3yIYiyN1wVxod19uQZ50wBoZ/oX/HgITi1RxewCLi7wkra
dE7pUWxoktK8WTRhZyNF30xR1sZEn6915UQNmgJdI/SG+O/8Yax+VjuT0Nv2xN3dy8YH4Q59Dunf
l4Gs+JDHVwV5snPURCwSGhJb2J1Xiode6z170AX3IwDFBl9Hr3FCn3FxKjEqekOA+bLXfDKXvcs+
Mden3cwwUKFCj4HWaeCvPxnvRAo+sCpmCU8i/z4rSOxQUkTGoZcLkXebWuhB136esI1e98hRmn8r
fkz88gleQddH4QATgOZi4yCfipQR0OQ6Y4orQYQbL4L1Um+TaZ0K/qiJSglt7vA3MMWwx492rdSJ
uH1029KSg4bjMPNfhq5XZTJSe+JqFRvs2os1aOLHxDm10fAJotHmfQ7pxF72kjHiTWLpBIkU1Ia5
eydsLg8UJdvFjIsCIsa660rNwQq5+49eE0SVCwmeQkdGzilw+ucAIJRO1ri7lBGua1bbb8qvUDL1
uhBnrHM7feDkUfK54XmB3Y+Yee5nGH/gvs5YJwxfF6Sa3Fj8Y35q65YdiMM2WNLlypNfmPU41MQn
fy5Mh1Klb2+lKRT+Cwbk+ruwNTYc+99qnh0IkjbNM94FM4ToxkqUZ7mPHqnUnH6skx3ipmHkLje+
hdNyHycVRIQIjC5GUdOhqduKSS/p2ipe+nH6ibbxt/EjOsAo8dY556Ce4AMHHzIAVeEhhLM0oBQ4
YDUoQ7WsKWE+jxx9lKiW9FnLRMugRwgXHyGjOGzSloqxPXOFh1yByWaK4078a5STJ+m5m7dObPqR
6grZ+/pcHkiuHe0Eu4LdTwmMJKJsjKWbr+Lp+dcEae8tTyO3V0b0MLxBe8o86vqQhpB+XE7O/NFZ
xPVF3xQBqB7FkpgoakEERB4d1HEfsjNQordCWVPn8DZ2sm5Vd6MflT6GgOwLIbyqC08QW9AfkjM9
BZOYZqPeZQfSRXFpfwSoh76r5lNYhTVsA8WggLpVwllwsvH3nEgRJEDSv8zyZFXos8yQvsha3nLi
0TsuVRd6946XN2WjyuO/Cv1RDVRbeN4aCXrWuTPJOZ3fQqW4Wvky+dTBmFrF4ppqwsLJzq7oQVUz
dHTKNBdtkar1pR91uBn0ffy1hfFCgj13oFNy2EH8S3IVUHrK1QtAgdSGcV3IsDdlk6DO3wteq0g+
uCy7jDSxkvGd+XPRFIMoPZApPAQnk6v7w5G5Excot6bDSGewfqqD1gDPXMlgcTChEw4U1HFutNXe
/DY37E9lC9O78gBpSATuN5SQGqf5FPjc2m+5+u9sLzsYewOQ6TTgcvj9eVM3589Ucz6Ks9L9hqO4
ZPApRmgSZLBUv/p1YIG8+6HqvkC86f2ICRT3KfgEui5k39K02pznyLDeZYi/TF1cwYXpozV7robs
CKc77P7moS7LRwxZqP4ov0Ddkf33SsWYB4tQqUnajmsRF/nkOR9HOVoIejbNnKT26Phu2m7ck41J
hSNEcMpAjIObdffezvT8OAVl7Unom3q+2eQB0H5Cd6YAPX3JIqCWP0jleQTVWoU6t/oq4jz/YaNC
SBa5rSvgloGwEX8R0rmF53jOfXFc8vD8uPq6qIsDzBYHUtUjYsb8oBKCRvMGKxGXfu5Z6dmRxN6y
9COYT9BUPYubp36amfE/s29jq5GN6Ip5yjtBdESw4zyXg6fnqUPH3iJGRvo3eTZUv61xSVqSwcaB
2TFpbyzeUATBBiMnEJckQGgH9bz7V5QHnhXRu4+VAibCHh71h8srx05VTgkrsY2DLmn0gsXGIfXt
cFwK2x8RBHaV3LvkMSMD/sEWlNBUlA8DR3elb4PQ7BemAkpKLG+EXWnUus0YvlFnz5Nezv3vTc6G
ekQwu7pAfCYXlDF0c43bmcukZbj1H4ar3hPgCmPRJYVSaA06L5tRfcG1FPhL8M2PykUA3jA4ED6p
QUXAwjbDUCbiF+kDnaRMGGG2UpOWx5zcvjcWkmkq4w8QWy0v5VJpw6TxKF7EMzgtRH+GLTeoOP7d
iOiBkCy4qpTol1GOTONPaAeie37dLWXcjojlWJE+1QdByemFlVsflm7Wrh5WEtbIIS89U7XwyDPS
KdJGhdACS60+HkjCy8uW8PV+ixAT89yeDYNvhBV3hmUU/3jNWMyf0dkfkMLjMrEoTvZOQjs9WGkw
+TJGC6BGQcZhsR9FHN4BDWPmsI02GCvAp/DlFMEI68nZJFfdiuDwTSunEw5tVSgzSsyVFtJ2Kdw0
RkH1XeBEqALHJ6JiH3/51k+5JJuxgnjtyN8PWXnLlIsSmfSnt1wZ8Uxo90gIiYz3FOxodqzkDLRQ
u9bytREvHmaLBZkt4lmqZcKC2YrrsqWAGZgZ9suS2xf24YqVtdgMaY49cPf6mT8AUSXcAAwnGPPo
kw9Cbd0zc4PpGMSgniSbvqKxhGIcaDK8CUXxbDjOZYqTi7HTolpwYXH1PZDgUdBDXZvZ83Rkhmwg
wbqAMtUFGqj21RJKORZBjvdmp1lIUnQa3sZ6oOYa0bgrfXMfZsvhgU9hN/4IJfXYLIOqmcPHFf5a
nMAgmlcV/W3kuepfmxuupDrcYuRhgEe/Bdo8UBBhtqK9wjLYElBnoRAsTp2zaHy7av0eM6zQfx4I
G6HqGaTNaSh/5VDN2TkxH8Jex9n2Myxq0e9uN1eMUgUowWl199jJusoH9YTwtZNe6nBg26x/7Eq6
fkDt3auukgbNXcJNiiFMAwtfMf7goyKlMIBcz+cyZctYUhTSQARDfHf5TiEg6taTmExLWc9p+Ib2
EVwPL2ZfLgwx4YcXQ+Mn9qZxN5PDG928dXuiKOFBaWE16s63Mya1cYtIjwAXy/hs0y5k5Rae2baC
igFcJrHs6+S4I2DcYLseqKXJY88XzX7OySDf++3fIozfWDRSCDQbjDB3ls93CVm6VwaKdevJDZD2
iCfVA5D6wBwcf/kWxEkgU0Zm09OCzdv9KB56756xVCdUzce294EqKWO9kcLREH5j7ilEXPg9vOzG
nPkgJBey9cmBD6dblpr5q6skc/AyRK7e6jlbugTcmQER/rlgYqRi0G9YyP/knnrbfNzy5PlmVfAr
YnrR53htoGR2WnlHezxvh9zeJOTqoXqRRjr7Df2OzFRflcSLWatxIjvH8Hn0muBCzAlg2qYeIqoY
26HVGlyQpne4iHozLrAdfiTlc2Ztew5Wwa+rfwdyA58Yy3uApmWF8I9Nn9ah7CdYCoqLgZ7BSz9/
pQPXSu12c2/W8SBh+P3T+GDdDb4+zc5lCnqsseU/rbdwnetJArVHH1jolB81cv2pSIRpPMxFQNIU
ADcZMbWhf54J9Ty1HAa3spL+98EfkFDhaRzl95iszr09TUWJjfUPgrOOVIrA6lJrJzYd+Z/fD/E+
gNXAMOAYuhIdK9zQTtJeHTqb8QaC9Qj8BouiLD95gWhaRcQYZZWcB6sRGIBjluXxqPucRU6D6M7P
n/OGAowezqKP6O2t5S/KRRJpqaDWwsXgMReO7So+9i/zseZJJ1m1ueLeulKd4XgTslC0eKv4zc8R
NRSVUTAZa1Iyw/YDpuS6RtlXHekZezNf42KEBVvsXQqUo5gRlEEGhEbBjTJRzQWXcRhP8651JjS3
4rp8HSH/xjLjVcGWxJLxwwjDT3CRxR4GeUQyJbOlxCCJSEaVyFczpAATQmAxcnpYWjpIB2ZB4rIu
QAGxpywNUUg/A2Svh/PZaCUUHXuD9Afg/NFbilu/FDT9lCpjzfryxCzN+mZcFa3QlHJaKX/sLGn5
BpYI0yDyblTE74mJWqVg6q5CTRxGJGqvm2c5VQGFGITob24YP01JIVGm3gPz0jKalhpqb+wOtbwy
itl4OboNDkMaymRGZ6Z2sDZrTenpcBUaTaxKtP/z+HLx911x6OrzA/WvoWQp5hdsp3LRizc71EIE
KcD5GcpDm7rhDfyHF1QiwNuTyDzJpzYwLgqOQmoc5pY48cryB3bm19ubmB7Iq27/3qrRvnjynaWj
APDPTza0omts2nXG+VHVNxOZDwIhR5NBQeJBOpNC6JpnZUap86C08RPovbqzdq42dCtOQfjPCwpw
PGifwK6eCDBVv3cmasr2xCi7A//NoOnEIU2wvhXzCXEgZsKw/2jvP0ZnpQx7b8iAzyocGI0R7alq
cOKDY0+0ddiN0AGTnesDMMZTgtHO77KCaB+IshnIX59/dy6Xg7F1LZshK/dvsTDjKoFazn55CrdZ
to0s7/A9NqJXr3kmpClzLx65NTAaKju4eQE3L+7TGeSndehIYMgwXmVWLa6VoP/+U0zInxHblBUU
GeWx7MAqiICAngPbrEs4JynJ/izCSOBqnK1m9PswrOgmffmmbsIfI1bfqlOiyLJwj4TcWWlIWdBL
PryS9+pkpZfYuFa3asW3KEO8Y27k5/+SITaLXpFeixxOeGhQ/+UYGJdNB77GBAF1+DXB+Z5Fzukq
3aqKzdXlETUuu4un342erMZQ4WUcdqXKE/EYmrmycIKnE1u9yX8SjBOu47+rGIKDmCa8zzvbVE+h
1yaWjEH/BdTK9j5dVERzmxIshsw4t6qOp8cq4bvuHqsHwGMlbPiTbVPd0OXHoPhRt1YugDhDg/cd
3viwgWzMz+xiRpferWUP7ZgS43+v1vdQlXbHjIGZaQG4AOsSjuemRfOHKMysmBPKJLDCwo02nEBY
PMgD3eTasp6JUw6B477r8q6slhy3wImGWkMijI68PQs6UjuIxQLnbaM7j6tAfqLjbA3jlQsMemoC
SmFSSfWqcMBAgDOxI/DyjIQ8hedHIoisnKdUoM2gGdjFhHISeF6mgYua51dPwqqfBVnph8OywVwh
zCsGjnUlkG+1Ysgdw1ZVx2pKRVLAeviwMMRzfRRNQR4Th3+9cnvkWAf6RSJdbF13OkdKYaHX/e4Q
1wdCODpMiLOGyqeR5YHv7FUPDMCoRpPK+F3M/ydEGbdzrcV+FIGEv+PNJdikcSLk+mDapmyRZ4IV
iXGPw/zu8Ef0fv9uoeZ8kMgEFT4jx+i5BWRFt3KOpb8Sq20BH62hSqj/M2OecMaDC3XzVtWo4X7J
KB9UTpppuVAtKjXFa22QoDwhJjbFJ+hJ4H5N/sNhv4G4gdauvpmErqoXj0y5Xiy/IfTQxEaKvTd+
G65kmDhU9WixhfKC8TaUUfcuMqf1uups7DVxctxFnV7Uvhe1FU+9Wu00pDRTdWqLy4ti+zuVi7y9
yIApm1UfWr8RhdpVm/AxmbPKoUgdNGeqD84JSAj40MZXMf2EBRsFssUcahZY3HMt3UEf5iAFB99Z
0G4ymgLK5EgdWfwwhL3ely8is9JVJ/BdiIxN5pI9j0NoUeJGGjEMXdrBHz9xXizoB5cpmK2wV/ke
ejgyotwVuT2Vw5DODpUsO4oX3na6eTgwINwV/F36UtI05xgHXq+bL88TNrzPTwzm27G6nZZTPDPH
9YTxPk5+WPfF/v+PWlLMb1lez1wEbKJLdxNLJjikEaANZniRMh+bGNUstRRedG7l7vBrNSE93kHy
yrR/AyJ3YvZib8qRNmLVKDhbpeQe8NyiV8JbNs9ybHjGiFirDIaWRX+vv1T4ixjaJe2JiBS6ASsM
VJSsB8aofoy4bZKzjXBNr+VzVWtIv5rq+ThoIfTBfAzXdTpZni3Sf3JjucSsefiiXR9+gkFfJYgt
xBtudKEF/8614IVRY8vTy45AvqVRT/W+qQCuA2COeW/Nyc4DPBkFdKk92A5dk7QdPxrHGgPCNG14
p5j2riTppXPpT2HDWOfZpa0XIjq3DlugmucxKex0eqI67yA85gIaCublk8rrDdIk5XjyxnqAYhJ/
MTIePfPVWWlQCG6eJT2YT+IpZGsWJ9fnR76X0k0FC/MdjmMohCzDlqNFEGLpcbK9pxmga9OAH5OV
97dY0kRRdfRqwi5cx7SBEI6Ss6IBNvHSiKn/QiPZ4l26FJEdbEHFEsLSkQmEyG4+AgMKmpx8TGdU
8F/wQDseh7/Yb958LXKGNn5D9jv+VTjaG2qOFYEQXglp+W84GupWPfRUzvT05cBm3jwm6UtfkAuO
aunClK7I0ZfHDX8awvRpUyrxk7woqe1tZhuP32UvE8G5lfIYNbflDjAEqAUCuffqeWrZH4YvnuUM
ECCKPNgb2Sa9IUQ7HLjdmgUGpU79vwrj3lObpj8dS6c7O6H4wM+80VcwYI4vEhMY4TlUJGJygcUn
ALB3NLPW6MOCE5wzhnTggqpVAJtLiR1tU3/WvmfnPL9XmEvlU1IGC8g901pKisEVjKESF7HRGFbe
zTw8I/isBP1P8D/8KWiBkQRUULOVCSWkZxDws/Uaf1Uo+qg4Y/+RCGyiDaOfSwXF6VCUzhuzsazB
g+vMFkBazh8ntBq4n45uh76YoXRGvBYRXRADWYCMyLtD32DQOEqGCiGUseyIIVzWtd3GvVMLvM2x
KWNlK7WoTw99+BaCBaM0tK1QdLjQJtchQ+oWs37QJVsvCSXkxIIwl2zdmxXXjh5IVvprkiNW2D7F
jePh7kAThsZb7C8swrNH/sqbSPyhPv85lFs2P2eKh1sTDW3KXpjUyE+3rwJgp9hTizDI+zGEjKF8
sSplf+69JKod4v2NZGOAooLfoGbUbjbrbB+0XFmaa/B895SomwP9dv6BVIZG7vT1xPfKG43NQqBB
1/UPBSGf0MO1ndg0g3PuCWyE1NeQqDB1Fv03rfBtoeG5gRAPYWv4xqX1bZnfdBL60DZ/ev5qmu1J
ctZp2WpqOUY9Yf2vWnqhL4b4DuChttkcqzPyqat/5QcwDYp6zLu5hVqcpp7gp00V9qNwQPXinV1P
YQZCFGl4s/Q2lkUSOvClizof8VcZKZN0KXxHIN6xLuqSpuN1VAsAlG2B0k2besA3tTIluq00iidX
6rARBAfc66iIV+B2eDguIxoL9ztE9yaPClzvWlPhYZKzjt2sMrZOQ3iSOVJjZ7Ha9HNfZL3pyor5
EMc58sw0ZfQ940bbE9GhcrTJSsSgDXC1l9GET3gQlu978PBGWa8U6F+i6J0JvOC4Vm4ykNGNT1S9
NPDWDeAZxcmEMwe3g50UdNUvlSaa8aS8Bql/CdRBqVnJslHhcY5xvyJNSCszig+Ji+Yi4sMu76Gt
zzxi9h+vO5mjWQbEFY4q1dR67KmkqrefDpvz2+1EWOZufofrr3QxFouhBNM1WCnDb3geS389ka+s
fW9IRNndJDJEbvqAvgvzrWRvjaIPDC1juJ3rh3pOPWAbY+ROq3OxoKa98TphM/RG7jKsWFMdRGT0
viP8oTxkwyH4qS3dKpb6Nc7C9FVTk2jY+Tekvx6TLB0EWXG2u/xlmNdQ0izD1VxqYR44uDqb4z9F
qsiElGvUpo1UssvPWE95/snga0q5XUUZCM4jN8vhAJyZw4Lv8CmhxyPtNSnqLK7p5ZBi8n152ZoL
HxzbJVGRLObx+l6Dfk41ibmOGc11mOSOkbSBR9jwf3PfNMF4CHDE6xBknRlcMpLkVuFjmGUd0VNY
fmVG3CiNjWNiBrn28wVKV9DPnPrxiy3N7bH9eWpApD0At+9PVCmKacpH0g+r8BUGR3/oM+IdpMIj
Bda1YbjohcoD4SuRjU0Q2M2l/4E4FmsMMNzjKxOp31hk9NYg1STOSvRvI0fKNXjW9aERRz1KZeKD
kyd3lDTzFsRICQaOqo4o/bnYdflOKcA5HsQx9JPlQXhUpCIfkICkLNZYBlTMu9+1ocHNpEd4B1Zy
vnn9xPIpX4XOO6uIJKZUHy6hDRlatPA/hQS5JJ6jKsw2eLjWeBi7ww0G1MYuojMsPDd9R34zJXTg
oTvCVUe8C0psrQidNItdwk7GQakW5dGZiE+3nuLR9Lb7sN5qCUEPeBdYW36asr9hzMy/XWHZdgMW
6r5Q1wpw1kLAHjFBpNGM04vs3tHL7p84Ji9Bm5eb85/QqGZw16PPv1kqeL5PZOJNM68IPETM/+OF
b5icpD2mHPFpL3/XYlkLiP5z93SiWn+UTJgocCeGfKpIOgLFPU0Ws862zuHx3ON3eGgMFyozOXNs
6yLkS1rn/bDuxcyTeY+p00n2a4QSXdXkF3604IsEkcqbur9GLF365WIXTZvEYhFQxxhM5j8BEKbs
g9kW+oNZywZXZbVX2lIgympEQW1Haui8vEc/DlrA7WMbgR/hWiUt1itKqjjsMzx9RRPolb88pdhj
HF8zGRYWbulchc4PkVBXDQcBXzIU3MUZQ2HHB6e4fXxWrzwFrJoPdtVk6/Z71a9Vw9T7zPWiWePE
mCDhZB411DlnRoxfOPM7884E1D30EtBgF0f9RBI2XG77d+FDusI4D92GGIV4DhICBhXdXpIKQfie
b1EKOG9VPtXSsoipM8P6xo8eCAuXzSJ9CRMRlBx3ibUVQOblDVXJGzrIJFPnhkZ2d3dLE4qE27yA
s9ChnCy0b4z6cfXZzD/9ru3qqUd7GWa8OTfGBXogLoeRAgwnFfDSg40opV1lGfLWQ6tYCXTAD85a
vS9FrKZVm8FYeNl4Tz9QovwiRs7RESM8hAVE0akf3vYaND/h26O10p48nLE8gKTJxg9cCy7HTlnA
E0a4UoaFO2+5PmDp93Mm4AhqY8RMNmRwFg8LpySoWSFhIJcVPXp9rHreZYlLaYwhO6jyrdwYJcsC
iQQSM55a+BZw4WUZcj25bk3DPOyEZwVFLSpiUZkMzlArg7/6x8P3VXW2MMMv4aqyCRtq5Z7avLFp
4Wwe7Dnw81vKMwOdmMgyXlV7l348g1f9p8cKExEQAkgzn2aIarPHgHIU7I3sQY/VSE2BhAZar1TU
zNkQfG1GYioSgAj6Ha0EFv6oRmR3i9ccyGUrAQ504WymE9IHkad+CWeXN40mgPDIz7mg5ks/feTQ
Iu21t+/q/qPubygvi0pZivQ19PkzE9p6IcN9c4Vuqwf2EXqq207RhrsK2sYlezLBi2upVQA92yGh
Dtue4I3TWE+m0diZXC5ws+eWsl57aZtnRCaAtC1oLBugVTTwW3L1VX6/HHDl1H8gS5z8MCY32ADV
MBAJbNJF/9VkHlZ2bBrqRW8LZ16X8zXhZSDeq0QzXkH1fjg+KzYSpjHl1H/UMIq5hWsCvgp7m1cQ
J0b3x6GFMmiOneTHTbPIOLqIYpzPglB0Ikq+HiiZAHy42Gh897k387r4r2YgF37E4FmfBKkeBUcd
CdiYN1YPG0x4pf/a077A70gXC3AS/nmX4WgJe05nV9idkY3AHS9ke7UlfEbep2L9GZiJqhVuiis/
a9356GMmmtFeAWzjIMjLP0zXRi99ddlhLcU2Jmoj828MkSj1H2MRyl7Nz1V5QFPljBgCK79YOVrI
zwnAZFpW8duqAgh2YaadcyI2t/kemjBD4o5kdkVCFqraPOKLYTXRlZ/zuiL/P742AxRJtlteftM8
9CIK20BtH3DhEKt4q5BqtstzPvc25KKam3hnJXruvqHVCztJQ3zDnY3FZRvKNkNQ3Qhk2OwSzToy
WivSrdrhCb0+mC/voW8Q7+2+w/l3ITRYdyScq0xbajmrv6mq2ZfIHR3AUVfs8TjrYBOoc6UhbSK2
/uudlkvyHey5y6gRJ8UNPc/CyZKRlb+vA4P0TeNC3asx324bd0BxCcNBsgGLqc/x8TtCT+ZwZ8kQ
fqImTPz/zhL41SnzHzgFczTGQA2fufjlPM5lbbt7SFGhJ7W8ImGq1m2yywMzUKWF8TOHIIA42fIx
BtLw7Lts+Zvy0ONue4UYZsNZMKlWbHMrsBPPXezqUgf6RZel9FG9hzlv19vTnoIwoJME/GcTiEqt
u40FKeYQ1Gzg1A0zGL18fwrVy8RkRPxpocuMehyeJ62DqQaxlm+SW8BkvF/umxT9VVVr2l8x58f7
Rcp/OMnJ3jQPEdnSDWctBxi6jQSFSpBNFd6GlxzrBZ7ZoDpjkrV9V77B+VW45CFpUjIHqV5h8iAa
KvFbR3VNoHaR2XNGwhOINzKduork/MZtEioX6cBSbuL9awzTnSe8iYMjnBNNNnvIkEHnv4zV60+X
0BZqdP2bE/L6384IMIuo8dDoiupG6Ld0kyMfGClP27lzm3B5h4EtZ5+agtHVhDc+69nwyNL1g/qy
fWELyziXUo+i/TenazoM4jf1aBO7qA6Nl2vmquCGqfodR63/rohTp8OG45F8UGT1dO+O5r4up0o5
yfHNPLMmZCh0SOZw9lOuFfEA7Zc3kSfETiU4JmF6FcWeiTcXUMhCBqqD1xlTkxcyNFxjEiD5PTTQ
lUJ8HRqyGvDh1T+/zvjlSS6cEWL47QWHModpK9FOruSd7UW45A3rvKj6l1jXNBrQ6CqBj4o4hSbc
HCN5RTX7dKuitNYJIKOf0VxmyxUDJ0PG0a91Mwx2VJ2gym7KuToI0Mt1bXbpRWXk36w1CDgMYVXL
owIEdgAsjwmtMRP4W/LDuEMBv1PP9EIp13S6bubzatwRnlZ9xO9xU9sAMN7pcL0SCtiUG/KJBHLM
ycDdxvFy96ALLH5w43H4vcfsmrEoqAZXegdHVT7MQiuFXlOPHK+PTCHYaKSryRDYoHE36FO3ciDB
CMVG/GMKxVtuYdyVeWP6UiJIlTfVtFGBxmgXTQeKHYzkLh66LqcMDG2vMsG/xRFjQHQvGGKhB7bx
K5RGIuasvdislcr7UIr0Otv7aUsfrIiU9x6tdFKJujzGXjQUpBEZFciJEIBICKlw9B2Cx5wmuk83
9/TDQNLkVtpvMNznJzAnpVK5XnV27JfpWZhFOYsuXqXCJGVdGHClEGU8dk+A+r31kWuwim7mXBOX
vHq/h3Kans2CMZQhSydUKaIcJTeJTGfO2oDnkYsLmOlyNVe2j4sPdWNxnGHYGRSS/aIe5pW6mLad
RFORuk8sD22PFYPPALaax0rnx+fj5gYjowCMbs+w21gG2e/padLNGlAikRYaigPOvyMpUy9Rwfzs
1vBhB3W4U4CjJX0iJhoYY6JfGmOMuekoGpLMoPw9JdeL2Gnb/U+stmruTGc1fGJI/n5eHtjupnkr
WWS+FRWTD3EilWcoYGa7xjzAaBXNxjaof+F3YzF3pjPegegDijKb+LVwMXEeyMYHht3YJSiN5fvI
1FNBLxgGzvQtOwBDM/pOjLBWryZv0DYxt2cxwVeSfa4dyrd2FYM67wmLVJCjdblmztw77tq6BCTn
gRZJS5ePl4hgKPjNyYrg877pkr+fS+jlDBUBvO+WoTGZMPrkSsPNybM2AcTt9h3jel3qm5WHP9NN
+Zupym7A0bPoCiq6tYL4GKk8pSw0buKi3z1rPp+Egc5z1AV0Mp9TKIcjrXKLeB8fnA1N9WbDf4TH
7Ut4joEcHtQPMqvQe4Idb2KEP3+ICq4asVtm+GL1+vGYdHDOUOyUFNFwGlTg3uXs+6VcGMW4Fz6r
uI0dE1W8DvZlditfBvLgixzjvwVTU9bspyjt2GULW015ugO3YbEnM1tTT4lQ5LRqxDNFSxCyjIJB
bJp0ZBJ4+ZaDBe5Bwhi1qcUpEUB2Ggzp2O3ExjhpkmZj/bikQHJ8thRT9cyEazsYqkIzLWarxRVA
DbXdHeu9NcegcT/V8xlSa3qRz7bxYvWwWuEA62/VmHEqJZYMa9OgKsplLApLqjfWjRBEmN+tl0cw
8TRTzYzSZ9w9A6/zxCPLvOJH3TZEhb01tC0s4gjb4tRKWw9fPX3Rch6HEXFM7KzR76PHAsGjX0sG
3wMGiF1uCvYWxBJYSY5PJURQqwfgc17XPByNfkUI+Ip7N8w2JAH4SHIEfHwXEm1eOP+iZqk7JqlP
D3S6u5LU1UtgLOG+h4S8lbRl4seWWwworvCi0lg+bXykZRzg+pYsJAHpYMXN+NvhU7Muk7QFJ7U2
K7vY8rcmDhKEWiRKMF8vIezYeGl0Tx25X9DZxA+wOuf0cRZ+r2FvQ60d32VdN4NAB1nOQLPxsJ8b
LuTCHV5iYsvAJsuGaUpyw+BvgugXbrDfgQSYiESpGTogv8oF+2x5dO48HE3VmSmimh7AeBksY3aw
LfUCdRS6KNj34XWt1eLxEV1dsEY7kowJCgsyAboX4h5La1Ue9ZaHgyUZGlPZwTTk9HDa8x45SuQq
P2eo6Rnz48CHBVAMx4gd1wIOO55PC/n9BH4pVnmPSUkz2Wsai2dBaDG7SHdjQE8bncvaNB8ft4Ca
yHOuWRei8JKEwRyT76917bxC3+wgpvHAbiO5h24nMPu5A3TtZdVWj1C6bJZtsVk42IqfTUZz3nNu
1r1atTeOzZ8GAOUqE7KUjZXUUac8+rrJYUyIRnZTiXr32U8gZDiHelyQeydvZPEJN3vr3HsHF2vR
hx13X9PDUS9JKdffNLYwRri0YPW78fNJd63FidBUHU/UrACqOEYjyVVcX/qGlio+aW12Buzize64
OvRDQY4EsCHUYe2aeOgBEK7lO4XffRnBwLKQ9KcFtRH5bwAsC2PXykhD4K47XituhRxDj8LsWqiq
T8EAKOVQXM4Y2SzHakcLQgXgd8jdT4vu4vj9g03EKr/oz7NBX8LiQGeQpij6bls+jZz1+085HzJv
e0hk0EE7S37eaWgGUlYKwLy8IyTxhsKhNSuDuWB26s+weL3NDk+96xWUFtvKjjTUz5mjSSaJy1EY
pDa42LVItNqt/0wwqERdzU6BNTrq91Rr9DEGexcETcVmf/EIQ9HZGb1Hk8jXL/23yXOgMqXis3rS
/tqqI5XmTsfJJnfj8xkdbrW/a+PGZchBUHF5qqlAuLsf/Rjrxz3ZNOFp5lhBoDm2aqvStK0pt3Sg
OZOaPv7BrljSEZKQnpvbMev4sG/CU2swHLg7cBQF0IVwGQ7VRIiO1MwQ/JpI/+5c/ygP4QYgZhpK
/OAcR4uQdcojU/1uOk/mXGgTBM6YP+ZdjCxFmxrhRWEcSMogg1SVD5ZjO0vWbZEKr9JPRnXCAc/n
Saw9GcY0Bq6VkBGPFZoHwNpF8550RWp8kiJLfTkltTINQcjB2qagMfu/6Oj9Xq8k2Ze3lObDGHcr
FALeXWC0RYa3Sy51A/6KtZrG5WaEDk85aVCnDWtQGDwiK5dH3j2pPYr0OqaCKjjY9R7MnYk9ZueG
zLu39j5ktOvmXdNJw6WKlHE8HwdivFWNh57mkUtKUQS80Gr4dPzNE/mcT0JFIZSMwgGwFMbOGeba
V5WR9eNj9ak6MXbkEkqTh9sBmH4OIjvK6HcH8wFLSeCMKU5HJfthnQJnIkbiuvPMunhW6d9/Ts9w
RcJK0dqXnvClJPT3GU0CI+xdljQsrsZaSfvx43gJOec8kLQliWt8mshujuRn9nOPuJI3QbZjJeBp
FtrksnzDCn/vetZYaqQKjruascVbRbWz8PtelituGiL3+ZvwAP5jNrLf+sgkgqVqLyTWN8dlzFle
vKuVO7KXPs3BQDNq9xxkjebssQ+DUehlfENT30Doo8XSKrFDPKfeNCpCoOI4eDUIGQ4Ks7u1iHEe
VJI08b1SA8A5gR1boHP5v00E5li8x7XXYNbJmDfy7Yec88yEyXvTN8WJ+x5hX6ohoasYDF7j3AE2
6iuk1ytJABEeLaSxKG4wwA9L5pvCW1AhN5tSBnZb3hecTtPCk+jHJ+xLJAqfB03hlHa7iREb10DR
caPw9niVwUzt2+A5TevwGQqHSIuiMITc8UFKJDRfjdSoZTY+YXNMMrLIoJ+5grraiU4ek9bx4AIs
JXZpWPkWo2EXhrSy8kCZxQ4sUBVp9AE+0fqh2BNoqMzTZvOdx9FUaT0vWdA9uwY0oH8KJ4e8JKez
AJ5H8BacfcM1mc6DiG31g8YqrIEykv4VlkiLeH5SHpFuJ8itXXjbG+37VNT779WSryUT5669RYz/
QpSTy5yX9Db0snXrFad8XgkUAFCxag32ELa408J0LyeE93yhCCfypXlfbNOP+tesKnC4bCw13ZAu
B3MuuttQCLVoGU279JUK+0NKy+hxQlrM5YL+EPz5IZwuP0ZFka0HF0T44Q7tvQ/tF/zfsxylW+9u
KOpGVTb/CRVevzEO1S91giczdvqC4M68MBRCqkRfUtRJ0x60c4Yp4eYbfSYNQYh2sRMenq2U01vf
ILk9pheebgxFoi7yr2HzX8aqmoP5coRU1suBdpAEJrB8HpCN3CdJyxJCx49T4SBadgVdXT3Zf6NJ
HcGX9E4Wwp6r0gPHMFGdkqnVGAtCWsWRWLOaea6tBGmpDRU5BKec6z2nPRhDTWo7lFr3QpqQCqN1
0gqpzhN2uNOk2cqr9vZ+k3WAI4+VuFIwhesbeKnsJORprOTjEZumEKqeqq+v3h3uY5MEicIwOLgQ
CR6jAZr1P/+LpbwI1YSX2f+yDJAvA8BxCaTFGJ776HWnGZlf/aC7e8StWaQ7MNFbMEiVIhO6a+Gb
v80rbyto+9mmjMGgiwLzgM3cIwXGp70ycy3rp5lKqD2+6pYkx9pUt8PQBJ7Vy3gPKh71naRHaxC1
UTVVIUHW8bdOu5EYmXMzf4oIQnI3+CAa9EFIMnvZ28pTphFBE9Sy5sS5cul8BeUJenmpcDflVnWp
S79GXEx3eqrdGz3L2Xb4SGkV2kAv7qaC4St0inGq2b24lRaNx70fC7od0iwc7j1okILWxyZyet2e
/yZbdkLmjtkn0eula8Jqrf0V1wJ81WWC2TbvmZEg/+a+VhdfIzbVJZ+LRqUcEtwiw3GTmR+l/Ml6
d2YSGESAZPuRpf9YobHVjVLnslHiXhj4k9nun0Lkq9AAY27b0lQBVN618XQYj9prEZ54hsQ2zBzO
huY/fBh4Td3Rj4wyRjxLESdwHpJb/c1yKgd63zXjEeYqsRx4wFijqfOImB6fSqy61JH5E4RWUsYM
1qHbTALAOHyUVdVbwoL5eG6buaZFD+3YteDd51cNlrWtm58M12vFTxy0mdMi89zfZDYKKA7b8bRV
El1uumQLi7GedYbaKTdu77Ki3mCncACyLSULi4vCrVzyLiRLxMblJS1nFZIIcFUzCwlqv8ExnHWo
5X5RN5Mo0UKft/BxMAUbmaBS4paTj1KgHJ5QUMAF4OdXdMtlGHvyPGfB12SzxnfMk6Gtf9BdeyRO
PZgt67ROZ+XqxtwQE3AKSmaoVCUj6RNLraf4Hoh3wif5fcI4RLw756olVRWKuaHaN1uOJeO+smh5
m2pPr6nT5pQXPyj45dwlXXPb7C03IkHhsez89SNWb7xnrnYxUXgV7Sdqd1cbkPA+IT7BKlgSQywS
pFDLt7SQpZd245LKxcco5BvY8yqb/5WX3OgvcGPr79Qr4r2Nbf0zEIA59Xqk/TfOay36XhVKZCOk
nH2pweNg4TRuXeYyO8Qff6hMhuVZuAHEpYdWBB6WrrxhLHX6zGjIwyjeUNjVXqjomi+zt5bDd7iq
NCKTFm8gsu5ujXncCxGqAOFuKgIIwkQ5uThOYZR0lI1gfqSANJbsAFGB1cgEioid+Kb2rRhtyL92
8T6CdgxJVzab1iPFY5psuAsjRA4Iv8JJvjxIv3d0rnjmPMU5lkF6nm7Dls/QZRBXnQqZsZvIWq2p
YtDofIt+gjP0et5/o41AstE1X+103k4GF/arwpie5aaX8q4rGjH0Qi9vGzP0EAVahFAH2W3KbslA
k4JK/NKvBJ++OiJEYIPx/6RESV8SaZHMroMBaLy/iJFgWeltID8Nm1WLN9ucMblt3Xv48+iCoAXl
hopV6YkA6DJ+yCqTOFzxK8i10B/5ILv3FRDdWU4fpz4wz2AX2StgJfIo8Qs5mNaKzCTWF8kM04k1
fR80jd6CeFdjKTZGhwZ9NwSlMXSAH4c8vKOj7IPlMvccmcZZ2t7nHHM/mpYdyklipU0QJqQCBjEY
vncSVI+P3nfu1mHzfOtqOEJsd3zs9Ql3o7TL57gaQUfWTTbQ5RI+h5tCYK9v4k8DFzaEzDjrcjfA
etz93+1KkKZoyYo9tf72pD46NSJSiBwTOU0dNv6cKWbzGm494fWg23duLclCKCmMmAZmiIlffVTO
dQAYKhwFk1eTU3UPU5NWKfv86kqZlOLDd7l4m2xx7GhoVA4QbQQwxJgiymaOOphCXBhcXwRs1aVg
a5UK5xb2/7v0BzdAKVDX71Av75X6/r9cEsJ2iYslfWy8l8r7nBw1DaywuP9AR6FkvyWW4U9fKJCJ
6Jmfl8W+wGqI2Bg5PaxbJM8GBTiIsIJwlJ1B/0SwmzSQqID2ssbCdQ4L8opG7Fselzc6cOT4dIih
uJ+L+WBRXK2i/LF1rTNk6Pd8x1URCZYxqK2sv6J7GXjBh05ebnypWBHuA/FB97cinEXPXeHabYAl
cqqe9SI28ZuSmMQyWEVwsPLOiz90SOlxLF2KsP/3IHRdIczAkS52li7xqvDxOVYqU+itef+oCOKu
Rmff+HMhDyGdheghohs+F9oYp0WQMmzwlyxNfmV9Kr7zXnDIlqHDi2W93vOjRZrYLyfo1prJeY7g
PSxN85CaAbhjZFwHoKO7I2LxMJSywvsIeVa8Icv3VKqDGVhe2WKI0zbnq1JCVmnLra8zQfMIciZj
rAj+MMKupPWeHKTu6xhf9oBj2I/Riu6RAgyR90w8aSkZHDwgo5+pZTNfX/9uWR50KGGwQGY7W64s
Pdo6dnZbtxyhQUxx4ILwdZEkAmtXSq48NtTolJZWr18uzpDCzWAKNFcYhRdHHhCAnPhddmpGZQHY
GA37hq80qj8OnSuylEMLxPkXurDeQmBV4+VkLsA3bb9AJr9WSVRGcaPcKDshqzhzGsIIE5B9bjlj
0m5AWDP97vsk5z5Q5zl8MAezy1fnxDDljO7XQBbs7/0aFBce1wcbo8oiDPMX0jn0bemFw5YvDpN7
TldEwuwijl9SeYRyDRWh/sAM07KpeU6Vtj8NdhYU+7lrXa/vP2pPY5PfXVUTTBhbFE/G0vscbLVV
Q5F/YcsabZrvK7rgVuYB9diIwPN7DZrsRqDJRjNowgm6741ImDyciYooBCFcOEcgHCKZeW918qW3
bCe+VI2IV2ZsRks8fn/WTfukjb3euXNVQzWqsv4Kn7p+YlJzouKkn/uaBdRheuX2nlpqW2Wey50I
no1pDFBU1PS3p7R2VmMoe2vUk4XtJAZDZ0B5nY0Z665C4t1hhVk/HhxMzTjU9Ln0L8gBII99UOYd
jiKXb0qTNLIR7VhO6dtRpk4IeZqfRIgXqXhXQB/LJVPCi1w8qzSlnpcNbNgk86q1UlXmVFpzqjPr
/Us5kymLZvLokM+Gd5G98p2n32Y/GQkJ29im+ROZo6dofIWvv86idNmEtVNp9Bvtz/dj0SmJ8ov1
AiVUYG3Y3XzpLUPygQ9kLwzn+FxbCqdFQS+qRJnHv1PcjMXiY7Uy4U1ukPcWTbfcGfU75NmIRHzV
wkOkTgd70VY8GUkuNq1cZyPZCTTY5dSvVdeVPkWdqvR4SS3V66/qFntklSKtUqiDflfUHdg5XNAN
MvP79n/UvzM+4kq9k4zK2N7dtUnGsOyRTyDeIOFJ++xAYjB9Q1st56KxOJgb7PfKEhxdUmbGfssU
s2IEe3d6VAZRsVTqO1LbP1gpJ+jJyOJTLzhln7zY3Slhdl/v+rJs/WtgeIq15qceFFr9guXBahRE
0Z4EFx5ie+YdRIswpRqeqXgrf49kfRC3Uj77vHnrnSpNf7QPOa6M23rd94xQDhlSROYYsIU/878D
3TI8X5DFmrvSFEoNCpe8OwLQ2nRyLZDV5R2XiRyT210TvJjHjojlt6mv/Zr+OjjTUOXTf+ta/Nnb
Am2/Lrub33IC8Cga+PakcShLNRkzwaFu2a/1UOvH3SBNj0mSY3SIagNUbootwkUseCHY+bDNC6Lo
O7I7Tccl576hck45FMYvkeJcD9V8nK4lL0aJ3dX67XBbFP/jEXLf2iQVykihhnFHrYDQCX0ypvhO
UmpZ78Oo7a4Fr4MwmChyUtGKRx8BEcZRWO2Q9x+vciF0RM7ACoCuRelCIM2y5D3qR4ABf0S2D4oc
vAoetNVVYpVuh+NjkSB5603/7HnxoYRd3kc0QlKuSgLh+A1qmTdovRW3hbDIaiXDCSjjLy4pdx5b
pfMrUVC3mPYLhjKLJhwr/Ucg0nx2hLbN+v8Nx2cCxc2/tpfcks8ynChImQiGnRVIekn7v8G9Czsr
b5w6jGALiewXnWrRyAH66jiSWLgpVxL74lapfQWdRxvYj7lTnIpCT5WjtoIirmELkQ6T6S3TbquL
zr0+i1HVDhjAHouWlN1oeswl/oPIMTp7bIW6qR1fJiaXYHP3SVGWidRgZ/N2uyG/cI+Tk3TEbdSG
YbIfvjxpYjaaDyc5i6QC07EilrjGYr3SQOb8G87/h6LUTQGvUbG6G0Br72Add8X7v2uh5kY5d5zZ
h4QDz1UrED0oAWYeUQOgkUorD9v7BhSiyatYM78eixqvs1P5UBfCVklAYGJnGwZkKYvnDhpLadTq
pirzsvxLUm+wEzqushGLa9lvoXYMkZCQN7pVaY8wyu0Vq4rD+mA7T9MDid2E+qL6wWczbHuJ07Pg
ZxsHXytNXouWzFxHOJCax7/wvAYmmbs8kL3eRuWFwKYeDG/0D5ZYrI5Z8mX6/iu2258+ZRf7EORP
CIqQEpX6JIlkiyol8kjc+XUvOeTHMDRTPALLXyzdOqIGrHaI2N6pPExAJI96W0Qx9b0HLVkfdVsl
M9Nvyi1CBpTvyLkWqcBRmdAl9GcZwvaJ8oB2q3kV38yhdWU+0AapX4uXpJUJ2JE24UTMc5kqM/F/
FmsRJE03GB9N028jIWdSL0HmGXqlpGfCJCVMXGxLDC1c6GfJQR0P/y+hNye+ogyxTuy3tJnZafmD
XnsVjO93qGmgoFqD1doPMUWX15FF+SiPEAvqA7LlI5pY80iSIMndHlVf725I3R75ukWxYEOHWj4J
Fk65QY9j9yc8Xeo9Dk1A6UnHspkXnjuZTI2rnz2h7xr2/28GtGq8xaSmA0cB1fpg9k3YGvaGnw69
oMETldrXLrY7h+O5EctHVr1vlAq3MYxMs63zqdl+8gzDK42E0Z4i6VG+Nu17KOfkJjSt2e+1s5FA
tQGoPKBDHWTTL/SqdeWdyebUMq87CgnT4Bj1U+rI5RMhEK/XQl6osxA/RM2PqwhFRENnofI4zoMH
5s7dNMAjvJyJF1TkOcMqwsoaIWa0Y3I4lAOoG6yuoI32/qKS6Zw7j7juK+b54QRr2C9UNFegiOsD
eXwTGJzPzk6DrXCnjeSbhwBfoRlXCpECZzDneHARbP3CaycCGvyBuV1+KQJfg5lHtgeOxutveh0u
iQyvrhi/NmJd3Xgiqn1zV3IcxitRk0lvl9hj/MMt6bucH2oYottwBsG+4F1DdUVZIfD3aQMADnpn
4r72TAAGXGZde5eL/yXEB9zz7TkkMjnbBvPwN45n+b1sJh6Aw0xDZ9oniC1bYdpRigTOPMtp8WtQ
g4gpuqV01vLiuIXVbfCFCQ5Y0S5iZB6Y1DEJ4cDGlBTd0xmvvQUSpuWPTii91fAuZuGloOBNWmzJ
NjQMBkFfn6Dn6yvt5tDbYwpdZo1xVA5CnYJVr2lwC3qqHDMQyoicLG2nyVZjtHN/ZAF4L5sR48CJ
70xJ2hX1e/3hrvgvOFIILI3q9tXkO1Tt1iG7oICdXEeZNCjgDW8GXFCAaguJKdC2nkhrYqWwCosW
5nxoVOkq5FA0XdU88qMDcYbJIM0uf1aBLtVhDS72kfCIg/O06ZGHah1NQtDrC0QghpT1Yg5hyVQv
VwZbjhuX6jJdC2Gkt0GOoWCTEINrdF/JTpvn7+m3r/AruXrRlentbB/fg76/JCr2sQ1qxbVWHcuI
vAGHiE6Pak9eESpogv2blDjGbzeI3W+emlcA6lvwhZbsGvo/UwXZIL2cO+3tDfm82ar2o7jUUluP
KOTrGXZnBj/ZZ0ab6VS2XO2jDOILZsp33CoJ3lObZbKMHSgo0UWNOA3J0EVrPbShooU2RN9wNng4
6J3G0Mg5Bc0iQN4kF3iXHI6o7C6Fbfzwpu9/NJYiolaWbVlLVVmuFvhZw6b1cD2vMQvc+mArMprG
bwPgB6Fm+vlTH01TlcyiqE/Uq2UgIBUuB7ESHNSqSS0OmSpzl9mfVnMadYBNz+xo+7to73EFQulU
7PysVJcFU7FUq8ocLaSh+HNwC4aYPpfh4SHqPUtBtw25I/ioLKqbCGPnOeJifYMY7oLXEJWAqpKb
AE4CzslDiL35TI9kNEDvnrRk7ELDbCpgjDMuPbylAkRbfXNX7UMD+RtkSVwlvEBahs1ymkvaduAJ
4SeLZngeng+j0aLCDlGbFVDADivImYwBzRmjNn7hG1GFgTb8ona6Ls+EApC66AaK/wtvzwKASGGi
zV1W3QVCLZsodZ4dyfu4cq+3sWggPOMBwhdXTRHpAAcnWoDZnY25hqm2YljMNpFDeGgjZj376Wbp
MTDjhF6UQqLztrlY82Altnsbfho91hskyH0Gk3gDYbGrMiXWt22anLMc5Zp2/kthQVsXhtVmRIET
qUiKM/3RNGDGJ9jcXZnIwdh6gNb5Xf8+9kKieoKcAhcsl46cojuXl6cs60nRvqkKgLdJ/wp8nnfH
EFy9cad3azL1pzndjeCzYOCrwMDm51VBr878X5X/1eFX63Kc1WXm3doDR/ktUAUC48A9dPuyX3yq
ueVt57yXOFPAqZfuhgEb6uVoaT/in8QLOkkJxSu5hvs/IEytd5nPK7bpT/MiiEgAh8Jg8PDlHOcc
i6A9DZlmOI55K+u4Lf99jC+8lPvOIMqsi8mBsnhEy+jvv3z5Z41PvxK//xJLQXmSlGA8VtgDO/tU
g3CSFwZGxWq9zZvc+spRY7ot7hr8XLmhR91gdJFLaEeWGngcRHCauc1xR5ITwnBTwf0klsUTwKYf
3gih8faTF2LFHCMdXiLGLFJ6UxSNzKsHHH79Guj3SoW+DpSaCshAnuHl7ZKLUfePk0JKHu4fN9u6
uFp7MmRGnYVTRv/0xoFYfbWKrqfWWqsvj/o8MvQ8b078DOLcwxy8DWssQ/4YrtAmL+fH5wFk7R1m
1yza0UGXKRCZFdoY+1Qc8aSLNILJnoix6JGQwcyHhoRJd7APhc9xrJxeGNI/PHeyTEjRMz94r6TY
2O2htQ7tWmU6vahK6hHDhed8PxkzeB7oGpK5W03gHrvzo+wJFMLycXm/qkE/4zCSalVYoQ4XKtuG
M6vpmKNAPhW1OaHgmD/j361FusN3qbzTPlBoNQKo0FfTeNT3/GFPXjuziXggganZpOfZAa0U6QjD
bOEFfHNHvZ+gYAp4001svt/CJNpT7XZwld2O4X2648wfpCgs89JDvMuUDZU47I728nOG769yOV5z
Th+OtxMt2PgPSvovwKHXglHvXsMvx0nF1yuSq0yD6fVh5G3Rlhral6g82DXLczY5G8xOl0WAowWL
mrA+jBdTNpjzqV1jJcvQgHFH4/qCX7hTOqW7W4xjwf0mPDQ42mSw1DLj7TT8IuO5IRJ29j/ezAuJ
7l5dGUol6OvjkElXQ0unGR03oVA1HdHnF0ztvqGZjg0DeeYhnOE5sdRy0lJs2CUOGPrkIjKhnj60
zgeGN/IiVAR84vslF4/u2q7CPMRGHKLyirBNRy6ZWpcMGijHjpPoPSpEjMzgxThSCU3g0QYCFvf+
8Ml23oSGfm9kbFO5adk10VzJri9yNc/E85mMeEykl8aOwG9p7tS3nnwws0Rlpr2LHQzGIlpDLcJX
9rdMuRlEEnp+ftncsKjknEFo3P4SPdHmih9p/uNHHkU3ytsRAzNftq3xMAHWJ093IXDL4Wdj+cyj
NoBCIxsVlSh9CDYX81nCOH+xgMH2GFO56mo6BcDNILRMjXlcnVX272rtrha2ZiVGmQSlv/X3hTPT
zHyUudUeAierBtq4cmn+EAHp0DBEzZwG9HxBxwzKEMI3ECtJywLcwZHd6JZhNiebYAyZQ65sngwC
d4dzW2rAr+IRyUPIacmsbKhySLrvV3B4J4k7Q6W6NCpIq9fghtWebzCZ+v+lwQQkU4WxZyz5ubZz
boCsbjmRt3mG0aomcuiQU09X3GczgzmGM0wJ3ljscCJNK2Ddfi9jaNz2UmEDHk6xOjklfKXg8Ayu
PSw73/j/7Y8Bk9Ej1CGJnbliKgQ0D3Mi2qtSdYxqzAUwdT8sVBpyIZK3knPEh2qYBX+D4+vsEooY
l6g7n0jA7q0lwq5i22ymPS/JDZIcw27Zc1+rvcB6Uwspuvhka9Nw+nXZC5Vfe67bjj6bx5P6dO1g
NLpd4nv+GLmSp/G0OfjDBstZqYp+ujdoSpO0ZrUw3EdulF5Q5llnzv1c+mLfivn9V2oAsWerGB1G
NDw65PuE30/EKXsZjQNct/qOhaEfYz0N6yKwT1HO6s8H+ZJSxyMtfsS3+KXz8YhO6soF3YC+Cl3+
hnznCefnrW/3HClVlNxNiJvWM9NR3tU3qYcgVkrpDEfOYPdwj6o3JVLbfsqmR+EyuC15+yRs7d5u
KAIV3KSczg+ny+hjfwtKU1RIIzzvxygdQUh1h9M/E2pPh6zmijDk2O7QgbYzx95TA7ZI5K4ssceT
GOCGqY2d1XKv2eUHkFL6dmI1IjfzKtsOB0bkRLTtrzDQE9kIcDFAOGSWjUp7F2gREh4EtjIAxMei
PHRuzuM4K6AruQ2XnORBntgQdzJO/cXtRH13vXlR9qhG43hRlAIE/a2lz941ivBrXNqjREB1cNnD
n3cL0+BRcry2miALiJVtlXEsq9H29Zyfz1p+BNB23BkqP1nbV5JJOGTOwcBeRWKIw78uTGRSvgjc
UCYyNO5YMI74gOoqMqHHe++wQXykEjII75zNdydXECPxhLRLZvoi87klcBGN4Tk2j3iIXISL7VQz
0EMBJgppq9hdpH+x5vd6u+zd5zoy7w4uzO9KqPItbq6x7N5W2qWayjyBqs5ktwEEA7VifwUzE2O2
Eg5nbzirAZk3WWFDkFVrXWEe8/I/dfrabUFxxO/8mwb24ugJhB2WRnQacxA2NJFPYZLkQ4CQexFc
8NIV1t//1uCt2n9WDOihQ8DHMR4IVBJWk+QmCixSuoO0/bvyGkpd8Sy3GSwqlSMrbmPKcX2vMSlc
V9+PFUqMDsFxL1jvwfjhZ0dvRZ+M1TmEIbx2yx99LWU2dlFQwG9EPylQUjFmyGME7BcGP92XaMCW
qzlIrUs7cH4sRBRfGgQXzt/F2qUxy4SZp7+DzYa8OIVs/4SmBJdRltd4i4Yg8ElUeYxCE5h5du6l
jc2XiB6+kb/qTACvJuOhJsBuPhf+VJiOqYCFXhBJsdx7MZK/kSIFZvxFhaGHaBLUro6+k40XsD/n
sTM4bhfQyOAq8fp+3u7Wq0B5s36017fde87FvD2ylGne7uevZQJQHCeZ/2iPzcgnp+166tnLEy5h
+Ea2sO5gY1dVWL+oUGqmACLJkZNh3HVFKo5VC/dkaeFgGUzSjgTJYuo7K1MzPsqz+hRbpqy/G2qL
PjCQ9QinTZsOyizhAQU23WaVf9y+akAEbrfDdk+B8MJTE+UHh2KoMBeFCrNXmdCbC8avry5YWgr6
mGizlQdHZl57oydC46trlXdwywfhR2sy/xK1jyjFoDmUMQSLTgY5RCoNFS2FJU1vkRx+IFTNWLkr
HgJlQAMSqADq4q8J1x0CPDLwJHIm+Wf+nbCVD//msPdkE3nlRe3ZF0mOPLcRCkyBijjC4K4F4Pwn
euT6yzGFQWvqrxou/jaqZkAQnSgw9vBvQvNd2KVu6gBFrL2gy+Zf5Z9cwePdpwyC5KYqUqWb9ULk
Ew7D1fJqH1oarr768mw60jiGuSK1M8H92C22AiiNP4DYQ+GSEESNVXWvU7/QegxvEGBkLUArQkTm
XgYIr21NwDu+wXm3bfWfEAxLKvSYyJQmUFGpmDIc0tpxvjOKTpCX3bUFptZDBg4jFxPYSGSgqFWL
3YmtBEHn9Qz7v3dGKFOFv9twzYKhGLbrNLMmXEmtHjPatHLpTfDNL0WVwYpTjkb/2Y0ayALQmzVQ
ho8rfCirHeAU6LeoQwma+oEq4+fyHB0YMvjrqpyUcGvM9S8v4C8j2LEv19RHgDW5MfJNfbmhHmpc
Z0vnxrVtPe4ryyJuYq9VrPe0sFya0Ad7aj3Hc43g7iDZLU3Ueu0G4zWJQteKsy8MvTM9O1qDXBJN
+udreo7iFnnXeHZfiaLw/WKD4kmZzx46CxzgK9s1nKIoXUTGALFtVffx23+AkACZbSgAkfnvvgE2
lCwBe4WMS+p5aO53AC17DRRrjkBv0NJQVGQ4XKrta70WCNHpdx5Hrw9fDZ0xeqp5k4awWs4c10s+
ZGS2xE9e69vtG9/cBwR+HeWMGOG/mUGhlrmZKHP1GV8lYfcBavUaY8MDw1cAFlBbKE7tdehIWm4B
j/ht4qyzuDjPWW4k9ORmBa+/blc2a9k+rdgL0KbnvczP/k6XX8nH8D5q2Xk+vcPpgGeez+IC4LH3
8FL8FUxeaKw2eoeubyzjaCo4Z8/vRxsykcO5lDuAsPP8pUwZctnqhhVF3E6ymIUvHQe5LGVJUFcD
fhaduwqtkHkBOWj+1HYoxApc+tw03ZhTFP9OZwmoOQvfonqUMMu0s5fpAHaOrb6G+SeXxE8LsNKJ
bZ9hb3I/0gA7+rJ6bkSmngSAxScSMC6v9bkP4plsFeIfRlmleD/K0FuPQJJB+J3mIDscXn41BOSO
sShPMGGqjD+pg32JRoQqn0JRaYyJEtUdS/wWOFOUTBeaS0fT3qpKNZWJuhtvKoOiTtTZwGysZDLG
HXwNCqKKh/CSxL7lmoz0CHgi6x0aAejmR1MQO8m8/khsaJY/7e9o3WAG2rmUnTr0q42n3BJ4JDtH
HvXbInsDE2rGE3l0oaNG83twAcuEjo+KLWlO2YZYCv+mz84ILPadN9Bh8YCUU4suC/Q2cNgUQGop
V7/QUZlojGc3NUrEaqND6QO9+CBn/wiHfjpIJc/EjAW6IROelUQ2Kv6T7orEdjBbPswZ8B3U1rWE
v+t/1ERdvIF+IOSS/MiTGIzYTQiAsDTUi51d96r+PmvQMm3kqGBweR+lXDZsLo9vCgR+TtUVXUW0
07p3nO88zo0MwvSvmvt/h8ZZyuuLTMImUqRzT+eTM0Lyi6uOs6G+HwM8Nol/ZO2GvmhZhrWNFsYz
VZBWm+Yl3Pjieo6p0jIae1QKNHTwLivx//Ey/P+8xkMcb6tSQeH8oBmoKuZldK5m85o5GL17yW3D
m9p7ZGijGA2NGVuLa/fclJ5iFg098cdmrGMEWZGJMT/SK25C837HT1jkYY9ZnyPpwi6dRu7LFrFu
KmQ8ecZKu9NeLP4Xxs4vaQmPeTPZHWq/bDYAo6qbKbi+pRJDPPqKQHuw86lZDiiv2cw0ka0HVlKy
fwlrCw9PFvFIt1Si1N1aUV1D2xKzfUoe44MGw417RD5WEshZkIVtXkmmqY8+hB63E0X4P5H0xVei
SDgo6U9czoyWI+j0BhysNxhg3skANwnw7wu7h5LsR12QrfFV7LQxwwEWlcKKtW0G7mmv61PG87QS
1fWtxsho6xdBqWWE50oMQw8kN0FZsdoADQjwUvYr7MjP5rCTaui70j2ixFjtHk32oBFkhbO0JNsI
0zbqXrlkcuTnpZPXNJo2Qxw3ZbwJflQpINyjhhhjWSO28FXL4NUNk37kYfGKwgforgoYUUF5/5r1
0aBSPUPOODlsWU5Sj+tiLA09eelNY1o1nmGM1tDN93G050HKk9OsG81+/s8DeM+cjy+uBJjAptnH
MQr9agDzzq04MvvrwIJoWOcqmtEZXZbjwu8ij6i4ZmDezN2JWLLj0iFsPeHDqH8GhmmMDrg4t2DC
v2wJFglUBYmStS9TC8qtkQcexLUaX2kEU7ZQMnnKjP6W/AGctiTV/W9beOtvp5ZweDGL5WW7I8Ng
VgfJloiYiO6U/ytciKxivX6hMp3NtoR6G1OfA3FZiSJ6bfnvNcEn16/oCD7DHbXKiiM3WuFFfou2
U1Gf0Wv6Yspcp9CR9ejtYdJ5MmQFz2YEE8A12XZ3Mh46UiQULIGXJ27zCOFkV9fZT8RKGlrVlhsd
O70KUjCnqYJsH2GZ/5mIoka8qqWc6l7GGY5OhgFRvaI3I5OWiU7FWeU1olLeGGIPTtz7luy+sU7o
gBz5ZhVsRzOIMlGf0S1XNXB67gw/mALZKBDeausuErQKX5Vd0sxkRWkZR41n+0FI20HcjORL30Zr
rIpynbb2B2oQ1uwTsK9a3R0CUHGw42dCfkGQXj2UVNuHdizC7k45BHQwL9EIpxcEaVNtB/JgsLB0
b5xkjVVZC7zQrF7HYiH/kalyqVCN1skC27CJHl84KfXHi5w0vDwMrt+Gu/bs2e7MXsA8ElPnu7xY
xiTd4HeVJpuPMaJux4tKqnt414i7+776f6hFCFN2Q1eCap7vp6YDQbu3HGSDFlxVhuA3kYFg3G0v
OFLdaJsIsp68ltokuNbBQO9tReDLPCx0wKuX4vXdvXGWVNj5pvSpNsCr2meoILxR42gAPBwKpjYZ
xlotncgSUrj+z9LhjHS5bJcCcWHvchOltWyA3ljOFw6SKppfJiCNLo0JGRTzth2Q2yUYjq1iIxlb
F7j9GNfA5vHBPe8ydpfMJ/8kRhWB2mPasy2UdAKqkurNTuYF+WH954CdWQ3wnvI8l7VY4JEn2YY6
+G7bwdmFEyG/FSi3hZDw/yya6m+7MMGQ0Cj4j11srjV9k07NYKv+S4d4l1jI+Gb9m7b9H2+ufc+v
cq5N6+v4MVjP0wanxBgEfT8RhFqvuMaYp+xQSmcyco7MHvehYDHbqMQqQgnW4y61OWawdqfv+mKL
/Hl01ZIxnXHQIaYOl2gVW99WRlWiu/+/eQf6FCXzbQCtKqhwKyHfkGHOhLlVNjXHfv1UqsQPwYOs
HHJlRJtXiV2PiSAkfukiOeG2l1Q820y8pTxJG43kMLuz1ndNgEqwTgPmodpCHL+TGaGlMp8g4B1Y
qdGvcJF9GbX1QLkkMjjHiIdwx7aSBJQewluLiV234v1IoAsY/Y5EM4euUCjM+P7auVSKFJC6711D
uVJ5gKKj6lSGCeU6hl2A0YHC7pI994/xov5RsPNkokvyK2qdZfn9MhbibvXo8hFekiRLJOy0gki/
rSPISacKKr6iqlmuXml9o+c2KJmTnp5gRLEX3h0GDDzpFSokpHa+K5CeQ9NlxG89zICxn3sd3sXD
yB9z7Yfgc84yfiuBZqF87uv5ZVfshEpssDcs26ZX7Q5wmfBwGArUjqBTa7gWAg+Bl+TwrsDEsixN
MVBF4TNEmwUB/NKxNqmP5NFPAt06Uj/67uaup8tdqzyIK7IdX6dN6zv7vv25SITzqSAc06jZ6JH0
UbUZh/SrKhkjzj4+1HriM+o6HzXrHH26YX0n1HxiRqOvnwI2Yu/fchrcL0cWGTNEnmfDM65r2+HL
3Zhc8lek6oyQRgjXXQZ9btlKfIvaXLRbpidGKkNLban0WghAmxb/Ttwny4RFDvgnbAYGkTgKwcoA
5sGUZJj8N9DULbxPJE1DH9Tw8fVMj0NacLYLL5X2ELtlpOCZfE/pnzsQ5tDOtYDk5LlHaYQhUvQ8
3nzrnd6z9R2/ma6rd8UQk3at7mr+97vhBbhuQ3xqbUKrRnNz8pqNhmTcqmE/4Vhe6jhAEvp92l+w
aQhW14eCq5n32k2dmx9lY8UcGWuTM2HW0WqmQnWmmePT4hWNuZEnk5JdZ8uehVFkdnB19DT1D5VI
4b1fxveiENPY+AFfnTWuIk07UaLsXFecAZDeOMUh0Uk1Hfi6Vh0fzska7sqqHPgFJpRADqVBg/a5
3evOlGOtcHPI+HgagixrWcaupIX9favU1qY5laDpEmVAwPOBtlhJUnRwUrRdmRoN7WWuzaQglg4Y
I1N1CmFlnkGhwprpD6Q/RPraQpeFPFopQDGN0Q3raRE7bIQ0h9F5QCpq4Cc62T5S2Xwl9AuaoWHc
AlnLI85m6ehb/Hi1bCQp2qToNfMbC4AWcpK2RV/xo8E9w5OjkgfMw7bfY2fSB1jfBnmJqJG/QDpa
F5iiiMAkAPBevO5Wz4sF2co/HNcRt6ZdZwsehpgzAWPvu6UusjwPQHy7ewF88/g8CtqNLL6sLadE
FX4HPbqqnf6FHToEaRphEMGlKw6vviNAQBObH4rsOQEUVy1yPdO6RQvLL5xbaAY23TZOU2ahRFva
59LKGEyzSR+yz5PPq/XhhM33xPGkxpr4SUFIB1HR8AMx3dCEXvmfeUSZP/+O88ZHiR0e9i+cQo5u
4Vtnwl2unFqQZhOelfq631a2dCmuhhmfdIhnm1ryTBE+nSMbjoIPCtwXdt1q8OsqnHHLswrcKIwv
ggegqfRjn5JYz3QZPKO+48Vs6ZmczfeRRn1JTgjZPmVuX3/BUP1NFdKNXtQIwKB0BrEbC3nX1C53
Naaofljh09Wi7l204D+mLeBUyZ8A8o+jitIxOqyPEWc2oLGJvd57/hyu4PnN8QCpJ9XiAvlURgjV
XwgDEU5Hz44DXVIANjsk1p0pCPDFTHbGfmD4mvbZy+J6FlXQ84KRmIpt/h7ZFekDjGz7qabGeJ8r
HlZe6CiaGXgXHAz2OrtQk7rnLjf6X0jOxkVhoHAwDKcfwNYYX2kPXM16kaNANJNBub5vTIr5Vnmn
EBovApjjrZ5h/4Q7FpV7Zn6Br2s7azWYd/gHnWPNLzJQgv94nQd0InoXT9FrILRWOqoIgVqmysGy
jyERCYJjx50L+zMH4ivgA1Pck5aNwLofFN/wbZNuEFIj3KVZPCjoFETfFix1tYfB6H3B9KGUL0AE
VBDgdlECGKRrkfhhxo7NXLqjreD0cwp5y1oz1RmEgRtC7JaI3uD09IHH5AItapenZ8hv0Ne/cNrp
8j2G2dcVHSDeFcH6J6ypaqs5o5m0JAtqcEHsZgFRLqURbXB3O4zM5UM0vwlHPzdt9+nrmbMkcGaE
+KMW5oq02taBlRSGjmoIqIcmSTjI5c0FNPL3ApO6a0sjEUjIH7YMRj2x7ZlCwcmbX9VtxNVUPPbg
NrncaX86kijkqNduxqxNCynhWO9VLURe6Cbnry4de470Mv3Skg2RpFT8lJ9YnBVNO836Nb1Zrvsb
OPtRNedZ5TuM4pBQxwg3VZDmsI0JEHAY+ZIxii6qCfv8+4/TOodFv4dbWtfi8f/ls7XZj/xNmtB+
mn33G8SaANJrVwgGLTAtwgL85MXqFMOErZ0aXtCcrtrq9U/NaShtVIVPRSbaY36+v7RPprdHdlQQ
ZA9bQBlJXOqMHyZMqXX/oV5/1ZiLPtncmEmshnvoFTvpxuY40L7QPArqyHe6Lzy0+5U1B574VSjZ
rnaZVf6KXiYnaxYBYLCdqKV669lJ0ssqlPBEs0q515ArKR+xpDjkuGpPCt/oounwEhn9lpVm2FH3
RIjTAEK5PRsUY1/A6VfFEZCYeBRFuunkxjiMD7hCwzdzd9fdm7LXSwJYoOM40yo3O7NVlulJc67T
eXzumBKax5nFiqb53kvhq7o6ErZSI61iuuP1LTOSyrYkGL7WZMzrNQPEaSFb0VeNZna4oUoqtvc6
+5RcZLjjRTFU+MJ2oBmfTHN1PkRiJuHEhXH1d2Bjb5EAWCX3cxgeEFOqiaslnMDiurI+ct97uHTY
dSYTEq7K8TZpa2BbyCOUYj/fJriEVOpPb+V2AfJBNdR1b+GAeKUCZozfBn8u5D6SqCtgQwg3MiEz
zPGcBxs0fdEpJJx27qhSPjxuZjemPdONj0X0JuQMkWW+CNiT7JOgCJJpapOHsGS8+LkZrynWqlNV
HmzeF/JaWqWkf9eVabnqIpCjrG71lALqIKX+Uuekl70TODsUtwd9t0wZlfa93NWTZfRFXv1F5mRz
KbRe5B7Rg7OOQkxH/D+3xJgdqKEzY6OLqVatMazCofxDlZ/wL4Fg7A8zx0qCeuSmSVekOyi93OC4
sb5WzNmNgqQGE/yLrEFb5L++H0GjU7suTKl7Fp5xjre8z2nip7x3lC29y45zmzYD2dB6V/8TkRzn
piEzqs8h09YlcdMtht1tU5GcEoNwoRhDCbRH1HBz7HSRfIeW/Omxn4F/SbS3NnTikVVpkWNPvaH+
GNbdOM9ZE7GBrdKwmtRvv8y4rTLK6NjQKovmrgCD57Kl7835LGdc6a4LiFOdOO7RknHEhmaBVt3a
/Jzy41IX25orCE4Xf6xdkwswphiaSCKPL4JkDvGVebxQ8yR2EpJ8Y/NLs0nMSfbOC8Xw9nQi6EJ5
B9vRUefRiksO2WfsbL9hJgiVFpvwQBiJUkdY6qM6DwYpn7lHzfvHGlgXhmzpR8BvTCnMLUl9gti4
E6kxjhKPZnt3BcE7/l8HwDdy143uK7rgtYi83yScHVuvO0VBE62CkjOv7h1qOltc1cgIo+uRbQt0
0EAdrvgxo/+5RMqOOT0ddEFnsxGiz/epxwqTAcaNZvuyViosRl51cdIRFZSF8OEPQm9K1eGDQvQ5
VS6sfi4cFu8d4gmUgifnFkY+avbdwn2V3RtVG3yOTyMbNpcy/BmCpEabCFSo4BPffnw+BlJSPnVe
1iImNJASxOMtR6b7y3s93LFFJVXz19aVT09VxjitSh5gO2K5sJK/KN59G9SgONwu9KKu2eBGf/Er
t2g8pF0zTay0ocxMDeAL6GKUcJnqsGur0cCa/LYelZq0YXQhiWmMhqEysWNCHrpJ1cB4n10KB3qi
KP5lu+rwST94CFhn38KtILqV+EMikg7G0CvLm7wcZloGX7YOn1Mox6QyWjkTMQqfZKt8FqBctgx6
VjFlu2Yx3HUydNCh8Fa5JJpSGXpfvlyFbSzgHNJQ5X/+pBBPynbCpmq9FgTF194Ri1uJRuZ4Z1sj
fUbI2nu6JLDTLTbkhycRbdy0QeTARGeoc2UgUvnqYHQmyUMt6TuLpEtiwYhqPpul6kyHUn4Hm9HY
bbxvyd4QqjOnWBPutucsbsj0CPYxdLYhAJ2hfxdqwW16tRqfo18ubBjyOKU2gkrYyjOoxBbYlr+O
5x/wSP2MIexL0TEV7gidMIlCAjdhNwAMieC3990CO8SzISTKqTH137e5V0jBxDJCILWoZHAxRBCO
TOpWQwfmOV1dTnkVtECpSxHG+YW2MkE8P0JPXPVj1R+CAQsSHkxm4qJ7lBwbuUoSfjm3VyaQ9QWS
ZHHLee0hpcOaFgUzyAjX2U6RWMsYsdYNryhpntxMPj/WCnC6vKA3tfex7MgXH4qN6ZNXR84++cm2
9yAVu6XYBOQ7rLEaywUR6fmQkm6DRQ3FC22/Uuov1oniSME4+THIoOwz/COS3/ZKtyNHdxAZzXZ6
HLHK6COosbmM0+sVBDTBzKLHI7slhsbXK1XWaYfr7dwEx7qisq73afEN5ijFGqyVrTlvRTTo4HMA
4+5OpyqEIZwizuLnNUh4JiUqfxJXxQ87UyCGcJM6sBOudg72U+SjkiWXLpbpMN3cAdVL9q9kAGOU
oOaCq8jvmx5f6xSEjWNqwHS7f7Gb8T9H29q02uFnMWT2JOHQ3B58LWbK2QfHYKwGIVuB4cyX3JvM
r7ceHHOQ9yWyZsggBSExWgEJzkh2k7KLatK3f5h4pI5tMpBw7dZzfBTUcGEOsN4imrXDxm4rdZ4x
rh233VZEUt+9jZqfRXZZHIf1MJuIhsh3ybS54bJtfe3CbdQh7hMwTyO4AYnKZO4vDRC40WeBeO1o
gpo1V7Ery2ZiMGFh5uqcENqYGGOUI2DhMi285tF+GQ+3cw5pxulm86slUt4h58avXUjyHZL71z/Y
QE6cMFr0dhtOoIWJi5I44OT/iUWCR/avgkGGaqO8JjkoefAGZG0XfBrnV5/nrm09IzHba6TgeE/S
9dtTBInWWVYh9Z9jgl8QiirI9cVAj/v06DTxj0G66oxBaU/8dlIBsny68GjpyIV7SvFKdu/Sj/mT
gF1ztZOqpjFOu9R9+erVXzq/WTf2oiHXyM+gJffKiQS6Xx5i0SLt2Iob6dMV6TkeuuoxFhizDDKK
ZBiSl2UtsTvvJd+D5+MIuHZQ/y7mzJqlarQ4hvSUmG9kab6LqBZsHR1EU4G8JEB6LnINg08npcsN
k/aOIykzqfp2n453hoWXNDbULjkMdX0VK+E2qvsRfvs2BSHzH0tPVI0BeVKf+lClVXOi0cdEREpG
61vWiyUqFnq1NtEBDMWu8d3fskoOGgK1/mkvaT/qdtqJJsIK3gumsBLAMka85xoHJw3e+0QyYCq+
5FWZknsunTWDU7IFnF6rBw/hTFhNOZmJcpsFaK9jOyv03YxY7UdMNEVJM6BKp4NvCT9z5Uk8ACFw
2vuXWNUvxHzui3zYU3IF4b8MSUazi1HfN9/Jw38mLlJ/C/g3I0IBkBn2ATpEo+cV+8mofXF5bZ0f
CBPMyNK1D1ef3VuWN82j0et1oYaUMNsfrHdYzYyGqQfU+iGcGFEqA66u1gTmBSgCgrRbwpUtjnr0
XW1XjUUeY46qw+ND+KeFKKLusKrBTxCG30FNyso/2pc2T4oRunLFYxIfovF5avylMiTDQwgb6HIA
ZgT3Un05Ht9Lxn4bVkERYi4By7tJ7dZgFmrZ6mqgzrnQRh81EWS1j37J5vbhUPYchvYhGh+ksyY/
8qjZHZ6bLOIcuSrTR4U2zY97zepnVjXgOEmtlI7kABGLts4tHpvzIMU5ESpMUYVKW/l5GqEdiwHF
tYfR8U4YcNpEI0JkGxwN1tRLMITo3ZN95lkFyRSib3Nn3GLMOv3Qkih95in4cpbr0ErlfqBdIg4o
EFSHZYHUuJRxiI0yJ/xfOc4lXuf+xCn658WibuW5Q8t6Lv5N/M5OBNZnqTKANvTNcbEAd9u7RqIt
s5OCyYFkMk5vyQSBnPzARVA84szLi23iFQ4VuXXv3Lcz4qWqyWLqVIamKYLHHw9A5Zq0CXz3AZNx
llYj05gqmXZAclOCzDsCjlViun+WkJ0C2OE1kyoD3qMuXw8JdU1HVnZAsKBKdDb2xsNsxSLwNW61
4WpSR8tQ7W38nRjhsJtBGKzN+Z888UXnK0fC/aMyr1o8RsjGHvlN0gqQDCzuZFGDHcAhvseaCE8p
fMU6M5gg8OqtqNzFgoex1YdKQ8Q2RFtEZongoMCMOW0lz+o0f0wDeYkXW/2/3L7vwpJr8acgOaQi
+dcDmWbdk4BXjfnr/E8TIyKM6mgV2gkMaAGB0A6dLME93EqKiXWXH+gIov35AiYqG3I34waUJRkc
1VzTDbzAHaj2CE22/3uJFel5jqGnmYQrZake7igKloHQhK8PZ9geyPiD/Ot+DaJD1sFtTK6RfSRy
jRLXdV/6ALnxA6J5kuSCjZXthB8ZlwOmRdpf1CwsPEYj0RQJANxb4Hr4JvshT/i5YwGU6bxIQsYQ
BrjYPEbrsVbgpVLCJPM5luu1S3k0GHzlNaYRxDF/RsMx5AW9NC2yNHx5GRigorsutIlsZ93TdhI7
eRrwAExL/Gmqahi/YYf/Mj+ugUD8L2SW9DqVyntulyfzV22/U1eZiZCo56tdhuKsNsT+s4pdC6No
e/pEgtZDW2CPfTi82hib4otmsKDKyTgbjMHfZRV6NJLbTxyy5ySddMgb6SNrJ//vCi2E+r/qNUJ3
1VRUtUPDj4hbmo8n0OuoB4RapuTPkyR5zAF92qP7L/XDB00wdAuWdarkL+dIX2oiroHEOYF+drks
ZTq+uFVYmqdHajr5d18V2YO3X+AgMWAleoU88rb2/Va0wQ9aHn27ovM0KnZl5K8Zbk7laiWSOoL4
yI3wd6e1go+azF0iJWEfeCCT8JcqNAmG6Rc857j1R4pKxuyhNSJ7/zzuqaSckSrzDJ8AmzY2KitR
mt/ReI5Kxb2xYigtDoSm1PbE1VvG6r/BiHwi9h9Id6GkTIfbGiuahwAmRkNfWGk+G3JBh+EH9QCG
RQoN+ES+T+5Yv0/QvuoifNf8Yqzl8RRYRFONaOwVFGlxIUcx0GD1l7ZRZtSY3b7QuOPspYwagCUm
3TYcR021l/l64PTJN8iiptWaSUVKHP0eHXt+psBO0xfMV0Cgx3BDkds+yIiVwJkvDlPCvLlb5oFd
G/kgOOftvt+cyEv1x8jBlIwAULHUVRCK4djxtrAY79o6gwuZYsmsj0Rz3gbspnJUEzCEjDdO1wr2
7QmLeifEq9kMtSvUmW9rKlcdKeMmPjuaOLXQatGfXhAxqyoMzubgp5fivO+y2kp3m8PPTKDagbv7
dz5HA8zP+Ulnh4f0/dA561XrkSqiYpwz3GCeQBwmgzGJgDDypghBsH8gzvaayrpx//oPekjunaow
CMZSmg29haBDemKdF8S61o1lqC7Fy1jDOI8/HZwcy1d1r2nYrmkKeK0PgHf7U3H9YymKA/eEc+VP
tmCmtFiP3zH1wrBQS3Jh+DYimAy3oyUqc6OInQoAVA7FZBf4K3b1vKZJ++vShpwCsVMzG+oUP92K
yQ7Ibzd2WzI9uicdgul9y2F4B08lf8JaYbQK/GbGB8NE+vfVBRBGOMvRMFi3qPgqBIGn7F6xZT7h
jD/IIG7UbQjk2mLdkU1yPNhT6xMdpZ/DzF4P9pgAapXodbRQ+yReIJLmrFT3UlEjjM8kq9ZMTv09
H9lXSzgpj+S4Oozi9HOFh7GVJqDK/hhbAQ7b+gU+kbsypFgi9Jg5O6PLn4bA/iUH6E2a1iGZkxnL
hmQc7cAgSs4iAmPTgDOtE8SyvJazlgOHP/YR4VFzWqr52frj02LwM3M5d3X0bDJs/UKylBWarmEQ
+/sozhuLKIHuEiPfI9dlodE8N+RbK30kkbd2PKYm+oKo9N8p795CLE+gDqZEi19YdUFEuRo7HmEO
I6KJ2xTVs5n3gzHXcwktR3G3KmlD+a43CIUVrvR4eolLvI++MU08HVl1N+uDGxvPNHofNl918s+4
v3scG3yA+P5hU2iWlHq397dSd4D2OKpfRWYshILK63A3WffeNDA+cdP/U04d41YFCrwkthXqygqx
nlrJ24EBL1JOWkD4RXFBVAFV0kIA63dyQY6rKhgiaRBaI3ku6eOHyNR9IkjSWISIjYyi55XM4UeB
zH2L0kNGEG9tBb3ks3kGq++iCwDuMzB0Ps8KZC+rGUOu0s+vXUZRhLTDwcMpy8F/0TdlvlXYKvUe
T9KialxhBTqr87doygyjBxGzXtjmvvxKEVxnky9L8Rnz9UaYhrnzvJ3auORUYbE4WfJ1+DjwhRwS
mxUasm5gX+nG8/dmd/w/L3jEp/J/mEwgzkIQUVKdeKVkxAvlxNa0CLOloiIcclcUOvCrkLAU0MF/
v0b97vH/H+jww98GVpQERrg81605YusLG42IixvI5HFhswl6J3kQoBf0/J6yNRp3gFCNUT/FDsDt
LsM9q/s2eVWc+FwTh48svohslZmZV57xqmdu2Roiu0Kbq47hjJ/G6zVwzz/yUswCxpiDoOkhIYGd
gRED+HEDP7ZZnjedQkrlun67i2xmSrG9oIINDE93pA1eO9QwnfavkYrnFNN8csAWzmKyS1dE0I5+
ov90UVpePoFPK2eNH4SOD9n3sZnI65qTbzhnFmw6TZMaxThSh53Fp7f8hWRlzePOGxGLXlESoNx7
dzBgXEZgVexGiTWF7wcfoDLGgN4Dv1k1R4xQexJ/ay7FrXwXWucDNZavOGCNnmeFDPdSPdLBFsX0
mY3lMGsIDU7jUIMUXp195so2n8Hoj8/eFCTurI9b8VO2OcDfe9n8X1OE3IiT1cucGEQzzLOQJ2jR
tMSE9BgZJY1LbsWgwBHv+QmevGdcN3ePnSz1ItTRhIHunEpf1k1s/9VbChmnxxFqhx6BYKiw90s9
+SccC/Qj/ZitaQJ0WiRvesno8GNegw624VzDBrV71DESRDyTax3R18W7XGX51GfFyxh4fSu1WS48
n8uY0zgPAVqfBwd9X3wzTsVaRgfr5hOyvW1LtvSGYlHT2voAiujicY5O7IWaAuqPHU/vkgR0B2ol
mcFB02b2SVaHHsKIBm3kxLSePUt33EyBzZ0/p92j6vKVSJUOzwEmgDpMfnhB+AX3LwFfuyskOuto
I1l16mjGQGktEXuVnkkxC7IFZdSixU5j8EGslGYxjPS3IL32eLAbhOqTX+zqp688PxTSyn9Mm2iT
wTOTvNg7y7gfK0EL9J2TXpvkiou7Y9jCUKlvxsyh7A3O0hdXTyauU1glviCiCqU1s7WWf84i0jtD
nwW5fPokHYKrNapVnjsia6VDyUJSyPvm4IIyAMMfKBI1k4ulKct7aKprHbhJfJyIl575T3h/Cien
DRdVFhCuRqG9h5e9FLcIUY651U5TpJWKCQQbs7f6QU2PXfVmIHNXduAoW4kB8ODAejQBXMNVpsDC
BVUar+PxW4n/7qtntDjF5QTPM2ITWMClJSJASyOxrWEfmJh1Xvlm4vUMJzDvVnMo6sUEqTmdlnWt
xkJjnAeqF7buExZrvzdOmNVZ0sroMgWOEhrqZ7FGW54Rf0MGuS/6LgeHPUME5rWLfj1KrjME0piR
sD4JnV3RClVeFiwop9paSEQ6rn/C2ZWDP3cLWqKF913Eid75NqD+kA4eK4gPIw99NdFxDPROCKFS
mu3tLzL9imkWtut1cwOrfg5SWjS5psCw+HLNI+L6K6BL9r81qThYeJd24P5Nv5P1ZmWKqmZuoeJz
5PpbiFnHbP+GJU8KYMNtUUHgTDotPJJ65L+muP5EDOcroJoJCieL4JYSBpu1iFCZ+1dZKu2UipHk
fAMztZRupEQ1U8fD3+5uUI/TfO7aU+NH2JnKN8HImE0lynwTSCWfhMsUNENcM5E9RrB7rzG3QjrP
MNBaqTmjhNop2/XJOUm2id6zRzkH8PUhDbh0rGynje0vr5hMyxDh3iheE/ByiNu7rP6qPcTbsg8N
ujNvY0N2IruXZYAZ6pSVrBFnuOo0SsVaXF5E9LZuIjm69qs4GMwcubFd+LUqFNnOT/Dcup4vpHfr
WYo40ekuV232br371q/p9D3sgqY+YWNspOuWLecWsQYUWWty9qB1ZwafFrW+uneivVSbW7ylQqJv
vwK6ly2U5a+r4XdD7RLSvXUa42Pq4Vv6VZ7HzAhNgtwuHHRRXYKgXXJ1OVZsQb+nkE+OkT8JGhej
K4dMeKybKm4Vaq7gP8y8RbXYqWvqvT0OSciVgASSHUKhCXQD3XKfJpumhsURp1EZ1Nii9BJ+Sk6z
QYstgxJ8Fv6AlTy0/8IZ0prW/sE+PxQ2E8apY1U6DhQ53kBshKZ7EKKgvNRUDeMghT1WTTFsNzU3
WT47XmQjAtpLZH6kPw/h9hgbj5mdodEK1241WaY5HCQ0PesYgD7ejVqbQncqUrciOhiTJn/RbJFX
amyeCd8ry21uZh3ajG3dtKfT/1/66Mydmtvj1yfVDf2mrUA+927MZE+1hW5sF09lkP+4LdxTVSFd
5FGWg920cJvRec02+8br/dHWJVBPGRbTGp9I8BAFqkSwJzhMSsDlep4Vwp4o4UyL/TZgeOuRKuPl
F3GGi+SUGNjlCmQ3V7TKE9FSwi4/5m9zYjh/eUxyD3YuO32pviH+CLYEllSiBjDbQZ5HbVG1L+z5
GXQZNYucbLhgzdEC5gMUcpXgqwO11YsRMPooX6o/dVy65/JAKWmLa1Cqp8ltjyb6WXmHhtC3PajZ
cmsmRPBpQPNTRiydYyNlU0w1cz7x3Qy3xNPBHhXi1hejSiviZ2HH9lc4cBpJJuhQtnuEegn2d1uQ
5O9eUNpXR4/YKt0i33hpZZZXbE+tl/rFgr6pobBqSrisR1dw+2t5btB1e84Uw3wqdI5HtK+bLNQj
y1nYk7VgZCLsfL4FvjkXoRHCXrKw8oCwZE8lRNExChaoqpw0NnACWPKv5NoztlD3xgFpjF1VH5ul
5zZ5qRwkH6sN+1ZDETndsZ9vp+lBcM+IKNNnxaLYS++8077N3v1pVQoefMRsi1rUdlXv1a+k192P
vTFpsU+579YzcJu0v7qwymX/1ef5Qp2GZ8++RN6m6LkCw1hhfQodcZxWF98S9BNvYh6UjyvBNvQ8
sxA+EGHHpF/5gYg9bICD4KsjZCUA/cmYeuPJdHoQXGkHSi2Xp2IIntNhygn6VdB3UdkaDtzulreb
5gmw+L3wDQ/jdoxlTjA4mBBvhmXOzWFl/FSznQky+gISuHxRjqnzRwKwFf5Kbxxx7fEQDcr28vzf
DLYPnhr1Py0qLqjHg+4R36W9UTKgEVhLXDGdYiX+W/K/c/yZ3HWY+EqWa6LaGkjMsLJZ4EFml15S
nWdoygTn16HoD2l8nueHBJyQQyOB5uAEyTbdyOYnqMQNSXDe84x9bsMUf/NQ/G8IWa0aK+y4qYYk
4XC0F9nRvLlgSqqRRkes1jU8bgotKQHp1JAzXqIfx9zRr/mA+joUoYYGyQzd1e5qS5XEFMt8O16T
Brin0WtrH8IhX2DlTR1/CPl1bZ08EEshaNpmLvV+8xuuf7Iy19Oy6DUWTdUprZty45lIhc6oItUK
civY87kdhDmWOIB7j3MOrou8Xu3tSGvhIhl/7h06eCGiqLE5fn2eLbzB3xVSrflQFNWMSaaT0ivP
cTFe9PRtcYCnxnb4KhtNoNLwbHTIBqW1T3vc/qsuJIk2n2enpLSCfvWROlYKI5mmsF3ADqx/gDY9
oGEHUodXoLhuI/29rsQR/EJpWpdmLT8hQeJtafxfu1q8ej+BxQbcK1sWe1elmC1LgK0NvTnTIP34
6lSCNEqjPEq1ONjlgoroIO32pWlsDZf/bVMaVy3vX9yDChvv0/fu+Y+4h0NMHt95pYhdcaQLIIdX
BwhKK3Vz7saZwUynd19gyKvUEWgUAfGmDEidcOsQXeBXuRdO3+TvAHhEBM4isIJP4puCqRJSc+S7
iww43M1eaLd0ti2HRREuBNbG8xlabeTIgE+/0bAyW0GIREZ2qSQdcM9FP+K92zclqETaiDILTyQE
E4+99c5L7v+9rXP4i+6xy7JtInJRqRNCx376lIeVE/h1E7HY1zIGFZAIsS8XjTU4BKjadZuySQOa
jZ6m7DZaRWk9ZR0JjBYArhWarOkYoFgpmzKwAKVkmweDvxwcMORXXgCCy+fRd6A8L2m6q7eDifzU
oNxVwsCGFXOamk8nCV4oDvHwWq0Nl3aq8E7/Gjq+xLangvVq06usMc2+elznxjHMFdxZLMSIEYn2
X+SPPnPiGRyuKTBaY7CqcMZhwiDLz/b8KMLihqTnaIlVo/304cu2tnJxbRH8F75IP6+sMqI2aThk
l10X8Rg3PXLJ/Gh7d8qt2RgEUIEkRHU3n8KfH9oIK3ZK7ZT8trQzG6eqUF2aTlZVu3f/z/YMqfRf
2XgihY5X31XvTq/ral8AZPZbGUP1C8+QjV6lsh6cVlrqlBEIGt1f+KlPTkhwkzXBO0/281jZGKpV
jGQTLAeBetJe7fyefbwDslOict8r8Z2rYcf/hq0up+q8g6caLPZ1fiVls9ilwfnKyI6pUAqrm5vp
Y6BVT+WNAm93csAnledcWxWqcqF2RcqwLavanA11jU+vmU14+OmhLsCWfB2N65R1WwV2jQiAXUpK
eRDquf7dlxbEyxwdYu1zB/VJ6zyCh0PvtQ1XbEsjvj1HYmJTrVRUfgDa7q7qRhaLFFYvLYhSpz3d
4uNvM1GFtLJEo0s4eQ6Qf6DVnfiVUkx2fXjHQVJwqGFKyjcuaP7Ep+zuCvKjxn7io43qyV9zk9dQ
pufW+knZ6jSxoTpvjOFn3wA5gfhIojIxv+NYMDcEGtEyvJrMnAi2moR+RsM9C/n0PxPMCf9doAEA
Gquwe0cO2NHOOFmSx7Q2zB/Tfe84Iavp5Ydeq5Ta2+b5AVaamt+gdiywqa5o7J4K3bgn398PwsHo
2+dzYdLkCH+mwqD2KUK4mIXn6UIbHD693iym4PAm/6B49DFPNVxWjnTEx2zvhUTinzBgZRiqKfTY
lrnNe61lludLSt6Rsp124EstRFHAn4bW9t1eA4+2XzJ4eIpMPytsWgqUDVj6rE3Vqs3bpLdyM0l0
vWzkvTUXttvdS558iv8ciyKeyuY8DBeZHW0bJJR6lnsLD37RGGP1KiBc66qY4OrHMGYF229mcGvO
zPZ1wDJDkKbo57E8KxOO8sN/xJneEqbd9mqL475gjoSRZosIdbGE5bQqlF9R+Sxebsw2sqxmB2Ej
A/iJ9Js4TiC87IdBwSP6mOC1vI4pX3nyH4/Fs6RAWtDfQEXZMnyfpT+5HZY25PMaSvnjzmJxGT6R
Tb7Wpk+AMPVhjCO1vebd7zD2c94SQziHi3wRAwbU377yRmZJRtOm3emo/UD5ugXDZ6ONJXxZjNwy
EtxQkkA+Hch4tl21LIt/Pw2WafOVJEb0A2ngElQZLNsGynaH5pDnNyMaRHFb45v9AEmRW0OMgVGp
rCyAT317O5jWvsPZfyUN8xK5D1PTziXSSCRajCrX+F8aQos5bgGhHgM19wIatBtvPWgL3zyjmWcD
sfmefwQxEQEJk9VEH4xlkkADMzNfpzBMjoULkLK5JftgQBLcal1iunR1CZRO1B8jiFIYBO96J8pI
h4DivGbemuZPUbTPxF1EDb7hCRYx0uXxgjfAAGJp7g5qGbrxl5gsOdE6QfDZSuM+r9hGoA3A97xC
zsuawqWlDoAC5xh2tX8vVpBlIdT/P8GgncbS72kKv8Dk2KBU2huaOljIoS3lSof2hemhZ+boJMba
hHTmvJtGd/kI9MfyPwKk6FXCZ5lvD0boRacMaO6g3mU6hMOhDuPA4YOGEZVFw0sjC51QDDqYqlHm
Mnl9ZKBf6gi4ZhxhVLrl9NIPLuvf3IDl6lAkJgXMExvgrKEvkMgw+Y5TxfvMq9ZFZ3Bk9mZoClXC
vYUTrlNExW4vEzVCwp3KmtnnLSwPOVyyWwYriE0z2DLUi2TdjtiVOS4rY25z39KY0yAM4Ga3in5M
A2Z+M11943xjuibhH8aCxVNexiaPeKRyCUeBL56Vixujzv4vCRtV7lKCpPlOINDbwPXPRiwmZD8f
nssXoLxMSZsAneQWQN0zLWJhKqV4/hK87Vo/iGtOJGQfCn7plcymoeo8R6T9cvmpPE2s7dvQFAMA
Yg5IHRnFMmOtqkSEONOBWRJISwqdiv6vuVKlzfT1EK0uhBcNqRANthdMeyX3+UWxicKO5ByunWqZ
NplVtHFSR79pUFQyH3ysnPlyW9VeYh8kiwax+b4htncX6OVIuUMyTgp23PL5H2x7aJhR9ikE1R/Q
Vvx8F6/hU0RSr9Sm8okpjsCB3rsd7+G0KnrIfF+XfWEjPgtcXr4cUYdAS6w9XwBejo9TqMKPdvOa
UQ2Tk6dtEPq1voEbrSGqnFklWNPdDQf3dsakSuXHYOJLMAmftCOfG2t4aUgZ3Pex7Bnp60FmbdTG
tk3LLIkHLZpVTzJKcpATUbDeSFQS2hAKMiA5750KXHFKEAwC9UzcY69v5YZGRalOu15OBGWWRymy
MXBiD2rOMfo19OkcKkj9NFYzOPDOF7r+PVMATrksIIgnhNf9RT/H1gX/Iz/aX9Hh/mm7jvHk6eqL
0W4YgAA+rRdXmT863JDjNDRqzRs2PVAtf/XV8jzFs16UsPoEgcNbF+IaMjjid0frIBub/vNrlGAd
TyXwZyRNym1081yveTS7MK83hf/m0XnJW5oClvxu84GfBVjDMhgD+VbwPzfVF6Bq+jD5rB16uzSi
cdOKKUNXspmMQkRLIgZKCA4gcBviOFxyWVpK4rvhN4/r4wNATNm+uUpdQRb8NyXiZS0q4w7XOP1r
Z0gUqQ6KhWTnCD9yq5ZtUpmDFO81+lXo4yQY5Os/Q+RjHEoI9DQQBuSF7iuprnjH4VRzeziu3SVn
EZo5FbZsDnicAGjHYOIIB1I28aS9Cxt7KUdf8W/QsoE6Wgi+1JAeyL+8GYWlQPfbcFz0VIInD5y0
z7hvxp8Ldqe725eYm6hp5LGGV+gnmnqG9Xfw6q/qSe4ldl+Vo6AuffgCo3hqJf54gjSHgAGHTZ60
Ecb/9zG9RfS8z8/vRI2ix/2wEaf+OlhPcNtsC8feqWE3hYZ0+6t4pZ6BR+eGm3I1kHCw//u/QDtm
zG5/gUpq4Dihxx63LpEeXHZGm236AwBat5wq2xBvPkBPnQ/D0Kr2j3yAIXdNcMD05oTI7JXgwRDq
MwAjQzZ//alZOUPT+JNNJfSoy0CcXNOu/7YohcNOY4sl/+qtqtNylm9uTEIy7/HxE/VKP7sqpRl1
bjtRMA5cJt1PDRuhy9QejC51JShw8/5tqUixXgHv155CxWd+dhzvTCPNYak05AEUkcvb+twZ/Ghn
Wd/rI8a2MQ98TlD9zR7s20/ySHmynGEVrLTnrxSwBcrAeNLNPccJeNJLQjmvUp5keWIkcDiVh5Oo
y0iF1jt7X1VKxk+kXeXDCaNth7kFcIdZypDEXOJFcsycQJTOhyB65WNdZi+yatbl8EBwOb8n60cK
S2fpjXq0sY8uDDsxC0RUlAqgVS8INXLMaM6Lg3EhiPIRfkJr2lb5jksCEX5H7RIw0wr1G8Z7rYIT
b/x+TV8BUmQfAzboPN41p2UXqD07ML4DMEI5//8hb3eBcDljbQZba3+tK7WLX1aWNtz7hgN3oPHH
nbJk87OvtQoIf4/FyW7Lk7cJqWfXqlNv+ozu5Yda144vgo1VrMD2v+wHmeihuXDvvrX5lFprcrEb
pDiPQK0/NknuHsBCYLOHhS6oDW+bY0Xt6aipHX/Y/3hZg29iAgNUAgkfxJEXPiO1a0Fzc9j4kh+T
st6JcDhi+KeShtqBZIc9ZEErZy+uj0U/9JudbVP2jSEjuwFHbgTVtoG7PLoFC6jBqpa/0zVBDV9X
4FuUz4okgNJ5oU85mUnLXAXWPKJv4wTVYEiz7sCd2edLfODGN6b/74jTyiE1FA1cVvDSoYAYn1K7
PhLa+igZwOvEi8m3OtgBKpGKorHCxOsD4DsgXSVIrDniCcar05RBb+wSbNlUbcA6DB+1Lsv4MA5z
Fl3vV+XH80dtViyJTIbTwoxANGq/Ig8Au2/7wIocm6NwChYcl4+d6aO09LT6M7KTq99fqkFJFQW7
5F7vfPwUmABfyf+uuUr+EWg5fbWiEKnK9cLfi5QkMKmd08eVNyRYNLW0/Jo5U9P3AmgjR/LTVNts
EYGxMJKmsZrkqtjRc5C6dQ3NcMj6bvu6tWy3Cy3TcoYHK3OAYHW4s8HNA4ln0Pt09nx2Fmc41GsK
R/+Se5RgQFleKUU4ArxUdY4N6XuuD+w5saMASybtCR3JruiA0AQwtqhLS44AVAHxy8wkwNF0x/rz
pUo/rNrho3Vxdu1bdq9lwRegCL5yi5C+dkSm1a9qrfZ7vuUmHfIlnmyhnGPXLXeIPyF00NlGjbHO
9LRHh6MNgf3ryes0hk/7/x6rcpnF+WOl4d+4+Gtr9y/w6dBpqo122LI6pbAErs0Otn2Dd4FvCl7e
mxHmU7TYddI2CBNRkN3agpfsbmgzpiceiY6NZKTABf5bN60kxB8aIE1E4AeKdZs3LQKRrELetUBj
kn000D2XWGz/k9Snyd8SGT0kMGqmZBEIhEhApfs0sg/xjTJv+k4Obf+cw72gRfIFDifG5R83B62M
gCJ1xfPUNSPBOYCafl1Vva0pbwW8srpXF/G7yFy2PuuWcRwavR5MIBvrHEI+1OdW9VJAFfYwfii2
0q9Saw2YFetXXQjEClt/wDlyyb/MPmnxYOe5us3W5CcZpYwX50Cx8xicU0t0fIfeF/xpj5C2gMnc
m9Zzzsx4AuBw2I6RgNlFZbdAoihhIa6iX5XTvuIV7ZSnymiLRLGDALESAgXklEmzBcGcx1EMku9i
DMZ8HPxDgx6VaL7q4nMlVs/B6QX+4OjK4WFizANm3d9hB0Z4c67Mjjdk2Mon4//eGIhAF6/rDXlk
TJrFqg2y2pviuTPF0+MCuQam6fXGBIqHa5pfd5HF1RleXy7VN7Z/ZPMuC+JMFRMq5Nam0YbgxxRJ
9mb5HDeMd+kORbsJoOYV73LfTLyY0nCSe/HhOsRSYiDdLcOMDG8XkDYoJp1rZ9rs6Wc9GX7nfWLK
nOpaatadSDAN//AfMIzsK9GVC7BFLwoDKTCcqGVVEFPkxZYxprACFvzWJfPz2bTCxUmx4Mj9KvjV
i/vi2NWyxFig9TyfZp9qz7BwxVMb3iQtIPNxS+ZW/ILHxcTKPdIE/+IuyEfj8QTov0TwCMQcPY6Y
oH9IwHiUCbaaU6HXsstMVJ7XamKokOHtfy7Jl3tskzgZxur/1qjCbgXmB3JO3p+f6H3Pw7+HGNAL
lFJW7E2CqFJXvneR5orBlDYthhqcSA/Q/9Jro6f65qkL54FDwazzhUa7flReXs37zlmUU7A9oX5k
Sq0wPLYdXaSG6wGC1RvwdqT0OUOOzWfFmh6wi8Ea7R6vuJ2I1Dw2PvrEEDa04oFkGkYbbsz/w0at
oQRHUoa0r12BTJ59/AarkYkzphl2QEf/B1n9heAzJeqaAxeK0p/c8UqHbJTW2DqhqxJep6OaOpIO
yZyF248VFvv8WavGqWSZ14gSZM01fFycoYb3aWG+zvbPF5kVRz77XCPQ9Ka9Q7fwt3qtuePR17bg
S8XshZfWvm+kX7hpPabU+9vDb1uoiHoS2Kwyb4mb1G7Gy7dJPzyHd0i3wE+lRWMu/ifbsCBMSV+/
kiIi9jiV0v9rFJxKb5k8RQa8a8wrur0ngVyxBCUCTmpD3yhZ5KB/kFutXbQCDVjnfxAcTTFN7v8h
x4FwSHWeGWalW8alRLSF+HURAp8OGMf5zFQOl35/RfaDGE3McWsXeIEsytkzt5UH7r+WIhfrBhpG
3gj7+4NKELGewif0xs0KHlb1FYH8AfxNCRg6CHsl7xsU+qpz8qLq5BN7zZg8UzWiO+OQUfMsJv0v
HtR1flWb8qxjSk3DyHo3FQFWLi0q5N+cGSsdq0UIKzmZHjh14baHQ4mtCWUGqxSSDnKEUQpKKAiH
UeC72s24+BbvqKymxzhRiaTUlo6BaWx9+uyrtuNTMMNsjIqL14YP7fv5GB9+/eyahtEUJ+7K3kHy
HcyQ81+wR5uYedLmOzbO5o4eP6DFcy4LixKl8OyXUiAb1M52ZOv+YQ3mQad8LdMdyZJArlY/Av+T
enJFd8/1fGjedVG0lKDUSPHGVYosFYlFm5CqdZUBEtq5+q1ZyB91pxDSFqpNIgwWir3sA0a5Fg4f
PWUlgxWY8t0w8bDTIroHNipOpDqK/K9GTI+IzRs8E+2cayUiuxzVVchO+wcDfqxAq8+w9l8Hj/J7
eYG6fOu80ZRgvxAFE5WNwl9j0MiSZb3nsWn1Zp6cilE6evzAbOll5AU4Mqa5vDg7nswHhFOx8+Dt
UDK/0kUmKF1env4b4XldZ7Nk4paXnMWApYoCQtONeRAQTDP4bj7/6KJ19IrLqggAc4huS4jkvD1B
mfZZlt0WOJl6ijHiGxkoYPeubeI8t09nBuvjR6dP/FTQQFq+PUwFZMCUH/aNLkod8bH5azA5n2ff
gtFq7TtOam0vXLWmI4XN3Wa6MvcJhOTv17PZ7FBqnWKhHeDrrZnOLtBYhdCg4EvcKlR9eIfkTU8W
2LReKq01r2j4cWagu5Rnij/k4mFzKm5EkMT6TMEm3lcQagq2GiRz6C0YPyegUos04uV5CZDLFIwd
Z3hAPanCuXXui15YPSvbIi7MqRtiZmPrZdBSLekcDywFGzpW03/GIapg2LMovUgbWNitTOmQ0Mc3
DPs2I9WLZ43vZBOrPMXLjfeHrHHmKP/+dJg9bJ3blMhkO+OFI4FoX4plf3IVAw6f1L3kAsPuezOA
dCZmnfFCTZwTZBGOgAoFuGyz4ngSkfEmsx9UmT4OGroxo4aYSeWm/aFflZRJOeXnl228ZNDFaZ1g
4NRXnk6KNvk82oHgZWu4tZImkWQ6sjqtRp5oBiB9+IeQusGXX0aOdik7NjDEoTZ34B30njyB98r6
hXFWw5sXCHzZfo9wwgJfIR8/qnRsmd+D/nEZlYY5a8ySRfWqPTiIq1+aR6DC/s1x8+tnDgAjA8SG
uj2E7/AJo+Q/Y1wzXPSpwnMK2wndiQgUbIat5bOD66PESK8K4R6juMag7fEc2U9xunFTwIlLO8RH
2zhjoQx9J2UOhRYKriey3MawoSLYl5j/IQNZJ4uZB3HYIZxA1YNV+wxQjSCb3R+y8WAVFfPOq3B0
eSdN4gY2o79IkRj/rRv5y2lGROPRThGm9XChQuFzgcpI5/0Tk+nZKGp4C2Ru5Dh5Azmimdv2m5eP
EyKgNam+5gZguXC7yDEFs7mnyUPoy7h2C++WtdinCzS74Eq1mFQuXIFTK/KJjL46KHMw30oAlHaS
nXqDKB46Xih2bzzLoVHgf/8bpZzFjJd5ViwbRqhrGExjANpXK+IhBqPJkarQpYC5sZuG8HMVYmAk
phZhP1oFksJgz3lBev4twV8LgESGsFjCLpfjh7huaLls98NL+ijEDlzLf+GU+9vFUTtjEaPfS3qx
QHx9WPFFY07MeVMknZc3r7+PaOE2yAAVCtSx0ykgr7pgZluixKcips0feI4qZHbR3yXIhZW/Zzcf
X6BxU1kKeAQdi1I9TVcFN+a7yYHkrm+ne5AWG7m3ZJwRVYr/A/fx2b8x7XHGgaH5bU0/4rEHCOf8
4Wm8JFoVUzTAeMZiFKolWRBVRS/G1j+11/S7qLzVYU9KEpWQl7Bl8PNMv+eVm9EV8RUwUGKU0hTZ
M6UeTPt921vbOYijUBi3t26hcJlqGGOeykexEyGvFMUnnU+VmeYJI8MDf1+7oLz7XFdRiXQRraf8
Ayb4oRPNeo8S2qGq7eTzrnK+m6XfqRogMHBocyLYphMX0v2HKLmtuoRHKdETV9eouMrGVJOUy63h
hC7vxcCKouy+7tjLdMNmdCp7FAapEc78EtluQTrbrMqzZrkihwWq27m4qtJG
`protect end_protected
