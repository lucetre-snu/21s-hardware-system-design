`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g7azmhtm6FcP7uNFjuXJjN8Z6yccOPk3SSjzvKB27peFKmnPmQmov5+YTGwYqqN9LpdyiUExk8K6
vPnJqontvQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFrqn2K0Cr7TmQ5al162oDGiY83d+AkTWOgFyXPYrTNznygR/tx44RAp24ytphNK9p6shs2EFMg/
Qqz0l8DCWiVEoJ/T8vMpnAn7Y+poGVGS1qAR3qE2njrl81VcGBZJeFaWIudhfr/DLTuuf2T/dWDU
YpelM3KbfYNPPiPy8PU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FZca5XZouG+/BYoQ8qrJTmnJanku4IprIWRkO6VciHehE5WehR0wsZJhfKlqLEeY1oTPA4bXaxmY
NjYkrop4EOwW8t47/hj2kFLI1OKUAE/TAhCGg/aNSOViUbB3dUomG/y+TBuDt9L6g0Arj1vb/5Pt
IChc5ZdEfRr1lJMTpFfP+5qmEH6lePPdzgPZATPB4Zrj0P6EyiEsU1FKBuAKd9iYNGiLCxVomaz0
3/RwK2Nl+/l4mc7PJt5Hso+4s1qHb4s2wD+OgbIwdH26ZkEnKVFpaLiuWQKu9uhDLGnsBMPf7XDE
p29f+mrvP9Zi/3nonA2aBKrTwR7XuH+ZYoakxA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jP68OjlYJglq3zpmKrXOhq7Sex8XNW8fQKp4hUNmuw06OOoKhQASNTnjtyVjAIk/VXb64ViBu1ds
cNMJybDSWBhnChfJq4h9PNybShGJXxSm3NDOo5wUHKf10Eti3fSotB9rVks+tNdTEZo4O97kgfdD
G1FNOqlsYcQiShEGLLiEQ2yYtgJBxJ+jc8mFjIEfPhAYy1ElrvtFEpnhkNS2LfE7xdWOQdO/XoKK
ibeY08pgncTI3pvO6TMbXushf0AX2S7hgfk8ysZrT+0gktqFrJnyR6oljS6VVPLtRNW2vo/cC8XQ
Bzvwwt4cpSo5KLS4XxB6qClZipItck2AUEdIbQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o7jAZIoXlFbFtDYmtXhfRBlb07dhBb6Wp03mlT4T0FXtvccSHWhWZgc+VUNwt6TohLihOwvSipPP
XVXpGL4pUVYNdQBCVpFzhMkt6jhyUgsF5t10yI5Of6YEfQrDHigceoBukM3+/zJHPprrPQE6FUvC
wXSGhBCXnHJs1R+n4l0714w8/WftPQhlD9QGQp1qT2VARQXUKBRxcRjxe9TcLfs0P4xnN7uHu0R6
JTmV+MHmhGpetSZGx+B2Wa1MQofUPURqwE70IwBoUhdXH8+39DT5I6x2+wMY6RcVATnhNd2BCgPd
RzAhwfrcqRiU9aB+eNNdFR8ve9M2nGMmV2JxZg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cl1Dz+fZIDYEIQuUd0pSg+5jknmtX/JERd+yOZ2SRaVra/4pU/eCTjEXMzhz4VFGYB6dgUxMsGBk
nL2WNdn/uaSPpi6mNF0UHQvZik4pUkYPrnRbFveVqW8i1t95SG0RW96uD19206lWrp5U1lqc4fH7
sfKHi8ZpU3MAg0DOO0E=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qqp76m2aV9ue8Qai7QUavb+lhRYdu/txrnwYLzwTe0vS0S2OD1vxr8VeIT3bF/ZuXlTGm4S/UCSF
bgOPp7VqEOeGNfsSPK+VpQ+foQMENCQYccwKquBDSg/sLjpPK9uuoGLBLxjw2OwsRzplVFXiPcRN
LYK1/FmCP7RJBNgmhh/ti99a+WSl6i2YIIRGocNplQlG8FXq8ZTTHd/x2Gtdf/zGvJOy/fNsos6S
Oq9yJ0rMmbGeWbri5c04gZM08pUmXBsivgOHm2IVEZZFM4SBqrsi0xa52hs2kelc3iKJcWiTvU3X
0fJP9qNFuIjXBPPZvEYwhVtIh6DwiIC2viSscQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
Zb0iWcIKs0k4nz4eYC9VsLEH4At7d1Pp17cCsw6OQVhCWHsWEKoXF/dIH5XC/saMZyDyc5K4d/Lf
g/wq6BiDeJ0OPnYCszr9FMVzjilUSOr/SHUL8uLqUf3jV/+yu66aS1KpM2yVKa3OaT1vGpBmGaBS
OkDHVFntaOmu5IdPpdGrES/UqLfRZt21YWWFys6DcfNdiCxDqC7hag/pGtMO0qEmba1aUfp9L/jg
ixNKZXN84qKl+NoO51qRV4m3kWAQa16LyeKHiwb4o4xs+7bmHJn6NOh/FDmR3qMhuM1sZaTGJ5I7
OqfNCnBJmUGozzGT1BwJfNmfiaL6V2rsGc3FkH6NyZzJe+xFzkbrtmcTmULmsujRPYnrO7W8rLbe
xh4KmF6JJusYsMAqdUqhSjIUmY2ykyYwV74yAHWc9ZfzaIhBBvl9Ll4PxX00iMwJaLZlmjjfrjEl
7RkrrOOfMAQl8tg1pPSGLa+XvzlVC4U1uydjpf+9CWg3TqZTTAgNTxUQjr5+BXQwJUJB6uWhIOUE
r+XCA0IuTgcNUbvsphB61cbCBiNVKug1I2zaLG4i8gzJTfLfYXalHxz1QC3qVAr8JX+lgdd3zmcP
EZBsOA+W/Zk9yA2CEz6uC2aGpJJZjKRHsGKZcTQCwVb6hnoXpXebUVFwPbW6ag0T76i+snVrclnz
XFv9ag3Ecf06CT5wcdNz9vywBt/FvsLzjUzpy8aoJBw0T+TGf30J8YHCJ9L9xVkmsMCSKstM4N0j
Ii8sajNb2mXhM+nEv/E6FaCYR//NcAgE5PtDLF/tZlxQZL/692mYMeEp9gSBL6D5Dg/+MSp6TUZM
oV8UMC0mkjP32TzYXDqW73+AQO5TlNtGG3RrWthy7qcAwF+fyKWUGHk+7C0AZRBB4y2N74nfB1o/
yl7osLFNeGY1gY4Qu0LhEzdng87q9VGON2dSCKeQsoig1pfug2K3v7MxCYwy2C4ZVFEs0qCUiszT
rEU7GO3meVnQFJf27bDSnzGuvuatpoQ/aneKYPAnBTPPl6ivJR2z7eDbwqeigBwrXWfFfQEMjPbn
BvtMG/UBnyCsftClL+qM8UFFAxeKZUdd1giBvJ6B7eZYEd3SIUoaMh+zAnV9aX6IMoidXcT52XAC
WaJ6MQCIzoUgooY4eM0pD5OXgeXHUsYezJPIciDhx34pSkdLmGGs4zDXFe87yyoYYYu8xiATq+4q
ZUO4PcgxmmIyMVYnVm9mFbg/HYJCOM834rXOAUlnUbWVypguS8rYTpNeBcHrSXl210Dd28scpa6I
RCJyMCEsf1jfovPqZl3w7dh5eByio7cZLaWsTiLdMRAkjfZ00vPwB2X+ZXpkTpZCyZwUIDfdmAYC
OBQfmgZm0LwaBJx2EIAEARyMY0Tp0yG+xZvlxbr6xmxjoKQpHYWRJXJxTibfV9OQRPpAjHcFvFpE
IoDm8KT6LaG0dbgM1BaGZTF1kPoucBfz6crQRZz5xCPQCYgHRctG08Q/gtOrQbx9zNGag58+4FhM
JJhhzddnDfrh92a2BWPkGfua66RWLlcTPQrus9Wyd/FHMHAAeZb0adUv9JpUd+rwOesbuQk2fiZY
7IL0IaKtG8K0mtqjKp6ogLQPu1k3cV+MQcTzTZtf3kXjOhId/Ce5Q8nkwF6vUiDJJke9EK4i8iOR
mYdnfXVodaezy4h0qdkXe3qRPwUe/2nSBE+YLXUVqaWNsTX9LZeJSoPSx6IBAwH1iaUh1/pe+rI2
uOo4nGPEzOAoHUVUuT7tgTBNjybWe01pl663+EonmtLDkNfGiaRRfcpmzxSYh3zWBIJUpD5qmtlg
OGUmeNZU0VFY49x399y14ZZIawqvFrWMARdFANWTzpMaUJiRCbLZoanW8Auy0wbfnnTQrsyGoZVH
vZ/KUn+ql02FeeJwnIW1kPQvW8QdUwrk+bMpf0tmTTqj9afkfIXhf1he1DwkZc/6eSvV2Dwxagci
9AUai1bf9khp3Cd13badEsv/VCCheQvnsmG8F1aZ26cHrTWzoAE1wlc9NTL4cM+kR8w6AxGyN9kZ
M6CjcQekDq5koaeNWse1Zujz0pe9Fd1/P8qcsBKgZ//iZI/G2vEqAy5j+5SOBmRUD8eGwqzeq7Zw
TyV0BTts9ZENpE81mXqoCCyRNXuPh0WwhQN2HP0tobws3+v9zOTM7qNAs8wqYjLI2CPsYKX86iFy
Eyob4sCXFzSEHmI3QJP9bQTtx9dzkDY93wHKHDReFiH5K2WvPs74K6NJdEbpQf/C43aMcHQCdNZN
KXGZvhbV5kehi2nrPgA6bpTTUhDwmCLe5QEPzZCGwMd+9ztpX1FwO/uA3ozh0/DCEavZVXEMNlg1
Y2/L+qRP7A1XCoSRt86BLIk0DtG9W9JLNE+TjRx4sBl8dQ7rLLIzyVFv5m4wdoPyqMWES0xeVHal
qpQhmbsTXt0zvAtmoWzUXL4+ZaiWgi6dfTlrJ1P7BAX94sGTP5/l70V1vGm3Eq2MmxWKqj54/7sb
N46QXSXFGWM4AozV6gI3cNtzAXVVO2g5eYPvtD5welAubfmbQfa6oVNaq2O4nUJxW42QzE08fNAu
Wst+Zh8aSo/XKhb7mgzivSwSwoaPQcuAywC85GxfWDP/fvay+BUmrFw97EfzMIAAwwkrbYFvYkgo
JfqEYpVfkrXrrpdM+5WviFTOxIclzX+bnu2hG0PHYCr/OvlnFnfb9gwUH9+e7G0X2WoyQWLMHMmu
hyeJIhsDIA078oPZ02knX3lKpx8xWNj33z1i8ypnoUbvqM94Ng2QVs36mKIGKTvyBGOSPUPh5vGo
gaziOfUtvTRd8UFBkBAtU9S8jcz9qb/dAdvhCMCyX/Hl4ZuJdqiuocg9gkyO4uoCXx4vF8py5iCF
blYoT4EslHNN9/rUzorWqu7ovgK92DbT47Xy+Bq8WFpM22cUBUyPscbpfWajC7hbD7oi/LbJryXn
ffNYcBWb0jCZNkoKFD5NVemkcll5Jd1w+fQ5cpx2/sEq3Sa2jpWwqJK092nZOYXM6anml9EN/162
8koEgo4fgUR3msC1jQXKi7IiwzmzXid6yOi0q//dWlGzD5KVKARgX71Lu2h0nD0etz5EBfwjmEsx
UHRBzn8NXE1jGfeTBFif3vXFdKtwf4OVwJzcNNlJYfarkKl7DlNuHQcdNSS/sL7KHOUQrLudf/Cp
gjuCi2JqnTpfJhABzoQ0qd4DDszuwPRGsACZba4CwB5mxDwcH8U/2/5OeGm2RwMiwUBzfc1n8djd
EDD4fQOB7GSJB7VUAI4F/UogtbQlJeoulEb3cfYjmlSReh2Orf6lJe9OpQtllM0fNBnECim9/6wB
BouI1YhGEFPTBfWx4FHH9NS6aHnfH9YkMrcrHPp7oxxAzUZcM0ZTaZ5b8U4V+L9BOCzSTyvq0c6y
Q+dYM6sXnLLX04GBM1ojJFnCyRv18MMcWLkKfQ5DxF4iR3oIeahuA7gxUXTw2PreiS0k4U923F/o
kDFEjXaL3hwKTMeObn9b+HKy7PaIN94xPuI6a7Zl33++f4mV01hXjuEWSz61IaPVjhPxWyo/6WRr
hDq3+weNoHCADOIdvOiWmrVzRs8rkzaCzFO9CnXQEIPN3MEHWDIx++AdsPpu/9NxAtqsTrGrOjc5
VTkD89p+xh+acuSGcgb3WWosDfarZ779kNx1quSkRR9Ge2W+k/C3ooRSmkt6dY891gcJ1mfJ5aoA
jujqEiKXuirpsN4PBkHWdwPykG6IZanULebz91kXPgz5+gL6JUs51riYmMHu/ahFiCiCm5dnDYyr
BfYcIAG8zTVl1j3ZsV5vlY8ixXihoMyxtsXGjv0YkaDa81aHPVcskoc9DnPluO/acENy/PYabv2J
VvGjtqww0uyfh8d6mUg0ayPvNXsX8zEIHEGo2tV38A1zerzAzCFoqGlOF7frkowEnbCGs6X56wAO
45twmVvt5gFLas3/pBF6PWsdDN670JPOZ5brOa4I9uBZtr7uGKA8fM561OBCGiruh5JaPMzaZJ8R
NcgF5VLTHnVbksldwjcKc5M2FK1eAEOCcOrJDfO+EdeGYYMosxr2KV1jxz/z5/uQHALRsbC2eH1q
7/nB0uvmWxXi9KDphGI1zUpsi33CZmztx9LzeAp8Nip0o2R2F4E9+SLMUomg6NRVHkff4iVqKrsM
l9TEqVsDrNPDr0CUdtir9RXdWxi5rtCPV8wYwwPiHt5H4bE9EEbqqiIOa0sOpzDPYkvNmPKpZLtF
mMjhtYYmsqVBXtslTFi9fzjU/8bzneUYpVI6M2rYbDLe3nDJT4knZ4GicH98gL48SVf+AoAlddBt
7s8TQ5LfmvJ+IicXowBVsagUhLG2iTYqTAmVo0TLWSXS/Nq4KnpMfDQldwLziOn5vQsNLFKjw4OW
UwTLSxTJs4hBGxi9iAYUnAY1WBVcqjSogn0T0yyTKkt4S6rBE84iVhAn4lh8OvRjmTNtycngcWuF
fpUogw0mbucCUL80VpM4+9C3cfR8pOX/QtrZJdKRE2aofvimvxDtJuhaATwe/ReCeEUvxIoxPArb
I8krtqw38rskS/wBr8wqmYHvqR8IUJ0X720da8EK3+XHB69W7YIWzMvVvd7LwF5vpBPTPKop1BNd
JxKqidQBhuW3CZmbkmsD73wdVFTZbFqyMcmR9DHhiNmV+Lx84V5Dw5OVIzQozkzcXijWHhHjxdt7
xWgD01eIC7dxmcqUd0FCSbA94xQTYMGAvzWRWn4DlDaMbt7K/hyM135i4SCG4Tp2jyKaiSeSs3V2
Qif/6/ZZhe2Z3e9pY07HT6F7pvkc9DxWfZ8ixyLxvO1o+GRWlBaGeCTUk7pMONbW0EVKA+yQlH3h
9HFD34+tPXStEE+1KVloyRgnQZ7bzh90sv91PZIqXqMWIIleW2jAuttkYX4HUUHaOcmLLfhLx3qk
HGCiyKajH1Sp8SY5gwrNELkLjHS6PWqwhU8Vy8fMFr6bjKfaeNMCVuMgzVnx3eSdJHNX2LEg36ai
D09BL6nDLouL+Yv8fxcMINLPdXdVmH4n+aOSij2URC5BQaRBXINHNDwj188u8+ynQF3Cak/+YSY/
/lSI3k0a8LgU2v9KU68b8dhxDu+aY4U9NJdsW5TN042o/SPVEbcXTEPMs0mZuW+R/e1DbFfbrLg6
cCceXTVXSAfoNBHjnpgLBJxPvW47vWogzR7jgZTG850KR7Zhw1z4p75cqslJTdII/F+ejaly43ej
x7jVV7jFPq53J+LhhQ9ue3S+/VDZNKwXj3ye79gmuAujHUhUG5BHwLcN5Gtl7abjGTV4cjD0/rLZ
/36KgTKpc6tHSTotcqrq817Ec16UsS3EBCFYGGckEJR9eLp6/nBtJCrZotvW7ks+/CXSoSfEysaJ
259E27HoMOoYGMIXRel0Q2TCC6wMhMF2968kUP0tnqsyCgKSkfeA8Rl4zRjfmdO0ymrOeL439Nxp
SmFC84h9TUt2RRqBRM9sTNlioZkVMdq2+xYhNmX56/8xS2UighY42S/zJmNCdeag4Nb2VTQ0PUpP
DD+uPFzaB8p40B2NxjalwKLnKG48zOvXWzu9dT7/0qJ85tsjKkcL/H3wSFDJ0MnK/YgdQZgyaQUY
M2vK9geuhR5y2v2044MT5J7tJLp0Q6ect3KVKWA5Nee/FxAoKE3t7744WeiQtfCHgNQxxYIqRcz2
mSy5nEGHYY/Y2iHBpIDoBnfXZKz7mx2kh2gZ+7jQBfJ75xcvuIk9i2rws1Xt/etVF4dSWlQtbkJX
QQdH25kLr6an0AiiTJNa+6sodanxtNZDaDO9clsMIlf0agydkejVSzfSUbTOOmgkshxdtLnJpBdS
FE7+rFjvLP+fZrhuVRjlyow2g3+JrUWzXyNtddEh/7RcbzqI01YsDuB1nJsNLbr7Zf8JtXLQedPV
pKhroKX1spGotRKxloES7Mfil+nobtgeo0Qo5L/n5jjNJ4VBjDD1hVILhZtfok7s/Lot/MII4OVH
+Xnn2wTjyxYJkO+sPMDxuGFiT8YOBXLYCIE3k+4FIQX2CyrD+2+suIgvGhYvJKamzN1DdJsbfE/5
jaXgHgdnbUOg0ooUxaklY2kpiRcJgYC7r6TWiooGfM/Qz9Ck+0RLpXyTZNzU0qpxD6Gawodp98NE
9pv/Et+J0T4HxuwSwy1KcHoLRx5PHwFJYHaxNMze9SYRl2h9pc/ZKkFd+XPpN6LsnKpukFWKP7xS
4lpTQP+JGVGuFKgh52j4XhD9BS+ggM9o6ujcnUPUDepwzDJ1sOdiZvcsfIqUOH60tllSMH/LplTh
lM52axqNiwZFUlE/eIFBFIB9KUS8OZT+Bgbbqtx556GWtfWjXuEerEDUMqkkxHaW0W98IlMVOgZq
4VfBWQ5qPqN4q+mIEJdyLZTANwwOKXtUTsE+tWiL5+NwvgT3vocgliL7Wo/BDGEU14/Jewt+6Gv0
S2h6MFd2bz12Th93xSnT1yerJCN3DaNC6OHg6tlq8gUCwvk0SCZzvU5DgOWpT72w7G+KwxkWmuVP
r+oaWAdUsvC9e4tYTYOUYB5ij2u7GntbrhTdqXP3n1jA7FsVyK/1MPITASweTw56COdZ3mCdnVHj
ohPr5CK8c+6qm3ZBvkUtS3s3FQs+7Ug8AWij19mGJdY74J6W91InLJp7amqAliGdTKf2uuKbNRtE
4edfHg9adOmbYu1fMoIl5BxeTd0v5RA/vjbAoGXlIE7MF+YOS86E663moUWTSEgv9dT64nB3zdtk
m4Lw4TGdDIaJuCxIrGwJmwELbjRjlt/mDtiRYvgF3qPhZ+B03TdPgT8c7aDnnu9kHCCiGKBwW9cV
tdqk0QXUIKgu1QYpiN0bQBwJJ8U8EY4rJjOB5KBrJdMSaY9hQl7Zxn9NiAXmSYzqmC8gLPgWm7g3
EzLMpiU5zK4gJ9lYxMFQA6H3k5vtdfPPjeo+h9Z4zJdsEFHizhHcIfYHu9t5DWa+1lrAVRxphsFt
c8gPZ/s0Eu/Ei9Q84eyxH8Dy8zUGvXE/hDbVgFwLEEh7uefFN9Ack9R+VMBhw/UhrxlyYm9p5jR8
bLMyzirVCXtqGqX4lKptsfWwS5kdi8NX3oIrbPiRB39neYy/MWdLQT8hQdMX//nY8t2q+Iz1sdFy
SibstFuEhdkTCCcd/orCbztlgWlsb0qr7jZKI5tKV9NHuCcylbbkwhjOQopvw+caB/jmjd5maiS0
MW1kRFmNpxfV4COK28b4GMDDOugwoQaXCxOW99lsb3gbu6lCoQs8944VfNdnFUQRLu/gEmoPyT35
VR0bqxkqrfijvu2DTwGfjRO9VOiQHTVjrdQAQTlHN+zHrV9xId0yMu0Vxm5QjYn37ThVqD0fcj8y
T68M0mTCHpcsvhnGCDk6dqd0EPPcz/pKawNxP1p4fHuKJBFkMsrOyUFuG0rr+IUbs0bDSFGTkPgt
GoxYPhHVnk4AOUfoo9HJVsPvV0eESADIadZ/JQ/F4ia/SiUMS7E8y9O7IrAML2H5DMY/QJj7WY2P
SphZQ6D1ROtRgjXK/VEi3pQv4AWSdUTxZJyzy0MVCkRYgEAaV0pjaXqtfmig7AoFQKsZoxh2KrdE
Ry2jjoSsEAlgwzwmTzdqMyLtN/MhuUaJcHLAVhe7OyeNKIp1TW7bVYD1Ufu/QafpUDuPsEprTz1K
vYPlXnZyDrDflTOIJztW2Nt+w2FMh5Betx5/F3Y03bdisu1AEacFQvEtWLVd5Cg/+WZe/tGfWEXB
bJWWfUAtKMHFWkuVLy6lPcokMblXSV5tz6YfZTltmfBQC6I61dbV3qAXrcd2E1F06wa/ddxoSzwZ
GxQn4DDhC1EzmnfptrMU0ymOw7IvAw86l+4fqBSdwmIb7tx2k6SWULA/cejTpR+JDgAJUjOdTduJ
jkufrFctq8pyB3YlOImNBQI8gLX94rkYe/QcLUK8KA5GAXJtz6i5uPv0+AzllX4myEHzoDoeVe6w
zvokjMtaUzpzsyv3JrTKwLv+7XoL7xpEKfrGxcf1NVXamZNtP2gvvKw0mtDq5LScTKa9PV8887fq
E9fwj6ZzEKK0p4zgcBmKZuXzYPjR5dA+CMPVzcIpBfV7OU/mX49x2V5XIj549VSfR5U6kpsHet/h
9axQtz5+O5Gzy67LwQ8JNMQmzqaHgHEhJzDGwQpEMzf3+I/W+pedIZ/2pXPleHCPzmW+zTTDTRno
IKx3yqh6lQbJ1C9UbaG9SLbxIl9aHJ9IWafRFGC/JvGkWkN2N94+KdGry0fFfYVyv/sE7tOQqtFH
49S0NDQG3HprCRZa6mbV5Do3ogPQwIWSLd8+2TPObEHtJmI6xAYpBQ6iT/AWjMzof8zeQkW2Zesa
johUmwvNsDrmW30mirf7GbtbNxbnE4s9Es0K186+KcKu4dnUohDLObQrxvsx4v7XV+Xz6A5E/OrQ
lva/c38Ctjnrm4YujA38fcPzHb4bOpz4C/P+hs6rvNVJZp2m9nhRbmVAwKhbiPbypFBeIk/TJhv2
+XnaZsJj+zif7yC606Xw1VV5ZcGMlRiUYFXBYUke1aX1WWReqZPEq3drW3XOw0i0bUtzBpI7wevJ
A5H+i24AutlVjO4qE+iiquPQmZ8Be9oKjbfnajd+4aZJ0ppJvVCJMZmF3MGLnP0ZMtGlflJ+OGTu
WEYaRG7+GurhGnHQpcs8wIon90Kg3eX3x1kC9+YIu+jaKoDF9lJ6A2NVyKRejF8lorM0s4u+xtDX
cxw5EbpVLBr5os1fHE/yoSI64O7BH/768TwQyDqnhYaIbMVng7ECSG6FE5BeLulJMRcqZq3LWnOY
eWQPUntjYL4IVEzQ38pMtnt/WG27BgvxvtjYAr/gfWuj8HsqFS7nhFGGEMVY6SyXHG2wNu8K7A5f
TkHYWlLsYwdirRxTFD6i/RUkjC51nlc1R2aAAh1aNpguXbCDx4fUom3vmZIm33X6xtmuawqxhzOb
1zroyEElk9EGk4N+Ggihh92TciILQljvrKSYwekZH4Z3snpjbIrLN8ni+tawYCE9AwMDFYXNAtn3
Cnc77b3bTMLq2FWHJt/6auSnfpw5ya2BFHa/59eVTbAk7jrBmpJ9LyaWLSlSNuN/4lp5bWtFkpyy
9ipoj9cYLHVCaMoWPIdENKmYFOr3L7ghw3rHd/P/eNbfdVFfKETxUuOw3IKyd06kqnAbL2pKuhfn
27s1v2XPPXexTIfOF+acBhgyo3NjsDhRvBQLoynN5jpvxaU9As5eDymfyxJ1Wvnav7XKbFQGw9rd
YMStBOg+mg3zCmKJS73OBQFUAmB3+6okJP99UyW0T9XB9/5QPeg8lt1RKvP0o3hvDIhLwIZGx1dD
qpG1RGrNrXqbpvFB2p+xHITexngc5kWLHQ/0dhX4X2GJkPkmQa5H6XdTkokhVND13LaETJmZ+amh
UhylPdha5CG2qi/TXUj7stv+EQdjqYSkfj00NPsn8KKKMKHXbA2rrBssp5mpOwoZg6FxfGlpZjyv
CZFSkQFj2CVeBo1qqkVtnk5FwMImWGvC/1wFZqnVstYtemqfma55vY9FekdX3oz1/CzLYMujx1Mu
sNR47XyM90k4+c9uOUG/nux00WP/u+w4PeCRDLPUDS0DkHt8rv5hf4/tHNm2dfQB2rJu9h6eWsg9
f0jbLb1VvI5ndw3DGbC6a6ZSERYkqVkuOTwI8wMglTy0bkWupcGmbCIpWhAx18oXOpugJeEOgcXY
1vRIZl2TjUmABuP6EJk8wdNTHEVxadeJJydOBl69/g+oEAWpNdbwnhnrOluIpTpmxpsw0i2WTaTp
0bxoxsL/OsrOHdxnJ8FuotMJkh+xNnUD9SVoboNjC1lNnEYbv6GUI66gWKd8k+DngbSHgtmOklYd
SS1LgcqrdlVDKBR5zT8F9eVp2npz+yQXgx6lmh3ithyNgKmUBhdZKyF0TvM2woVm5OnXygCkm7kH
3Laf54LFLzqAnPs83zFxR9kKGwtXXT1uPGNSv/i3Y5sVKsBwmUNcQw1KkJPpTgZL2o1/eckepm4s
t7e3trCJa3CeMzhkR2CmdW+bllennskTepO7pZjTSnNmY0SC/ALySXFQt6dXKnbaoceh6f9n5a+7
jPeU2yQe4epbU2gQkVM6bSSRpbZkCet7egAsviudukktkgfzF+OKPpU6+4pqzIFcMBwbhb9ZQxp6
d4tv4qb1hSmkVFYm6rFYCLuULVgVbQYEj+Ug90r2b34WI6cBewjMZHr5syOHfEHXPiDLlJ1Xp+Wo
wobiGIVsqENjVvlXUN3MNU6hsYsg6CVWR8kEJtuoQQOp27v7VN0npKis/nuJS/o7OlauR1hmhH/L
PRmpIG9AkvIR2vbyQBkpuxmz8Ic7I+DzlzzeU+tbUj032oN9HpROEGIhpC76xOHOA7m+7nTMKnv4
V0BoTNzNUJtnvWi8gjWGlNCQji2TaWH3UAz58t3zULb1Zh7weYzvCd2zoWBbeBrrjDBaZKH6XYXn
UaMxtTrXMs78aBRXk4b+wsRKF8RATSz261jeBKXp5kKIogiuPP6B/Ew74G8j7FKjIvz8dJMMWfwp
QyE9Cl+0MOoZBXTNF1V6+TWP/s69IQnEiA9j7f/6e9DT1rxbGPkdWQE55ygaOSdIauutR34rBFF6
FLyd3TVlF3xynpb6jj7n49EZuCXfMHSXpZ3kZrIWzl4nhcuKgqw2gMY81qW4wgLLdPaYIDGSYHEA
WY+Nby3rJI2TyNctJX0o/QUwXqw8AFW3Sk5/PIO1j28hbDRghivtDiGXpwfVxYcag0Q1A3W/+HyE
o5zfDNqdGSne+htIAV1GUxIestD/ofp+sT35O8agxIeL3Y+xHJeiVrkF1pdelYbHO0aXqEG2cXpp
wA7FyRt0Q/CTvOYGa7WiW4bECAFsaGGa/rDmtAFokCIfGJMsvWwjDwpljbw0C5b4SDMPmktA7SBr
3Q6ja5HI5IPrNuBKtHDO24vJ9k2lT/JRI99F8PAPyktKhgH+PRBm4B/sU/BsfLcuWHGN6tzFXlJn
3iYhy5qMwYZOA36FKX1KifnsMjxNR7ySE+xgUFGYiQTIxHZAyTCAMNNjHVn8aqO7kzwssb0c4T/s
KiWTvgE8OlnAupcOJZtwRQr0F0VzbftdsJBTDOQDk/LBfOhc1tJlQHMmcbSGrtbklvlKD/tJoz4r
DWhfYLH0X/ezVS7VFDMiWTbS0kn8PES0ro+SzB+LogI5teT6c1HIxjwr4ZDgZZ/x46ptE3SUSPFz
XugxXLG56SL4b/Qf7hLAvWKzZ5IsRhYJF/11aBAngWLHWS22gfaslRmPdUn0L9xX+PxyawTjksq1
Wxdegl1nadwrO9uGbbxdV9CJXRskKQqbPg80zuwDL3F7bNVb9XnuSPgDR+VkdUA0fvuHus+A/jNo
LW0ommzTzeg1dz7UQZuNxoVjJsLXX1q4bO56Ahtnxo9LDC4ep0UxsJWF0Xw8FjKF1X2lR2HMAMuL
4Y/5CWc+s+rAQ9Kkr7JV0MjgnexGCgXzSZk40xvW672AEUGG+UJsXTWYsPsu5yyO1dSiyOGPO2if
rKJysX0ccpSRGBJtIZ6WB7ZI8CK2KEsXh/P5M3NFA+xU/wnV/a11FpH5mUb2yPUJW/H82KFly1re
kLtQrrnuTXOkczVFVJ38E0qtOYHNXFMJfxcPVUWRZQ+d+Rx4fuykug/LeOHJDXZyKTTewgq4r0nT
a0YGVwzZ/u66Rl4hcODp6OtvsYs+Iv80DyJQjKA64lavpvgiyjNm9tk0dKcYtjCkr8STCR6eHniC
4AQgFueiTvi8oR3KhA2ZGNPO4klhFTkbV+Ev9QTNZ30b+vRuymX9uEwNM071VFUvpaChpcv7PnRw
t5apgMbYz78NlFu8MJw4zUOnCFixDb4kNVKR0hxZUwRYe1GF11HhGX/26reeZD/qCRjJVqRCoibQ
a40owdzSmwqyP84yTeo88F1W4IVNbMYcYKTUXwAHHp+gPP5GWcx8uq5iuYmU41fLcqN9LFatTcw6
oBxHbvUQoa/qrZyRHmzOTCB6VxClzDRSzPF+XlY0x3+6y4pepciLvozjI9MnRaDnW3xROCuk4KRz
22wQSjzg9EN+ZDzzSRR0i3ZVxgu3f3VFAQ54a91o8X4+wpE8jbQ9PS3Se0QqV1IqlWa5X9SZAkmR
vUTA+20AiRsnmqm18uLDlesoFPAfli9q6/vhpC+LeyK30yv1ruJL00KX8MGS/wnvIAFqjfNGDbfL
Rl+Z6+NV2yZEJWSli0cfbnS1QohFyrIWBusXxC/Z1spVQC0Gwy+B3Lhgb1E89D76MjHh2mLBy10o
sll9IVLmm05CPsXlurrec04I3K0b0KLGd0W8BwfRhjIn0KyEV2E6UW2ldh1NCK25qWTmiuqvk8U7
g6yei33JE002qRrF+39UAeSXt4WzOnSOXm9rtHQ/TOKKxwWVDEgu3wEjzp8JV+SqnLM5M16dKKqT
F8JuGK4paKNnewdbJFBpBX04HzA8Mdty8Alhe/2M3YkFQECjMyaGvcf+ecv2B+Y4+Nypjcb8e091
MinbddEQ9cV5+AoXOpZtUY9SxqiaRqikBy9SEfc+/ED7ie2MuqHPor8cO1xaJo+8Ajlkf7th7Tes
BbeHpuKQbg/n1kckU8PUxpM4ccqFRYfJfx6B/llEycdEtqb5lMj4BsVJovVElOtR/vka/ZYwNVuY
a+X0Y/jl5bMTRw4GpUCCc6sYmd08Spw0hDYq49u2P4MYCKeewsXFzfYFiqEF4/OW976ApEQYRCAu
OhJYlXmD84hiKJ4k6+32LM60KZmIuM/tQW34M9SY8sehkmtCfVBClfyYQgfCRgn5MXn5wTk9BdLG
7YFxc/D5i24tsN6HAieTgDGDOAo4aSj7h7S+LYb3RZ+lonebJTmiRnz9xZP+zYu0z0ECDd9UA2fr
jowxxUvTOzBiL3bFmnGGaWWGlL+coPham5x5v2t536LaZIi8vHR9YkZjRaCLFQPnLzN+AOEpYhY7
eJTCXbEXMDi5Pqhtsq1y2lGKKAVTr1/IDmQjfsNA2eCItU5oDFVCeobm6onCg1tkDBupck86aSBo
+sUISa6RSVskpXc/0VvqSl0h4eac9gYkdyBkxmskrxM4nBfcfdywh9XBj6KH1LP7sPnba5Xo7oOk
APu/e+KutLpCdQtah0jTWiqJ+3O4Nq51QPifgU0B5rA85Yk5qT9s8ACGBDCMdEBR9FW0x2pNAL6A
YQ9WNV4INXQ35NyL8MSdjAYT6X0iufjwsqFGo4supm6Vo1rw7ECFKsplxVOmCp3gSci7b1tMQqC5
7KqwB6Vbkvn/aCBmIOjHi5w6Kzacsi+r2Do2ZnEQ4SysAfvpEXlY+qarP5R/6BGqTXHubJbGctOW
7+/YuLgbQVEX1PbEQ1uDlnGfRxNHO+M8lmA1lOH83b/hAyyfIDiCWTJDh5YRE533Ap13/TtX0Ud9
ECmHTP6waHk/cRTDH/D6Y7y6iFG8niw3XfYXWRXuQh2UfoegmLo/6XPxJpYqVgYydKN5DeoaWyUa
Vf/Hkk7t6/kLbJcz/Wrle8EcUh+79t0sFdO7GGwf2Z4J3DLyrXf8QKcQ5341FZ0oYHlwwJM9EGAW
szuhGsllfOITSVRTJpGZ4pkPQBC8+eYlnY24x6Q4Kfsj1T+CBc1FQhnI+ZkDmid8dbObmJYjHZuY
dRn4wr9saK1z94TMRiq69S2yynT6pli0CJTXw6iVXdK1UxpdjhS9iUiNjNZQxxqf3WcgSQcxv//H
cgr2PxolHiOVz0gVzBbqKsQO2VZyU6nfez/SpdvlwfeAsKPNai0iSH2yVo3TjAU35BodTlrA7sMg
CJe6jJvBBAJ5qE1gFPAtEcqzu+WzseeVjLPQcBktP2JeqZm2/sU1skDUlvW/2qjP+XUdVjIsEEV/
BeAQ4l+LKjuBuS9TQAdcj45eHHpSCC84RtFjJ1H+vsAtfGdgqESmpCCj9iKOLNT/8z7gQR0xaG4y
bsxfigQVYiZfuR3YUxMpZKDm7GsW9EZvY3pZH6Fgwsf8TgzqjE+wZ1ksQg8kUaZXnB+dMx1E3Ba6
nPEr/SfdI8hr1Z9fFWubihhpBFOTOSyEtAgNlLpuTwHPsYbqV2fstOHEqJGvo6jltO4Me4PHP8gq
QgSNvXHV5Ng+UrZX/6IE3YEDnLi7oTJylmoQduH+sR4PDRx/cAqBOjUHAZZvtjhdKVgTGUA5O8bU
VO0to0fKegyFrsydczfGsoJTzgA59FzfswP7knt+slWbHeUxwqs8KsI4/GwMIOHGHssQ52WxOJFy
7JAlaMTdC66WjSuoPJg0BknhyORPHaP1TkN7zNpB3J1w1NEpNAcMgRR6nk7S0IHv8INNLXK/s4Rl
0uIsBXfCP71HS9mTS5tOsyWMLeSfHAQNiAMsuH/vrOEksMjYkSIpAsJHmAG6Dso83ZtUEJn/aWTu
/g+AS0YrlxM3iA2VV6cK1iVesclvRM0UcaKcDn2sUtytcYtT3gxpzRVaWw8/ox8TI0LnjGpU9dHB
R9Bws4lrwgbmhsKEvg6/YNi1hfKF9QR2Ha57jzTvd7VoosVnyDzXETnFGCCqmRJIugf8ihrgla/x
s4lJLrB+2okG6TIG4FvPyJHQi02u/CiBGhXx+X6EY6H5j1/hNMIevSHgOtL+d5f76157ZNNekMNH
Ji/jiKFFa9h9jVk7n9kSedsTewQPzV44vqrKFcfxJWdbOkfgzBbvQO/i9swPW+Bhqyg6kwm2PjG5
YYOGvxSxZo+WK2eYLt1po77reSo0gO0/ejLKTFvQdyfvDVcaYWvvE1ZzmimJH5FuMqDwTIgvmbon
qhLIEGt7iVWvTcqcr0X8MeY3ZkarSAL40r7mniIbQ/2pWy7y+QYba+knhmfdWogVd/YaWNcCazmD
2SObwIlh72KpNca8sjhExzTngxy0ELCH+9s2CnlpBNPzGvteOiRryLIePZC+/EmZ/leT7W58IDIl
dQMNewp/2cEvPGi8hKJqTK/ZqrYb7FllmtEI8oOPeLBiCr3yJ3mACbQL3fDEVoTi45tWNEl8P1Rh
sWNcRwZZfY4LvLdUwQnOOy9IzlUj55iV9jjZd3FazrL4N7SFAGRp6EYhCsbWdC6lVGdpZsB1rgwL
WXm69O/rU7K+DpEfVKqUmPMT9tJkT/UL1L7Fq3/ckMIQzJ3ZZ253fhxgBFOPddZmo8mX9yCYND2b
PlA0CMvoS9RslcBGXrV1b8cTpAotrvy/OW3jbb4umtxx8z5QBjWbRoPkMLC5jw6eK4bMYmnCEcaa
uWw2G4MRuz1+tVWUf3nJMJgeMK4LWCW6R9nN8VsdLAotVdRrnfG5ZjC3xCuAALI8FI0D+/rsBfFe
RUXELgl157ZgWjCrUPuusemgGSECw1PFum35flggenUaRsP7eQb11fuuiGlKmhrLADWvqbemUcgy
XfezucCJzsIHqEuzLX0gsWr+WwA9nDVRVtA3RzQi3o8WAUYQjemCf8pbyzF4hkTKbKpG/5p7Z5zf
42TvkgaKvNZEoizYHUQV5a6oVYprwfkYmja2tX+x/emmsAkIszoAeXggAn80tmhMwGnMqkDetdWz
TYZxz6I3EX4T3mfG9R1lNfCCAWKBFHA9g5MALjaN+8VXJMfErF6z7YTBH9VSOsaqXhaac/blm2Hy
/uDJTqm03xvCFiNJPXpUUe9rF220+VDiax6Hs4+FclPr6da5C3/WTfGkhrvK8FOlczUkSxwUeZvz
dbayBPwyJjCwIGmLhqrwbxNlyoxA7oMS0PFB38X2KPXtuyquD13KspuiKrYEitCCbKgkA1QAwXoJ
CQo2AwsQJbaRt5/0/xWj4z10s3J3LTMT4mOboCDZCCSFG/lK0H0Mv/sZ+hz595VrpIVb/KqC1bvC
e4k9X2Jwa03yLUEx7t6gm+nJhJexUzDRFn+Wkqqh1t0sowLY90UNRwwH8T6DpVJROXnP5CIJWyB5
UInJRJcrz4x7t/X2xAV0tCuyfMVn+c89h21BLLsKXBxKM1l4Iq5mePmi+U2yi9cljyZ+twBwLGNt
B5ritfWYWFCzectSzL8xV0bmlaiy63NZAeVSlVEXnDBLlRtxvc0GaPrS7qf5KgNhNpWdf5QQ60CU
ZEH+Y7TeOdVi/Ix+a+3C6zOmGyaVPGpU3JIlSS1MLqmh9wjCu+6ohbmkIBuFxhkk0SO8WkK7K1qL
LNie70DiBeLaBp01oD6RBRd3hbCw48rdRyl7Pd6b69s4hgF5aZQ96o6pq2SfV1R8iILq6MhjreX+
0/R/qPc+zFO8JDk0Xs66G424VS8+5w+dhelAZAkr3GpnxwTkHX3Y7F0PotS8tHPf6aUuZWW7TfcD
khCcmjY5ZFGwgDF/ESMf1X978ObfC7CHnm6yHJGM6LwV1M7vaZobGPgdSKYYTBdQxa4sKOB4MkTw
FMTt/F6mUycXgWHxsxPjIORyRM7uHEvlwDtVHovBEQf4TI6oR6RkR1XKNbwjN9/gWwc41pXb35ty
Ea64gD4B4A4tn6hSUx9arD4bpzlXfvxVDMwsDRibzdqe7UqCUouKtLxK3TubUWKHwfNJ5+opSuav
i+FHaT4XeGCVvjYK0TYe51qeU5ugX0NxhnfRBkxrDLU0p8oTdj1k+ji2GBbQOVIzo7h/hE5LgcIf
ijsW4HqwG58gdjZTPeDcEcCKFFzN2HvCfaEXKTeSnogdhHycKGaumt+hJw7I9EVzX6Nbfzql94Jz
SLiIUhoZfGG8cxQZmKH4KrdLy7t5395nUjpvsGheevabMowxBjcaK2/UbIEJTFoRwo7ci7j0xKKG
LmEhK3FdSBNwNSq5jjyU7ksOXkcyYbsB7AVgbbGLkdS/vdALIPldmqweCbTAu1dw9HZnek+YQYMW
QsRKzbcJyX7tSwgdGvzxJVmQRaEpXdueDjEHskUCl7v4CJ+NAq+E+xq9KhfLemfm9SJcEfTjyuqT
TtUvIL4+j+pHCA/CBDmqNn8qul6Nb4ffetec55gwGF1hPdPXHjId3x97NMh5bQzGSqYU+HOtBqjA
OewpoASgAkrOfYlUFmZhLay2nIQTTY/BlKw2uPpiyKHlY9UpbrzUMEiMFg1MIdkoiZ6yeIlwMSVv
ed7oQGLa5a4+S0wqEHKSU6LO9NLVxNMCFxfusXmayYF1TqYl42PDQcuBa3ZYHf/no7fpk0Bl/Omi
ikJpFGqFyOmdodf0pkjZGuZZGtMpye0sC0nWde1VwRXAw8WwmJPN0BToltU8Nzr3UOpSYYp4ywSR
5Ek+bMNAlFnS0AQBGGxFJPCOFSrzKL3VI7DEkrPqXWl/LHAsgFrsRnlfQXx2Qhcdt2ZjGrqHgfnq
CQTRrd4FMnCp8ESmsgqMf8iiGpfKNAoJ3SSOU6kGczvq8WsPSHxpRuRZUZx2tedY5V023lUbJadb
QDPhtaGZJehVyYWdOMBtslN+OW2N7IKApz30KIXH/LMZ0oaVQvfI1IGz4gr2JuG04N4F0mC1P1pl
Ayk0jr6rSq4gi0/WwahcO9vnvSYew3XsTtVS+l1/FMfPPwo9yWkr9Gs25zI0UNw/izSwOklPDeq8
jS7MVFB53fd3/dBH6jWd5BniRpUt/XSkZ8zMXzDVoYE8kY/nrXEE6hp/usrJ/GCq+YEY9z/LXciy
NDEBZKvN+4quxysNlEMJPl5Wcq0kFYPPz4KoKrZvNzLTwzFtl0AiLX/yOHkazmfK5ivrVmGgT+Ll
g/nZary/ZWyCKy86/VMwEJv+6x7zW0U3Oq4iJtmm6Hc4kQADpVN1BhvhsfyIQK9Mt65s+/Ty7fm7
TRhDmMOkVkm5UUR7QYKzL1Jz2PGIPL686ds0/h8nnZB7jXQIytocbuMRwca5A9OqJpbS5jbRGlx2
y25DHfy/OG3AxHsO6n+EXvoBUvgN2w8uY/UTOV7lLmBTtAXnyyn9Ji4hPCMGGEdp5dsI56o8SXCi
qoLCr1iK+CCE/piACgOKWT1lGnBc1GvcYBMeWCAsSUP5XoYgii/h3+dqVT1lZkt4kIyjvB9R5sCB
QWNroZy8w9tCynVVNMbsNE7Ga/Blm3Z+obQDFhanjIrJ642py6vDYeuFFB6iSMAa5lZAxttQtb1T
1cdSn8tfhtlVIYWIasfJXtpkfXnlQhRAOE1orX6RoMDQCdPlrBxji0e2bkx/Z326ShsOzI1nIYm0
QzXL1e/ReF9vvxbwqmZ3C0XjJ3VAkUgBScU6GF/I/UZ5Qu8WlU9mx56nS44p55Aif+DUcgTf1Ktp
2XxP8W7BTNgTi9EgV/ZSd9GTZXDXd9LsbgAm8dmOnc6PkihvLJmyCdSHlpolIcRuY0rkfSeGWSPR
efA2QgfPeGju3EyKfDeqQRNDUpXqCR5ey0MzFNfxcHygevqM+vx5Y1Tjj1V9Rl1OvUWl6WdLVLEj
XTQ6cAdKoQzNFvKUsZLLcXJdFjfbRuex7+gIefNSsl8OSeuiHFBcCEOMLMTzycklimd91kXsYFmm
c6fpVg/G0pGB9B7stPYuhTXNJuRTPjmcMJbjXukx8cPdBr0KseqSCz0iZCta75bL+5OZ9lWul5Xg
zoLOVxVrxZ0hknWcX1Bz0Izx8yDPXqcVATTawsXO/D7UfoMeKWEdIUa41l10e+cFXNV68guVW6U4
kxuPO6jtk2PvGQ1+Xu+t8naOIgfJdDlOiKiPzUtZxGr5R/dvd2pH+bqJRgTs9rLC2quV8rxQ7W1M
qRrtgD4kW39BofLvqj4tXPg59vKZjHfaVpHc/1ouhoR9V0opxIeFh0HNq92pMrqujiTD0IpaotBY
2KF0/NCOydpuoYzPxAHri4xbVqF1xzYZogKmuHS1BhedWoyRUMyJmmUU7ih6gusU+64oyn/hZ/XD
vyvctB3Rq2a82VkcBF/Zo877oaAjWuKD5TvWNL/J/9LOmnsShXIUMHPT1BL7mW0GgvDWImMr6bLa
FDzjvtQju29kLF/oYrpn/CrvDKoCNFOSKxltIvK6Nobs0kiMyo3cQ/jY5aZrexZwjqwgG3DM/oLc
Kp+7EdUHAdhOWEA2WdRTvGuYWNkSl0snQN1uJ91qqrJoZ1NgbpqL8LKxLpeZSa5HGIddUaNfcNLB
NcBFMem1/gzKN6rpLGWiJf0aLX3lRMipqJ9DqsIDW/A0/x4Iiy4aTlo7cHFattVZz4JHatTu+5jG
i3KrypuzNKOqAc4UFT8VpkfMHSKvsVyXYzm9PiFU18wqXOJK8woJDkpO38Qhek9hDNsbXUvBB+Gr
nz/OxHLixuk36Fd81DEcJ7sRKk9y1ohYvCkDb/V6F8BTfrGBbRNbiFm67cv8JpqdnibmXzCt2jyq
6/4Zvqh9YdYx6k9Oh5XsyUYtG1UpJzMHui2JGNKdtXQSN57Tti5LV9lx7G3g/OGzR3ZZSs7bi51P
3MSoI8a/tgOuHCY9YfuF0UD0bqccu2ZzNQwQF82Q+U9p/vA6fzQeg5bcGFUXiXiMzPzhZgvLHzBa
KcD636eN7IkLNoPLAEIdykwMCCC6n1W9BDmSGAKtrUYwl8BI8dkMzBQ3Toq5ZDngQzteZqel5bSt
JLNTsfG41HOmENuQWcfL6VmcLqXJk0QWoRZWM5Hc/A9IUckjdWJOFxuVRR/dzmATofFteXtctBt6
54ZwriBeL8DLUTPn881jlB6AaUgZAugcD2xZ4vwiOW/ea6vq5d02gCz2NLU7s1BzRhUzdIdFLG9W
P4DOAqjqNlBZzdiNuYEC1A241L03/ZUhSWjo2YHIJw5OHIOX4wx7JsULpHh+jo/mIeQ0GcmVpYz6
jmt8NceC34sxwTXpMn+IyBYfQMsnPyJgfaqu5PKUkRlCtGDdus9Dgb16/F3FaP9CPX1Qowp1njZg
P9JRYVoagEZI8Gq2QZyvtoNaia59irM130c7xOfckpZkp3GNdHyT9zCHmFf2qAZ3h8/cQbdq5Ry3
ltR30mjUwr5oHFA6ICf8vohD5HZBFYGKubyWSPDdG1U+mbF2hLxF0w1/swnSJGfxZ2baev2QETLM
NJ8UX+JgnOgr1NqHq8RdCQYIhZi39k+Kb+yhuXYVm6EFUG7qcUqczOajcF8FzyXwv7gyuxCbIj7F
9wYaJpxjoBtOJDG2eVI3vVjRongWkyV+t4beK3u97VRmhLbLq1HPEWYOuzy7vytk74dfuUtAcy+v
Ald0TK0/LxiipkAXqRDkT71i6qD405LnVgFFEsyWHdsFxiNrgnPVj0Xto6W14PViVdKCLdjhWCd8
HPdCuO50kUAEPAoRRLYhkqFhZ8wRdj97KhOytF2IuSMAoLT2CDAQvr7hHNYur6ZAqb6I/5ddV92e
3KUitAkvdzZzy5Yl2tkjHavvHoeguDgmUgDUImoZ9ypi8ODKC38Lko4tCM59AZ/8Z/ibiU3sBdVf
mzJtLBmQAvVIy6J4fu+9R2xnVvKUxA8d3CUe9jwS+awGgbmxAstMrO821ijZThPqRow0Aj4FMOmO
CbBzqOsk0vXCNO2/3b8qYNcQ9J+sE/EShk1eTTyBFlIVmXE6qiwc+GHSz3BTBQqRI9rrwZrEkKfd
HOxd34jC/ZZRI/Pa23KDE3iTCG5krQL8mest5ds9jIR6FzQ2/GbKn88za5TNqTIzcplCyFWMp7Ph
JLVq4OfMb+LtYJrEi0tI9FhceQXzi1JnppJ1U5D6LqWzdvD+W1ZgJZGQF1/IbTsw0ZE9909KXRyT
61ivWFtbwwfwbHEmh47ViDvnyoHRidfj62DURRiNfKfHxY8VfDWlfnQlvwiuHpW2ecLDkvFOgGAD
OURoGM6JOsMM2GOtoJT3X5xakUJqlD8Sfrrii+4rVrNJaK8PmaA1IzGAKD5kdCcOIS4ePDC/S/jD
zPcbadTwkw8ajjIOOMVREbx3hTo5ust2au6aDHJa1xPRVXYQacOOEvk7FeyKxP19bsBISPAKeb3Z
5Do+1f4/3Uu/FWoG+mlhjxOtwHLzBffUK2+T3wOHaEBXb/Qgie4W4GnYXv3UmNOJbziSk+ram1Bh
T61vx9nLGmE70hkW7peCmd+6RihnFyEtN/n5S2mUQQUwngYb/cZeZPX90Wef2J4teIPPp5Z1DGb+
ea60oKKpr4Mmd0aYiTBOuqEMEjt8sBpq0irU4Cy9soP9M6aNY5Cb2Dqs3IKw8dRLrj1CG5R8F85U
dGQBWJ/B02+fdaxRxuzDSs5E/0ov4Vu+Mj0X9faDhHo4kAmB7Deg1ZxvaX83e1jZoRtx3T+hkplq
TWMWaewvUqefVZ/Xf1crTE/6JBzcS9UlRO90VTzX4J+kFq5PafcdOfYs6iY6kp2SNNYRImZ3HN9F
Ldp9bPEcZUcUjkV9UhKv1IrB+1xE+O4Dkw9ecmSjKcIJDYu4R4TrJDE6pptNla6ewfso3eKhWW3+
fIijnbrdASz8ghWGXtd9DxwdsNt1MkuTt/D7fpzne8MIcR+Qq0mlDaTGBfr4BpGCoMADxd4Ksfvt
HR1nu7FXE2TZaoDKVr8YqAgla05TNEqe78HrvCT7V8jxihpSFhLsMIZM7xZrY+I+hS/qJaxnCTP2
A8XxkOOMv7jcyndNDGxrWacTEcG4gNbhN28qW5UdvvK7SWA3IOtdjcCDcuHnEPnuUvCKy/dyHTKK
EiAHwbucKVCy5kjnhWZcUjs5kLsPZhbsLGwTqwSCE7u9FO5HwrEpw+SGV6xw7a7BU9z3fjTpbBx5
lq/UDWRZZnxu7XuaD/IyI4kA7hxgFQgoA3pCUIPym9KbT6tYm/tnYsEjoLWDHncBMjdwmYUqgKr+
OvjmyZkzMBjo2ADiCSuUkMiOnFgXCz8k3BmvRfkNiYAXaoagzetkAnhsxX5xAora/3cDZ+94ks+0
B5fiqCpL51AmaVn0ou8/2hWYKE1nW0RtjosgoUliLokiIiiu63nUpomLzTbb7wTvyPQy+kKMGGAh
uU7Wy5cL3FpzlqBDa2rpkt/oUw4wrAZ+QFCBCPCveUPy1KMB7UJuEG+kEhDIh+N97+KHUO+4g57z
gV+5nsGY5ioVK0oxbFXS7jrIb3+pNH6XYiYhHiifM1xJyeL4lJkZ1m8wMvOCMBOcfO73hlHViaXC
kskSCqnQVobhBnhjB+qhQ8S3cBPhOYrIk4Mc0nVfzlG2AiH/BfFhwuNGvcM9QexJ9NB8MhUCTwjc
wVOc24zC9uWzR4InEi/lOL6a8RHbdKvkWZ6Cylln8HQNMyUOHVE+NsJQ6vaGltHhCFXohswv548I
zgHNCtO1B9NzHXtqaN+iFvWBJnPF9YVWPM03hRUcsaUNWwG/+RSH7WP3aCMDt9ZeiMnnFYMt6D9W
REClfG6WqiQzn2fwD/cNZ7Ycjcx2iRklYhRp0CuMIE1Tg0S72/8wdwwS/BflaKLYtdzvlbXnjTuF
WOJ45F9rwL8rpmkfCEt2+iNQRVtY+s3as49U/jZeVq7/UYWoWEar+/jva7Ec+3xZZZMPrespyiuJ
RiwtvNqR3j5dOd5IJ4qEPKJ0WovnGUHlsRJJphziZT+tFMH0sMD3e11RkFpNqvpqg/x6Ha4rZvDV
75DaS1nXY9KArocA34/j8EVZht7ldLhX9rB0YLMA9YS1VyLxGuWSkWiUk7CU1fCnv53dvKirme43
WJsiWcf4Yrh5pOWDhNiVTBYZppR8pVcUNuRM/DABNsfv7X9+391D7pSj5Y/SvTbTeDnL+Jfn6DhD
akmmY4TMSes61w+SAd9Wsfd3YQewvCUDblgnBL+d/8SA0VUgVEWDD4HTxJPyxGRG0v6DHMvhZ4w3
vuTCszRRfeJUlJMoMC9jB6+TejvWiJpBJOu7zyPwLDsFMn65Tl8VmP3l2l6QZs8N2tubozM6GLHS
5pFLJYsmZAgjHC8goVx7PcpMjxH5ApUkYohmLLvmSfzoUOBsR38uRvc6OKKoOpeKVDH25So6CNN6
e/XY0ujkUyE/p/5abUwd1iRszPh5O8jW612PpkYKte8CqDYPQG573l0t+yMplJkxXTus9su2Y9vX
rvg7PG3d/wFYJWeeQxWpIP1VBgyekhAFKeXZLUz+Tsulaz9+x9ZpkUjP8capRbG+Z6/UeHjbNKV7
NMQTEQnxieSLe0v7YrpXDchCwytMbXXEW/benMRyDv2H/7QzNq3UAkFO6gGyvC6NpHuTxG07SBGR
GUUfeVvLDlufz0Xex9puSDpEVsxYYmY63QDypnUsVAU6+h0ZwYVuURTHDkuBidLRSqd2bIL1SI47
VaTldOdv1mDEjI7evXkGVojmnq9rr0cPy+OW4X75unu9UL6lwJvlglnAf5aZIZ3TsbacfJMx76Ja
7TA5XHnuOsK4KrxIyW7O8qtwLV5Yhll/xU06h1kC+UBqzY3lJs9LjfQn+QBV7JF/ARmctcJTR7yo
aIuLuk2cn+RgTmjpX2Wy8VJ1IbzTxPTNs1AeqlwX9aX2P6dB/ny/95KSs6iTeOZpDFHdlsBTW6wh
lCEoQR5nRgoljNpvVDo45yYW5EgV+8dCUebh3T66RM0PXA34JrvYzuOT6ECChXSekazlYCbcEqxo
FwxjNIc9rpPriguqW1kr6QidrNAg8yiRQY4TaqqDm0SiifLnln+pk4i5exQNwuM5EnhQ233EuIip
M35JXJEGX84L0RFKzpHG8S4L3Q7vzrmWz5NqCpI5Dtnid9MzqWZ1JDALGQA6eEmhJGa7iPTNtFvc
xxx+bQm0AMQYIVJMCoU8zKCV7fmmLjmv/Hv9Xz8DM/JCXZr2DC3TMDNS+n0NrkCUrduSPJDRuvkA
3kGeY8n+jdgsdNOj410KFfS+A88m2OUVYNzHxzzoQfSU9h7BZdXiHTDkDJLEQD0NUbEQVd/zvS8Y
LkrR6/094tEdNGY1HF3gDBCn8u13swAEAFYGCYG8dCHMjGtlX+SAPdxdPV4Em90AP2tb1OQTUI2d
2pu0GiDIMHhuNp0IRvE5N5Wt3I/br/hdtsy0xoGiIotKz8FURE61gtNe31WJw4fHR/lqHH9uQQQO
WtaBV9cnxTeLNBVsnrh/jJyXFCYyE9QStFxhHDnArQlWeiXAqntktW+okKi5Fq1i2JaqeQ0bz5J3
o/RIcbBDSn+xso6I/QiW2RX10Y0RehqGpedSx1mzr2/j1gZS3bNqPHrOXpjqi4Y7/XxCi1H119hT
U9sB6pjb7vYqrbncy75+rTwJjFK8qms3mSUBkxRUADSLIQ5/kjMm5R5ne/PW625mcgLiVImQjEa7
bF8S0iAywOwgwO5KN7HIuG1lMvtOloN58Vl2l2+BAhadbNxU2V28RpSrNw0roiCtknq4pIUk+ql8
8j3WoJyjVXTlBSvSc/pFNcjaqJrPmbtYpxmytD8G+2//pIhT4rURl2raCH6n19JmsWSaxZl6Yv43
yESnIoAAItWrD6GiCSZ0RGMGPQJfmduTrh11wuHhjctOpNqWzaHQS8BA6zTh9jVS0Pyp5oW13aTs
J8BGVajT+lBjtktcZ36wVOYVADjorZwtXLdFEEm82kNZL+wvX3vdGZ1OHHkziw6b/tzpS/foodau
9wjnNFqlTPHL3vSpsRtAFbSO1IFp65mWDsy2ZfN3k+j13pdmg+NZfXloTcF7eeFugnSgpmb23WL2
uL/MEQp0mp6ooaOMxq6hdnp89YzjIo0NXQU6eCxG0BOdGUpEwklLg9YTCNfygVHkNu3iLzbF/0jq
Ca1Y+nemNcHztCbtbddRoTThePeVRTFGftXfbOPcMhd++xOBr+aKKtrAqXdyRfs76c0v1w0kjeFV
qfoOip4kAkw6qXmW9fE63LyQTED5bD3oE1B+YA6Rblf3qRmeQ+foYrCfizrM0Ri+PU+e0vXCF8+F
GC1y7BQyLdQqskpSdvJQGBop2olma+lbLYOLYOTD4VPkREY5qlbhl2o03njyQ63eGVedUtiiu9Ml
1fI0iD5tBcKCK3WNo6rH8/6Q0UnVsmKE1HbpoXssuZaUGckcaBdpZv7SxIZIGBameNawSxoaOt5X
MPWztxi0tiQ1O1YpG9ayxJakAYEbjGFt4Cow5zNhDRficDTkluWigbXU0Nj+7or8hZUw8CEtHkKj
Ay60Ts9qXE6mk8fRuyTwITzf2/s/YhYHENt6rzjbL/xVaF/At5AE3Y2Jt0AtFhgJJwFncNJbaLhX
ePEArUa3Oz1hZ3GwgQKQeveAHrTmMCnuEHc5lt/Q+nsC7r38sNG7k8Eg0YFPqCRVgKFaOvv0LE6i
DSypAy/GjeoXBG24TejUzmmGNiJawQSYnyty8FqnJubkr8MNH9yXB/MoUHGZfn/t6J5AKx6S4AMJ
/gTEqwe/jiXH/GI/ZirBam3UmXEMMwvEnmmRtIc8wOfPrElR6dZUMz1rafQGq5BKf7vDo4uFUorq
TjY3aXKI7adyV2c8rgxa8sH99UG2o7F7uQj2HNe0upfxUJw7PjnhXbJz8t+p8IIWDr0WBQvGD+NJ
yQpu7Ipc8jc8hH7JkbJk3MCDVsz0XUxpbjxYanM2PQUWbR9fPSzlTRHMnAbCEfhZMl+cx2D88MDV
/vUSIJRO2Q5JXCo/vMPbhGa6XqVahFBDSB9OeXRSccW1ZFusvVsLCISnkbRbUJkdPlEH0h+5FOq3
R0zx+UcRIljZbN1uRKW9wOex5yjVh4CW/0RJJzSaY8/+6NN/cSIzDTw+gaFUv4/I2oIneW4/d4QQ
d5CaTH2Ed7pGN0rZlD2nrP8NRk7FKtqWuMsoIIIgi7KiYKnpj/fRhiZ2PwEFHXaCf1525o6joebQ
acYXZu+lPGVNQsEVIUZLPhz7K7diymouoiULUkLL8Euiymy+8r92hV8MsKBcuEBgZYVseXt3Bnoy
Bzr/vUyGrhjOxW8neN8hb8dQ7hMntESK+epk3crnIiUkP5M9MSfIrUpzf+ZeUzzYk+22q2L+igV8
b28YLcJrAre+5ZDSnFb1tv0gC7703Fru03MS6gSSZe87Gbc4WS9lJvsb5LSlU+T9x5MqeAptHzxf
4HhHdvgFhe0CzDa3y6jLW1VB9ihcPA/Y68YvgULwfkqwdAKgp/pPeRh9WihNzjn7gX41M0N4kUE3
tqy3BXQ0ZlM/HvDS77Gomo+MVS70IG88kpKqrNg7FzG/nY9KWsJJooA4RPjS6o377KHTPgC7noZl
VDVd9pXBnx9MrTbuVPuTxNo6E4AOSAxxErtI4Of3/YWnv5eKikh6hWkfoiJ9cAKJ6SN7nwamv7iI
RK8LaCEiYfIFifoICkPTbZpW44tDK3LRfg0zNcFeTSAGeVVp/hEpVRwJBI+wojZz5pm2cImsah3E
J1wptcPTNSK5QD4wdrkdrfymNiol9uxS0bSzIyleBFoDb76s1wJ/M/3AvEr9fRSndpbaSNgmiuLJ
kaSlSJxZ8RibMeLslnhpN8Y2SrMxsG10Bb6V+Pnk82ho2Vlt5sz94uSlVu7l8KxMjyQASxlQCSRx
45GXOdNglW7RC7CFIZq9KkCPVNrp32WW9MGfp20fCqvNIByb2vBscNw62JSpwRl9CCp/V1ga8TfJ
KM5g2KPgrWentj+eNVU57EvpHLdTnl62zlQ1ZgP8y9NqSj06THFs7vRZaeYlbScXZya+oPlM2OKK
ANKT+jlJLuAb6QVK9fLGsXCqbJ+HdyE3d2m5FLPKQBBytBa53vKGpVf5twSLD8t4YmksCMvmyRUN
uVCFaMopXDQzrcwoyeeDyhcqRqwYzE0z1xcc9jhnZsD0iUAGgyRJiWYYXelNawvPG/kLXWlRH38v
nxSv370CffIAjyaiNrzDkY5ajC3wy9LC+PL7DPAJnRxHcjZEtfrmT4Hq9v2fyGbD+wSxPOQGd7nw
166Q5B6cqH/uLrEy6Jfve5/mxkHau1b7X9M1BMh6gHNagBhY85QvoEKSkhxpmF5LgbZoKtYWnZul
iPl89IugyeahcW0ehqt746ErFGGzzfmI5x5Npfegz53+NRhfGFPK+dCZCqop89J1A/hnIyMDarjG
JLHKQ6xvvnK6p+amqz2s7riwUQBVrYkVJtqOAughEI/zZRJIFNQevN8SDTtl/AGDLGp9I5Zldkre
SLiFbesjZylY8AXjrS6B+nsOy3QYhvbI+we5GMlEeBBqfAM/Z4p8IZ0ALPaNBC7fejO8/lxbKDHS
bLLWZnYdbZCRk6lavjZWX+OQeCEN//BgFnrbIxeqphcVRDzGVFxqMl4ccfwfx4Y5+ksx/LwIvZgt
GheanzBkF6mccBdKVXroXbtnwDya5MgIwzaON6OvjRMQQrEo8h+AWLStdJRjgCleXycVpWLbcypf
XwCCT49MZ8J2EhKvL/2ZpGZelHgR7x7WgePxbMhJq4vhuiHip++LACgkb6y/XRN1+rKC39lcGPyw
qBf35I9cqTagMDSLALAD/x8mrI+Dm3CDg24Vqhua9nCRWvpDeyzC9xQwFHrUJT+AXMZRe8W3utlk
cpu8I8ENH/sC1ZfTLfZfZDvEqNmIzD0rsTs04fR8waZPH0bYrfPeo2bquYzTFUyaLC+U0NgzMPFy
MiPJoCH/miusyvuvQPjcK5hBYAupPdHb2doE+7c0umfedqky2EPtz/RmluFvKcD6I/ZH/wpsrqRP
KfyjHEw8gpide3K7RskZI/dBzu+UchMPAlMjJCFT+NRJEfbwVllE88UAG/NlnmYJ6TWwjgkU4M7o
zbLucvpVVVpkHKHWWwJlfSo9cRQrEEyeibNECQp0g8al9b82cD5c9Yc2yKrHfqaqt4SYUhWPtF15
zZjpDXGNhmpo1eCAQTmpa8zhRV7N+6fJh09xP1xaqW00lU3hE8diGWnegX4DkiXtkMiVrRgJWsRL
E5hr6kfKoxuucqDeCqdL/Yblmw+TXbpmWX9a0tH2P9R2zo32Jg0v8zpCqi4VWcetEqnJrbGUGIUT
Wjrkz4UL+mfJOXxSYk3B2u44YnNe+Xi2npHJ5HXeNAIHc5QbCaBhMtunbwaVoSo+j+5VSypr43zQ
rZ/dzsUVzvjqoiog3YSTNSY22ECjhKM8RpUCrpDKMGF4HWnBIwZloHwLDI7dl0bIS1VZPqkkOlrt
pJAS2hviVpP/enDxRIh/Di9MBCMMloFHNZB77Xul45SaDiSa41tKDjcNAxy9C7OloNZ+k74QnvqO
3c+eXm9KpP7Jc/0siYUG5+QiIluPOHtUk9zOC7nAv2Bn8dL172QP68zb951kBkUB7XzyFx5yJSoy
jpBNSWcW5og3IeyCYnPVopiVTgqLBoz0g+A8lUj6A/0H/1zJZ7tIK3QNlyeNGoheEwSdTLGd9kt+
k1NGdBFaqS7t8C/Ou6aPSq3wa4FtbSTJFYb3i0UM8PwNPZTKpKnTtd4IlpIk8PsMG+3deKMdRGh7
2pYlRkZueiT80RPCjM/iy3MXoBFKYi5l1sTsOdbP0f668g9YutioyeIcD1pDxgo9u01YHu3vOA1R
cfuIHCtRjLQ3CGgho3Ha2gyhqJapjbk0/OuUlPRKuA+pNGlDSwNTsgK5+wfn8FlbsTTuOAvfMIg9
32PiuHinAxR+7/qID6BGOXRM4DBppDLE/ZKqs/MSDvbezsgAL3ywS1SGLE57VtrA35/PDolSivnf
YzyMc5psGrbvv9jWhAZFEFqqel484EJ+3n5zHOebejOK7pDu9V/v022jPxBhqXapOR/CRLr6dtZc
/sbhyen3f2WyV5jxcx62lqkY5Ddoy4JpHd+P3R1Et/P4BAoXftblJ4T8rsMUk3r5Hnv2gTthpUxN
C1ue82kD/extSAMbyhVewrnyiwyTYn72Qog6jCpV7NRSaA6jeOwxOaV9UpN7J9Dod3VJ7sHKhCzD
pgNpwB8dELmMsWRWIqbiqN7HRe5zVCbPa2TRF3taPjhFGHHu3dNySKaxYbmsOhaN49Dg+l0dIaIu
dGXPY/Zo4ZfVu0GHluTb6/kVJDnDki+Ectdzp0v8F2xPfmhI28K3R8Q0YrnSow0KI5TD+0jvEDXX
exVoMVacNYPTnftp/s5bWlXggQ3Wrn/kDhH3k3iVNbzW0QFp7O9FCQ5a2CTUOElGEWbs/DMvMwHT
dbQcNcA3a5WNxZY9BGWRxOWkkSvrPkKwQAn7W3BKkRACSa83k+UB5Xw0QZwmoQb7vJ5Uh+DdtwdG
wLmmH8DYprnfxKajoIh/dMaBlbJFuxTPJNJbg9dIu84g9Yt7A/6dQWv2MP/BreApIBpMdAJYcTjT
8xR9Pr+CZeiq7jkPa9upkXpxVzCPvI4NP70s10cZQ1t3iPcCNCVoEvVtS8OGD3fLjn+6faRDvZu+
v3d6Fhs1PhneRGCX+v3fmrz7fx7uCLranVIR9BOHP9xkNtJthwO2SrV2DDH9xkLW7TnpEfdEXIED
XGiR3JcfgH/StoLxv8r0T/W0Y1UWptGfT96t//DJlW+6wYvEuvo4TAYymLTt01x/vNfeW/GsV0Bk
nM5MvK6FFaoECxYzcDYbbYOsYRX14Y4s0CntR4/9OY6tKte9fnVqtnq+9acPbqJDyxIZea2BFsaC
ApRDT4MfEyeuboxtFU61NE6Th6UQQ8DQMan2qiryqaYbi1qi/o/yvVYYQwZl/ewCGF6AZEScG80P
A2Do07izXq2NgFb9YNiCJW38uSi9mKeqlRv93h29mWKqrU5yWDxwfoYueDv+I1feQPDWxTWx78VX
5OgR1VBDoZzVtwG7ruboBpW68a5MnxGeYVqCLUzSSlmStOA0OIW9IAjsrms6gzmBLp7WTE2nORzJ
/uwFSfWDViWQcgQn8yRunwdcLi/CG4NQLitdVBX8Jp57LyJ0izbdsY7ALIYg65E07Z6a9sZx9mGH
xpHk6NvAndepILM53gzynqZWHArTKISPycURgZqdKjP/bQSo5LRv9Dpc3Ot2KLiga26J5Sb+ueyQ
z/Faq9n3T9175gDK+AnzeYOQy36RYdp508a44sdlmiiIyn3txmVSyO1ZTuGgsiavyHzV46r9/+rm
56aBjpuzEYyW2kiYDN53Kc/KAfb+dKst2rcKExSd6PasautORWxfyGXpYTydAMVWII9C0zfczP+x
PF24JVT3b0vnw6VKJ8QgjvNBH5vFri8ihGBwPgQ+gYVD2I6BjDNksFAIfmXTlzw2GvR7PaWOvbGE
llXtA6JVg4LyF5SCeyCxjaZKrUF/fLKbiNTQjWYan2K1qc6bkgheT1rgncMWhjlxXi9620HzgReE
vy6dBdsM74Ppn3/370j4caRqvRR/fcHDCjxksWDNyp7mMha0mcw/AUxOoD62cVqai0sAbNOdsfP3
V/1ZtwSLg1v59oSS3FjiKOqgkX51b80mHlVdn+kWQm3R8DaS8VYS+NkG0LsjMiBVO//vl4Y8yRkD
vYkfQ+MCeC2JyZOpeykJg0GgvYJVB2LCw7INf/X0ZcVaFZtDgTXc6rcb2MSfoToVt9/kCfe6bkFE
IGKrdL03ERDs01Pyv+QZSHKV8Gnz1gLkU6S0k0cBkTiY+sme9+g9tUE9fFAsJ5oaxiyFog9yf0Zf
hO8G7bYmOs/ESui2cSM3umHkldFHZwgN+gFwTXgJggEAgxZOLwnjjJolmGgHrIoKpEdR2T/EIvvc
0px+OotxcYLenPvE7YiDbltI0JVo5gzQju9aVSxAOyFjsfaHav2vbYgMNtJ8fVlWsTEhlj37UPkG
vYuOKZGpNqlmksuZV8lOCy7E9RQT4rJzFdCZRUjMxgfoDv++HrE2Mpc2yNEl/AeFCnDt7alZUG11
wWKQSzzOHqDWnBypoezyYySRpyOJ3CbRGoCsB2gYxl8IZsbrgGKjkAFkkoZRXLFllfNhrVDXtw9r
na+q7yKwzjaTKekH9lKYSGGgaeswWj/Q6dvV2UNKdnj/xc9Qblk2e7UKkjfOHS/Y104UnHjsaJif
W5JE3brBU9e7frW1BAGoGtwzuri1Rrst5ZLng8tXyH/EZFbB63YiAQPlc5JOqSGgxAaAXIrZ08b3
xE/oz37z3tcsgRLPWyjnbVGkzWb4/c5OL8pE0v3jRRMcmlNRJfo4uI4ojOw1NR9cv5F/bPuLi+Ps
v/pHs+C5xtF0Q0vO6/XeHtdTPARsvjfEkhqHNaVDjyviC6FILxe05Hdx3phcl56Awu6LFFM4E+qv
U1Tnu/jKcskZA3Jjb3wkDSfmNDcW79+DOL9iIJXfFjyyfN6mHcxUZNBikSVTyXmrbZGbYFaBbTCC
/O4aOlWn9zu1+mW5eB0BBI9tgkyxpBFEJJDoaLzNbiGoekzRvAyS4F1PPUqxSKr2sHhRvCRBAsiz
ExgGt43lybCxKBVsS0vy73gr2Asc3Sf8eCSpxG5N/nKVT7zcV5JnWt3xuiRFznmk4DzFphoS/SSH
Bq+GdPtI1/iVjy09eLWuPdlgzjPUkysjQZMew5ibV67aSOtWyjPFBQJ/W8XW2ad1sU+rbepKiyIw
OyQZk0oDxRK6Hql7YVFqRzMamDu2vcD1Y11SF4iaCcjNrtgSSl7gKjFX0DBL3+EmFLMguxX2vGgT
lH0hWCZ4+Dw3t2fZUNpTyQCSbiRIwRVT8eTZ8AeqnonCcONdGZM9N6ODXZjOSJqHO5/L9+fSZWdO
9qZ3+hcN2qoNgNnwp5UzaPFVFI9NjIaayo8Fi+TlspgGT5ROUJMCGV85B/mqne1FTqWILqwkrdrt
bBG34tH7NVDo3hu0mKdW/c+z3wlEOvgixllYsGYWk95c9cdEJ6cTsaGaQSeaq+GathlSyOvnK/R9
RNPDJnILOCwWKMaaTg0MI3TRpQ0wYBgk71ARqDbqhlytr0bthnYzIKnMjRhj0V+XZjUJOPYOMam+
YNi+7Fku0r3ek43zfTJLeAsbv/pbWTf/ZDZVltw55teeFb0nQ/W6ElJGbFn1LgNwn1Mjz2doIH76
SxOMnQcY2HOA2AXCScmHSK/U2JfokJw0FpCtGQ1L48INiidsZ9q/kznzfIgVGblFdqBLg0H4OtnK
dIfi/5JZDv8R8Wj/g4V0X0t2hnzb5/HadaeVuxeQNk81Vdq8FbCjqWMR99hSXMSiXVVjc/Ir7rfA
UAnVONEXrDDRZ9O3pjAN/DaBOYarRorsoCg13zKzU97AB+f1TEfjRMRSc8GsijQgcCOUVaRNEsmn
ZWbR/0H6kNzZznOzH19lpJ2G8Ra4ii6piJmqrGYEkVcrQq/deklf8YIoCwxe7Yh90D37IwGNryo+
fwIzJPclh8VCJ8VF1cMrn9pXuKnWsyd2C5HffkqaIclz3NjzslyhQitiTY+9Os2ussPCMpevx/2P
QbfmWyJ6yC3nPN5h3lwcHQBmh+bAYfJay+SzuygC83ivoSJxy3HnXQJJTWsKxDtGGGl+4FOzsPjN
YsIVIFE/uEWVdbUuaUpQXX+FDrnlAeIdtaEmCo0/pwNBNcWm05ZShqxAy14lDt7vdVkFocXVsD9T
gvV73uravbPvxjJXb6RZSShvvOA55I2v1L2shaLMkTuFKmynLWGlwCy+I9Rzk45GmIvkuwFqZKdr
ubdnZHCS+wlWMb9mmUMVqsQVhuMB8qrWWTVN2DKx+DmRsrVfk2Ha0mxkf8Bd+Bb6VyFv5242pfkZ
2uq1p10Ar+zqztAfyR9mJTrsLrZBXjrO5AIcRx6W1zQSV+9o2YPwGboxcWOO8jFqsHju+k4/aJlD
Uqhi6mcFYdWJp0grkVNsv4+poz4g+euHfI5UKw2G97+kWSxlYGAFHi1FXRo3tvZGDBFM5mlHugSq
cggbYcIw+Nz12dgy+bqYOrda4YvO7cbVa18pCZR1IV2fWlG0vfGUPIc0miUS2i/PsoHEZs8zZXIB
TcDM9eb3Wjy6NI2LhY8BhSWHpyw8g0c8grhle/BuGWB7hUPkrqVbtVrfcZooFNaRq6wYalgkQ0V7
JlHfHb6ktYFGok0aQEAPs3YOo49ZnilQuf321EXaXOqL0SUDQGG3HdTOE4lQRuSA0qtOKlwCVHt1
YSrVOQDWa0oAA5JL+E00NlYlcHZfGZOSQyKKqYaMONqvrf5PTSCIE8q12JKAt7s1SUMXwm3JIr/v
+szH+VwRxqR6HWXZcEoIFmPN3MrAcayDz8D0diXw6cxuDa9oFoaeRauyI56FibigbMcFFK+AM29q
ONIyBdYL+ZvyG8s6+QAXhcbl8LNdSPVMV7xGa6A2Eom6QlEY6tTPEU6M+QH5GWFwqZUPfX0MNwqY
iAq6loBLCbhjyUt9CF4zUm0pJ/dblqazLX0e/O9ww7XsYJcefRE+YjCuIpYB1zXqwI1cV+NkZMeh
tzrVYIt0+ZKf4QiICps8CIYKb+5cmhCsyFmlEgbQ/lTF5vr+b7gPeoYMTdzVO7ZDsCdZr0HEJjpa
rn2ZS6ZvkG/mjYP6kwUvmTkg4OiLu+EDqDuonwe58g6YgYeyIXaC1TTht7bgRz/opxVp5aJHojyy
ilC3e75tzfFOi7ohL0Sk9DQ9I37HnhrTRECSgTrBfxBpqYIRCTuCfX+YGdRQu226/09MwkresHPY
u291zk5rQKz4OsKkO2jbqv69tawGwjVtjWPYj+FjeIZH6mpp/cnqjqyY9yafwSpqnGVe8SFCBAWV
G4p1aVqCn4tzpxTa+skaDlz7HIYp8i04rNe94+b3XURo20sjA2QkyY7YSECqaUE4aR2PHJmGAB8Y
ZEc03fDp/Yhf9Mx9v0PIQeLb/Mn0U3NEvsiFpIkG3HkfhcZzIMiGIVd/v1UNTaR4+piIXv/alTxX
2io9+kGp5m2/+g1sxDDlk2BElJUDKiWhfURQfS9rMUCNRzlwEQFT9PQDTA6z1MSd6XVZ8Z54GZAA
/2Uk06f2zn0QW+9TYFenKf/NtlGAyqtX/ygHfrzXNZlBwuXWOsN7uCN73sxEyLuLSWqT9vPQ+lvA
XCyODxJmxPquNc0zBBPbriwk4pp3zUqo4Al9mtsUl29Zvo+WC+GAt5UWQAtcY9kh/FYKm6rttI5w
XB85KV1YCe8iL15aDGpInKAuQ4U/S5nzT/2qwsmtMMKTUyqooKyE6/MeHbFXf9DZjHd0A+6/YI54
hfETHKeqdoWHUyEbsRdvF8nOggZwid6ZuIkGHoH3mU5lnUKzPX+4+lxfDXE7FgWQ25tvH3A2OQkN
kDzyK28BkpzHnWZ60lY0cf4Kgd5h0CrVyCOiE6319JVtkdycvzxhbIEf++Xb8bW3BPIiAxkEc42L
6o0HghslKJOA/ckj1O+JBHJupm3xXJfa4+42/SPqNCU91+N4Bp8on2Y5rZuWoqVVgaDg6Jb5mQKf
IkRsG8F4g47kJy7uf04UaYM4TkZVRIcMqBmLJ0C8lC1zZZdD0tqSlhhP3jYmK3SOchA43IBGDJlL
cW1eE9+74Q1xWOjAJnYOGVTNx9sZ4swfrDj76+9Qwmhxz8Ocvo981brlOkk4vV9WTM6Urjo9n3aL
Tlbc0+HgM3bW/XrGhoGTCRGK6imLF7Bf7P+jQnn8vCpFKAN+MOpR/E3RLe8IgHOEuyxNxma/+MxA
WjlrrJCN6bcu/UME6YGVD5GLcTzyWJf+K6tX1uCZJlvn0810JdM1/xv9txu7g7gj6gcbPieSg8Lh
i4isw5uH3bspPNfRI1Ixd5BQP+timhi5jNC1BeZjV0TNGWAztQRShsvh2oEWdS4c7n+w085kNGEQ
hY8MA88/nllylguzyR7elyh8SFiNo2Gt9YcslfE/rgwstHTYuUyeBpATA4MK9fJgSsiuyf0vkNu6
TMt50XEBcGKNV/KkZxGjCtD+MP884nXyEoO6fYniTL2GgprU/MCZw5X9Nt9n0NzTYUEZQbFB/FVk
ftivngHAIIoBPfrf9xfMDM8a6DjRryWnG3MIHEHjqMxNkqleIREfFDqIPISqM/l6kmRcrvYYZpED
EZe8mKVDao+Uha2H5OcSXELu80/bbizLbGufAWFNZVNk0f7aLlHMq6xrHQ9xDnoiVlraLZxJG4Yp
qFSYJyYq6fquq1G2xa4qyQAmB3C2Me9D5sHDnv2H57AAvCjIngQAI/Tf+M9yoJ36uk0KAgxEK49B
6d82c0z4B4VYzDwHS7PYZI7gmQqE/ImdekXxCDGkVMDjcDwzFVD5cqEUT7Hs/5lwIo9d7XRVe1JE
a2Ni7oltJ0I5ubPVTAmosvgJpFuHUfKW0GEfIgVQRZaoNfWeTmvRfMXELytXiHmgZgSO8ddDYIGg
EsRAUWDA314dZFQ/BIwd4NczyIe19ly8cxUkcRoeAedwiVoRFXKY02zGCJs7ODQVtrtYgK83WlnD
YfCvW7ChPyYENIuwiCgkdIbJE4uRaT1Fp158FOW4cnjzRLDq6efom+B188NzgppMVsfbfKsD+Xel
Hf+Ch8YLTjRJ/LqqS++s6OJtOfJafs1Iwx3BZqhsyX1oxDM85k5kzwHpjfFbO5xUqnGDgytzx5Dq
pFt7jaFryWnkhdDbxljX72SmEXA1NzpL02W7kzGOxs/xSuugoTEnnzclMLudMdadnj9OvvpOTXsJ
W7JVCJutmGwfWkS+Wbb56zm23xsAJDKNjhBg5DO3S19VMuXDdYCDlMH8QJzNl2AgGrfr8jUcxBz8
xuIJswhK4MGhF//m6QPoTPD20foH74i0vR/8KTaJSiGtHHux5qkIJZ8fPvBrjC8VTF93NRIOsEws
d5M/MMYe6f4p0xnBKAQOQtuwQlacE2AXbiGUx3UEkGVBLoXYiNp4mszYEFslquYyhntvc9mkfmpZ
HyOnjGei+7c1DZJ8TZEZ62X9x8Z5PkCLwVb+JrCQ35y3+IK1q3GuwIU5da0Ztld5IaDzy5HbzNn3
p9ZOfV61FnN6jDnU6cVlvLtK04URnOk2y9F262y1K9he0p7X9eMNtlH52oH3HQb1ZQxCbwKcmVRY
WywUDnrihpGPVqWqoq49We283ZNFUMG31tK2dOV6Fnd+EZcYCXj13v0SEvz5+qcAPyBPXkwmGo+t
lGbyhqyh+nyWhwjgk8xJ/fYqISR4O9F+0pA8ObRG4suMz3Y9xaOYexlZZaMV5jJ3GmYYHbn30JP6
G4j/+/jHsDvp1bREkGJ3k5OhaLoyGVVAwFOxXJSZDA/PRmFZHrxwm8cVUlLsLtkWYeHP+4AQ6job
m9RCZKcE5uI87yTLqGTfk8DCkVnptcDLyDT3Y1WTW4sUnklBn3S7wedOb+2o2EwM4cj3G73d8SMw
iECtlVWCpL+mr1wXnUbG01WfH21PN1Lk/uzrcI2zO59DdNjYx2FbqRizWTlYwqsv0pbZUUkwMH8y
Hh93Vx6B1quaG6zNfQuTq3fSiCVX8dRUuSbKkn0JpTPl923MTclRPIYKOw66EtwksrgcThMhmsrz
FlLzCzw7sFjma7nDlVYe7zC14BA//TV6DyMfzw0uEmsj+swIad0ruxLgLTzvhw24lGkKlIgMIBg0
CJLjs+vbKgRm8piGoT5zE9E4pWUGc3NkoiuBNh67OleCDknzaptfOwOe/Glf9kq6GMP7d5L7XCFY
p90azh5MPoB9YR+iABsslAW/N/zV5y+RhVWX4Du6YJyYLzRDtNauXz3TmB4nXB7cMui5RuYl2Ci3
CH2XXWTuk/K4tBEpsmf7ap8nqdeP/b2dSS8fLmXdxJI9mqlvQNKhJGr+d4WuUVkvZsR3QWg3+u30
Vg2y9IZMcNugAadwxBkosJqW8L0TNWseqV0wfbKY/ZiJ45tP3XGZ6vPJ1QBO8Bqa62Zv22wp9Hyi
nC30kG3LCTwKDlLz9AwWgT9hjjQcVQ2SztIoDVy05rgH0vQ0I3zostKS9Q3EC/s+kC/f4EvH4ELf
MjeX8p5v+cEpucfJnPD3o2uxfwIzgtuFqUTGYRiY17XdpdhJruG7F2WCwJEd0UqoZDeVB2nq5Vok
zXF3CNUPbDp5OiXJOZAH8k5wH8qU+2y2zQ3OkLpBB25su1i+2/TAuCNcnzG/9m4l1jgJBsKwm5i1
+ColJqTQcC51uo3mVmG7O1/JW9YKq48gV/iLDMGQMtcganR3bC8867ZHLmd8XEbV24gz4dxklyYy
zjYQYPGmKZTgGahTME4j1wrGQPM1kRQV/dQM44INHCAmQiWuTpOQX9tYwMYGvfP9jSu5PC+gPx2q
QE0BZtxCBFUEjDYfWRyYi+eFgVpKHGFo+NuO2b6L/MLQS1bBmT51nOxQfkJTsz1MlpYKv10MI3CQ
3tmHu37gXf5/0xfRqOFQ7ptd1DAo7YPwu0LkeLuyOQWNCgsfiaeZZ705DpCjbz5NTfpvlP10Ss6t
O303Y5MPs158lu4AAS2Sj2eoHZ8kan2aTSGPuFDf7v11IJgz4xeysdEkgQFgP8e2+km+nr05E1/E
Z/RyXaqquNN2cESMEAvyQryENerg/6R4tG9ME5sxxn7mNK6U1g7+Efjo8q+hTWbsWFM3rDwhxkoB
rPsULYRFkvwKcBh0KRdW4E0Ah76pbLn/x8HRsnyOXJhLRnOIrgzQF/St5lqLvvRxggDlHp3rmT5X
MPjMu29lBxk3VKv6AxXGUM460xdvoQuXnxx9S6+DAfNIUfZqcJ1kTrfAwCFNNp6YJVqloGBBXpHh
YSVox6WeGIJTau+AqKdCzPW5AnrPqQxMrwe3pCIznrJ4c01EsdMCjHDCpsrtibUos1UNrYMH+TWB
yZQ5DsamIsVwZU4Vn2lV9imUEgSkoT/KuxLdn7NwcdV+OwLV25rz5PjwhI0Zv5ufaWT6hsIcbM84
yXAdyzaQ2XH7Z7a72MeBwSKj1nclSp3tUlgOJCRwk3S8YVveZ/xPvc6i3ztVswhaVHUppRZK7wZf
oveMcikuhDfTEumjYtwNmE6xy5kLzDRSAh/BtjOuqBpicFeMEDcemwypiynfhgOKdE7IQlrMZwr0
c2WBlrwY4sJJHpgM2pHuvPs/9j3OTI5xl0trp+9JdeO25EAvDHt6Z4KhqDYnPs6Wws6A5aAfXi7i
mmEXjzz+lN8CMfW2bIsS85Z4Az5AKvG7TpLTr90wCu1spbOPT0jEr3Ig7kwTTfUa5+cZZ5zEbkvV
S6CwONdqBHoLFjOD0Cro9uatHUlcGKU4qIL6Kwom2jqOhDGBma1JxJe5h+FraN21eV0Sc5TEPTUS
N76gvzM2/Nh5lONDRFL1Rs+roRXfA3JD+8VEFrCqtCfY+J4FICrmvMw77F/MvIkUDLvD+CzXWkIm
fGOKq23rHvSk71xr8fjxaq7+B2VFHCZycJM2A9l7DTuZ9XRphIs/kY/LmwtI5DbY7/Npv/zCIG6S
ylFAimwV31yK6BT6LvyGvsdisuizDKi9wX9dKMcIDuqvCcexluBnq/IHkJr8JS3blVYdabfEspza
shPEXUXLA5qi/PAlTyN7W10hjGh7ofxuFae2Zr5jntaCxExRDT4tDdWKPFHEsNmquZitPilgFkrm
3lsUvIr+2ZeHIbsQ9Zx2f/33S+drTDeMJoKUG5jcSsVa76E0829wavEu6MjXojeQMZrAwm8LC9LH
yr3/ra3uKErL27ruzOi9YY1Xb665xVdBJv6YR9L8drp0tvN5j44iHzCIuLCkivdiZXm1/09l7lHG
eSzxNDWE/u569zBI82PKkudzHxyB02NkDRK7ZAHSLoog6DPO/J2I0Hm4sGL0aeUCteETAEwEOqb/
jXUGP0vymI7gGvnWe4M1TUCVwE1gg32+HECSrSN7UTl8JJrEaOq4h8U3iyyB9YuonaOtqZqpyqGT
lDPcVNv4mvSF9GCn0iJKmDUUQnAs95SaHu1c9smXGQooABRWqwmUohqSUfA2Ke7zc3a2fvXMlgF8
n/w7G33JG/1dEHZP+iM/0XgRkDzNRKF52imVoDiK/01yzT3NvuicTbW8gMZRmx9Ee3MRKW9Ddm3q
vua2h/ydmcNg+qnb0B/B7maGM8GtwfrX29eQjAKVFtwPj3YyV3jk95F++isxpNdu4Ws7tacp0DHz
CvmuMsrkqGam6I/zaxKMjOeVPKYdsZKgLtFmb+7x9fXA/uIvQGTKrNI8BhTH64ybbtmeEg0s2Rri
YbtJE182tUnhnGTW2HzW/lMjwv9UuR2zpL7z8jaasT/o08kpzSBjJUQGT2DpseEpigVpKNWZzpgA
Otu6pdW+79sRSEjXzR1tHyhkoy3X0WPc64MxVWHuUf4UYLAa39aszcaHHDRT02HnUwB88ejP/Pb+
1O+aX0v3Q8iZBne4hOdDou/oLNMoy6T+GL2OPxHmCTQQK8qOUmbpegfq985MM3warwdXL3ddl6W5
g65gY78YXYSjiHsuOGfpKLpVKbPQC7xe36bs1TZZfH7gw4dnxJNNlcAhC1LMTDEaVUX1GrRXoL8F
aJTczPZviWTCtkJ2gr1+IMy8QN/6yngC5/UvCHU11YiO3fd4D3OsEw9xA7C2vsBh90X8UshFpj/B
WuDE0E266UpAKYIjVkBqA5AcedtkGAG9rXIzg1mfi0O25VUnxKla58upIu7SnvmSa+QoXzR5/tfe
M5nm8wK0SGQHudlnn9DVRHHu17PkibVlrveclnafKrCk2dWVp095KX/IcOb5Ee4m1Z1QMGsIYgvZ
VoJ+K6Z+nGa0UvnmpNIxpvcgWkOcSYxkhycXnE31Eho4zJ6UbjiGQOHsnzH+UqmgAF9CkAyEWqq2
m4I4fa5rGGc9I2aGj+m7sOVT5PtVR9WXj90DMoVzl3MvHyz7GrAnF2R9e/HSHfpXd/Of4I62y/iO
vC8EbWw1RJFQ9z2rg+v5UKYSFyIfJ1FXz33MiKqFZTmNddA2E003T/1/pguT7zEk9Qw2kUE0enN6
/iD69//xcbATHxtbrayYS4s8vIIfxZnKIejd/ntyNi2+P5R94CTyUs0ZjlYTKiD9kVHlCJMu6xy8
KeoDyY+Naf+CyCABbeos44LcYXiWl+2kBHBRJL8ReePwQbOWFFr6wpu17ZASqb4GbYqgxMkwhBfx
iNUmIzlUxyPEwX3oqgq0HGZBVOh+qF0qLmFSBvPEyHddT9VCo58J+GO02ZkHTlvPWuj0ffS3MaaC
wJaa1jxBPIK8SM8Tad7mKokD4kCzXKkA9fSeTP/Z5dbCc2bDbFplbLDkWfGUynUGIOl2U+/zttYg
yxKhLEn8+EPpANxxl7cmkzzNYquY/BFwdfcW8u4T0nGEZKAUQNMBEeoTP6pY0kgtOQCjC30xakws
5+7M3Hur0DZNXY/+JpKkkW5qpSYDvsZxU+wk3CAO2IxHvEvSa5BKe9UvE0/8nZtZ5coFxApkiZXz
RGXPzpShf29hlVTJx9xotIKxFjECuTfRpN77RqKxKUGONiSonHnPknlT3+fYnh0XBWJmGHpfBnWw
MKjhhjPEnEJ9WYDMd0VWBUq+u9EinNkRd+EMcU2zxalQK7ZpfYsMuEI48UedxxpEliTZyTA3yfBO
hGFxN2JvNlKSIwb+kieywmpwWqVv1Cqbubq6nmJ7yMzZIvtdXHETcsqxNEE1LyI4c5+jkq6RDUdx
z9tw09EEa5J83wvkQSultZx/NTcpjulIwWjo4ndcZmPEbQEWnA+iFqkhzHng1kyYFKPRYoM5O5pI
8HwbZqEBCcoj2nYdpkPkPzbHUQz1H5OiwcGBKVBzU0NQrHwJQJ10HFrn8x7qO3PTGfST8Ul1d0fB
ec3njT0ZmmKo9PovrY4HT44Gns/ZFPI068ldgP2CK2EuFYOiMI6QYwLK3nT+Y42nklnXT565ldqf
CsLOhMc9+oIoKSv1IPcPTNrj69VWwybaK15hXxtW/f7OMZw0+5/VnsiaC6FyO5hSIMd7NOiomIyz
sQQIDGVf49VfIy433bEUSVH0WTlHKJQactOSK4XHPEmOBLqiGQ7lTcKTI0q27pM1+oOYTHPv3GM+
t5U62r7aoIyDJ/baTKchXIJAnU9pGhcxXrkhUwk2Ghgs0HUHZtpV198zJo69b+Tk5MoLxWhoMgPV
CJ30C4GxlpqTQdnPo7wuZGjodL7KtipMoFSqWpT8VLzYqLErD9Gi07wNohzvxcc3Zcp+7IehaHtJ
qeLCNLZFAPqsh0xtzaEgD8xYFc4cT5/HkYEQC9feakF7/ViSN+x10JqTi9imeYsBjsiTlXlUPUXS
JeJNnVpBq1tHv99ajvsGDniwd69Om7ODSmARaNUvfjcTAz+gAdCWGBM9/FpEjO9F8w5lU0jLjJTB
3/DAh8uhkivylbH8eU1NxCm7/ZnBAZF+vXbOWZ1Pw/ZGe06tnRCa7fMqCWJ+Bgcb1TIL2OqOf2O1
8ahgFSBJaO3H2nUwH9nTAOimkQtKw6eTSac7xFDQbYQX6tJYN0FyjW7jygEIhJJtDJ/UKVL4Ufpn
Xls4f3xPSwsL178wiOEWDQgpwrcaTTqZT4mNC4MXgV0TgSUbYjnhJn3cmAp14BnsxIelQKztugkG
mKPPKimp4mjgMi3Q/qifeAAl7twpV/a/tfyJ9U5DwEh3sIL1sCczjmEuyk3kXjpsN0qhVO9qDkZr
WgXU3U3qMz/egqCIGwwAaqbfTyUyrjWnxCF10v1zbMTQGrI20z4zunGnvIuf1mTxfJnVJeb7+ZmJ
QrCR9CBzzGmxFaH0u7+NLX4gub8Gff7ObWedoWUUmABHjK8KMyimKUi/feQ9S04QJtVdWXOesiyu
mOsFHWCnYCGCaRfcluMXRpYl8YlbrvBtjpsjOV1pfIOAm3QCxnoInWLRFJAOs1S1VRj5h07S/Gs8
YIjFGDKMqokjGFNAxXcynYuqCpEnSkvkAnYcWDIPURJmfOZMwXGQeLHHEsJ3apbwioGeLLXWGoKL
QAmLMffth9t5KW8qOCWOGsThGmAT3pM/Nga9tl+U2N22e6aQERFf684iDOVfx4EqqgE6Oak5LRXG
CIZMZeMNkNIx4PUykwUC8Ju1uwBFLQ43NzvFiTw3Z1YA+ClVRYV3JV6uwhGSToP985+HmVBQEpI4
dO48qhrL5EOQ349hBm84d6FLbXreYPR28DmP6hL1syg+3D3CUwXYOhDhSVgRTk3MvCcdqLWJJjWT
uvGoUVvPz7afGZLx6HHqZTWL3TMa4OzOAMLO4LgLoKCwO3CwQN4FuDbxNSW8EKCCj+PsqBTWA1KH
OQ7V6+lgTvbDyZ9Dp5qWtX4FO293VuvHNSHa6hqVusePYqw1kTib5mIYbP7H58YcfqRCre9ayRo+
8UQt6nRRtZnU0Zh0/Xp3+ukCj343+QKTGeIckQzE4EAz/Bnrz7M9EPaHgghWlQCeSOJ7VQRX5diY
ipe+RK9m/YqM7UXrfGLUrjJLMwvBi5bR6G/3aSP6gCRs4ICCdKVPyQWqCmOXDuhHe9IggBcLR0o4
ElBT8IzIX4nv+VUSinPqpKn1ufPo44op7pn1RsD1bWQt4IGxLNQY4m0X92B43GswfeX2j/+SEs+h
srRU432Cq4+aphU6x3cFT5+26+YIWpClgCljg+8rClD2kca8XkVyztyp46g12uL1BTFwlg5RIg9U
bYhvKk7wVEyuQhAjGiKsM2eq0Pm2Iba+h+MzNc1KjlFP1G/HOBdBdnyNv4YTSd8tBOXEsE+epMgF
FckEsWRJ86L/GRsVdTuiSWkH0pB3S6gNi0mmMh0TAdlwNjMqD0HNWz0vgpXOMakPWumHaHKPpOEg
43C47M9AGoSX9dqpTmZy5pbL+/cBNmC3eYxhuer742TaVAnO/bTgI2ZGCLL1NgNpmwupgiFf2tGK
RZkpOq+cauCGWaFxiIymREevqB8xyU60l6W3uOHtbbepTpMDB4OblNr9Ic3iCgNOmW+5n2mtUGwa
aNnWyXtC23P1NuLnl99dbYE5KewMlaeNBtO9rbcQq4I18gTcfD/AAgDSYymcgX2LohGraOtYOE+c
T52l6Y2tRGxhPUma+dAEG8KGRPrqgJkDhkJpjb352lRykKMLsbzTew6rDBGKe1Vt03/z9UZBNyDI
mrrtlizmGWr1/o0Ck1M/hAGfkxC9Im2JfR7vu2oFOFjZkK1bT8AUa5akEHRlDz/x+RZgad823/od
vxYaPIXttC87Yz9r9PsUMfwgnQmbm2bgOvjyvA69EgCPWhpwYiBkEuH2v81B/A1Kd1hc5ykwWJ7Y
umIgYHBWZvH9K0e4GFffLF3bhjSvRbdjegdQ8ExIwbOH85IHDAT/Gix43vFP33/HDofaiJhwe242
wwOTREVRXIaiabL8UmcxeJvDLHXeJjX0r2/HaTFmIPL66OvtUMJNfnqYmEZ1pr+u6zMM8HD1vF4w
aN7hYpYatfD6u3uZAD6ZHTCqNtycwUH7L/WDINi+mC4bT0htF5aooRz8UDTo0pqfSTgMw5tB0ANC
m76qNoqO/bBewRKmzswArBFS+vZOxIN8OBsR3zl9rGP31qYCLuOqUW0gOnXaWgk4RRx9K5VF1uPU
7FnJ6c7Pqqv0ZMf9PZ4ju5NKCe5TC5MnDPKLtcvDNhEFjdIPatkq+9XOcYfXpsU2jlw8BrQjU68m
0NoFR2FgfKL2+FjatilKGwGjwcfRLMYNuRTeZbaCqYL1tEwe1TbWCiYia5fLI1XgBzsvBEFoGCWU
+JFiA/312pZV9Qx7++GfVGkGkz1aI9DUX7Cafq5AyJPgKg4do6Tb0VaqlOe6ddqA07DPb5vWrEj7
vh3Cym/813inijBycUE2g1UxqcK5Gup2fQaZyunKeW9RTAYm094q6to4zAVSF36TiEQc/q9Y044g
GYkffymbHbOID75sYKqkWBi7a98Dk4sIwODeulwoJeZRxncBjkZ3B/7RoYBN1EwUY911XjBq0Roi
tXYf1dLlVvFXMHDVFhfC5CUy8o1E7w69V/iHtn2a9jED0iAr2zy+TcM6+xJOLfmhs7pHHeujs0Rx
dLNutsyPtBIxItTldFgTY3iRMv9/t5sXMJHsrKWHUs4ZPpxmmY76YNs4Az7hNqqzW0LaF7QtQm6F
j9ChsTMrnsZVgk8noWS2pGwC+0jRyNBrvyViv8oHKHotVmMx5ebY0Adv52qzYy144yJyGTjTIQqG
jgts8Fj8Ai1QJKZB8rSVEpTK6WmrOnLiArDo0BuU2Vbd7MzsjXn7onku6w4+5jYfbXTsOXtyRXJC
Kuq8EYZw7GWEKkOLG0ubdWSu1Wop/Dvbrgk6HV5/QL4cVr+nPefX5JUpG6BFfrMJ1imeTgvGDhhA
uJIF5ljsZb5dsvNgykyedHaZ/1knlngRQgfbfntFKDO7GRy40aPcPugG/jYKfqBVaJP3K7NKgEJ9
Bp2cicoHsOWe7pnzAQWxxsVLICAbwxdrDYTQEMjLGQP21V9Mzdl9TSOtbpGhqxytEEuEUKVTML6r
eIY+h+0C2XAGQ3aqKD5NmrHZPeOF3ndt6BKqhvVfacgPu4BbqfkL1jlPQyxTiPncvfvPOhfI/qPQ
ZjfFEDPpELifDRDp/ipkBwm4cbXgSKZUss/uamqp3+DsVTnYTCXTzfHiw5JqrmvINHosgYLcANf9
1QnYq/0fIEkyn8M0mW+eNrif0FsMdmZkbWDxQgburYAvjudOKP3p9eenXIwos6TiKQ2cUdk7CSSw
9n4ECcquNNshpJhj3L0jZf2OLZJEN4L6wTq8DZx5qozaBvgnt393iRaWr23betnoLFzpZVuDBLim
+7TP3bXU+62vGNlVGtgLOrKynd+xpXzu+U65VHJNrWGqEgw+2vsAxb9oOmyUoslsEbxErmcqBG1F
BVm8AVd291key8ozT960sP660zs9l05NzOlELAQSecDVqla+IVMNiDHUPzwcsrYIDdqAZRinmjye
Er5s6/hnop1D2umgonv335QWYlMAuaZ71yeYlFWyXY3d2odniD81m+TfyRdYJ/Cx4+xUJIKxRS7u
5bZdG8XhbCgTj+ZIhhc/+RnVsGaV/q9OZVCCiRG8EMV4K5ha/TA0xLxqfBtxuweYMU3dzPoIGfQ8
xtBMG5SNO3prrGRlqettib0ReEt6qC7aawHow1YoBOp26uJrUNrENA6yZTpuf9BlXrPgcNTF8MRu
G7eERrzQV8ci/QGSIrw27/I8kcWD+fQ0w+PRTKQUyb+UfIwIHa2L1yGHfJSZDK9J7gRbc1dmuCNM
Q4nqqQ2+CE+Gt0Yz8y/sIY8YJRCylmVqObKtBx1UwLMLlbSxuN4XTUd9m6D8GmQ77/Ci39YxELg1
Ne5PPBjjOwNq3K/1J721QwIHqZQbWIm56vclx4U+VayFEfTcOzB4cDEu4FlkW9163bYW61/q6wRe
zXwDIpbfkENWywJUy6yVP1OrMj8KptCaRxVYCdoq3UGqaWepOsmTWxcmbAWpozsedeQjr6ZNp5Qh
I+3xfzYlzQEAr3cUSXkzDLb77nbsDeabczSKkTcO0m8iS634NVuHN0LRT3uRdJbTDj+CnzD4vh3m
Q5Q51AZRFgtDbg+xPo8zTOVIpzzeaCAymGQzrwpmYQG6AA93kRhnE9pDv6rr6HVp54cGLMK4VODO
Gk6HqIDvFmAwT0i7TktzLlR3Rr/3V4ftfr3vqqSeSNjLUotRVdD/PTLlATZJbV/l2GvJ/+RqVqC1
THbaS3o2N+amp/5GwfHBFhESgLIeNvpKj4n58bT79g4uv8lbePNg1K+ZGFpHmFdXOuiPrPIO2p6E
QB1QbJqs9tDyPAKWKdGiLPPZQSrcqx2jRny6K80DtxCkQL1LVeZuNZWWZ6Kgivnq8q3WSwjLX95/
xusyfWq96gVmF6sTC7RPlkvTul2o5GYvfB+6x5B/zuHRKCWs3v6+pWcG88sUmZyI1BKtYpDRIC7W
QI5w5q0vuJP0L0WB4u1+dcx7tnBsksR9bOxxTAxwgPGMnQnRN/nra3uYSmtOPcB+vkjJnnvfuwCZ
YSXHWRZWzDsxFV8s0MSqVVFmiWNC31z8dPoN2XpoFUlQoVJDsMpZP8an3NqUZkL51rNgw8WU28Be
wDdGX3kWTBfmd/sDbbAGo3rjFiGSnj7j0hNZNaFNKVkeQtwGLshNCFKfRUcmtq4OkZT3H96hbV5S
y/FDh/vgR69PraCgQ4IJ77xjQZLb+gz5mYN42jbyEvcuqKb+lMt0V/k67pDLJ67yEanfbeV7ZGqF
FQd2FPdKeCpy6tpW0BT+42SxQWIH9SGiEfOR3hYBSCc/CH3P9K7XB7NuHIhUOoewJpOnAj3ZAuXy
otaQIR7ThoFoEEmhMWl7S0e7uM21xw1hDJnpaRQjBsVDnOduYAuLzEJAHg9q6oo493anaNseHKwl
EaBu4f0z/Byw1jw6m06Oa9wLO0BLYA5WJTAuUB7ZbrxskoDabYkYV1NvRYvr4bDVht9e455JaVEh
4RiPCq96pbv6Hi5DIqPDQLMiac/CZhXu4R+0G2YixKVW5RdH39BSGMAnqnPpbxuzVg1XkrkY4FTm
0VlAfBoJi/RU4faKnloipge4LcpP+xLcZvlLgzBxN0jIqsOihTa+soFgMoWQRVB5JNiAff1RpWBN
yjawPn28gSr46wFl0diC75oZ8mVc5ANzdIFstW5Z9zp+yKIwTTNWaYy1xqwtfQCthtaYhXNWO2rQ
mFuo8ojUiwpKNaBD7kHPj1gjNSYlQxGyJTROoBfm3ILyQjx9E5rpSHck+3StbP41mu0InUM09r6A
NaFWwhL3PemiGHXM8wr0Dcjaxr1ATNOhZDQPGYl1hwtAopa/RQgzX3PjN/iLhBzquPBd4679z6Kv
S6YEH7MWjP8EEDDSaAX2qjlPbyC0TkUwv45p+MXDnVzClmTM2M9Y9evkmqurIlflfrNMpGDi6XFn
Vhzo5+reZAgnS1uUzlU3uy7jONzewKC+D483T/CtZlQFsSlMVxb7Ixk+dHJEL0UNZOkQ37SrAjvC
734bGqb2cDWDnuji7YMhCZybGX0uE0ryWqtzUintLi8FTahR8usyUGLsgE+u8O88xL1r2Ha3S0xW
haxD7jspPhthzc8oQiCls7MysJBwDXeokD8UaRC2Q3WvM9mryugDpTtjMcoEsSa6BrEy9w6prpGU
eCtodoi17ziihumFHHS0jJRCbCj+uqYBrE4DjclA8JwP9Byw6/Ra+wtuBMCIXO+7jFYWJ7zRT9F/
nvSAaMGHrI9ittrbX0mBeRR00OsYFj1gRAd6ZZzB7o0Bfli671tYBXFvNMAckkybSwiJeWAu2fhJ
zDcjcL88MxAZKmpM5+VHMf06VJ6Ceb8vzFtdKZPkGlH0SXMgdzPouiFwCcu4sifj7G5AoVPzEhmX
1wuX3k2/Km+t5UofcQnqcyJHwTKgpu9JevHT7RxZ63bInU2/i8ENViqaJpS3jZ/yh92mQnKDimTv
eCu7Mw7x0O4Ez12AG/FE4E7eWAJ4mq6uBKuNge9s0NgdHoxtIY7QceToh6mytjR0VI5/bug64ohi
wfDuwDZ6njwaPItCEAxysDKE2QwTWLDscJDfSV4A36q19Rqg0d0oZhzLPn1U3mM/FRp9WEyXgC+e
Fsp6yjp4N4vq5tAtrSx9vt9y3MpxzTyDi/yypR8TCm9+QQQTqwN7jqh4LBpVggFmXcV8vIKB4dvW
x/gyjmtNEzLCxli/5kkKpn0dFNUdk2q0h1Jv/MrFz2sJU6vbah7ByplLjGDKIcKU6HCvNeK+XHam
HrC41hpn8WOP8FbGkQIz+Bc1oXKtK+9VGq1WhAPZx6iBj5ar/j223KGD9p748wra/qxdxWCWchhX
gCGEjegRMpLGKXUkr8T6KkXYsSjy6f6Q6TTATx4amZM/zSUWGeVBTHN6VEqkIyrDw99oXiABxMKq
rTYwE2lUNsQ4nqdKAjuT2Oxv9BVrMTvoIID/C5eQKl8qyo2RAmqP/rxxRZpZEFo3Q4HaPDo3m+nj
7zJGv3QzaOnjkK0XGCRXPmPrfDirZoh2fHkJQaBlHF8jHlK0gBP5ac6m4e6ezOCc05DYTF6yLOHh
9E2FeeSEmgjRVJe/jKB/iQ4dg4ioNl8Igy1kVS1Sc1LcccFFkPVUInq4Rj80RSy8Y82vlGL17c8W
sDPexmcZv1J/ibKlbaJv2iBZY2KtvMs56PoyNaMvY2Ke4LjPs/hP+4ztsehjn0cTdfYeuC0+pZna
+ZoZ0CPYCw1GzzIXChnC5I7auT5tJgNXyZR0ZcacfM3V7h4QSORk7Vm36YmjDG5C0U0dS1h6UNaV
UH2E6kPR2XrV5H4IrCThLG9lRC1JMUUdbEW2rzoLcE/9mtRyVZHaq9FwWXRn8MBhfkNiv0Uvtorn
8tykbIYjwHdeRQta49BUlZSfimoTidG0v/dfd67SYJQ2FOWRej4YOZqPW46wiQ0Vhds9oBDDPZ0i
imBVPgV+q0Xp/ATOnUgJEfyZcgJi4wc5MkuJJOci8pGW54O0VWbsovAD8x2X41abZWN1vQ3OoJyB
kXkoMVZ3G2JBsAgOikC7B/fLmBRPwOXQ+DJcx7kBOE1TuYzTFWRcnFRylv9gqCAUbQrmFz8h8iZv
Gt32sgHC8mH47OWes1XWkR0mNX4sjgC00ENUdWrL3kcqTq3FUNy0iQXqic1fKUEam+XZrAN6tFl0
Rcwhh7emEiuxoliGU+CaGD71Tn0we/+a5JmtjyE34SD66kXftSIVtRm8iqAL3Xe8SP7Hy29HSATC
LVzkIfrJzsYp4SiyNg9DfA7/j+1UMlhcuq5Q4xnWH0ybTXyOVD9o7Gy54gmVUladJXwZzSbyU7eQ
9w0RBX/QgzOlZlSeFu2Ygv16wG8eDjbIeehd6SAwrOGroD/4NXEg4rh55KUIcaIoqh0uXwUPmgXp
GD2uqkRJr+FzPhQkBcKQrJdpQkunCRBo37gyTI7XUaDx6m57756I+trwhvHDZfBlfacfvlv9wwGh
YyceSBFmV55S53NnyPGV0ygdqipm4ywDH6G7tvTd5SnrjAUrqwfOwkzXjaRG1bnsgT7OTZHn4Rw7
h5bSzuzbJybEltgH5K31pOUy68W0CAJpwnaIxH9AS44vQNF+JNcSly+AKg6lnaffVxuxrMRkCKZs
T78gsr4EUPtKBut4TuXkv552LLooViDbto63Hm83N6Q7YYWGlUIpXSBn5Cn0djL4U9tyPNsftQeR
5qVgCPq+xrhHqp95JMTPmO7PqGwjBmtfU/Wa+BbRi2RVwkICVLp9d9E/JJmjirVjnFP1VvVMWXoh
SvM5r0HuMKtKYiX/fQiPbDISfC2rfMZ9zyJix8nldNRFzhPdKfeo7HOrTDYO7HtOcsX9qEfxPzfJ
DXL0eLM398GxeNMXSV5Q79UBX9AMq28a8uGEJyeJu6tKbmDFr60jSY76ohIMgjX9H1V2OIIJpb15
la/m7v4o81P7S0a21HvOeYMKeFIL+GtvtEXck+FpmygS3IMgDlvj+L7HV3p26D76+docvpj7J1Jg
ykb5X6Ti4+7lxuta5b88MXY4v9PK60Q4HyhMSzwDx2h2lSXW3Wd8X9v5wNr8QWqUXzw4Mns50acD
D7lqS1bQ2xuCb8rIPv3lNCk1Da5gcYwnJrHx/GeNDV43oVpAyc15pG21bM0e7WProK5qKoqLd8j/
BY4d2KjNNa/MhxZoTCVOyneTiD1jUvhjhu1/HVqgT7c3ohsqHu9o6aaFQpbJSbBck0Pnxze8XB/W
Ke9cJfa/ayOJZpHb5qwXD3k6uucHC/Ap6Uk9/xxCpk8+V+qUF6meypnibN+3lVMaMgRQzu9U8ITh
Aispd64ofQLeVJConCOt/MAzLDfqpJ95EwOPqZyrAFM56icTQPjfGFz84zAW4XmjKUM/hxknTNUL
JwYb9Ayoogp3RkEBq3mq6P3/jdHkX3C21l7U+4cxbNvsnd/Ai8M0/kR7aiMvtekM+D5IJB+BNVoh
BLEKBUGe0L58oA6Cf3OtCo9cbZ505letT8KR3sK3dom1gsXfygnB4NbfgxNLuARcRX+FCKPSqLAD
i8/6G2yBwyf7rmC7139sdQKTG4U86ooclv3GLWIlPYLe6ZD3NAczd8LpAllcmRoSoSFmV2byMov3
CoZl/oDRq4RbFhwOEKBChUS3kMcVpZHtahrJiQwb8t/t+FsUz/vlkEJy65JnqPxHJJBWaxPnDjom
LNccUcisAP+bhOvZffSgBgh943E963BIdKRXGe+L+Dmz4rqr9/nE7DAjmh8BT0FBVcDXb7gl2caT
XBMz9tBVVyJYlfedPZIWovzGR5g80riZyoTf0SylA3QmpIzNpMVKzwSqIUcjaAABiqG9Tjpaw/Y7
/4M1pne9wquFd7HavIo4fVM9468d/xMeTp5BaMPuUqR8UQOvezgh1m1b80SzMiNAhR03TvUjL0Sx
IQShZz/X52+jDvG1UNmXyMs2vqcooziE24C4Jp5kJk4PZ3JWe3llzAnI9Lg02fzsFJKIrvmjc9uT
PD5oqM6zXYY5q3zi4oiWro15o2hJC1Cdob8omrgZfABDa8UKvyIx3Pa1cuQWqPHVeZSphUtLcLBq
K9z/zMgKIAnnMNUlgWBAPOPaXP16zt6QCWSPPnEhA5NxinFW9Yo2wQ/6Cmr1cm2e+06a6dVKKN0O
WtqHcz54A0p8UKXdu8oxzkWy7CxPWLwHPjAid+jlFCUIfye3JprOs7dAtKUBANtNBjrHSkdYzKS9
UIAwmmCluGK3nCrNsdN3FmOhU1cQoohct1iO2yHFz+STyEVci/EJVZeTA9aLqBpYaeJ0o8Wlzh8Q
Dd8j5iWcZH3lk+6c5nnzhq3E93CXraegmHc0zmWXp9kqzDSSq/6EF30/KkHsbwI1YIUPfdpHSFxi
cJI+EVysJPk1lkEmVvEoD9Kj/pwv/CMGEE9nxtAmYNBILGiKxYgD4J5CIoTLuQfSLLT88mDMf+pm
shaqy8H+voDghF+cYZcv1xg5DYycG2LhEtvGybmJISxpbgU+x89rlVKLM8vgPfY5dG056IWH5jgA
mhR08/d4J3TOm51WQ5/MuKKnNDVb/pAszZMj6l2Dlg/cM2Gk2zST2KV/EeRDIVXE4zbajePYb2K8
y//8O5txZXuSFy/SYTZBGh+2126RLtjJGuyebJbpHLc1Bq8vUi7/Q6yFuLUTLaMiQIDqbmRFCh+z
P8as+Dk2+j37YGNZGUAviTWEAmcd/Xf0+cce4Eva7nZDitcoSC3YKXY7GlMrn9Hvdtats0DaqY66
b1Mm2fo/lcHesUtsfDCw74Dg/Dmg4Z4NcUmO+NYszFRxqQ/01yQBzRobCBttFabUFdx5jalWEOY9
FcrEkF2TQVGdP8H7Rg2W2WqqFSFyHnwug4Oi1wi69SCgui7ajHaIbzlvo/vQMi2x+08aUYVUTckN
vHezSp7kEIxUsR52sieIhpCqkKkrRvyWorLJoVqUKJiagUqBabzZA8UBoSpXAyxwu5oUoZiQ8ATR
+kR6ttEcmd6zAdxKZoME1jh4+Lxpk7LYUf5f0Pu0ZYrByINc/LlvRiU12DOWHZcQKF4bSZpjMwdv
c6wvccoNXzQP1Vf3XROwk94UavTZworgNGkL5Upb7PEcU+B/zGFrp1EA9GQJasIOtHU9hMk6djW9
t3fJ1IkYk0AWTU42xWWy5FLQ1VlBeLh0c4kuAzf+ZWJVdRqbgHUTejlplUq+6lk+oBpVFW3yeQfm
jd+udrrV/mHExGtjXbcsPaWWaHlxmryMaT6/65uHUvQ0rr7ryXVaBIBWVdSoKR2e6FZmFlBqybJ9
EIhWtHn6RkAs1AmovjCVKbYnMZagyAJIRmFvv2guHKZ1vNQugCcsGaFEChQTZUNlfP1sC6f1s979
aRofmZGmNZUOdFc9ojGbkRNgkGTqxUELz5LNR16TM7SMYZ/K41QMAH4NgoobiE3aM39NwwhgtcKg
iCLZ+7eCQ+4mJI+6Q/LYpqBBrKZplKFr2gSmrDrgQaR40+DCSy5chCVWnAVE1h9Pr4VWptMobPcf
TLLiyQQKjHXN5wEvFhlzpsneweQkJ+oUuk2v9XKLPjYEcJBZgoJeFNgEGlisgOAPMSmOwo4E/VUi
cBml9pEyVr7R0befqPPbg+WoJ01MeTLGXCwBL6lM/kjyJPaqgdHlIe88jrkoP7FdvBDwDFKfvBe8
oAMJXC8TpGUOGMdinal6Qd/pzvlJugNvNPhJPl+AUUdI8z1k5S46u+BM2x0YBtE/h8hzJuStcbY+
RJ1Jy5ZKaQoInWaBTnX27N6g5TctLecSOhW5N2yn4q4uOsDABYQ4qgjqp8piUimv57F6xXmB3BSl
c6Nsdm/nCvy/5SoEBKEdaiMOG9mXyDNke0Ysa12o4ISkxSWe1ukAC4WxfgNWAg6b/w3gaVU2UZmF
3GAjGraO0cYY4c4vo5dbNEVoGwWKai6K0M0VmcYkSyIJoQzIdkN7XgFz2KHxkNx/mknnqFRQ0c4v
4ss1BdagtKtrG1E1GyMnQRSR2A8nr5Eo5WorX2cUHeC70tzoNZvEbWjps9JHkPujX7sMh0BLshKB
rys1inayy/cH0Lb0ruUeIK/FxZ/XyIeI7Menya1WZPJpINl17BRjjRM6EwF6huQ/hgloIEiiB6/o
KmjzKgTib0tJaULtGSDd+5T5ba8WmruerwXgVLFkSu0nVGroLtUgeWYJYrJQ75jutNV37oacFORH
djIi/iIf8JPux6PHEo34/bPC36sI+oFwaBEyxyczkMJhlZxq+kHNG+zP3G5mnHqsPPk0qW9vyJXt
vDh8C1Xm7JXdI+2rHJ7Z8223E6AtIjEu+EH3DBl4pMSgNuHgEatsxR7tCS1w+sSR6/wYXM+CvVM7
Vs5otoXcYiIzbGAMYMAdSKPhPjM4kRd9gI3/PP6L/dw+hjFq0p2qtoKH7HpaVFV0VHSsAs5XzNYH
niryEBOqGQYKmPHVpWysqpMlXG0+3guGYJnREJqcuxWBk/WSxPEg15fSZJ00aNd7nDwTO9f23TEk
//prIt2dKQ1Fmsw/DiJ7dy492DlwueaZga8H5jD18ja5vWy0EZd7v0jqPhl7zy5OkcFwIeVRpTjM
wuYB94eyrvhFGvxOQaNH2pnCtkDp5cn4kfCxYxqhslq0FPy3A8vuIXFWZk50/Qw7MOw0DrK7DW9q
D29awDAikDPEVRpiz5xzCpuhogI8vNBkgB+lz7a3gAwDueEC6R2pKelQmIrMuEAZua37IcCouuGR
5kvS+81Amoj5fadzcBUq4duBdJzuD3yzUI+Bl0nxUiVOS+T3Vci5GryNO4R/KDeQg76zjtJjfwcr
QCXNERW6DKCw8Q6MJVvlnF/CZXW7qXq3EqJfav/xaN9kfc3FoAzZxlvXAs0KSoW99vyiLvSxL5sq
mCFjcRCN/14FlU5rhdYpDOOE8+1jRt+bMzfwvFDC8rpVhvLwFaiC2j0jdM6tfoOahztoq6Y5iIwu
JcQE2Uk4HmMx6l2Na6AKhd2smj1TD4muJJIg3waet23D6V4UasZ6TFC2ktKnW7ShDLSPB5bCl2gt
q3Bu1659qO8Z5SpUsixgsn1ESPN49zJBo41yqHo6eJFf/ReA14T+Yh17wXZK/Qfz65kfDLOfZPvt
w0+SicZ5qzlqWMpIk5BjljquxgEGwRXuW0RiQh6dc/u/kglL3CIYYBiRfgFZiLds/e+OPNH1q62n
oultWmpE78Eq1OMp9LmWLquoScZEQ1+DH9uho/eZ+PgSs/21KTw9vz8qe7DQd3AI6auh01UNfPky
/oQvKgKcAq36UAMgF9/W7kpfV/WmQUWF/Wh9FimZ4OUI3LRpVUUVWNtyZtQUAgveLAcCqcY1Gv8r
2934x3/Muh8b7iDF16b38kAM6+7nCWtcrUBiWiyAupSNlUq6qmk9eMdCQW18fMxzv2KAwaCKtTE4
JmId20u3TZxhSIcSVu1CHmH5krNTMn89sn+LD+DSL2oxgbNVJY/k0OJUyOODh5zmXQldn7y2rtk3
cnQY2ZvPUPbrmIx7H/8gYCKTPFJtgrCG4+nA/0DrnuxtlGjdXWva3PFl21+LgZ9f5xHVVfeEH7By
EzhemUpe8J7Koo7omGqWwbHR2wGEgp2XoY+tHJpVWCyylsrZ+/gAQwj5UjRjj+BAodR8NkYuOPgW
+DdyNivzlax2JdgAxptklprfr8U0jQXuwp2gNTRbd0IGSjYCt8kNUYYQi6A9ylmMQX+pCypQdVie
YdocIxf7unRw6nAoov10h5OjvpwN/tRYYy0hqP1xoJL2+tNvsAxtBkvAjyJtc4NHZQN29OaeVoEu
rV+o9aHcbxro46TTsBNB6yy7nP7Pyzh7htNl2einGcSAYSXZr+s7VVeY1FKDy8BTu14DY262p7pb
0OqPeAdT4EkquxI4xkhkNraB4Xemff6c32f/o2OEKS047QPtFrW7F49Hz19TX0/T651/puDgRuYX
3yz4vzRLI9rnq7tNdis3cpgkgb7lh9yD3xLJxfMKmM4LxIBtm0QlVZjaPQiAa5gOdyVQVcUAq66X
8L282Rgq4NPyL5JxbVzI1zmt4LjxKlDPsFphI049Qla+TVWW55Cf7u7Vp1yvs0v0uEMdfEKC+yMy
zmu50Cy2qiO1yI5XYgW3C3ZExSJxALWiqhlc/uiGQRalVvvb2Z8aLVq4exneI3R/tSbamnIuNL3G
AE1Q4oPb8D8sbF0FVc63QIXR5RVs1Gf7niiMj3u+PuxrrBiXoPVV27NbZuy1Ai30pUqoq+sshJhs
gi9nBt7mCgf3hPlM4KGd1t2YPyFEomgRnGkLpKuGcIk1GI/qAfimHeOUgIuvq6zzNE1yhaHhNgWR
4ZrM8AOxlycHPJUz9SQINLuFpXqcGfglQdfybRHUiZDOlizpr0i0s7DANntPfQdclGRgwBTHnpJg
z0/T6hipfq++DMK7elih7HuQqV/xbHjYPKItoLaO+lYiMn7GQ7oIiQgnHaJyVEjOQ76j+/wW88RR
FGTw9bkXfPT9VuLcdaDGaMe0t222dgfKV+y4pwy4efx54hMhzhGMpawwOAJmWMpxFY//aB4zICeQ
E4vokgd5CAFzDr6JHuubIaCI7ZjgnRxrFjix+ydc8EckSOcVnKOEj0fCOLlI5TCk4I+NqfhMwPF7
1eiw82pqjk5XPZFnbIQckDJSXOGqMnpyDa/2ladvUQjed4NDTDtEtpBWFzsmyblcJAFk7dXjTEBG
6jv6nEZocE5Gb8YdBEQ+xYkc++BTmU7K0eK1Q5QEufKjJw1flf17DVNZJnxppl97ldcTgPJYv6z2
1SSjjHbHxQQh8dEQV3tk8RgyC1iuPJ9mObZ1Jb0ZAT/I3wRjWzzxdjUqv1okduAqIGVvBKbZLCjU
KP6nQvqwd8Qj9MQLT7d4GVH+kuzL7FmCPHzQ0jHAS+PgVdy1q9e2VqISY+FmevZ376G7VgmURpWW
InRH4NwnYYpvQEIGd+9rMRv3nIDzkx6a3lwzovLMWvPyAvUgdAjvZVIgUXlF2A2c+8YII8/kIRUL
atyaQKyOs/qpC6Fc/8hySNBQFDPSU5NUtWCe14okkuQ2Q7AjuWJo7o7TzEL2+rm/WcdVupTMqLqH
GtM620Y++ReSsDDW04EYGNll5WX6Q7qPGyoMgq/PWTrz3kaeOWDE+4C5AIVDzMqmFfqZnwTpyrcZ
uXSoWacYch7K73jXTshvDhEyQ/ocjLCKgcwohMw7ewlHvumZCIz3bRXR33E89V2LHeSF/Vx7QwIX
x7Wly+Wr/TVkOc2TeC+zqUDyoHuz+tYTjKIrJpTZeIJLdSxXIxXDbODIFTMr7CYp6ghyciNnTSK6
+dd3VL9lP48D51YiPKWoMN71j16C9ZtdDIkSlAicHwne0I7v7/Xiady4EP1esDuntGBqm0afCym7
iyH1TXQx5KWtUNAsINrN5mKKhQs9RKMpr+Ipb9Yuehfo3MRRhOLTKxrJD6X29abmBON+n2XKus8z
rV1LoW6BF7D/TIrRohGtQovafu6nPT2B+zeFD1yc+gIgbjqUq1e34JajD/yFFTuEi6uKS43+aGvG
dRrkgGV37nCujBed9G0MwXHnfHKWdrjztOiT5+ViqihKtwMU3FnNHd7CYS23LnDrk/eeIjOJsE8L
CzFqgQ508ADckxW2+V4N5qryk00Xn9Gdya2PMYQ4aRmOJiSWLHdQm7+o3Wp8tGQMIa6yqdKi88du
lBDdv0fWyYXPojCD7EAxuoK3FA92GJRki4I+PmeCcpIA+XOrDkdiFDs0xtiYqAUM05fXmeNZp8oG
CR/rWST7hdw+r8Ca0p3U/70KdN34X1nMYBp6RwKxglJahxRZTou8JWVmgHrr6z0Y9vG0jgo7xOSc
N2RDW+WAAEyRBleEaoQca+bmRcfUnf/hGO8HRB/GjVK0eDSVNfnsiIKYzgR5Vbs5gph4Icro26yk
HKDxsFHC7avuyLZLD+Cg8wMsY+J8vLLCZEDtOsOFSarlT2i7k6c3Zyn+6Y+Ov41O9nDps6nyiqSM
qA1g3tG/N94Bs4wLGxF0DQky+GDNADZrPAFQVjnOV9aFeLHYrsJnSrbneSIkNbwkDzMkG/QtaWz6
tDV577uC3+SgpidmxrDzzOvCGNo8unQ9Ti7rXsTd+wC40fwxx+mTA/caKuc22Z8/mgmr58+YOVYN
6NhFLHkBQeSkUhuccPRN/Sm/zE5flpALjcPJmh8XMchkaVhRYPgt8kH85HNcl3CjPUHwYUErydNw
vQByP4hA96Ep9kFRcaEi5gG4rdZAGUPhJt65W0Ow7GlDQ0qsSmWk4mkN6B2ExYjXbHBZU1mfxexm
Aen1P25xbdWm/frUxYX2p+Xpxlc2nsKRVaX+/QrOsee9I1WzlKLkr+myQi13qwThnuYSYxL0k8ue
3PHrfQk3NUtgeEcgohloO3njdqpXSYXDB+fMLF8jSBw31iVeTnCL11iNAEtFWLoMrbwG2o/Y0qOW
BawQaiUcU0dMu7/l8UDgxU9wuciabqKQhv9kbKb7lSd4TqMlXdW6aW3gR0F796OGTH0v/YZTXfPX
ogt3W2uER9cqRmKnAbQ7BQxvfNvhrp+Xe0JZzSe83xmTn9b0RfQE3bSwqGKcYzUjBwHJAUruZKtv
WC+QoRiW4KZ6hc9sHTq6blS4u4LpWGifg/8gEX6gjctW8P5tNPjcd+uONykXqM5wKeV0KxDqypD8
DkbWxUXTnfoKHHK8NG1+4HC4txvJ+KX2T1XWwP6LG42gJqFV8gDtnRCM8uraWmnkIhc4yuOE7hOT
2r2H7XhxAyk74ya2YaYOXQg138Y3FUI/0BXF6J6IM7pokz1XDargnf1u3z1sQfUpwTRQ33cxxUHY
fYV0wR6smpC62ZgK0cCb5Cu01JpiyL07TjHZcWkaWinwNcpKmmETmDprfJcwiHu58v+EBINAw2xZ
rt6ikhszxX6quRON37kV4f8nFFcDEcU0CfvYK3k7K3JiFLUkKt05OkQdWhmt2E/oh/MLU/9zkyGw
rTGuwN4xVRrefwLCIl7je8bklxFsxZ52c8le5skc8pROZSLbMRfxEgIZKd73MiuHnMF+2DB0W8VW
wUtB10hVPg5cDk7zdqDuR1nGJ/yEAFKjo5xik9rzKiYiDO+5vbklILIrcpFaKAYT5r59RxPdc9qB
y3lCxXRVo/BPVYRxbAD2vBxoMvxxHGzRdlDKfcp+4iHvprNu7Q2HnuLk8DlS4LaXOIpVaZ0B/xHO
XPoF4ngAv/2fdWBA0E4bCmxVJvbqgMqEQIDV8QC9l5l1sacFAr4pXMK1OgvRuduGR1ku3wMeBeyz
tMxST1EVKMB5y35gRpZDlaVPOlAJNsc3gVyu2kr1qMFHop5886SOgNJYC/BSGKyP4MDk1j4dCmUg
dG51NtGMi0kw0IANuIqVcqRIgowXUiBFA3ySYdyuMoGwSnMGj/NtWRpQxbknEt/+Heg+hFXpXIax
EzMOaO+v8lP6gvk8/YSH3aQwzJTzRnERa8MYQHqerLm884Y5GwDEv4zKn6Qeg4loIgbjp5XOTdU7
oetJU1G7dAw+ufreZP0AoJLx1B1VpB9KwOI0a6NMDdEYCLasXX1gblme60Pr91gL6RztJgIpPhp3
iCqVA6JEDjr0MISs9hIoPZS3AAmg3X0nbEb38OLOAHmz3pCHDjyEXtsPzmQ+HwpRhepH61onqaQI
hUnTJ33Ldc1pURakr9VGJBAQ3P4z8W+oQ5KW5AWPPErdBGWd630gQ5EuvEnp0aEPhgh6dWYaiPr5
TKSIURiungeLWRJGGjWAY1Kw4bx8bIOpzFYxHzsZzbPwL+cQabhrgfahgKXPCjLxCOb1yoHHnGjc
qSNPzQWKnxGrhujGxNcn2n1I/OgqH986Dp7wfsFx9W2cfcuSZ0iMkLY7cF9jWnnrzDLazfzRn9Zg
vsrlGM4FXKNobDjEn8RTnK8Wxql0ylOo/+m9ilmx/3xUl5TTp38KFNqpEcCGwVo+L4f0segGi26J
r/gnPAxMxLhbnyOp9v+SpNscVnLJ5XGCEhUAlsFgmOde0eJtApWbPwL8D0Dj/b/w9iMMR95xGlxN
LwcT8dIow1Zs4Rw8x/d3yezuVj9uJGHu1BoU96brQK6LWC8bpA0Yd+TH+iLkTRlYfKTL+ADUt6zk
qgoOslZ1y9N7iLReL9BJhAKW7qJJsfZX6UHv5zLA6X5KNwtJ6J3iaG3eHkFfQqt42IYX3FFlxjm9
oPUyPvE4TVctKyXSjm2nmhp782GmP/aJt4sSNwkLou/sDc35RJyQCQa99fZE3qZB59hcVHEkxwWp
cOVhU+OMjtskNNhPlhCEEEF6Qgi2C61UiwoNskJ57Ea59TfwKGvBOyXsLZfEYgRhcTIeXbHWsRZD
qixcFRRDqo4DysjFVUNn+avcIf9IIFgrtAuQGJK1jMKWuGwLGzwZs4J+vWNzKs8j9lw43tCk7EGY
s8eYJQixDt1xN/Flk8ED23XdgdABxGtmiCs+QqthSOTtZPUg8jQ4FEd/VNAQ9AuQ03+MaR06x37X
D3P7QvXtOUuz2eOwwQaxc3mqNbSfekK/9jhqzKxZtnEJmazpe2OdbVpnr1lh64hNr7MAbSP4+0UA
TZabR8dsgNMtU3SO2+LplsOrqwvYApB//HKL7dCZFcoTP0u7544JZieKDKK2PFAomcOkfTQL1OJ6
lL6ZjZRFN+ou1EGms9i3GaGVzT4I3pBpF06cR9Pq3z6z7Sf6gPWe6EJQ3QvrPJOhRPQKSFhK0hkg
bV9233J5JpPP2CPI1IFUqvuikST6DoVqxMZbnwl16io0AhPSSoLySoTLG/KazQYw1+1ng7KjOcMy
OE0RHgLpJ18QeyeL5z24qj8kaOFpN6RnLPTEK1SjNEzOXJK+Zr5RpCl5BFdovCjyX2idfpMyqlrp
5aFmKE30NVm+SKi9OgD22FGYHdAH42Lv3p4BJXAVLxP+j1HmlUwchOkyxZU11GSm4ZDseIuk5WyD
k8FRUx8pGOJ+JuXfkeGJhVOAKZiX+h0/lp9J9+pO2Vp359jw/gS6UgAbXrLS2UsDdWz4QuF4IkQU
joaNExXLuSHklpMmW0DHcxwDIr9lIsqHdmvoo7uFg1eWRmw9T25DD+yqNtYeW/rrTbakLRYleG8Q
kAcuzqW5EKRpTVqSiSul1QdxmGTDE38IP+/fZBgJ7jjJEjzEgHetE8jOgPQXF7FKOSl2TIU7Bqhu
F5aYt2vAKylHtcI5JgHZgCK4vg7VZKz61SL+oqJ2uZwyUVihn708EUCLNQNKovu2Bkkq0dbWYFel
tON/+HfNHQFY+y5gBpyBruBH8rIWV6SrQHAPkqc41NyGzaKauV0W144jJCgQXYr7djZDiWpU9YD9
QUq7CRFpF9yiO1Q8/tV2SF/yxe5zPDxjP7RhcdgcJ+s5n+9tUhvqd29CTN00tT86PHn5NpjpBgrU
UtCWo8apIb70iYSFIfZ4uV0qC7oN3o1O85RyLTonc/ryGxBmKk+vM7SgUtU0RDgB8dDS6p08Gt56
ZteV8+7xwn49cx4px6FLSsM4TxiUsQ8AhhkTi6s/ozd2VZSQISrhAULwVzpLiO14HAi/X7MEOm6r
rpr7AFiw3bSzlEwBDYXEGb516n7QgiJo/tTv2SzxXvQU1BbsDlcuPmAVRhPcMXZY5F41cY1th/Hp
vr4cwE2/c+yQh0qAgre0FsyoFs6qliaRb0kn90W49BChZcduFDzxdY3979f0H5luiE6TIlvoY+P+
xWTxrGJIOEE2oD+TGZR0MpAcXX5onxrAN/V8S4wtbxrCpvJTBQwVAzDHe6XRtPU7Ueycp870Vd67
FLNdpS6fmipnHJ7PZbBLmbDcnzSXrFCsZAUmC5aUI7bexXY7X1qMPciiFJqxyGXZT/Cu30Q3R9WL
vwSMxcPvioki/ZNBCzuZlOULsTxuMJuWQDwXxNU1EFwMq88tV7yoci32OLR9JWfnabLSOyGT+sZa
wBJ51lomT88irZe5PKnFs6mkW0NRZME9Mgp/AUJ/rEa4FmKxXl44FegGffV+dgAYTFDQ1E7Mo7mt
7KMhQ8fIvBnE7t7YZ+YN2DWcR2ApoIo3iyLjmdAGQek5hsN7md1pC3q+nWDUXvoV6IcgpHZPNCXa
ReBMZpX2agqCpWDXM2lVztt9lDqFkQEVGDRBSxUV1aZhfSZYuV/MjGq9bOhl8bZf+OJ6uhr01nkl
sQ1IHJAeeM6cjpu/L1e/rzpeKRmgA+8xkZ4rl8WCmjJQJEBOJgid3TgabNfP9P4uyTFYVJYvY/Z8
xRFZsyn6lLAlWX1tu0ypiGi9n4yg4u5F1gFBFfAx/XkRlU51xBQ2XwSw2JTyZ3gQf/HLMJmsrpQ6
ofnfeiMS2OxMr3f0igzA7aWbCDe0m6BAL1h9Iv3zg3kAAY+1wvjNKynx+xzVnybjkjElua4Bjiz5
M2uu1PRODX3f5QxXu5/ecAHIlUjOv/QhjZkFbScQZWq92EGmc4pDxfh/qZ985BIAp/c4M8/8TiT8
8OrgBQBPM2tOO2IkakH1X73kjTxLppBEZqqKh/AwPjLQAxa7/qq2BORH51kcolgpm7Ypx8p8Mjqz
9UHx6lDpDXJlYkKhfkwSONmFv/qey0BiEtlcpzG+ta0Vfze9jVZ+f1SYJmvm1Ch2WJ6lP2Moavpv
0b41hhn//VD8w1arJCdHxnYORriX3p67VvOHQ2nKQ1NJJO3hTJLQ9dRyM/URPWhJH3iMMskvOg5w
M85nzOWbralqPnLZfsZ/Z1x+xJ4NOH4SubgLH1c2G/WKwgvhd7otN7v639mzdixugxk4+yS+9BtY
SjhCu+8FsGCpWKvQDuDyZKQHUa5HoE32CpM1MRd7lHlyI74rtBemVHMg6ULszHbP3fPOdMBkwprV
4Vh6KNiAh0A9E5HUhjVLpdkbULNWeZtxpIWO9XVrNrYp4Gn50O4UXoyG4Pr7rRtntxjEgref5cZR
fkmM6XxSiZTEOFPoQHhL6HIP8KRqnvtjjtGuzk0V+G13iwaCDN6myo1CdVAxLsGVBNdirovJP0cF
p4e1ldnK7SQvTjdHxo+dsc1LPtdTBFdMSZdVF5m/YM/SNS5MjaH31/loqnBQdsx8pj0seMWcctys
mfWbSYDU/J1xcecGZXO6QGuOsVSHPEYxYd3GbHh/APdirFx4NovhbXYyz4U7a3iQMunixwVmbp3G
Gx0RGYEocQLAdQyJF/c6OQcOm5c2nuuJGS+J9iaNqeUa3sezVSL6yuh81svYuUTg8WJx+rFHigEX
vnEbBp7AM1GmFJC7RY6asSXWbb1HwIYSmb66lNj3bepzJ0F9ED3LZfvcN9xLfpiig19//AZrxolw
qoEWuWagDcNMKjl9y/avcqmWAGhrwbdNJMCj4tK7Bcan+9KrJAkv6JIAQPzsjyRYoKo30QVTeJgn
UiyHjLhOsjAV75IbXWkTGfu30Z++U448RnfeTiSjkQ6pWU3Bs3CnrNEd97ITfOjrEE69YQXgsZP5
qvlT7GlDfCDMRXDdyskroM7t5C2Gy9Vn+0sFMmRtphcx3a3wppjoevxPOlZDjvvAH3oMjIpzGFs2
oKUAEaXdqGlsmmF2M6B6kbxYUhXmVWg06F072iyssL88ihimQEl9LgEh5rrv3y355f6JY388uuEO
Cuq8AAWfxxxqOUcYKRZJR7ZQ0GuV9BTeyU6o0XQ97F22JsbAAi6sSUAjxjtpzAVNvRyKZm39opVY
YKXZXDgqW4Juo4Fu8BWkjhy2U5D4KbW3q/SyOmDu1CUHPgMCu5YYY/ZMMHAbtW+AxLGyxObDE6qO
AJpuH/B2leiKmuScY1tgHhZKcOL3KipHSXo1XT+j2zNCD7HS1xHJ7P13edqHfSyLJKw9JtSPP3IO
dMGOaCtcdD7nqDIyap+TYigSAfgwIMcy3g8IHQp5Ym1RAMiFyt/EYKIC+wJOn9N1MP4wfbnYz074
1lo3JNJ51vlvejqw/JfLmty3i+6KxpnVcn8qVJPpAHYacL3daycBiEcNkVZM6AhwFypWzhb2+TyA
MCwYZzRFdOvWEU4p0Cr5DVzaxux6tceR8wD803dzQKPQX2j3eGxnv7G871g0YeCUO02dE2RzjgQ6
UaKKYyhvL1gWhxpmmpL0U8mG1zee8F8S4FNL42O+GpPV0fOwZxEchMY2tssRabhfPEqGc4Lv+31e
Rpm/BuuIEHKtcgqkIa8tUsKNpUIwgBZqr2nqAAap0RWBPDm5I42eL0Js4Ug+/OplxhoY49U4vTpO
izxAZKT8cFJ4n1Gyr1XnA7ePSjJKlRGDa3F9NJgoyoSOAqf1GbLdJ00dYRvaguUVKhaMISv3IGYm
H0LXL5dWWvxAr9Fn4GtKQ/bt6c5QY/SVf0XpIbcxYQWKJpEb54xKvhuFRpEDKla/eWxQwTwIAZ73
rKgwKzNYCGsPFFh/aHdzDNNjduqCC59g5HL2F9qIu1nPDf4w2eF2ssTcz6ce5fbco6LpAzCEbZDU
RhxLwXdw4V6GF1FxZmHRdOmcirBKa26wrR86XSfTh3NIMMK/ygCB3pg50doCiuGGVb7gTzR8ORFw
QAP/OJ6stGNh8crPaiQsCHrBy/zUcR33opD6EHRoNLuwjKx/p1wJAsu5cXHyDufNEIpxdKdsb6hV
nZ2YfxaBOmsbxOZxbIKR6Ei/cWkLK13s4irz0C52UWlq6VmKkPAArd6xGDAmQRxLBhSrFPnAQdjf
ARCfaU9IXV3QJkr2epJ9LYo0oTSG0Z0ue0YV5429eFVn+gmvuvNjqQ+2OBZylrYWQGHrz8K9c1IN
ewumEc7VZr1IyzwG+omiQPghgSPrZC/hXOPARfUnn9RnNOCXm76orss+yRTLUKCGW7E1hFykAHnx
q/WkyfuxsA9G2LLlcyHSxez+9sHVhnz+RfjSK91DzCMRDNfRF1BRc51o75k44GJX3O0NsSfDFCCg
8+P+BPklJzy2TWGTgYjI6oUcnONoOvHNftO0EAVo1d7bg+geelBq+7zT2uitWAPj/BifQyMbo17e
T8qmLomMGvgGbDXWz2a+996eg9VloNjxDzp8Gq1WyBOVdUWYbqy7w2NeL/Qq1uhYdY6SPpk3gyOj
TIdvYzyrTiXo7ZGIfjmc+GYCEo+tVSxDC9lcy91BLfbHgbUnVq2L+xZV1BguRDxS2S4zLzvIf+OD
9SKQpTFY/4scFG1R6B/PbdNQ9xfUKWxYYpZ8YlKetJIK/3YkZmLxubCWNKF+G26ku4t/sDl67QH2
h738o35To6v/gz2wrTAyKbOIXMA+IsbOnXfJ4AHedc/w3vG2zf3J8Uglfwtuab6QAYjNJ6ONvSgN
hywHhvxUsM67BgRz6XAUXT1lGENndXB6AFbwp71FfcF3/y3L6DmkYvXbgBlT4bMORBEBaLcGYc32
okBb1p771oZ0uEOaqpBXu1nJzzIyZ0E+K3g/2h7Ck0wVl10qv2kCe1/hmcMrTsr4Weg19km7vHfk
OVliTIEmJTOruYG4+x9Kig3iGeavOofr5ctBtOhY5Y/GplGJAMgUFgM20jFWe0q4ydh1N7WC0V0g
N53VJn56yt/7oDywBKRTNRzfi5uz27DzMTC1Bu6TqKjX15JHwJ+8nNA4QZvLK/sr86xtj2Zx8V0m
8xfRN9ULp0I2F0l92bg0sA2lWECfSqR9t+WP5zYMy6AwwJryIGZP+sL1Bvsva86Aqljvc8JD4Jjh
825oVqy/WjfQl5NEjc757mWIsAGXdUNP87GMmytZyt2wDbxyP6GZyoeW2V6hm8gJ3iIKiYeSeZQG
9XsasT60rlTo9EEiBfFXC0/r+lrIKPp2UvEF8xLSv2oz6Im9LiaLNW4308CrJL+i0wvJZRqdoc39
znlvuyfQrS+W0boogzm+NHsUGJ/QnCuYedBqnCFYOy2twOwmoprXHF99RazDT/m/PIQNDb9JYf1I
cQm6gbtMGjA+bUKmcoN/impqE63EX6siCCgkx6sP+KUcwE+7bFIn3nqpQSAmvlB02KV7Ax5JGO//
KiNd31xxBtJ2dDt0kbpl4ntoPddNWTB2r9ZhvPUJsQu2GRbDmEO+ka+8JZBdj3/fRH+dCAJRxtvG
FvEFWt4d8cV0LpYgwJQqCR5EYm9Oi46cpAaq2LvToxpl5bOTAKyWMT+bCZnySPBU/exjqt66PoLa
YoslSngwAYwnUUgIau6Ib2Khp018ohC/7sq47bdjIvhOM80HRn+nYyN3hTjnAkZ11goYJzGpBl+e
4m951OPDfBhJVi03BUOG3p4yxCnmtmfhHrn2Ot5eMmBXUgJ454r5o5IvfmcQMOSwEfcNSQhW0LDz
ahF/+NAcvEZPjAM3gjonQubJEFhWPmwd1Fbj/zKzTRhxxZXtaZ/fH85Nsx3vlh8XcnUiiyrIl1AS
CdJKgo/u4OReV8l5Ia+ZL7gIjEDSTYvlg20yGanSBUN6B6byxNeLPbUIFdRqAunFBPdqBWUv2l9i
RJCan16WQk1diakMcRAPoPreTrg0RdAb2GaWqQHSDgDBZ/mnIfdERDhlUWaEhKBLb5qWFKZEG1DO
gTKKDEFtvNwlWUOntGoneXD4JJdYKC/Rxz5YTSnkGe6VpWW4flKIED8f2+p8lZ9DkM7MBRTZNG7P
03U8W9Y+U2mGvqy+CyVOIYXD4jGyu3rMph0WVg2ThGcQtMtEXOcstDOdiTzm1+zpzgz/5OvgSX/1
OJ3IV5K0RRkFoBb7ggLsTZ1TGX6BgzahkD2ta/bm9yAGQjjshXHnDaxe4YzRJhvVHnTzQM1O1hqv
tP69lkv7HlqaloP3qGmPF62I5HUL7ly5PQFcJWTBO0TqEqhg5RLGYfW9oojgUHY9qcusN5hDI7oq
MmeWXG0lMYlMLX9Fp+4r75l4NtGihzsvxNZS7jwfROBORrZy7Q6AyjAwhgrZM0cC8yOcj5uU6CKl
DACKcdK9W0AQp85hSlk6vudaaHBnPPF6hNoASY9vTqVDVlrad55sP1K5WV2Tva+X0N9lSxrtmOIF
sYOhNr+r5aZ5CWSKzKP1a/yAz+7Xya72jF1yrvg1l9FAKpaJKJF+cA6A1AZBci6WDwscuTJIfkAm
5FMAWmwHkao7m7KMG3uraEYmStniibT3m36mL/hC+CqSWVZbN6TBztXjALwJF5+psY3PsNMQc7wC
Ky8JY5QK/iO3Z0A4asbZAZapuM8gVE5irvt5RiABJMLcUpV519BRvu3m1Wm8LWOqRKqCAuuOaZw7
cfrUx7jXSHpJ3ySJboDpaw7EoW/uSpp7cUYhXsEhM5HsQr+MBl9PxnjAGCe7xSmfUY/6zA/BAnkE
oJrFfk0p/DukDOah0sH2q4U9wguis6QjBcikQzivIQYG5ho0lGzIsWN/Ee/QpmTKJCOcG5mYjrJv
us0XBUJ3NE9Krva46FTqvpsYRFfpxMjghHAO6uqDgcHMc/NtZKQ6yc6ZLR+xip/Uf5rywxBz21zd
qI3NJfwBVQse2wupdrV200tmCy+Dh8t9jpPdlulRt2xXob9VwMm9hrr3II/Vru2sBk9rA5Pto/zN
FuQ1e/WyctvV4olOkkMq/2ByBlnVYj1TgvVjtKRYZv1joEb6XueUBk4YlFwszRRAwIZoqUUgIXUo
lP6YIFSK2uO0WARbs+W/fYmNVmqH9Shs5JnA++mlSR2yKiTZDvzvJtad47whSCF5U4GV8t9SlUCy
zsetSjtuEJEX2JM1VXwazbC09VpyJvI9+sOavex3r5mkVbWDOajLqjHMg5QTrEI/+xgAVcNN4SDU
zsAwuwJ4zSYYQ9Oo98sUZAGybFSMlFVFjQMB+sJH16hc/JI4FeFj9+UMoeBLqBcPNudmIvW5T/77
O3pxagBssnVImckV0X86Bmmv6cci4ixZAJV0MEB53LaFUy9e33Es1U6GKyw51Dn0AJQ143gEb7wJ
ptyvTTJAqlIsZ1lH/kwP2YTk+o+Rlz3yOb92e1fzQHP9S8RIU370H0SWE1NeNfpYuCNktJv+aUuY
iT+14coyVL47i16kMK/rq0w9YLTncteDMolkynPGf0Tko+SP7jMBCp1NcZmrej3d4+fizkhUXTgT
s6Vcu7DkrmHnYmY+/HYd5vZiQmdpjsUSeA62GCrmf9beRQioxqcxRSDD8ALTELuG1w5zH1iX6t+9
MhZMEUkEeZWCeWeQOFGQmstgknDX5r/1ZxJCXYcXmmlz19Z4ZQbnRHWgJM5Gv2mqQiP56AF1JlS0
KBa6f4ZWTeuqDbkUtNNahlUKZd+WHm92yxqOXHGCghggI00ygO64Qs/ce0Wtq0liZz8cUwo4BY8z
D9MTvMWqAfeucDuxPksZ8KjTdKJR1Wd5V6WQWhhPt6IMjlzVzx9FLsHgLPC1IzHduhtELrDX3O30
nH9RCfq/8p9zIiCpIb+pdcJ1akgx/vb7nGtaQ/iqe0TQ8XNtbTQ9VEh5kdXNlt6zhNWm28z77XrN
/0jQhISZywdUrunRGbA6mExxh6uqpwG0CGCKhBGRnp1WiFKdF5TmOnZApGY6JTERSajXI+Te/+N5
HXiEFbxRwy7KaL2UKNOvM95rVVS1wPbW7G9DaNFBL/bovr2xGKOIZt5MdFjXqMzOhpj5LSHMgDDU
KcsCLgMKOXXM34h/1sTztPZRmvA9DHhx2nvCLoyP9AA0JL7M3KWOaFDOcOMMV7I8j7+R/9zMnUqr
Y4rK56k3bbiXaHFfJNDG9b8edOnZ6yjJT0Qq/YYoLB86lrKomenENX7ufUk03OXUIkA9eWb0Och9
xRRtbmQRRDH/9SLzrGkP/WkiSgjBhD5kqng5CwJ8prdrJRjlS8VjRj6TVo+7hYx2VAcffBHh46U5
n9WOfmnylPIvZrjjDXNmZPFAZ6CFp90FZNikw2CR40IF7dZCkpWVKBWzSNIzATQUwJWhhNWX7TaK
ZIEs9WaB/xMxibY7X7DHHgCHuK4LYxwLTJRHrB98C9N2a1AS0fXxp/Kk4wh0OH0s7oc8f4wsogWn
qhd9Dn/bol7iYszZhSb39eS+ENTBy/BCQav9WX9z4+Ex6NSn/gbmIyKIpch9YLBIFQ3VhthhcwCn
3fOsWtDSnQzk9QYD9I+H3dngZJo70jD43O28aU7WgjrVXu1/jti+ZbeyVg/UcwDqlJmqwr9S0Z0j
sR9UquxHCJxFmosb+45vYIgb4f86vYGk3CD5wdPzF7Q3+KlJbdelxnqzeGvxpod5h0aHn5DBs0Wm
TmOs68xovTUml7lofOP0uriVxB4TK7xuVQTk4g41ikohf+9d5d/3y/ala2Joi27cmWHrOQeapRmG
Zr5pwdt3jq5zRKAqqz2HgXNBLpbzJ09GXERzQb35CfBryk0qXVaPM4/3ILNBFOeLVNDwXe4UTUvi
96CjoQFyIewtDXAcY1qjhhNH1uxx7RhQrY5Bbmwu67FNRBjb+kZHJ5a0n1riAaAdVQ5reh2k4K4o
+OwJHiSWB3fDq2Kv8sE/tokEQx00ois3805kifA2ShYMz4MYfr62BJ2RurnKH+OgttITmbL/6pb+
w3X41V6jMIU3X/ZB2QcABnBwzVdNpy0mqJe+GVNcj7iIy+UWFfcFFwmj5dCu3TZs/5Xwh0IQ1ABC
lih7Y3tAdKOjONfvkncgHeTpgGmb6Pz2X5UDyCHw4p0CMwGglTpif56qA+3AycSFDJrdBHFrf/GA
V/lY0wXr5dLJPEHp1tb2gmMOtsu+60c4Uch3F+7TxkIRoDjz8ngCvQ0P8Sv72Rc4l4GkfYJpt7FU
zM7l9OdyyBMqM3w4UzWnamDWaY1+e9DJG9iGcL1kzXGuLifoNlfHgCMHbar3sY5coWYzGl8/Gga+
9mFd3aiXCRC0VEPBtECzCx4sVT53FhBlpDvTguevqfKylZyRQPpGDqthOxV2KcEp0NxZ+buBgEg4
Y0H3aH5GrSluJ9tJD6VsGnQl94rA1J9VI+9tlkuAVqNKK8GNdTERrdR/SKe6ScTlIkTymTJ+2xKs
O9g8rApWCuh8ytcZfygPRDlCmWaw+rJQAilSzCMez4CbJe4m8VdQhIMJoCRLIvkYYfzAVVqMUJBX
0YBnW1AVgeUPu/JgmsHbbidUJGgwSdtCx8Ne6mBN5lkofFchGsU2Ntky5hSnAa3dh0s0m4O+UYeH
lEkmZJKw/x/CsFPZX7VGkHEP4Fcgroj1EKh8tD4lqvM4jwUAkEY4cvirBcdRUDzyPvjia2gE0P8m
Nkn99INDaYeSAqWN5ILATkt77KpnCEGCT+UQrEq8hWD303I2YVvV7rxVFRVjQ3K0BUYKI3lrgBJ2
xQmhjzeVxt0ew6QNgSAV1QHcoXAflTAgg9NDptEnU6ICs5UzZVC/19U/IZofEnEDkrWvOs9Yv687
fNx7ru8j94jA2YBSs1eqRIFlWMNfdHCnMX45GD062UgRdOK3t4VgjLaqqYHC2T2Lopb+EE60/uga
d/WCVpLbV2ERvlv+Xv3qxKkZbrN6kqvX/1WoPY3HlfF0DLqFD2pWvXlhOJ/Bl0/wSe36V3K1Hl0Q
2ehbzOfXdwI0HNDJaHmGziePwEowVpCRrkI1Zw3txv8vx3hNBPG9v4UmNajhAz6xGD7IDdq7pon2
YsfY+j/G7IK5OX+2YtZ+q7IzzG0pFYQ46a4l5hLWq5V81Hj9Psow4I1734Sb3UFBACHVrYEpJx1o
7MCTasRFLrg2xmX+otLv9k1Six78+rTfE6lrD7AktMwZSs+ZgHSnSMe3tNbDxjZjloK3ZVgcpJPQ
/WfoM0VtPvoqD3bLlD3V8eg+D2L8w0NyXGOaxNdiFDRbKDCh69Yu9hfBu2sHSjWdIL2L947AuiYM
pObbEzE4v3QJ1GHKS5ZripuL4uJ08gytbBxiXmcBTHUokqe0r20dItazSrJp0FJhA75HHkpq1/dL
E6o3ATLOvZ+hUQWGv9qlGtjv3ZkM91W6eDCeiRSlWnOxnaY6TTn1euBn4n6OYG53qzOT3RC+YA1n
2sbW5iJDBTMzRkMeuMN7GRApcKmvJk9q0l7pu7p4c+CuFCCYdwn1DuT40LOIMqDQZVfGeB0fhvvH
Y9g10MiVPva6xlh3v3Ipc0U4t4Y8E78XhwyNdY8XBoa9Dz1KI0eeV4x1vMVhI3FyfJWM/+3Z9Y6h
DVFZfBTQDKCkncZAYVh8MGgGGe+4tLjKCLFPyRchdsVM6ZcOFu77iNr7f/6k/WvFI27TL5YAmodw
hNicVNlLA0x6uoWoRGLb4S+ioKeggFrt8judczh4uDRD3/XRx0CkqQZfaBtYa84rkhGtAwQSNt5I
T9hfUoun+DVpCfvvNY3zjnidAEFyFalAeoaPxQrCKR2bgKkvkZinEv3/QD7/zycfs02tvvc236fN
cd4v2rbSforbcu86LmEg54rD2mo6IBlUg8R4clBWkScY2CkckSfVF/tpIdGvJ5HTTDtb5YgwB8ua
63VQgYSMXxVFpnllRGlWWNLrB7ij0whXJrtFPpJEBpcznzLZeuQ1jRwU5IwEYyOCLj3i5BSaIM9D
9KOs+I752ymtrbYCLODmgj11cH8Z3fZsIEtOllC+aEtWTabRA8ebc2i8tSe3YRRbG7PO44BP3BVo
7TV48ZaTREHioIolpXL2YzPIJes9LqRPtUdl6r2PODPJEQCbNGjwVILgBQ7ALDslcKP6dfZeV2Pl
C7oRm5wrxSnCgpqPboKudY71eBNkdrNsHaes6Jf9TZfHdJQEf84AA7RpMxoS1OoFc9I8lnM75IAD
czoaDb0sbmToXhWH//SsV237es/RITv6f1K7lxY5wSmtcoKONAHE0wSsgZgvtVSM8OtVYbPjTNxD
3hvVRJmz0VwHHUCP7mEwT1jkcHNM7LQiKinddIgur2r+OJ0OHVLaoixYmUl2EBCNVWCkFiwIk1GM
YgG/M6S91Ap9uQsMCZLddB+/yhPKAxgak3FCfpp1niorXzsuSv5CkUYDJZ793vmc3Y5GDQi2/Z3e
KKBLywD+hAU5T6CQVxMQOYT19Q/lHXA/0MXxq10bRwb4TIDT2HuBPt/YXzyOiFrKhb26QOpTRLQ1
RdTCtbpCPJcteiv7TNw5673WH/0aWCIvFHqV+GaOjaZmHiJRe9b2iqSC92bH58m+som/b4ssVO0O
7LVihVdvjZ45r9gDu7RA+Dzvw/RSjFMsO63ufn90wntNOZo9dG06/TZmJnOcCXFJfRss8e1x933z
O3oUTpTObPzWLVUwZWR+vSo1tO5lhNCRJMEOz3FQnMSQLx4CC7NjsP37k6huEaiHlzyUQUQ6kjrC
R0gw8EpGiXcQFIi9wu4DXfbQH89i+xHEYRzNkmwl0kl49qZZB8zaTDI7A50llKzO6TYtIbIy2334
pp+EITRyeMrlTXUG+aopkcKim7cves3p24riOjsbMWZR8W+VZAaw3Sy/ePlRziHn/UC6NOTXsG2R
FUi+sK2jXL0RoUG+NAsTfnxjJgBS+mdzimD4Ne/YRblEJSTj5Lt+xwN4565kCUYGvhAnYPTS59gn
TNd3ico1WtIOdwm5ZObCUAYfAZvzZ8M2lkBpFLkCKqVBbqJWgewnn/ninLPi/07MzefB71Lx3Fu7
Er2AyAJqTOrssa50UiOORv7nG+C3bgoKFK6moyxFs1+HRKn7LUHwaIc/v1gPpYnVeI7XZBJQyrdx
QiP12Kj3++hOMABMaZoJogtZ1x4BGeljBq7H+qK7hFBj884A09i/ThjR/2o8TLI5gzMWl/Kx5RC/
5ZVcaJQlqybxcxTd13xAfieMw4fBH8Wg+i12ClRsc1sauGEk6x33qFqI2uwgRRRlm8iWif1uDfRP
wxdik3N3noSoVyINEoXbKc1ASyK9MhNOKK+QI1eg7zyNPpwZJdP0MJSNINynxXODnKMnH9hQUwAK
apGt7Bkm9KN4lGm30qp2Qs3/DyO2R0U28gYhyoxMO/y9rVGo7nc4P5SYgdITTYqMU5h0cul+2rbt
0Zz5iOJ6swZoBoFqstzeYZiub17+aQym4Qmq7aNQ1mdn1R2cRKSlPEpW7vq0JTqg/FJLE0HHl7Hk
3S3qYukSgiRGMuCGh5Xwl8ZcIeqr+s4OSO7feTbLHVZauVPHYzJaBEHFFD5CH8OPrraMJaDNnhFU
mftPV+qjWf0DUoyUg5HkAM4nCJRgtdwmo6mMRGQ4rATeZ7uRKJsPqez/ZgI6tS6gxahDhf7V3jBX
ZZSCf4As1TtuOq5/7y6247f4n6tA0IiIp5stywNBpHyuobeKs6wKBJ6lTM02g/062+q2xWAjk6zQ
Q0pxdzCA8jFmx8aTjQgrMwyejtjXATV/DbpooTf7YxW6Sh/UwNqQw7/PlktbNi0RvioJLdyZNGOY
p+NWvqB+kF0yj+VGyPPoYjNCsBh5v6Zzzt2wXne0ldXWaxGI5sBDdmx9/0shF7FQe+6aoKX1WnTL
zZM3mZ2+D9w/3IYbJgVlKPZRpzdM276gnNn6M53uPvVNCyEG7ociZlX8WCJ8pzBVNWRYk47xPCsg
er37uJGArgBpl3zeGMieSICESOhHchYpnrTHnAKBovDOPmht1lAKTsBKS5BrebRQEuUDXIf4iW5b
HCck1S/6w9F2MDFNWtSunTwHOPsiU9qtLy2u3CIkatUEuwdoCSno7t4HIF/qxdYbDOtscMU3Vzyu
u1cMnajRKKFYTph/ah8RyqgKEt+N1MtqJm9ZPCa4xNG4vh9GNtgRIVxYHDQ+Yfiv3/BdF/V2VATo
H7kbw1wUB1HI3k5kWiHAZOwVrvgAPDXbE1oT2ID79XZIHSfPdszxTh8WbbkaFCGhzLI1CFWwd+QU
527rFoPhyJuGgljtQ/GMJ85mkXj1VN9GDEYZMzuvKOgrDy9XRQYlY+UtqahPoKAzgNksCe6qzBOY
WIRMxN0M1cWinVMzv86Z+rPur9qRZnRPmlyBplIGgNU5FhGINIkOzYaLqp/jOJk9HICDeBe+jHDn
bZo29dxtPBG7qS8kyQ7sFJJeoxMydmAKwmKKa6kW9o13db1MNEYnPZMsjLbKNCLX3cH8FNhf9Jfm
OYhAIpPJxhvq+jrGo6oshmKBMDwvGJAKW5zL+S1BEIiREG2QKUr4V7BR5DBfCwKv34NZL3bR1Dmr
W98VRV8Vh+Seq3yyzZwAVpb1DeK3Jfcp6fwYPmtZ0gaSYQ+SnLWq7ray2Ju7YkdnXdzvUEHisJ/c
k0TeBSpkd/NIqr2nRcggqNFmwou+8XwsM67JoYVUJ6XzKPQ0y139evPoFiGZ0bZy5mhRWqBW94BF
Eoq0UiDP3L+C58/kcOj+Cu/vqnu/UnavfsEPN+PFj2TdRAM7OPaUZMjdETm/12c5b5cS1qbS2uVz
bIh6r0F2qnWxCh0tzihNJdEpq8Aq9A9cprAZnGa/Blo5niSV3XPsgwcZZhi0vUZ6qKDEj70RLhQp
0Z3r+7XNua9f/UT97uCtVejEUFdtLSw4QiHEbWJlhZYttA0/kxZ4gTVgEUVc9kHuFR4g1mQ5YuMk
I+Lz0MNXwb6VjSlvbQ1QRcKq5+/HwKgD8hrC2aIgGU8Ktwmx+KNr8H36zhfNIxuTDZKU+YovHiTO
C4ABXgtbOEqwCApiAXSy8cTEFbkyZAuZOqHJFokUzfQro3CcYYUHH5d0S1ij5uOib5iypInR9Bfh
VtTo4LGAr8l3xBu2TSLJ4Vpsi1C5n/aEZc3OGQN3fJBLqgvi1T1yj/8neSGvP6CtDtO0GonIg7H7
8i9qYlp6iVDX5WGsVJRT1Ts6WLTtdt5CppfJ1to0ejx8sKL3eynAE2fbCLde+4X5lPOggifUaiTA
DvByeg3bQmy3he2cLP7NoMQ8P5Ydx5W1+3VjgLioYNs/zpXRYejozAKKIlhQYq0mRm+m/DIzC3QN
b9TnhpWwSrDDT+ht4/vGC217sElTCGSXhLTCkgARpDVDXAZy0C+i92ZJ+hWk/Vyu1QYLvIhbZFXN
L14t8CXPMFkqhB2iGvwXJbjAK1exeyIDJKH7MqBBfxBqrLVI68CJblp740n3MZN5YXa4b5/qLmm9
izAzJVuaeJqlsCx02Gnum8p8n06feOZS7eDMTXsKH/mZpwgOvrSgN+76ZjkG07C4Fyou8pum44fF
h65sfMENK9aFygpWM6mx+RIGWl/aD2WjaRjku+y5poYtRKQPkB+vPfVZMl9kIRviW21k4mwWdv4j
E56doZpBf3TS310Czy6ZzcHTYV5ULzJ8IoueDNx1b1HsOJDT5dxruHjhj/tLJZLqI/aPjK7+T9Nq
SgJRump4UxsVI9F+AidbjGprmq5V0GTlFiypWvI+wwDCigM7IvutMx7ioG6nNIscxzNG8Msg3QOx
Cvtth2gJhTHCEFTloQE4C5tBAJRcBPZ/Hiv3Z0YiphcHF5BSIjIyKWpsKkkuo/MF2RGzO4vvXncA
Ua00ct+nHR+cS7iErBUN7dDRcAoTgFrn7UQk/QcH+s7GZqU7UlFgqbkqxcnQEei2TLn0WsONQeXb
DcdPjNcjEDhRjFbcUr1v7AmwBQkYOlKDfJlMc4b/FOewi9s5Htgk3c3Q+uoqKOIekCPvBSgkObw8
DsWCX7wh3e+jVGtBPEBlwCiCZS7y6l8eIk088LSs17wFpCQS5tCpJIeCDPvzdS3INcjckm6poCoz
2Wqf+auTiIPIDyhb42sX/MrjygfAQvRnQRbg4WtCWZdJnai2flZbNBuZ6CxGSHhASvPhvYuPfwqs
xcoZG+XdZJwJPZ6pmkrMpOWzLeYq6tlBXu0sbcGn6rdQGhooXa2TBZmxU4lbi3TuYY0kMtw5IFUZ
HdBr7C2MHzYCp+1YRn16hGa3xtwOQZirweMZ+FR6hAgX5pA1nK59ULd3uTHzCb6td9dc4+znnK93
vIi086mHhklQ1KyqiOpI9eR86Lbie7gN6H/o3uJvNzqOWN5cztoXNHqVTbQAa08W+kYPsdMfznY5
DV0kffUtCyW3FsV/NZVIWVtinn7YLonyVJokU9umJWMNKT1+5OX6F0yT4TWvD0Br6eoZelFoc1OM
+AKglTKhKvDR0CUJSIoPu//zEKYKP+bouGuhcpEC+jn0v555or038PNXsJyW/DvXC6PXBCH8wW9n
75dzZ+6RUOHlPmG7X7Cjf8gPxvmOATSW70Cxfq5/2vNpqcwURW0ZEVU3QT2GJv06AKgt2lN8MTyA
VyXZEh1nrTwjitJ3YtM9q3tfgz0epB6LZewdhnLu9GO72SuudxBEbuy+bwIy6fnyVCCc3UgWc1qy
YmFLzStuw5tJoTXC6iYXMVcZXF32A9qZ4XPqhf6nhnu3Vb1OqXfZ8lhZYkodCR8mYsfrWHFLjVnN
J2zdn9zZhyWJv5/jn544vibK/Qei4iDrqW61kkZdmX5e7wmqYFQtuDwM/PRWI6+5wuEQnSJIOXw9
UmlKQQL4Ki41KeKqiJ51gT5qcQnlEUMtlDl6a0/okdT8GaUpkf/DVHt0oDdyrZ5HiiJOGGC7wTGa
VKFKN+7kEWp/4jW4KJJmnBIRMU0LhHDIZ3cINThx2uKy4pXzq3hhH+9ZoMKyq2ZMQ8M6cBkwaJkl
91vVai8DqmNjG4t7WsOueJvSH2X2aBIwtf92hvIVa2BezOvEKkpixykqQTcVExv229TqNdm3Iq1g
i3c0xtx7K6ITYfAhWBz3AP9aTxS2V763kiDU3kzlZmZ4eeBNcTdhQ0X0zmhaBBzZHSzR3SALiMNS
gIra6FBF/5729bAxb+gHoOjOpXX9YOoz9NmWkmNpxFTedCnUqszkXQVoEbJFG+zCN+BZb88f6NSv
WYYqhWt2XATCEOhIZTT7ploiJvZasnKkTCDX+bA9xzYIWrfpobG1H+XTAa4IJa9n8Zf41R/KZ3h3
ErSGy9qY/W/I2dLarRWC71OtxIthnm85col+t866Vp9MajMLnOuQUmsLtCDR5CUMa1wQcE1Pcc1V
/tObrXYApQF81dO9AAnwjD7nhn3E8nJQenmaSpuhJk7sEcokL2P+QqB4+LpNc19f4jB+wnxM/O9E
lKg2oLKW58Xr7O4On45ILmD+A/1iYRdihctKsh/p6f0tTO66qx3ngbomuZkruF6D1WDBW2y4lJ01
7JZ/t5hktQWmuUlZ7JjBuwJMzvMEQ49THfnJwo++4M6aB/NrCNfaRNk0ap4wEgcNLksyNKASA271
l+rH+HTJ6zOmTFdjS9G5Tp/SARVJ9yuyvW2QnMYjrg9ogOayyySqvZcFNTMjCNc6ownQDVD6+6YH
/NEpt4w6s/tL8x1yhd2kmXxXzwy4Xzd3WKLD92ATLqHe3Mi095fcQRanlztPi9f8AqSoOfW24+Xk
P1L//PJw+Dkb4DiW7ahR+EN8/2+DYswd/Qrbv5ig90ZzqzXxRX3KXnUkhkRzxG+et4SHJh3BFxK4
awHQ37ZT/qoLNpPsZmrLini7OResR41+aS7N5o1223evirKbBNxZIGp+f/LHWga3uXiM1hrtHUhY
RbLSLZY1Aed295UUO9QEcPDBQ7z0IZnHoEBNyz+Hu1vW0HLz2Rtvs7K6CeWJFvmoMo2vSM5Wuovo
2ZGYrgTsvtZqP0c5F7gxXhl7pQYzkrdyAngRHu3c0mTUCeNvChxarDRDeJ2oxDAH+msc9isHoEeL
XthfQ5qVH7vfaj0arluArDyDbFCjiOELzMHFJVl9PkcLQhG/orkdz7Ap4KFfO4/maoRfxKW5um9G
3Bd9J8vhKymIwy6JVl/SWdvzFUaR+34ZRPsp18iHrmueKIGmayP/19aLJ+ypm9r/aYQtwsMFhzdW
ZiEORldEoFKt0Ok+umABHzWmKpkJgAXO6447lQcwFdkMvsvwHvp+vl0el4byVzd3MC3XnNL0zczc
GoOe+PgkBb9wedYiQr9EB3XxUavTNEtBC9ERN/qSjZHhPKupeu+3idoEcbm37b1dtAI/0Td/kiwi
VK6vjecrDf/J8BO8VjzV/sJIs+YIl/mgOt1Arv/pyphXejov2aJ2HErJZO4PWQAlEYARvEmLvW3M
WawSOij7VKc5vdEOLuajPNWA6geXwVznQsjMk39CCNGnqprdFpCh9LesfIqlgQeyg7LoWrilyV7y
NSZynV9+xFPb2zFa2GPNnMuvF7rf7VqZbDp3wg5Jd7Wy5XhGBgZaeQW4PIha3L9Wc7cJmgog3FkO
co1Q3ZPAzcOMVTfFTm3kLpDCcnu6pMil3f0Q3dAD7QJ0oaelZl+w11wBp6Iesz/DQAYIPrTZwM1n
PwlfcOzIPYxFUPdr9gvVXH4KRNJTKMjsns3SXDYkHUsqfWr4O9gx89ZQSIuE0f5omTboYjmXkfQ2
2Y9olk+DYBYoSb0u2t+CE0M2IB39OQdBKEmMx4NQSVyGeEpH7mRPoeIQfP9e86HR8jxVLkHwzj4L
OBCyzukroQcb5P60t9rvkSao0PPhNYc5e0jXJk3EcuHVK1SGKZALcpAvTy3/kc+9Zvz0pCZVNYcx
BCHONTNmckUc+nRU6Yomp0MLh231sgGhaPfSAdr6025T9SoxUZ9ODK7lJ9LOfzXDzK1mvqjHxdNH
UbKSziBH/xCJyW27spba9M4yWvQNHF5c4jgFRMi0bwg8Jip6H76zr97BvaMP7+b9f7xXMXmkQWr5
j4fQmxEnM0CUSaT4gKgxiByiGWO2b0Fq8ZlV7hQAb84+UKzb9UDOGLfcTy/1/Tk2hyO3HFsbRnG1
JRTra/Pfh0JqkX2hG8QnYDKqM3Dvh/sfrWaZLs5aiJsBOTUnQmhAl0UjAU0TvqI0muY4KopXEbtf
B1hFTbJ5DuCXAV+k1ipNXlgX5MxLk1PPtgZxwRaI9hk60ZIAMRWA5d4OhNlO+Mizx6YLcMhYH2SD
fbDUr+m541aKI8uY95LBRF1IGTpxRgeuaBne05O/OqJPtp1odY635rYm9x8lTfZQjkfb6UmWFmZu
wnSy+0ffWzCRKAmlpDpMFfHON02kEFeropxRY/QKND3Tb1f+uyiZFeRpp/gjwQwEIh0L3YJLuGR8
mhU64OSgAZHWFsNLSta5Wu9uySRhgkNmISe4T+T8LNI/pT7c1sNESGcNs9RBzxexujrO6JRtdLwP
HwMq+QXATaEEzbmD/Ay4AFYKD4tEyvLsJnQ4fwJW2ihHqHKli/Jm+B4ZGCg4FMHdtbUA90VQz0en
JbiSZqGK2DSD9trzmlhXVzZvBLyARtHD5/EEQ1pV1JVo+6nSL34HFuZUVhFxsW0t4k2JSPwd1o6Q
mbb34ziWgEx2hRrmpLVUwzcs9u8S2BexL+my3ZWAT1HKFKCf9s1dyR5jCYi95xE1EGXCINFA3wVD
QQJCLdTW/Yo/EaaKWUbDjtBusytWkfIz5e5tKfu6AR/pOO1I2W7qcapxVVSKJyO188Kb1if+W65k
6iHUhi3/MpHwEcCc99afajzHG6Bu9al7IojUuz4QWNwATsm3Q5HO0N8UvxiALg5KyLFef8vEJei/
lCix6AJAThOmN4VFzrEy8t8lyF8yh+4AEfIN6kPjEEihX+sLXyp7H3hQAnryxmXnUAEciueQgOLi
fNrWrJHLy9PjYzUreoq3HSZivXlMuxZk0HCbQ49ZFd6ZnFcXB+64iU/zPLPR6XeDlDlUOvn8zuKV
DvysFmjZ9bTe6viBGkQaktyacZBOTdqD5+7ISPEaBcNA3HtzPV03i5NI1CyUpgSPL6bL4x1DOh25
JNxo9ea7zmEcoKZ24to52vsBKge52DsIkLUqFb912ZC3A/hvWZam3xiQGWtBudMRkv3w0KUF6hZR
06MYJe2KNjU/E2EsqvIAWHzIRVHSnybVH5bJW2JfnqOAhEyJTYNR788CsrOr5LKKfCX4E5wb9Vse
jcIVUu/yJSDV9sU1tr7i92lANrCGG3t44DN9M4FufyGXYDcTWo6VaJsPGTVHANWiAdIV/Pi3aypi
CoVyUPgBr8o2WqxqsTY7Gusyqr6LacUlceiSS5h2JQGXljZKfdf6MR+mo9Q/ckXpxUgo0CV3xBdx
A8AA3ncfhaIEeZ6lVDynoZgg7IUD7jir3KtRQdisCFo2nPrbIMe5Hy67KxDOv8y89Q0RKRhn0TNR
OrHO27s/qu+/SDMccTIJpKjMQ46bPCjWGcFCLqiN+3DKcvcBDmPOyLMaozB05kIJL7BLzgAX8ETY
pEUdJBe/+zUG2Co7neGyJc7rlzGbUCt7I5T9YqXlbaKJQATghAhYYa6Vkkebuc1MKnrSVhvYwQ5C
H+p2hq8zNIH7RrBzunYNG2je12paWB6va76MCe0ODPa9KxwRTzsDkd6M3vWxLLsvM5J5XvMn2LjT
0K2ZBAE6P8DYiPKkPtpBOIn54y2TZb+cL7gJU2jWSOcaz193iUw6NFMAL374rH9XwHVNsB58yWCH
UUHYAXUmm0BmS5pUZBbyqde0gaQQChI6wQNSqwUl2FaOTrOtgGT9AOVJoUBgIjFATK8Z1ko32ibR
7CyawcccUQC+vcAG/6los6FXejkudvuROe7+ksvizaVsjXrXk5plQ/u9CTznPgDkXR1mvvnEkB63
ESW+lS8nxG/q0E5uRfgcvNXo0FDlT+/wrVrn94u73/GlJmuoYBDarnhXvrQzVhQJLezoS1rXdqC5
o8ZJIGV42SFFohYrMmI7EEHWx1Ppve9ww/Rv9dDmakjp0RgUEw0CK5ai45yWiFbHmTLoz5xJYH0O
2JjYOnyVQs1mQuRHzyv5g1CyXK8mShEbIIzjkJNpzBsayLuqk0nFGNkaWY+9qmWL/ZTNBliw4ZPZ
6BtoLjDuNWUI5DteK42k9SOvpHdpfJU86+/90BraCos7On3kglp2PhxZfPTUxeIYceoPmK8N5ia0
ILZZ8OuHwRtVMtD6UJQrBRMwB/28y8K9I+5mTbdbhohSF9zJGziz8t6dMhTBthzBtdWtYB/QHp3E
LRWNAjZuhO+rAPQ8M6ITdWJuIgnpz0xyrRGWRS+E0U7h5rdAcfwvmGxdjXX+4NcT233CC0ma7IXO
0WwyoYJvH+CRpCv3GlZ4xHaXCO4OnGGN0TcR5elLNdCxLRL0JG27aTu4GpsjS+0oqm6CaVRGriEm
A5W57duzncxm+v08czXjn2rbsTsrnm4/jWeqrSqaXYa1g8UjjENV1wJrbspPT30Gk5KQjOSyzqLY
/tP4K6pldsLCSnwWH4m1OON7XnRwwQGIjIPIlQ8qzNjLfKYPbRQs+1WvOkbnoY33cqERShNS10H/
ptwy8syum7oJqBrn9JJuHjudUbcsJ2dek7oRX6pt0zOvkfD4mg4g26Fiu8r/arPzRMS/jhgSbkks
EV6tD6vX7K13ZJsx5Cxs6A9X0sCMMNiDCVG6P6xJBy20riqyVLDDZDnSW7sWL/8BahiUaLZncsU3
tzRss93rxSYEceZMyMEJAW47Lqcy1aC8YUXXSPuoPz7ggcLNuHzc++D4GGXQPPqjy0Ml5BzAj8lU
fMSpSrpPHVkZ0J71cCOIaiUPk1IdtTjQNX5je1aKpmbY4rsOSHA3oldG8yZeTD4t3oP7EqyOarpo
/x0/2YPr2XCXdvdPpGzEqWzRO4GMKzh3/gmLI82R3M9MDr7iIqZ0FGkLdpmqr4yYMtnGfSyPK/uO
j9XjB+cFcmkekbWMgmTBqksiHa22rDU6ILyLhmZRWVj2F6k6SVLfWKMMPCDP/DTYScIlKreO8TOo
9MZ6oYgSjVjzZ7L6GaqRt/I1PTF/KVFso2itjTAHHW/g/t/atZtCyKxzdJ6Yno68p4GjcF65yjDp
x2DvOBvDVWVLgs6EtuO9N052BlXPpdISWnMXPA8sgyHfVvk7FkYsMvfftaP/JVwL5ktueYMjclZT
v87lnnKmmIEKLqieClqm4D8hfhIVAcKqSfYfzHUmKvbfh1nu8mXsRPJ9ti7uxKugl/upCWGpw163
R9qM44bW7zJhPTBxhVPjk5RcWtHXp3J/Ppdx3+mZLyWe6CjCeW/KjIknkkYWIulTH6FW66RKUchU
nk8sb1kFqdNFcA4/SubSRK2x6q9OSL3Uvp2wP7R+wDznon9M21TfddBVMuTJVblPi4aeaIIrt502
b9B3M0yE4MVml3YVO2iKqpDlEL5ePU/lUvIqifPGbHWF7UjoDXVthJoPFykgJ/CoApj1UbEq9O/3
Q0kONMYvOIdXgF6p3IUf5tSqzr5KZYwqu1MfFpjWfj+I3OOoTYvnz6VTAQPjY3GmZ5iLwyUL6h8T
peeasIK+bkHMJybaO6x5d0m14dxT/YZVGfuTn7tO30TadTgbViik+pk1xdyMY79aKP5/f2K8XVGv
3WKNHiWkrh43xA1xSldi2NON0blcnaevwaCNXpkOtmKlk3ueE9lkcdS64VG3xTv5gBIA4Dm2fYZa
LqGznSt018kXN2XY/ype6TnDbIF5wiHPejZ1HkXklCUu3jybq77LAckgEiyt6+LwZ0p/EQOU+s/i
cwsJ41FGB6mUnUFqLj3jN+zkxp1+/SW+IW8qaSGhM2164QUYsHI+80y8cxLaX0F2yqtFzJ5JleMR
Hb/gLcSMl+qcTxsJOqYG7i/LiY5Bqvry3ZdYBTXZmFVnBSJ1lXiQkIdIRRQfLirMMU6jqEMRui0Z
KkW+dNICVT9qbQhUn2cT+CZJ3fA62nyYGzKifD1YaKe4r0oyA+sbcONs9zOnJDKPdL0S3ymqeX3K
NYrPYlc8JXcP5THcXn6tYdHh7NZeCWUXyxd/OUn5RwALF5DejlKcma60Qh3pFiSe6xr81SGq85dN
PQZvXtYMxUV+qPaCENE0CBSmXF4JZAYIZ50p7+piauJUxRYqpJx911P/uLluMZ1nB8aFDk0MvKPV
4HSMh6KedifFSZi4LFRzUM9BDltYrcujVAxowfnnOBfUtocy1kHWzWT+4sdSfwBGKjiODp77V19Z
yF6RO+j+3ayxJ8sLVTt7pR5QuqyMTJFJD4DgHr6sxoFyt33RpWfHX814qq16ypC+EnSy8zpaEUZg
IM2vs2L3r07GJ2tbgQ/mCeyqXchsGQX56l9rYxzOG6z30RE59cMCbh52yXkGwFc88O4ea1WIDrNU
I/2VPtVFUyh48LAWvxDlKCj9+41AsDfgS+t1dphsejUBasxFj79Y+By82mdD8FMyaTXNAOwPrdmB
pv7dGM/DISiMNKQXJYHtXtN6bglj+acytFlJ7rC5rkuCA3+ss/jw6qVJ2tuAefEQxFX0ezOl2+Kh
NDB7QKzdwCsnYxXYG22VMk/J+BupqRi4hJd/H2aHBZnwJcTm7cYOm364X6C/eC8ZcAUYmvjLAwk9
/AMq87mUVvhRrsB3h5ZTNkBq3yuhD93BOdw3wj/As4zWITOsgMpdnn1OnxcWSa688DKbHVrcDs78
tw8OxMir3cuM0a1cTTkClvRSkiUPx/IALIo+TJIY3oWeWNlKIDNeYSbrZvnkBaZl0Erlg/LYvEuR
Xfnx7yHEzBk4WTBZKjMxt5NoqjMgohV6fWTSxC4LwsXcnRYTDwhYJgdKq+Jh9lHA/jkXZBzr4n/m
RxhugPsPzCQi991koZOh91vo+funstkpRwh5DsYDadlw7CpkMcz2xW6BRkjn1kNBZ0OWalqcOTXy
uLuoa/TkUveh3PMpH/7TR+YA82lJjCLGv3rYo9DqG6qGmbMcpHBpX9AVDBK2D7sKWqPZiBDpgFVG
rPTwwTbrdC8q1n4ZrI9obczxjAU6oqclGlwXEQZpIUpStSbCb+uuJuM1qYAOQrZBDz/uKWF4XGPl
+V+vePWtzwZnwfb71BaGcfAypsbRTEpwtJTSpWcGe8q7U5BbQcTOErwvbQMORDV+OsMLRD3AzxV5
Dwu9ifaWUv6I3Odv1yDAVM8itafbEmMu92CGF6jG97sepb467e67q7lk/NqqEXJAa0nPldZOW7WF
FqM0gGAxFoDSIX7hZrYAFLpSBL4LPjsu+PsPW/Uobi0HA7vqdh/xjTz/Qr0MI743mBFA6ZBifg2T
M26KvkT9E9UCKuY9EmzipPJVzfcAnQn6OvzWuK2141yvmP45jSTT42Je8f/4LIAw0IdJin3FnUxQ
MR9Rb3dAszfppkjJBpSRB8LJHt7E7fQqZ8vYV5e3hDO2+IZQ7D9iBjS8SBKRPH2rptmyttSxmFJ7
EVmb9fy7qrQnwMne0e2T/dk6oWuwloZn6fS1+WU2/J+IEtxPJSXO5UH+VVQOT8oPh/IGfgLOqYOS
4flc6Vt1mKMjVGCa71SxSJZl35zYuAVSdJOFOtgUDJ13GpmLZqkDVDzA00OYMKV6TpTfcmHPdTDL
gt1ptdCAneWo7fBG3AFORB/K+Da5pb3xhuBdeiGCbMJ/YVybJ96AoQ+u6pIepea8sSfdOkQgrqny
jEckeWzPWrGhaxxqgWeOhGYT1MyVM1RWca+sfLOxDZxNFDoRc1owcByikfAiUZjmWA0QWbYJsgGD
HXOXDX9mqMDXcN5rsCzpuqVLlNPgZnm2AyCEXFcop2GRGGb2DtBaV2iGnvmZw0ohoD2G72/ZNzpl
5TPcwJ9MWPYS5Sw7ehXejp/6+dD4/p2bkBXDRtVWHY+wbAyQ3V0aZO5eYFgF5IWt42donsY5Qjnh
rarUoUaWxbeDr2xIPP2DDZR5QgligZ7ToEAgGZRwYiQY3ElQD5nFTXyGIgl8eJ0yaygpX9b9jGFO
ur14/L9zRP3ZfoT4SlmPOVofp673f3dDLoH+KVfzioQuKWrSCRkynBsJj80FrIh3UjdA1iF670HQ
vJDwJDIaH9ozBZXsKtBS+3fI4+rOnQOj9kig4zMZBL6ge/uh0rZRoihuihpcvZb99+IbwLacnK3U
knpdjwvTWiLdgXpxUqRw8JnfgUrORHYSFEyHnXQPVg+ioCnaVskUnRX4l9K5eHcguAt3kN2O6AbO
0Gpgo/E2xvTvlHDw1rZTtzwCSQxKeIWLZWa0SAS1wBc0bDGYSIj2sRqRlUzkQKIpOfZo2xKJWirq
h0PvcYfRcN5QhbkVpOzKxEy3RpE//rl3ZAvfVgqV6w2QMXlI4EuQSVCjVK/UZPq7rMgkbslTlGAG
fkxUhMZybkoPpppHvclAVvn3GXM6n02lIoHZikDmHRnK9MwGgnelaV0HDpmPPAiW9LwlPtThx9tO
KSHV7fC5+A4W0mQy/DMWY9xiNeLNyY2kAMMuZtrf25ydjTaPh+gTIk4bZbYrgEROneNNwmBjg108
Csg5FS909q+gnLH5ix+2Viy6T+1CGb9250FgaNQziZ7Yu3khp5wBmFFPuwMiPCtprLwqxQeoHppq
J0snQX0o/a05BREKZAncdt+GqIDs601z59TcRvmslAlfgmvSE8fMTqHYH60rkNjrsF6T3PaiAZT4
3M3dZCkOi9Q534Oh1NY4oyMV7ybVuNVmz8KXFMaS1VmbYOvrnmEkMCFdRyByJ6jaiB6z79v9KB2G
7Oam8rAHWY5QT0g/45H7hDt9P0tqBarZRLAlZQHFLi88bjB02RAU5v0UaFpcLZVFwOtu4BKFCk9t
GGjybrOb8YwGsizGSL033dwidVFY9wFXUlYLel7dH048GQIgq8gzfCyRUXcUkSGn8l1b/BodXkb1
APYdR0cyZPzYNp99nyYElH03cLY9tszGK8edq7wwUNFcz0zSeGLZjcoikRjuXYOkgphzTDwhRHQ4
1BlgSOVX8vKLUBUAb/0x59/64W6Capj/672k238QMBEJKD+e9eHaSOQARiiVdPLnj35ipC5hyQ4e
7RmnHpVEcy1aacKu53LeCXebzXDpZeaiNPPVKJzbMldWwXT6CnX6wERFduqaMFO1T/iRjCgNQgM9
smcIqTUoLZopDTq0xR4Dg1RUFMJPWoWV8BA8NqHj7uCGvXyJY2H3i42xmMp48xw0qITbSd156biG
HzV/GxqHjQTvYPRuBvLCn46Myw3rPyVOoqjDzAi5fmCLz4nrcOO6ZbGdwWqD4vCUpCmd09yFNH95
GpIjNuCgZmm6iQQwnhq95T/FXFXsxyrd6qOivv9NTypjQfCE2xEu5vg5IkXT1fF5myHff0gUYBQO
LSsVTx+YrDPlOv5D1o1DlOyMMNui9Q+x/geEY7H/fNwQ/24lWIEFpAszMCb4Ug8TQjeMWMCIMdQF
Yq3LrOIWtE6pSnzEj0q20FZCk0B5SsTugOY2ubCBfctTp8PIHbuiaZIiWWRM/g849n3KIQpBHrAD
wTSQDRwPfQEkdFkdrbfS9R7MDaMMd1YTtd6zs1wrIN6J7vsg3QacPfgvQ05rtP3SH3mhnCL/iiiu
OWc7q4Qn64pgZ7dStLzvv0qUtaeZBKiT8i4SI5IjBb8okGAf6yb616628L5JAjJK6hVMtw7ghd/4
MZMJ5N0S87vPMiSvIWtZ5KVfABsRi9j4228wgcyKFbbdJb2xknBEtHDrDcs8P/xPVQSzxQ/ZQNEM
JzpPvFc3etY9bendJESujYhJIpVcXYD3HsljLJ9wBtP1s7+xfCvvnx5JNYgqSoyEEJGnRayWG9Bv
The//H3PQsBiliPKrQ8Zq4PBZ8PCgbiOutJYQJ6uG8CBqo9vWi1FdFT9KbYnx0UJ2qwjLPBXrJiB
C5CzvA9NP7MBD/jIiUic4oM1nUgTPS+LQwZQNwo8JujnOG0Vi719YVuXkCwZLVDgXwchj899NL3D
lCA3IDKPNN1Y9WrZxeSxeEHLOSh33W497Rrn+itCFBNyRE7LQRXQduRP3KPUgRWSP84pVopR3oVR
2hcYs4e4bOOSsqd5IWIvAOfJ2EgeNnkvXnHEUTDd/wmLHp0sZAtudUOhpTJpQmwVo9N0RkayaYwY
xeZJvqkP0HPev2zragdzU8MgPgb9tjz73xvk4Hb51QggW2w8u+higTVF878CHD59uWkjVdx0j/uW
wxIoK/fEvq+cgtNwjpOEvDmUtPXAKc28GsVneMg/DlGCP21GOgC6iQrn0WXlYg61ergNk4C2HjHA
9JDJANG+7eicas5EHUvEOPtcs4BReM02S+36pp91v8b17bKEFhTut4GtB0hmbT+NbAuomstmXHIi
nHJg3Z/bQxi9x0pzTyaD/nGezOhqynqiQsLCHPJ52ZjBP3SCsL06RAX9+2deapbwuJiw0jM3fcFS
0pAAfMoGCe2p+OMo/OIdVj4WVZEbIOEnxRwCpBWoJgnjLsoz+c5uMgnTTK21XH8UPfGSE51IqM8Z
KaUWta5w0n6vj2ZxWoAGMv4aMTpnFEz5mKn2gXPbBt3V4OaVy0Hg2bxum4dOO6MkoqJ8R7XgBuw8
RvlgmCvBMjVFo8/l2Wmm5jg4Y4/HVOsbQL8j05sgtBMJIbYQANXanxUHr7GL4iaH9aasEM5/+0NO
L8OaER2vjFC5AzjQmtNxj+f7IflfZ4vE9slBM/DDCrN+x6cH/07TvK/Tb8HBUqAX/S3YZ5pTQzHQ
87oHDLbjkoMRp8fi4dCHhBobIuGt5MG3F60x+RUIroMudDds9HMB/KueUww7R398N4Cx0FIEECgu
UpQ8WN6jgsx3d0Icp9rZBu0H8HzHCCkCtV1tztSSNnyMutXG3YtiC4kFBmLIze3rBdfQf4XxtX7o
tS49eGP3Fwyi7cPaH/k+/mRXOswIcgxBIBGgj8GLG1SsUFJ9Yxy/9bJ+F3m3UzYuQ6bNSZdQaFdF
ZBurc10tnyqYxfFWgHm+odTT+yE0oJQNhjJTxWEm5v76MEj/EzaM/CbFWI0J9aF1K7Y6QzsG2Oub
hg+60Wv3EpH4+UUHQPxAYf5lyfky33sX4x7ZNANb3YF7gWQmL/ulnuwnYwrcnkV6qMWDt9RUSqbv
ePGGrSHFsYhTLvoTngPU5b5uzEkaLi6fiB/o7LufWElyjxz0t2f/6OPL8bXPiNQ0GB1Zxmpjz1io
VFZsY8ZrHrBj5wvZeVgsk74U/+BXBASKL2dwa/zJTgMAqqmaA/IE/QaEBb5gnryGPhkvN3xSwNLC
INe79flWmJSVBTd9nb4u+nS3yfdaem+f9Wrv2YuOPOLSFmHxwJP7WR4EJHWWrwU0CmE76vHcBKvR
78WAxJ5hGVXY8OaoJlSUs/u9G6OUf3fXr8/8xNdTnhLSYl2VYhTIe8RBKalC0gKdpcfcr13/r0JP
cEBZD0HbMnOdsjQbyZFaeh9vfnTwThfo5KZrzmEbojryqaCN6I6NVgQ2hp8/l8r/u3jdMZVgxRlf
TtGsrKCgeJjVRWTiS+35lrqe0/+9ifY0Fjv/JHFMIpje7cLr42s2fyVRhiwSCthmaRXF9uYMzOf6
5jwhWc21jXcSf2RNBut9LNv4ys/q8VR/jDw2dKrkvrsepKxeX3idApK1LccwY+zV9JkP1BcqcK2h
eDUL24+keHnQN76nkayVi8HqJjr3gVgDw+nieRzKG3gldmQnakvEVoO6l4Cp4ugd9PYq9tEFAc4P
AFxgEoJ7U9NS1BgIDC0Yj/X9MmoK0VlTZiYwMsenaKnFxdCC8I6wbpC6jXKdBN+VxAM6+CwS1Lri
UIc3w2Nl+lkkt+ZW0SWTyr/JC5Msj3IlYUGX1cK6qRf4SEFqpiTQ+a5jqUDzzgTZXALxQwMwvxc1
zEK8uaqD3IhLFe5dyb+bBKAgcgci0wy4XIEsUVV6f7ap4fgvkvzaJR8pwj+EXw/hr/cbSw1+BlC9
+AssWd+2x2sTffT264udP0BzPqNTuSeZwt5SaHuaN2bSA/ql/RsjUpbKkKxWp1Rhqljk5Y3OVqQy
8FmT7LjhnWx7+4ndIyOxDk3sznkSVVk8m0SsqGaW79USOSRVQUV2KhOz+T+C6DFWQutHp53WPlqv
XhSor1VaTNOVdMypJf3/0LO5KLc/TxYPP5Z4UQ02MmHSPczLnIZBqjNjVdr4ulsJkdla6HJDeKvk
qkMH4ENKLTyGDm2MKJHwf4xiejDaj82XTDMBwiG3K0ELwXVaeI8nYKVjjb02Pl5vj447vVNJMpVE
m0cwWFipam7V4K/U8xaj/ECnFCmQ314feQAc90nfHwXSGEVkFK4+1iaAnimVWr1aJxKAr6ykhcfU
7XR6LfmPpiDA5Wz1M0V+RS1JkryAyr45JAUBVylX/9LkhPstvcSN/hyyghDvDeu4G5SqeqJZCv2X
3y/uK3m3mbq4CN0i8SuO1efHieUHe+8EEO3BUJI9IGprv8oxzRgBHeUhX2ctJbcxytHG1LO0mL75
bVOncxkfps7S5P31FbyQxDYwUx3T5SXlNAFOkWI5EYUwXgZ+3WE/RMNzTm/9+up4+ozUSzWLq6W0
uO86uPf6l5a+p/bgp2cqzzBcakPHa70raOQjDtR8Kd+vfrMBn6fYhiH1LuVnt7mwj8Nr02OK1NG/
jfUmwAx0ecST9x6QlIk4riZXc0KgFNk2ZAHzJE6xA1ipAqRrWTK0r2NnGB2SgXM9OTSMlXBrWpVf
s/fDFwt1SBpt/xuXebCnlyUPu6oYevZ6MuXeRcq/A8LkbVhwNEu7ESLf2H8WrpyPWGWA4uQvWI5I
7UemonCQrsrdwKg1d15bDE7KsVScs0C+VzmANDPrMni/MWopFRChDhPBZ44Dxw0PrgpLDWrYtbfw
a/ViSoCZ1UkKEWYuiWj9Oxip1L6t5i3vgm0A2zsgl4yQgVDDDOOwVCsaCUR768o5J+WPuz52AuzX
uxu2rOuvocj264ZdSi6U1hk5LHgIcYfYz1r2tOCRucGn0VDwI84ulx0aP+8ts+Y+dlCpqV/hdnBN
mMOE/tK6QgXGUNlTCVML2M7I3TPylnJ0mrtaohTYFq4AhaTjjbosAdsli0iDfZ+MBR42XNz0oAC/
4IA360tiNkx6KG+odeaihyKju4eJDWpR4j/IBYZOHJPfT3FNSKYAq2vq/jbZo5ptTLuKomMFkAg2
b8gXbSSPwWfYLQ15Fnb2TnPoftQ1SDRtPR+cg3A8aTe/wCNXt5TUYoKHDpvofvw+QhBf+ip07x/Q
Nvdklrte6s7fGjcDTX0FB9HdEBmynCRztDSByhDZbGGikklegbMytWOE6H09m6lKNS2pOcu2Ess/
bMHwal0SJH/+6oq1tT+/s0gIEOvyy41PIVYeW/tH6BOXFFeh3ktDNFmbkxKH6O/vxfTiMS7rDLPp
p0sssXiSPUV7DNB2UxOdn4YbNG1ovQudInu6TJFBZn4BXY+lOh+VeQVCk8M/26ypHrIO25XfTfTA
Lp0bCRjnss34yOGpZDZAK/6OfWa/NNQW3jvEoB5JCaohciS7QS8KBZPPjYJPaPf29Gw3b+kQVuqo
Zv6CysT1m1zjLkcug/IpAD9tq7u2MzwHO0w6k0DhdtPMRbz6gp42rdSlHc9+dmfw5iLq9XjZ/SYv
JNgopXpaIepBbvuU8bVrVD6dN2i62Jj1K/K9imzCivqNBlLSuhHNYStV6XHlktpGbTcZj+PqvII2
t33ok+2oyDUwvNidHNN9OKSGNL9kZmP2beYLUOmMrmb69svF0nimREJazilCWTtP2ckNm7EXQK5g
h3g8MrszTFRpsFlEIXvL5pTC9Bb+LB08zBllQpGIdKhzrZ4j8wUgoGymyRpIc2p+gy8ZRGUOl9MW
JQJpwrs8gP4GYo4FmAsHDFrjaVv4uXHooc1Om2em0cfGETUXfPuJ3kkPSGfc4BnTFxCHTBYHeQRf
94WzbrdA7JKOi0jvZfrDY8afX9AL1OqM0DBwHhWurWq97IhFlznbV+BTvDhYjOXufFCJcUoz2Z8c
yrdXLwm92i4X6Bdcd6yMDeT2N3S9kjNMZMz15BZbKyyp2k3bW7/mQPgw3d8v8vLmMvPUjURiidC8
BxsNbJXIFNxVsEyKjIiIXuu8duO8+sAIyCdkw0F1artFVupW00ZXJvE+CJOx77dSxYKOC8Elelsa
VeKocJz8GnX+fsSzZ9s1MZduz2OKD2HPZdG+/HDkNUMcmPWTvD4OR4/uLUIa+Q+03ZmPy6u1elix
IjlxJ4dy1euFDn+YenzdpHviX95PQwuKrsIOSgDRDvRij0vDlEJfKCl0OtcVr8dqSR2CQP92497b
boQYJLwPr4qDiMcAORgDm/50IlzV6ULZZBB4K7VPJt1HppolBwlp30SZAqlpi3sn5MC5eKoxpj4M
v9H8bn/8A2aj8Stngnkeoaq96PBzTTVokqCIKhIi1Q0jGvkWSQxB/IDEEmsqW5i0XJzUVesH/bW0
uq0AJkMFMReJCIYls6bKUk0Zc5NQ6R8ByyDhhWJ1rsZFZ30WCSLBkbSOZAesRP+Ppz6R5KwETaMP
1fH2ZlELU2y7i+6Oq8cjw4ot7B3i1HmbIkvIO0pBwATe9YfkJbbY4Am2WKQ0JWH4s4Idj2XLYx+n
L+z84jmrM4nvDwFGBuroodcmQGm/S82G6rQSBA9snnIx6zdVFfl9D1Y3GG3CeNRqbf3na+AmjFnn
7SIFdsoljhLy6W+SDDecd84/1t5hedPrUtpRe0BYRyDKfz8QrbqnRZDyDro3FSmaWDOmS1MTmtii
jAbxWXH3YgCVkkQETpfTFpGLSEBUvEEJm7sPzGr+Pj2ddhNXjmie+g2ljg6Lh/Ws2bLXsoCn5KiG
7R1jp8fyD+6R5H7s47UZqCZKZxxHXf/AENhKhR3UxgXlVvq508akaJX96Mmr9hGgFPViJH0DFLUr
2yqoz47YKCImV+UsTSaxVH1AOU1+iGaMABgkee8to1/J5ARtCj84eYP+9eEbOvkS0/6l7G5zo/Cc
VpkPRmL1YlGgugPqNfN7zwmvRTNTw2q2W/whwjCpmtcLFSKjDEcACytbG63ra4NtvjtYIXYKYdiG
m2mpiO1cdMRiCkMIMjNCI4VeWhxZH+0tqfOjpNzzAOKjU/uD1ImRmQIucBkRBMAjkHenucLU/Ej9
SYD3Onbr/ShE5SogE8B0AvUFWpJxA/qM3huxZ8NZ1Y/bwkP8SGAybSMZA3tiGzw1KoyhYSmNmZso
ZpXsmqT5z4H1ky2/t4a1U9qKswrqy2LNtHFcszl6k6/yT64/+pteQjA1W9pMV1SiTtkBoeoDB2l+
ftb8eKxLNRZV4F5Ah5siKrjnl0gZVJzMn3pX6cdZ19KHgrW3gdWwO+egOxrW52sMZUL0VCAbwHCf
IKKw0f1nZYGDpWnOBt/Tlbk3THx8BQpdae95Vd+Ip0M3AlVC/17g/rrQidM9N7MgljMs3tpNsEXO
LcbqbnicRvvjf/l1YfGoXe+yoCIet0TWGbi1ECTkHCoCikwoKXr34qO2hQiobKg1arnyjyjnecJ+
GiW1z8VPKL6Jog6uR/xTa8TICoVxbUIo2iwKfK7T/WeKkJWpYDMKdDNv67bbnZb+8bbbUrwmUqA2
ySv2EFTLs0kxtXGTxr+R0/hDtxu+PkAfo8s3sWrqIgee0K9tOLah3Ms2hCTowZFe/uoJ0WMcnVCM
punF/bxjhFCy76oYazRdA8WzGoFTmOrhHDjrfQ7jA16a9pcwMWZpTNrUbrUks4iQg8r9fILATICz
/uMcEg5QtciEKT0/dEidsxOKFudTszEBzuiLZNqQUDt/eDEMErbBfn0X7eQeoQh9ldVZyNc/nGXP
7Bp+jlq2ejhg0k+fgjHhWww/eoryUzDB/jx6EZTat+vdEHfcWYK8zJlD3sxJuJE8eJALCnZXf1Sf
nA6bEjFPBbDV1oqI7eWX7YD2oA/lN6+P6Z+mXznFnyr4Ab2xhm2Xz4nxYcOUviLU/71bVdJnk8Rq
qbUbxIxeOYRX9dMeXRcykJJELSMJAO7u8WLKkigg+mwHv4ikOkEY/tLBgtbsSRlJ+3ctwQWjvRHw
ClCRiOnBeqikYu+0YUs91YqBTI5qYWPUb7c+1cb9soC07zr+u/YLc18g6sbhz/uvwuuVI7J12Uhv
vtBxtQ/CRMy+lKu+QkVavGuVMrzpHMBy09mf9hd0Sx/ee+M6TmP658lr2qR8ZLBgnXmvafkWglxi
98WwkT02m/Z7X3avIxqsFJG5opN5kjd+fnih+uZdCDo0cJ2jAN+DpsjpIzPVhrpUB4p8gaNKz8eI
41QzjCDls4B5Kx5ROSyufSND/F34AjNhf8XW/V+ctDkrmOXdMKF4M8JkDFIauuoBo+cLQSxs4lW0
XQfQ1NYoZ5RHK0QnDCJZdYfHbz4EVVzNmpaffOJj0Hx5DPVdxBDVJ3fzRCeGh/IGQBD+NUweqLhp
bZoa7l/P2z/xcmZGq/GNlSNkal3BJBrL7B5D7aiqQqfzVCKsgMKIFfnleeSRi1/smcsg6aB0Qlb1
HgBuqwuM97SU6j4QIKttyFAxGLMr5GJSnQTFhR1i9ZiyHrbVZNf6IbI71MAamiet2L/dc2zss7Iy
YeD8I8kHEcJAVm4iCf7KDTnGyc/ET4kitpSh+tPxnOtUfv1/L1I0HS+HWB3KVz9I0+zANVOLydY7
SUBroMiAVP8FQy9Y8cguhQe/5qyqbX8FLZp/4pDRc017zA2hFPRFSI1APvS0y6lyxwsz4/W1HdMR
v293qyyFDKy2iW+rzvyHZW2iBocYFgWM9nXbGPk35YRv8WGOUs2jZNef8BZWaFKgYhYGYf+5MOQP
HMjFXuxfoWG5wZO6DclCoX/e2ZHOoatNddYgGVY7iyCbzp/kmFdynkqI5FpNSfSpRVjHaZyyuYz6
z8peJBkYPwUVBt/HXTwAT388FDbZNtFWu1bNshIbNSvi0IDWeLFvA7EuomUIKThl9HbSYf9jLrPT
tJArDGT/bRNdIWzyo5n9DRV60qxiqRctPAx2I37PgV7OW2pwd7ovm6NIAoTuFe7Vr23wVwt43lUq
4Z7EuWLDy3eMU9XoRTWVpFiZnSSx+HaB402Wr7W9qLaNXSVIyt6Sz5y5Uc3Vecje+u2voCxGP1ry
U7Jegg+FMgsuymcCAYUD3F8+UrOqKrJ5XulaL86liPc/5koB6gQTHMxAtJZnztfIkogMFxt+wFmP
UfCoyRxiYaujO8KoyYVb4A2FoBbdZvXa7HSev5pSYV2G4SN6IytVS7zyrjfOgjvnT7C+uQWPtk9V
b4FT5lGaFkhemjucrI4mrxmqWGd8D8u145FnnGZ0uOckl/CnA+CvNKKQF8VQsf3vNC/fCsG06cfp
sT7bacSyENJZX32f/EKjopfwge6wjraEHxZMJLj0PAJlXejhvXE/3cyEMuX5t1kYpgAvCPPoHQKd
i/1cBdirtG6PP04Mt0NV65Et0tFV26ybx3m4mPLfgbK/mF62fs5NN7vvrPWKzMgaGsrwVq1bqhVn
lP7n4wXMVJ/3A+7Qj30g7O0VianBNa8MqEGQKvkW0e+/Q5TL0o0xiOZmf+mZjzGrOk8cDAoZBY6Y
6QNc6ei+TkcsfNRmwMg9drNWwVVhUI2hdMW5jHuAyqvgenOgHEyTYq+swc0x9HTLZ3dZxoREq1vP
4kwTdW07Mjf++P6s0UVfzNBf/pe7n7a4iOqaoHMtRvzIWbSY8D6C4sMcBlPfFdOv6fqi1JvcVGGX
AflfHihSM6Rf7GFdXdAZM2BDGIcDcoXKDIBGqOMCqZGtm1aC519tl83BA0D1QzQQHdno3WHbYTZs
T3iM7CFM/TRUNJ/DdGANh+hp+VeVDar7bizvO3BeMUf12fhAXzSzOzBNmrLeA8yl+Z525VukzbRL
g6PHGMwcJkLF2+r2KK8vT5lx1fELa2ZcRHYSB/Jej+tz9vP3pDn0r0I29OwBXExh39JWUbudsVSF
HABlJf5kcLxEHMYorM5Xn+LGnBhMS0d2MBH5QsCTYXWYUXwn0CIJN0JnwdbJlg30cVU3YUcO6D6G
McogT/D+zzGlHlFKZTCQFq9Hj0wG2rVmByRXiRWLC3rOQn3Q9LKfzjQ8k4uHUs3Yf7wH0zrtCeh7
UiyhOncZCjz5/CXMmmJMsswkpGPVkyKYfg3Bv8FiptDighpn8ZZpJCX8uS0HlGpAdEL13haWPXGu
a+d7XbGMihE42sj1521FtVbbL3iOiSD+jhW8aSMPJe4pcIOjus3PJ1WXOjgQe4jhtTPn+pE7zKfU
lZVpQN7RmBxAw+kCo3nzChHWVbl1Xeyxvy7uSlxxlnViDTvQTATw2CQzwuT+U3sv+hbXy4HwoHWK
jsjf2slwI8P/acAUXfRQDzAxW+VtIwBFdb8Z5Lf1r8S65IdTRlg+tgNdc0lS8l/nTFsf8AQNqPrf
eo1MTlXqQ7u7M8y0qr2oBizIYnCjT93COm5y3dcTacGpeEXVyRwC147AKpY8p2WH78vHO6OwDvEC
1qp4MKdORLXxHDKEyNxazmoYq/X2zr5UgExSNNDUMTv+5WnZxYYD6uJw1H7f1ZmA7l8r2HZ9ja4D
AeX7afwZ5ukLxpmSE0GEXsaOXnMqd+tRZ0/2sMICqbDt3cZuG9hxFBpyRwSX3W01dXrvFA7aD+Lr
kzNgtK+dqn16sGo0EoT1z1KGgwmL3ms0N8lqbFvXhwcpuQx9bOUENy/Y2QGWkwMCeVtoPCfDq8c0
/fBHwC3tneuNMLztzs1EJONtWQzR+Rn09SjHBowHeRSlisL2ta8s3A+xPEZc2jRVbKknZydyEfGC
fem6YVDi1XyqWYXUB76QvZLevw8nfW6W1nHoEK2x9mb/fLYwuLWo3Ln1XODs1/wJekxs1CvYcLVf
iMlR5mFdl5WRr75RvjfhYkNKQBg1rgtlp/otjXfWUSeMyjO9XtoP9OQZP+oP59D6zCZlJa/3SF09
ObsSGuzEdYUOsgT3wCatqeZnY7gVzfr4zzCFt5v3QucXJGfXChyShm2qFwayeeQYsms4gtWz7nq5
uAnrqcROm2Q+sJUvOV85822T3C3QAbz7cPXT8juCEWLmtpdc08NvZnt+OmS9oxcMnaxy/rTwwujT
YGVJY+iKPK2ALqBCFhGvFuJlbuu4HLQfd+42EnmmG97MU3AjJ+U/QGT7LZ3DBZh1PGEgWQyZP8sw
Zuwo+aSr0/qC0Wah8TpWXHi57mZgaJSnP6RFFa9ZNREK+aUSEcUpzwXkkfpUaqWameBaxIMAOzhL
p8raduUoCjYKFZ+80Z+TBJ3OIofVvEFTmZGQpRTzJLQ7f4awGTPINzQO4y6LjQwjuz0bMId3QPe4
qAdOWa1yqZRBHzpWx7Fhj/ONHBwTDfjJ1hzRo69MS1Afl+RwttdycvivXBqTfL7cDJHUCzA2whX/
BLTPIUq149MmRLHsQ2ZqVnEfImXe3jLQAoH8W9AJJ0+H7Dph6pCrr/hOhpbEqORkAfvlHXKTKhEJ
PeWG5B20eERrFN7mx65MxuFSbLp2z6Kx8OKAkc5A3JCMd7iuslJwV+9N83nfseOP0EDIbDRHlNpM
0YndVLjHAGPdBaghk8eJ9bd6rezwwoPKxP9u9BTa3WU8hzj+xPu4eDgr9vFZ3zp7fd9xSxNUfuCH
fXBXWzBbEikCdMbuUhk011CCB44aBmwvzTPEF1arf+LE0lukvWlSgztAuJj55LdSZ1KG5gGsreZ4
x2QKfvFa1lo3azI9BM3rblwpQGYxnzkS10n0S/KiNacTSIQRfc0nGdgBP3NhmL3nq3W5qqeTj+vc
67RP+KxJ+fKtpIgqHhw3qNsY07STunxJwWkwVkaPvdMW1ZHNyHGShng4fyL/BIYJLh3qoH2H6zdh
4sXbBCapF4f9JBjL8QlmqcDMZ0TkJ5Qxuyx5zG1I49gRBmVCkTE39hE9yZS+P/Rqm0eYMOK4vL1q
R/lAtodKRpAa9roouAlmS6NhzE4vR9GHzFtBmwtbiahEdIGfJz58m/IupGT1C7ykrBk3vbsGpUqz
Uk+rYx5qeeqT2SSUyEjOrxU79UbGwT8nchPBT2JcWwpQflIOcl9IduLbqtjECYFT7JHs2Bd5KBhk
Kdw1EgtkoBhArTvBTSBiDUMeuq5XbBhjLiwrUUG9CLEGi7XvCZflIe9wPjFBEBdH1a8rpVrXXnRr
ISIJlahVlm31Wod9ZkbvfBwbMDV9FL5a3SoUfBoUyG4f5RYK7HwGadUR5lH+R1t/FQJZPOfK/pMj
F64qSm+ngwICG7RXkLsyCGUp4ePCppx6K9BRuBWQ+Mx/Ghca3sT4aeEjr2d1SDSy+wfTuC0sIlkQ
Htp2nnU7Xtk5odFIRVsoKIrImsy5xWHvwZWwygKghFdGMFzOSQXgqOkwuJASZTHexwRj1hJPyOKL
T75sn315rJSanVlptreEamqW9XlAQuLo/LUfaLBaimFy1uKWQ7Vh6IiEUJ/smU0BmxbvGKOOB9U6
zXBeReRC0EcVwbLXwdHHkL6iWNEj9QX/BosvmXY1aSzUPSGp32Z3mvf+aiMBFBqN6Tgcwdtu/LVP
DmMqb7+Jjd7u8GAHebl13oqMzAKyUAmlNd5x20Qtlp7x35D32IKYH0bvDk8ZHqB53GuRV09ZKKdW
WmhYAYv4SB26v4lcUCOifCtO7oCjdvTr+bTtGU8PV++kYnesfvMjtq51B55bl4WibKv6b3+H48lX
MpsKocmM4QoNZqJuJczw6C6nBBJ2J8FH7UqQpLknkrjW1UrYQVKgJnPoohmrJM2hZ3hmuNSlB1LB
Ft8m2qzaKK9svNIQ5ktQhu3S3+WGzRtmnUCmJ5C9+x9lNQSPCwsdUBauHE5BGXMEdozCcgf8XcMI
4bAEqt3xaoCw8Xu+OzDuM41O5ZP90uYGFfTx5mxNHbPwIBOb+CAp6G+lalWeIpbrO9woRCffVQNS
EbTSS7A1b+lnXXbgH+n4lvuf+SEgiu1GrUhRbjQ3lXFF24XJnoLXTq62EKIffiySqA7X2NAB3iTP
rkeI+9EMn+GVfmRgjYAdHbT0iu/22v4ECG8OHOoWT5hdroRfitWzMMD1+FybkAfPEWm5BnusA+qH
sMMhB0bAbaB8D3DlgPPrnN2T3WtNF2M2/xx6PRc/IeHSW66Hn8t0F0f+JC2UdWMrNnE3ciV//FMb
WnEQShA8GQTeP+PSVxOjI/8f0ocW6+QhwAOKMEtnwBKyA8T5ZVmwiMuQobA8iS/PezzMgw96VuPW
Tgd3iYNrCSMDerRyrJj2goTRl0tVcjJzI9LqU6UwDCSScILiG2reeh9YmWmWqO+E9xHGSt51vdcv
/yFU6FRR0/Qwu4FqUmY/SmTIwY44MYF70SW14XlT+yefk/adZGemM2zHaJPPjBn+vhJV8mxWulO1
gJecb/IWbJE+Zpe6qSu8kVII/kcNccn0d+fRfyzTOy54ATvwayjgnyl2DHS1W5/W3SJ83/f4s34i
7xjIcHeDFuFcc/h7kN5h2GANRbdmejvNzDR3xwRAYCQQUuTXtQdF9TJ2ImKsCf9N1H5e4RlHxKR4
tD2rdS4IwiW59396/mx+WmOaEBjIO0MXsjtvMraoZewcJQ8jcv0Cghxi4ROAwd/u62RFNBIMfYDX
iWZshFuDeJnz8QUqP/LgINAfwkLBqu3AR5bKCr2Z7zBb46O5u4q9XXZnj+E7bGCABR0x2fEcb387
gsV6t3DGYRVdMNMUXGgRKEdjhlq3DkncQtOAvV6WrpT/0ow8k02OoCm5qAKOajVgUFrXGbLZwiU1
HiQo2PsyDZlIw2cjB7Mu/qovvRGAkXFTLfsXVB8o6gj5DppKaj1oTduXyibK9DULXpv/qWtIAZWS
aFv71dTq7xjApo25dcods/b+GssoKg6MYw95h7kNpOpfy+wWhQeSQM5gOlKtp9qG/t5PMxaCChk9
C+SCiFNoUyYkvM1w79rH+k5ZyNQojNslih8wvislYjri1hZl9085jt7WIjkTa60aZ9eSD30y3vFN
EBX409ndda5lmd4CyafVyC+v0iGLseQxtOaFqSWSc08N7MnXcH41BM4tK2vilzlRHV3wUxPoU65r
Muh+AyFWmzmBmkieQrDKUpL9hPQCP/6+O+KvqX2CzC04QhX8wT0FMvMVcGyP3MljdAQ6ng7LKYI4
SJYPc5mB1yJ+zaYdcJehfErSuYzVsPPfJVAKl/Fm882XUIz9QBXvULVfozVgPjSE3uW5ymteT7Pd
J0WMrNfwTWI1oIAbQlBjK5S/CgPPJ0dHj6DHwk6YfxVCg5dxI3LD1Fe7VKuqlv2l1KVh5WqV5AeP
9y3zwjjUcuqGMjzgISwF96iUDFGTi1ILIrIlJI8r9dedttq8QgL60+zcbpha9t4T6UzRtqMJtYgB
bt/ZMDHjvkkEpvbiuqLTJ3AAAGQ02tJx8XMmWIkwGZM6aovc6t9iqSCbWqMNhtngHCYYg5T0zLzj
GlHeQW2spWPWZ0z2P7k12pRPftQKKBdcYhMRyZNV2og7K9E8/5UrRXCF9aEwTzwNyrv08r670OXH
oOw+lPV30ovAIQGyWIR5x/v4nl+IeVcbf4Y0PuatzYTwlHhg24uHCLhLCJNImqXefj9IgUm4KJN3
jWCwQXXdC9cZqtqyVKllZcVy3E0CFppEqiyiB3BKthrjvq50h+HIZqK99kGsH2k2vDkj9ktIM3kh
HgJ3vpLh1ayH0k2bAHA1g8sNYEAi3lf4lLV3J76BUb2RElItSIU4qmjY+MpXQMxq+92P26IDXv1r
3wkhXyuNmb6Fl9pxjteivc3a4xjfe/tTX27nco9sxi86AYxAdgajM9lsTgt11QtZii/cMT1cnSIW
ZU04tPYHsNYlkg1Bm6rZrPua+YLuQzzTL0m45BYm52i+EWKFauXwT0dpD2JapLe0OoKu8uB5u7/Y
aykwzfRLmuSPjx27LuR0ocPPlS7+PU4GCwYZKZoXYgi1c53m3/Y4b+3wenY/liH0KR9F1kSCht3S
9NId7KaRsDUyCXkNux++G0mSaTJlPTGHwK/zmTEYkK8upSchPca/ZN85eqrf85AGTVeuf+wALrdW
yIF/Xjekb7xjgbZ7mtSg9/1gmtubDhJq4VgItWvTLrnjPmAIKBiLxL5sO3YPzSmcd6niK5XcQz8t
1i68UWpCYUa/IhgD4uV3H5anj4L76EoFw14hkz/Hd83Coot/pX4uS63wUPEHl7LaoExn08zy/+FI
/XO3oWyzIybR5+Ng3slIor9Adk4kjrZs8aUQOpVvG8kp14MipmDBsVilshgorcwASezXDiSJSptZ
p0hYAytaTebwdExTB/I5zDgU0Wf7OvraretlD296Gv4b1M65tLJZuZT4aNF+JZ3UgI3BUdSqk7gD
7MwgPIX0rvXuUs9ElNHQPvf9HHIQUGVCkK/okVCmZkAdsJq5V3e/fDIdbLjuLw/z0Wt5pjQiQMA+
Su0MnM836jHpdo6yx2O6Dz/ePM36R549hIks3ipmT248VvD2x+4k+X04yGE1Tu0Eb8dRNpqv2c9F
a3Z3M7X5qxVClbx3RpjfCj1H8QgVPmZdnl2sJQ1VAKpnR4/RRRIPDziasIFXsc9F8lFeCcSvzWwv
fPM37/aUx1DLmf5H+UFshjYN1OoCOTKythpDYDgMsKzdhKG2h+7CKSRB+9+qa67ul1iUC0Kfr1yP
UvivurI/vIpuPOGzG9h+eJlL95E/qXeWt949POiJSGEt8wCh8mkKtmACm+PzuN3diQABjNxUUQRR
PrDH5wncudNUVSnSlVHJDy93PZvfn2KtqzYn1CTqxTVDt5fPKjbmQZ+gx5jPOl7fYrHj2ZfZ4dqR
s937ugzY3iLj6W4b6bjCPnGFpuEzPJHMBoaK6lp7i+rKWgV7oKQ2sz/yLIyMOLsVKif+ML/ePeTj
mhHtbWHue1teA3vjkMFT4EKNguuxQqXVcPdhRswGQakSvMSPk4JwBaVfIH2ADJBRWtmrbZLirmfw
RshXm+am2pfCC1fLEzskNcB3RbGKLA8gz4jmSDlD4lHASJMndzeGleorq4f+T5yqDB9LwilZI7KU
8nfEQGHTa9YUquVqiM8YrLefxs7yA3D1+w8KOvmjdlogINDEGD3S5anGeE3ktK+GzrL8CmhF5V3e
C3qUFIv0crc3y2tsn7zDo43EwAMKMxi3Nvhj1S5Cbxvc1cWaZyYN9NPdr51sVo9w/AU+9w2ept5f
TN+nKnX5kXeU60Eu83SjljMNeImqNpCCrh+cDSpstp3Uvq/KJa0iAH9ycPyyy/+zrQRggRxfCVbo
+flnoR1DLUE/f5DELhdePUXnI3euQ2w2Cg5fZD4s6Os7Jjfn/mvA2OEtIhbWa0B67hN3lLllW6p8
A4Q14gT7TDRV6z7vFo1/GEA+SXGLNjQnIPugd25FwOIvWx/c/PS2qSGz3bmPsxVSb+aw7Y0At0VD
Y+mUS+v+GntqoVZB6k/se1gLHvRbhvZ41wstd6xy6OyNDHH43IHfzlSXSwgzU9rFMv6dUtaWKPpY
TWIIE61+CToB7gafv4AFKYIKI5VxhOJxOW1K/vUSMaD3Q+DC6fa+xZodhQgk9FeN6LvZn93yYn8b
jHI3a6Tim0dNSzFp7mn/px6wz4gynC5lybOzF6cFHCiq2l4w/kxzKJogJ4sMlLqFDmBKHll1mjcz
tPSUydfvgGKFgFsFoBqg2xQDPGDaofwWm01ql5sGkrfh+D6uSrFpnmXcjN1heXY61Mw/wY7L/aKb
A0mZNEI0GLfbr+SGKdIlh4S8Kg8gh77loOPNfdssqzOz1O2yEApRUhbtiXhNVlx8h8o/LpT2hTqF
TdwOBjV4vuSjrEZFo+TZi4wq/TdK4Qe3mJ6iyBi5z30iecDdaxXZxtz3eZBrn3Vqt/kSokQgGz7X
2f3G9L9Gmt3paFKRHe8b3SCZHfy9KRdOQOgA9r40q5V7vDSRScW0kVzzbvU5JG0mYcUErx2hrgQ9
Op10tEsJSECdUIiHJmZOqw9E6YWPf1WMOd/yf1zEesU9Zun0MNjEn5Cv/8mbitNlRihLmu0HkD8c
FxTeNSkBIfsOCVfb2vJgNnzMRuSt4NIHMBHHDUjE78BD8Z8w09b7eGX+d+YOM+/PM+VLM7pNc5MR
0ww0VLSVe7GV+yvVImvusnoyHAes21p/qYCavLZb6GVTMfaEoJWQO9xr6J9mX916G+V6fij0Fhg0
n6Qu1hrIAJSsudCQ+J8X+IyO79OmCiST652eTVhEvqXA4/u/kZ1DVQC2Uv7tquGtQ5XHN1IOKjbw
EkLHnnzAvWyVmWlmCbEO1tepjaieuu46tdzJR5PSH8Mn3joxQg/Jhb3SZ1iCrFy5vslkbx+ayWzN
PL+qU5HJ6ZFg+rU71o85CjMi05Sp8TXkazEHMu76MofBoEPgR/7MNADdj45fuww4obEqgzlb4ntr
1CxSdD1YdiVWWtlVMGsz3FCAwLu39Heu5ZschRQJw9SX1V2rbsrFSoFwsj6nJoS4qOZmW2Z4jshm
gdivedRbqrR0bJRvI7ZB9G60K0qj0W7CJ2jRuzyFtgS5lh44sSaWt5FHG62zOhj/ekIicGbSG6I5
Vqem3e6tCW7IN1UasbScUg+HJ6n1fTA0QQFoSl9uxsAbVUC9NthY8rRQ8oE0elPCzlrDaQYihk1Z
2J4cOQDvfkXAl28aZXHApW5gOPA2l1jfOhy0LLzrNHOj4+taUVbULJITPxQ579GRZS2k5O+9zMmv
uZZEiK63X4xaXvg4rnPg5MZfwHsUsNFMY28diGHISqkDN/Do0OXsxuE/sDxSNIyZ5a+IuTun6Omj
Lqa+NaPz7lowvJwwOXHwCqRjWgmiIRnAmyazQQIRFqvMLR82n0mDZIKD/aQrd5JATa675HlEEtCb
qyQgsuK+4fJLZIG2MqPzEDY/pmvodTTponQmqRMqLiXvTWnMODGBfNFzotHRdOnBR0bRsbirq3Us
yqER4qIm2/9fhLsdn7OYtt89RqFRNRZo+ZJTQHkweH6Uj2Bri+zUOKrHwdj2/EwUsUDA0nKZMu+7
5j2oD2f/VyT7n2NWaQjnBECGa4gMbGFWZEsQBWGzfMGHW3vzAbY0iPcxkph6X0lq/FOd3c1CJ7AZ
icGlHx90HwBP88hPnm0NXMBXC1oIBu+wDABbAypDX1B+noiQdqnEHLNYUlnMJh5Diufv17t57Rm0
GPVTwFuTwk1b6CzxD63UGpeoRGUYiUJKBEyBa42Koy/thb4QpbtNuq6PoH9xdv/ms/i6dHlV3Qyq
wWay1O90clL7JEykjSe61S9pmCLDQCgqJupqTVgOq0164JRTAAn3HWCas73+cUJiSlDZiNXuxBHY
nGqF1OPyGPgQFu1aGoSCFOe20CqMKuaxVUJfsNzBagyAssuURfsEkCBoohyEG8tjJWoMnlymbvB0
qooc5sPJRxH+Sxv+V5lNBADlFAZg51+MfMrmvgrgknQL0klmsjFrOJt6dgYejKG+p+lx8rXJg2F5
KTs84espNO2BWZBAzgNIDx2rN2sWRj7ff5bHMK1EevJ26i5ib2q1hgBNIsNMhdvHfS0BZnzDuwak
XigcXaZlf81wCy118xR8Edm37nNKuFWtaqRPgbfCUL8tpMVzKlknpBYmunb43+VROHPj1HzN1tFD
/WXSLlNmyOkEzwXJjh12kU1a5I1QI7ms4KM9S/q7WniN7njCBVbxJ4oyR7lLzuO687Enn0Ekj5Go
BXj2z2R+/RxOHgVj6HVNAOck7RTm/UTB796bUYnPRHTgAGCtNRTBMkX5dq2BT74Ir0n/EwiqEdGs
ldj5rjIQFNLFMKP4tHyYsNhctunWAkYA6mCMhKJJWRr5wKA4/Gzig0FrUk7XElCGE/jA4gov1L1U
7jcsV4xzAsfAKQRVu/0sMoZqya+/HpXvlBash5Y18ryVUpeCZ4l426lvEkVoDSc6gj+J/Zb4DXcP
QYb4W8MovZvRPKq2mf9vnVSbRBr5LbZAL5Whk2qvtrt6hxWxziSLJOtc9ObHDt0MOEr40Urg9yjw
YUfeImBMkVMMy7zmnZ1bz4GTyxfNKtaoOpSOnFWa1M2pNhi7mn/BYlSXVJkx9PcD75apKSBejiTv
1diV6LVF1NCsZGED/mWumokUVjT0QJh/qvz4USz3Ka8VcMaVY//pjg63GmYfL9isskQFn0wxz304
KtOpdyqde/w5tycSwk66icicsxskpJs7NXXTw+ZyJNgzBrT9s1EowcHF+/xU9cnpG5K7dBdCMr5h
23L/hY0oaV1/pBNgtV/xYRI1RyLISBx4TKZOod2saBc/QQWLqayfzEkHpCCdznd664xHm53F/Qlv
XxdHQTlDiB6IblEmkd/L8fqrBPt9fDjF+LIx1ZTLUw5SfTWZXdUbP8j5AYH9G824e/thSGEC6Qra
8+ToQcM1IPrfDPzioK2PR7qkgYdsZonCFDFaKP2lwKsejVQaKxpqkOEa94iH3NhVUBpCNKqC+BeH
TUCmqzfCQDAQbi5c7cgtziQfUeyzwrdvBThDztjZFUGx8yVRuELtlmhfb3KFG6SiI8GKInuOXawk
2pUhKaNu+jiOuAR2TltNs4+kjsrQ72EA5FA3NYdXnp3OtgQtoLACJ5+6Vp8KYlmVbQ1pagF4mami
PqoHXZvW0iPBYwbI1ryxGhgQp3spdUxMikUHb9SDdhEbMul66qi2AHb0jLj5Zj2dozKubWypxqYT
TYhksm2ebd9R+YQMqDZW00710xpRsMZqK7cYMVo+oClc/hfDjXoYzjQaqNe5PKpKs4D7WPUXDLws
8MLuYj/ocgvYQBwCayvkmS3yJqpBkqzmV2Ehti0JZKUjGWSIBxhOTK4ulC/+35gYjGDEMqO6AKm3
eMQ2YORWWwRDg3pD8fvdwMfPXG6zUqSTIG8CEKNUhpm1bSieXHgpjPpq3YGx87K9LOzdbVPvXU2U
1rlsiBL0il2hVbRYbEVFPIk6SsR0leCDS0ibqhLk/I6aONPE22i9ttQouHNyg9dI+1y2Ds8VpiVC
6G33mOXFRnC3GC65CsuU5yaPuixjuCwnJDROnhfJM9N9T+Mon8nZnirBMgEMFC/H/8vqo6/Y1LMz
osdnTfYEGslpUbPpD/9RjTZDaDEPYwNYK+urGnsjGKwFXKoxauHi8VhiHss8+LXswS87LH1Rsbgh
G/QcHReauNa+Z+MOS3HlK1jbiUU+4adtTbgDrTG3/BpPfAJkXgfQU4HIuIpOhU1ow3Goerp0VvSP
SmbO03Vf7l8LPm1LufM9AQkgenwmJ9aZGkh1S4QwkIrLVUsc/hYvpaYnCu5QWkMc9ve7QPag84b9
PJ4ul6nDplDkOxETY9Bh2qn9HE/rfzLN0rfH5H+6qFjpCYQlByMx2QLfhGQcBchjDA8dFzwIshOC
aYxTFDfWWZ2KK5Fgf+YIVRRoaLt6iCE6+ZQ3yX59jSiVxw9sZBGL9G3XxPQ9/gOw5aniPwbuCu7G
qR1HzVJPS34MgTrWpzpjso3PlG6Vkn2/YON2fHg6kqxf2iX7I3OA0N7AJr6rZm0AKHh36RP5LXY3
N3+Bq4Uwg6PetOjZ+mjaYpxQ6KT0bNimGYCi9YqdfFPZx8AEXkLzu9NmnJhTN/KHcvMFKfWOhvev
CMEXS3YPr6xcGrfb/cmVi8Isns1DhFhUc+8QXaoBl8+TyGLpyYWLp2aT8pqaET1rEEMEMV7sM1Pv
sgEJNfO7fCA3N7PDcSXYtrNVhvnGLiPTphldY8UmMh/oAfVAnYr+5fYjphq/JT86gdIKVIh0q+uL
33ePk4+6bw93BNFobJsgACLyzg0n0GQK8L2/9lLH8MOfn05DQ5SHoYT2j7gQD/qs4urJBNtWTu17
gXNoYcVkLGxPfuhPZMNed0khSYA4b275GR8CSpsSXCRM/G+qguoPWZjxh0a25xmdML4hj5tVTWeP
PggbaH1WxvI72ratUOTqI/pEbPPwT6Ir68eu85N0IvDgChXvJ5oflU0o6rWStKp4NOA3dLyrWE6r
TAwUPPHPnycQf4wz4fxn9Re7FoWBCEVwrwMA7l5ATFVd8K7GWWX5z/1p8ya3khvt+gW6+Bh+0qIm
R4A+5pz+//FYOE2OfaV/9RkjHwVzr1ErmPdSvu17I6+u3TiPWTES2pVEsLWwYMuw5EMxNuCLKjXR
RDJ5P+AGsEHTwkplJ8XNqzh6z7u7dzW9oU1nxT4ODJTihpo82+87zzIhmd8LPnPpFEQWA44X2RaJ
sW2FjAR1ejgI62JxARjfYJJUe0+ykdjWAKI0KgcCKkm3R4+sYmiCN4LNskp7q+E4YEgPopWD1Egv
ZQOHvIK6aOuINrwqGT5/TUwFzyweGg+RtCwsalPHBNTSMb3jlvjJhAsXE2CozTz36wBF5T+ccV8L
aJbeH41GIzWSLYHE8pRvu+fb9106CbLJf5ks/NKGxNfOKEfvmPtNeJClRlRJdh2aSpVu5IWg/HCN
W1yIRjwD64HX2NkHC0J3WeuTtnjjbTkRvaoBZwh3sBerssIeyKvz9427sd54lgKKnshCaDl1Eu7a
VMJPYN36X/mCKJPwpu0e1RvCFheK+RuKkkuiUdCbDIvburwkydXB7v/wbPKW/QJHA/ue1Bh4qYUb
5Po6tW4ve3MzTZYDXjTyKL3qoYlqKMb5qLFHMD0hwsy9v2o/swxGUJYFKeoG0MOWhs6lYm2PzGQU
qfmiCoNyG13rXI7YnHIOALos+We3j8FzDGB3k0FeKgm18jxvY9jxt29kjB5QokLL1vKEk4tJ8KE1
o54vXTVPnrDJF7NB0FnQXp309YwuP2TrGUH5kSCOZXDkq2ieODzGw8PKsb9bWPBA8Hd0AMh/wD75
WNbCy0wZTnZyOWQZF1HGfPCGiXxXMYC87MGLQT1ymtaPLRFhKJVRgL/KuSrPK0knzhaKCI8sukP2
297qUhD7aeNWzfCPpLznE/jHbnz821VeZgJsKCaDMdYq8j/5Apv/6eEq13KYeBi9pYfb85lfvcjC
o0XPvBflyRCm7+s0m0DPskxOY2pJQN6g9mlUdwcCQNoO5MvcU9Npr03md0hDj8HDVby9WpqVM/Vs
KTyDwEIJ0KNadAtkTg6q08ETn0Fs/Q/s+ZbJA+KkV9UgS3HmbqEhdszTe9sqi3BROeXTgyhp7Ose
E6kfuaRe7wilUFKIt3gIKkqpmPzJYRE7PNCz30VrBZzNDGpljjmTiS82XlSe7p2jeHTaUCEefFaM
8zpwPY3ktTqML4nXhnA2R7xnf3Ua3FVAaVx/0GffitaWdDWbcyxK4z1ozsRP6nmc9VPyjI5IMzsJ
7udZhcqojRsQO2cokCmYRMWptJj/By+BEG/drdrk3cd4X18RjvsvCoLXmfGJi6ld1WffuNg6GU0k
uQO3Jbf6O+YTwDbxpxp1oa8cC1HXpjEG0qJkYxkyzo9NhfkB+81AqeiIqZzmd/92gsrLfX12bNix
b08Ol2DHbHY2wXg7hNCCW9ZoR07bKUkNaSUKiqvnfjFIFSJC960mhWZYmdKfCmrMgui+NZ2WJzv3
BVWVHlKKc08PUquR7nalGYNsMG3tzL+BeJ/nU1xGCGbMtHgyx5qPO9gvRK5EXv/u6Oy0nl7Iuink
i9UJvwtr3dYaMheWiTKYNppmLyg6weH7r+gCYsQ6RRKV9CxG0oxVE93DxDTOlkPJ/zO7kaPvP2xa
zPiRe/3NMfSyLVAUR+mUNV3WJZFuYkaHyzja0blFKd/AR8aXswF36oFDE4hz7ldXRh0tDqJxbiSm
6TKQ3lALrMUu7oe1oxpsy4VFQDQVjPQfZkcipvfVqzZMRKS/B++Qza7XGIwoyJS4T5FFqGZrnDc9
xpjPvQOSrBuDQH0ENMuDJrKxT1ZKtLG/73aBoP1Z5rS1N7zgi8JtWScjYduUQn2ujuIsjovEwpY7
K2/w1YVrr3sWITImYV39Ecuea5s0L8V2R2JILaU/kVuexu86w6x1VSXmycoleqIWPT6b83ORWZjT
Zr+MHDk4BQ/xQOj6B3h9wRSmL4ITIlnH2IYoon9Yv5TMa9OFXLbWeuw4uvIk51TYgKdF9ndRuFYC
a+eBOj1y39yaZfvOMSafcjC9cdR2Hd/wzCth7bj6Pgp+KswdWobe+0pdW78FxqzubvBfmfwth3r6
uYjjadPaau+LBr73sH3DSbDeq+9p8IZegLb/Yie13CG4SX1Zf/L+5+0MqOHezGlRk641k/M5N7bC
o9AkfHUoMu2xjN9XPUQbtfHKQUQAoTCkDbo2nXdAT52ASCr7GaC97XC8Io2v82LfNYV2K2yI8ySD
71g2fWyZJIYFPicsKfUjWyUFefTjXLCk4vv3Kof2lbS5ucmgdFsxZNBcpbuUlK18efHXAIEBgLeC
e8Adt2PKrndoXSknNz5AwN/MfMycU6WhDGuF3Q5oRYZ+bR05zavfC9oKwN06BZiTc/6eE5DgorUn
q5oB8EfOZFXRsL2KEwPSX35bOmtmLl2nhl3BrX5eQLXgylb4Uxg2DCV5eqQWllWopck5G7u2CBUW
NajEkfp/xrAcddEM6xVYOQcxaHImyvtdi7LFFeU16HvLW3FVqyKA5DTtOMmncyyozousXVM/w613
sE7IkNakrqbC+6jkwyBaq4lJoYeV/Mg1ukYpRcdxKwKHGupZ7B7Y2FsK4ZqckABYMHz29R9pXMbO
QJVfYLBWvVEZPAg6zbXYuzv6qJtet3PXYfwD8TsnmBmKAONjfga3grzkumCU+AtsK8CMi/pzXuxK
jBnT5aB3QFLiTxtWdENLAYndGXwdq04i5M8GkilsyYQuFDR9gC+pNdkL7GIg6ERzItJSDCeg81ds
mU1RCTLMwPPYsRHIMeCNrxUqnPYdvdc4AgEF54B26jixWZgkPSzc1UiPQQUL9d79UZUtWgBJZ5s0
XuhBdm9ldVLLOaXVadbqqEV+rjI0n8bVhY68ghb8Xn5CZ4YP3m3xXlp2WMOLsNMiLxx12+Esx7vn
TNEltCoX1zTUfNa2fRs1hyBoCcbDu1eSTXgZHpKzOz7nxKvBH8bwDs3gfOeGKVgyyQFoPeK65AkP
cjifNSQX9hi1Qn9kZ3TTlLroxofJFKnfQoxI1sTcnzV0Svyp6yuw4yvs9ySTxC6Gw3m/d12ARkMw
aplawmONU3z9cRUS9X9Izw/rYzHKpjrSa735QSGvdPlIghhRqjG2sLOwVGyFAdmGjM57qW/wZrbk
8Zhx4MXc+omInmror9tcsY9ah5xOMiOPLYsoo8+g63nqOJFmRi+4TiXkN1ksR2epRmwh7zV0gNAr
X1bh7OkO7bPNEeDnry59kpMeWtlsckiSchgYevpeVscm8xm/3YgfUz8hGF6MKq3q5SpsjbVfJXEJ
Wt/2RnrOU9wjFs29guC0dsshTsP5np9naWZBR2zPJHcCV+J2AAm5dnsSvSQ1p2Ntljpd5phdUuHR
RjsV4BdNxyYx8N/1z/5b2bu5bcQlB7DULjiKXos6uCBQsW3b2zbx/Pu7w4OZZjTyp02mdeiLkuzj
oN6DT+R2su1Tr4sBOLZ6LyhIJyOtejdvgs5YpfrtAYYoR5jjZxSvAebvoFrJmvURzhtQVtkEG+/X
g6mxG6PlXLIVRmgnvoA+i0PskaaEDIETTYfPr2VlZriZa/YFUcIrJqIgYdU/03hYAQ3nxNQpLz8t
sqTKFmHmevfOE3VX4m/1ePwMuQufBlde7BGHGsA7IpOaIk7sOkaTIoMD1SN7qYmE7BLg5TvJG4lu
bVUSnzcu2ptHHG8vG1HujLEFsQR0X27WiyQR0KgNJvkyix0ioIA0wO41U4Ol8rDsIcn+748ugrZ+
EXNlrcl3v/01XVb0RdzomW3sfDgqnoONtCAcJl9e2xNjxkNd/KGtFEcK921ecii0vionS4bptiLW
NiY1d0yj3HiPcfJZ7PuT1WnXD8N3lhaDlkM80IAz2H/x6B/GoXG3bSZB087YvKrCXxKqmPp4Ahfl
8l18xVokl9XKg/I5No6foW6cWbaagb3hYmZp5D+PMnfdiMi84eOckB9z7aPgLOPveTGYiVH65ymi
+4obhym37HzetO9FyQlxBwVF1nTs8Htp7D8ryVEp/AvfxhqYf+pJ6HXeXId8hM04nne5L3joIzZk
uvpVANeUNDTJnpMv2HNs+SJcQW3CU3IU97VhvDva4VsEMamoAhj4gAR9lGzmxCyNKJ2jyZIPBHsd
h0I0SHHUoGW/UhbC7CGV7xXZzwc7nQnFD1wdiWuv5s9iQ2shopOMptSn2XJ4hnMYAm0C2Lncfa0z
jgSCdTG0rSl/rQJ3EZzDYxp/rGBt34dXeOsWn0KoSscEfrMZrQrSWbwZ2A27gc3Rn98FNCdD81jC
ae3n7eFbk5r1QsJylCnPdw3O4urITzxtvLuUDVixR00+GUhAIttV12Udd/rx/IDGCve3vXF5YHhm
1VMU0TVvY6e4JZBHgxzD3+Yz0QXQ/1We+UsRz99usr06ST5i9AcY6zf009IevTh1fN3fb/Sc7pBI
iCKuOUhQ9m9dq8BENkyFuO0bk791MoSXTuFOjGgOuKvGiy7KVpKaAJ2opFJCC7cxv3qSBdobNFZu
BjZUubrL4DgXyoRHuc7CBcAimpVmWGvxvoRlbfJTqAL8Ey2KAjW3OwzOsQgI7TtA7PnVw+6NizCJ
NPYmdNK5mWu2Zt8U/KkcBMmMcXfHWpLRHmu2yC+2V7dU/LXqazVjesMM7hf2TQ+mNPKEBChv7cnD
coudGAhMB3g6f2L0Utj5tMr1yaO0kozLRXvpw7reuVj8HFVZ/qwclBLtY3MhPDAesmeIFiM2YINm
4F9NHHIqsfFEYo2mi/kXI4VX3g21yCX6F3GdIVmKbKVmpt5UvVeaRD1msMv+Q7fiY4K8BCyjcXCJ
XR4lBLqRHom8k3E7Z9LjKFmNyyqxlPKV3rYsCJ90hmLwbDM/3yipJF0j+gNcCf9qTk7FRejXQ1Z3
6o0zJxi4Wmvi7TFeZDpraTGzM/eQJHbVXa4gzX3JaaKHC/P3oBiZZyYZMPANU2qEX3548+QJxElX
KytZtHP9llyS0CPsi9oAUxJI0hU78QD2HDCqd0p4TeXxCBL3YAKpGd0h/7P1p4vZBzIrm/BirWqF
hfXLJzbiiHnbarI7EmxDmu+0Mbvt4B/V/kQrO7uj7WpFwmmC2NlSedmz4uj5+lSkKEJvMV0dcDKL
3QjHB5eoRCweZ8k4BOWXKfdN5rTlCBDmAzYdiieDk7ywDfGZYp2URgHl+wugSbJf27WZg6GNOVU/
v+6SDjNbXvf03Rqf+1XQTeldpriTf67+TG/kJql2cacWY7ldQBntOMDOayJi2oZA3/UvLrH0GMhf
9VkuHqO2vSdaUScXpPsxEGuFfuRL6oblDAX/aCytDR/34brBqG819M5WfvTfc7IVeVmNEzCnS03g
gAqLcsMHSIa1NCoMJJ/qFV6NFvCvS8CQe4DHU+baNCzocZ7WOtNNxKKe5DGKPOzAhxV7MVb7hPZT
bYM4eQwSkiUJJmfZiYZHxgDQUjkHbPyd16xJTC8W4xhGhHAoZ+JnqajkCSnZZL9bjx3GE0vOSrdg
q69NkTQD78pR7xIpHzHfYHXOhS5rKkzDXKsjKOwx5nSu3GzC6EOb4b6EPVUSJ9u/ia7IlTrJiO4z
pXNIwOdDkwvzP7iA2YS9MrIxxG0VQRXW684Ja6hH4CwaahoJixrOc1GHSZyT33uBoJwog5Z/5vZU
58jIXX9eCFfVCqXT6PFnr3nLzBELoWzLOu1rLG8jBy0tLsvqBLdLwTQO+3pQ9I/5cjRwPzWAAYM3
BlNlM7yLQD2rCHAUfFgsAwnFDJUgj/Qki7aZootvra1UsuaxM73uRFKSFwXvWgRpsfYj2UIUItoS
vvXEsVfcth8dMtTMViopSYEL7AhjLdRGzsh0XaPE+CrLwSpk4Ig2OnHVmI4EfzeQGSima1OIRZxg
2JvMXtEKn/yQem3wO5tiFXcjH95MJwWzANKUy3RoRYw1kqaKumnmzinvzkpONc21JpnGQTEhfQHB
VOIRGROOKdxcsnr31m4DnpfzNEh/pXV6sN5uwYxhDSmhFJl76kdHGw+SqX4Dlj0z4KZiFPKfZQtB
d5CohYKTbmX2W1B0QvK5Ok/zuW6y0cecc8pA8hWhGf18KKbYbjWLj+z8s37TxGugPK91ErARo+la
WRo6f//l0sHhmyrkc9AL9T8qa7Csja4y14h+JpmmpKjNp7dz+T+macL8z/dG9BV4HiBkg9sICvzD
xzFEHFFFQQSGbwoV4ReqTg5FRrXWaqtR7UB5Rijv2/c6AmFXR7snI2iH3C3JQFCuuOu8afhfe9IO
9bjbzgDJtpOlgTs32TCGujbpSsdE0b8FVi1IGrVGHk9Qfcvgs+b7OQrtkXAH7LW9hZ/xeFh7pLGQ
f4p0eN0DFbqwNcuUW2nUIMOMWLb6bv33ejptwYgqZb0IEWGTZm3Q5WgdbNc4vAvWzPVCaOAuWc69
zTAHTphN/WBjGu+17XkEDWNy8bahzo/Wjbjs19gAgj6ykkShomHp1X3r7Rv0du55DfFLNxm5gkwE
X8vvYhvf5hGrdab+jS9Qgx102zW3JSZeG4rFVSrxVlE+JikJSY0xtuX6Oy4/s+M+yhrEUdFgjY8j
7BjESwfMoRYAGhk5A0dVIGpBq/n3ddq1oldiaWDgROxUs0Kz5g6UHOSQCj/QWApMHLwz0/vZcyev
IWaSsoarfBvaRz5ttfAOqkne7u3PXK/okzY7+yrNEUbMlygYa1jnNLET92mypnbfjpbHddvVrcGQ
9i5C9VrAelto2Bl9qKFrsBjZF25knvv6+UgtY8Kx/fd83y5PPsy9M8JyUaTbBkYZouksRIzEbEkK
vYlA/Qbxy6HwxYlelYz31OsqEVD4UtXzC+yCu1M5zBRO4lgcqN4Zlj+29qiUJYSvCFlUEg6zpPVg
BbI1FwoYr/ch8rePeBNeA/0C41U9QmlilfTxfNgduFeIXuR7aNGVcq/Ag+J+IsLL/gBNPGfz0MHh
h6Ko8R9vVMiQtWX+wnFJyBoqE05bo01tjNyEiZg1Ijij+v0qNXZO82EpRdAL9o9xqGC8rkG0lb+X
2XB4mqQuX/sejT1UJlzpMQzZ7AjoZ6DVYhNOG0LgaRlFIhO4UPYK+64kPvXDaPfbs+LlCu2WOGBb
Ed7KxMr4WoQvFnrjP+ZmInQyhnRviOEknNtaWOgAlYSpsgBAmjH+iN4M6+6ex8TGvsZR112aNgIW
b5qF/1eSY7VCWXX5aDJq5Z7cM0NcQI/iuIteczBSxeN7xjXzsM66iWnkzxLexDRlRVbPfiXyBr54
k8WXvaAOILMe7BdDAj3cAaqVFuL4kCM9XlWQ/9ivRnMM7DowuKjdSgBA1mjXJbelpV+SaZ04xnp7
gIf7wqjMf+XfXwJ33dazX4KdMIn7eiumVWrHCBhmONGQvFQVKDhL8j2SUOHCNHJUWRrpPt47hIKG
9b3cfBLNObPdTls0uC8IGJcSIWA1niDKb7x8zr3YLln6b54osx5Oake1/0K4mgChdvTqhS8QMiEg
7ae6OEPiD7iJIakzMY9O+Ix/S1hm0UX9Wf/OdH2buGxjJ0LS5tSkNHnUWRPtoVMNQ8q33yI9zrvh
FZ3EvkBSGXK2lp2mBtHg9+0vpBRcBLar52TUjCY0YpeGGZeBrSBQV48pks13+SBR+vyx+m9wrSf1
NTfedCF7EHgO/+eOddfWzZT1+aS++0mDd9TVA/Eb0YNwWOPLLOWyhM49kjbqSDibAQFExS83tqVa
3bV+Fy2qenPp3Y6mZBNiJrgylMUCi8xGw0MG0veAn9ZOTsiDq8lAr12oE+DNBuhnIGemwif77zy4
oTS7cfH9uOPsc1HnVzXsu+eIeXNznGUD4y0ZCbPk51ahdcp/6Bju3HfjS9kEFIxKFiqIildC8fkz
id/PoP+jhEqBMTaFG/Q/ZJ3s9jsuejjTsYr9z0HyPyW9pQJlU4ZVMXkwCfHvj+ssg/c1jkDEIFVn
6zjk6HPW/Ocbq5njRNR/q5dYiQVDRCVHbChQOCeaFv1h6MVEJB89cRXtwCJsAGQceNnAt6QZLeFv
fdHRg0dwzMCRSA1qi+Ixk9K/G6/x77J/uK0UVDsEg3R8uJmIt6ypn+pmB0Xh4dNUTOod6FK0U+ff
dwK/iD+QoPVESn1NN9aJRGYnxy9bbp/ghaGLpOZWhbGtgDRvIWptYsoKD6Ha5zZklpdlO3OlN8Se
3yVhBZJeBL4yhg+2H5I8lmsSD4OrQBWJBLC/QZndDlH0q9pFX0gjGAE2QbUB/UdRKtd0AFtRpLDx
X1Micvhp122WIQqT+Cw1leoaU0PQR8HycyqzVlnZc6szM6GYssGk/VjH6XI4q/NUoxYS4QUHvqdX
BKWECNsCKlsujjJSuxHSiuk2q2veLPANToSz7n9F6UNa2lMAfg92XSHuoAuwGFAXbmrYnA8CWR+a
pRv2skvcLUVHL2zftDjomtQ+FaFx/O3MHoogBl3dOKoqfZrugffbBQ6zbyVvU7xPGmyIYWRaK625
nNbEAXDFhalTPQZ9LdN9KOAcO/NRaAiMUj9pjkEl3lKySJWnkgNdm9p3cLFb1eNI7xQ9ciD8xmld
hDFz+20M9UcnE/JwIk8FL/xbB8Y8uR/92UVfv/JK0r0suIbaIB9mtVUhBihFziAOURNXc2V9fEgH
M/D8tOJb1NyXCIXj2qFvNNrsWiRe1R4YLK6o6zA1vzanYU1p81s+BO9YZqUqUHfyybm3tEgTs4Ht
guTd5ZgKAdHg70V+/Yuud2PgibFnjKy5jlsn9SOx+J3p4vpWu+deifjx9WEhOCee8H3RCrNJ7maR
lYp/t/ADwzdFa/A0UPdPhQ1EGe/UdvGOWVb0ae5eO4TFhDCKpf5gzV2v8jbUeYD+CoNxlIiT/nRd
q7zRrUJ+rEjJUmwFsjaJe7daQUmT6T6JYMsRzguxMQ+DsUW0uJdi8y624VkRo6VYqszK5FGNLb57
VWKoXbLIkmUg8WJex6Is59m+z6ZmZ2GE3+GKNJci8ZOtK+GOtxfDWD/h2RWLZ2m2iz/cz8HpDhmX
va6mnkOZSXfFZ+aISknSeOwycisUL/lh1p4K4buuLjAuOE5r93tUs7coiIhZH3uPX7UDYNA1OnnH
LoWl0YYnm0WVteEifNQ2kb6KU2KsleB5Uw+bOD62Q5+jHCvXhusxDZgssuy3LN3mp75SlnjGvUqV
FzdZ6LSH49Kmpw6/t8EzgW9hGBjmCn9G8e6BhAJxOVbjYC8c9c/gwDrCsw7gzp6ney5v4JJ6ySmC
FUV/fRswCMhZheum/XVtejwJOO5st+NHbBuv0Gwluaqlk3LGOsagfVxj+HYjUxkFswJWbtTeoyEp
nNwNwKgba5UzgKBowkJdmgKq+0Z+yLSGYKQQk7VLoiF7byFjAlFBe6jr3QWuOsWCjNho2RW67Yk8
Zv4teKTnfXW272VGOSuC1ZtzsbpX2QkJ1s8NmpXS4shXIPL4YdTXtXXbQT9kz86qc4XohD7K8CMB
ZMWK3cAKmiRt/BU9e+9E5GW/eczR0VBiXOZldo25gwXz4JIMBzfd9umwTkMIGsyMgcDUAAOyjqkV
z1CW8ibAbidHK9MtbLnStUhsIoyH9eDLN6y+pQcv3V8pC5D/lEuo68JdabrtAb9vdFCQ6lBjDsgy
07RZz2U3bszoCNSsCSbnAhQhWXPXPBsSf8AYJhev4pxxxLne0AEbD9rBoL31ji6dS6LnlvUHOkp2
EYSJ5oeU+0yhUGD+hbaJh0+UoRxeE+7UIhNkuw0OFbdllBjK2euwW1OEQEQL+1ajyUhjshmx9Suw
urlsYe5DhviFDFd0IigvHrkI0+eBiLjoRTqbxIB25epM/mHklqA3sxkJgKyNyi74eL3KhQ12rfS1
XSFerenWX3eOsm+cDjthaF8chymHR6CccTu1JeW0lrO/b+hIUp3tJcZDmu/cEDMNTvmqRLZWge8d
8JIFFo5IwfanPWnn90O9JX1vhh2eQ3MGNpCFDQxiDQUdPGMpUxE1a4PS/30sDdxKJajNOLCCFZdU
9svpCqFtjPaN4j9ISJEHyJPLHMW1n8212nOofKUmG2FLmYzThqFTyjKejGuoVFuFHXQabPB0vWLP
o5DRGjxa8ex4Vw2CrBp81UtJdJIssROqrIGXRI9/ZqsEvgezsOM4T/zl2AT4e2/3MmyqU70jgtX5
Tu8ljRiHvbg0j3F5Uulq/mW+jHb5jp7FjZ9vGEdIsKjGfQ6vU/I6GfeTyvDMiL6SJD5UwGEhlNtW
cgspASDSDkmNzYjKyXzMi/UFQgDidh4pBqUq7TFWaBsFHkCvEBEzS7+TgdURibXHOU/9C/FcOdYO
CkkY9q9Dvl36NOwlZ97g9DqMpgU2KgpY4YLRjNmPK67P7Irz32sidVUxmEZh6i3wyGj5Vp2EK4h1
VmrXD0RuvV909KcXso4nhiPGR81B1gkc5YUmHB81lkDAarVdWEhlVsUksjGFhvHOhlOYdOeG606b
Tub2yDJFznvltIAe4zcVLXuqvOqFkj2I/TxrvAktTdhMO+bZNuQW61kOup650YvUY4GQv0tEKwzy
T24LPfReQX//8RSsZSW5b5LHz1DLdEAPBQoRdMPa7V63Kd21JKazaIt8tPel4FcG/4vWedqZGYoC
3NmfCXK8wEPOBvnhVFoDV5IT9VHSBm4sF8cvMp5LQiNJBLjsPizdqoB2MWYVbhtwBMZ2LJ3wGxSH
E59ucWyfcoEFDr2MIRlAPtJQ15TgPwpGTItyrA1I5VIjCfsYzd5GlNhrF/FIrTSP/06WGWQaO7Gj
1CGJmTc9UhfJHn/CMb4dsp8ykYfPoEHNN9aBQ8Vf2CPXZOh6gj1OXahdCnB3UYgpPN+dbtthDYiS
u2WvrxC4YHmabBAp23HnyUsLtqQny02TExCbleIafVi5MbBDDUzCEA+17ud/YNbZ9AUUbCW4fCTr
MXrHVuM/HcE/KHmihNX63UNxQ/Wmh/qP0zpyQUpe4/Zut/WUPK/kZGSg9cR1THbqPvWJ1RGuJmS5
rr9WCjzctHAMZ9PrVTm0pl1DYHU+r5xhu7edvb0u8PTMtW8GWtmPQgy3+q+ltlp/sBJiYPvuHuxi
LwHRrGfcDyiGNTlI1q//0nu7GpL2LxL+1FgqD08v9nzSAPOfHjbjl0JgQ5Ap5c06jQt/tw9wYvNd
KIlMvBSLXjYwKuMaxPaTly7CXzt5tTqo6VqKa75KeY+D4cJosmnIsydy05zSUeTFxTgdy1pd0h2q
p1Xie7HVeT+qTFKNl3O63fD5iCDryrI3SZJC9iSuPOOaW3UkRoEl4O5lvUuCq77DUEBLjIWfDBEm
IZ8CMLDs6OSStgutACGAlqpak+WA66us3mhYzqrgMc/ReYxAw4QjDn4/ua1eDWlVE2cncjAHTi/6
Ox5i5V1USGTuLrI8WgBgeFLpEH7yMPNyA2ZNvR4nta/VI9CAzfkgKNRnL9Gjva7dQ9a759sicool
Uhizn7x4UZgMuHZPjHssSt31Hn4v/vmYWM5h6PUAGzWT1xfKP+fKvqQBj1jUpcmI2ha5tXUyLOQJ
Hw/obIvRkGA8r9XM2b5/AMGEyJg6WlQzrrtswaaERzj1avMUeqs//n1EmAKgXssNcc4Hwa1nWG9r
vfy6vVyMTw1dOHdFNB763YE3RO8aQBNN56kpT4U2F5YsQEtgB78s7ObUemdRpgDGDrOEFwP+mbvW
9J9A+H/J2Yy/qLC9WVU4VhjjIn3FwyIwoNn6QOLxgo7iiDv/r8z+O6OEsMcwyrpIGyKrzmV6Jhmk
OODsT0YKBGO5Hk4NVfenaWjb9/Hiy83gpHVTamm+48fWhvfAKapgNBjQrkfxD+FINf3z94/E0dln
8jlLL1WJNqKxT2b/0DrZYhMdIjE5PMT+z0g5389xUA+3KTsHGzGH+n65THdmRn60BOx29aiy0Wj2
dugxjJ1PqIkSeYnCeawpUyk5rhuMiSQCx8Be2vGtI+CJMRveCIHPvXG40210kBEB12yvJ/Qu1I4p
USeHhhWlaovc2UdWPDkO4hsI718/tT3uWh3llx6de7zqxiSZmCDnK27Dxkxw0JcL/MZzjfMZbhXb
2eF8Jd2T55bU/mqQbPSN/wwONFmtowVg9NjcKqvNmxwxPKuSzivmmxz3Kw7E3+rST5avb1tDfvte
lcuDaEP3HKn8iH150e92wO5EMlK/zCXgR1u2yEoNU7zUoiA3mB4VbkI5ZC/NgJWz87vf/TxJJWW7
VhmCZv2JwZ/dw1KWMUxHma7zNn0/Rcfa8ldozDHWYjO9V6Z8nzkK0whAVDBXNlfvctimShlOERpK
4AqyJg8mjHws+mJdz9FIWm4tutylcFvL4zsjwjvv3nf/DHpAJFusA23HTXaZ4/AcVfQxVv1kXHb6
Akl49gF6e7i6HmnTy17t40TjaWrL/Ofs7pQP+m/OYdDgXv1COCSMCJz/Ln7ihR+OLsBkDKhUgsos
JbBpSJmS3tSDo17t1aAGWD10NK5ZTZkVHmhYfILal28I9in9kcBKV4bStfI9IXyIM/iq5nwsaMO5
pnq2unNMg+vPQnViu7qj2MsgWz842F8VeOYe8vIO5+IMmbHGm34QI2wLGc6/2j8TrZnZWzuIbrdh
lBzZyVNgkHr9RLY3QVojvtAgTrch8bgimfb7WCozqZf5UW3+8SpBKLr9TvvSnD/ajJjy3DzAbYiZ
AQpQkHvRcjtjbC0WxgpfYokbaDx/tejBrVbh9jgpY2u89u/H2m/+bsSkn9FZuVmlFW/Afv4gEwUz
67ykvM6PLnuHhWS/tSZwl1PcDfZUTzx3BOfJN9AcFFl4W1mbdoY7ifr58IBg/0B57/VDHxABajzv
QQaPQB0S8VFO+MIbnN89d6ESd2rnRE6h9wSzadKzGCPDjIlgEUPo9kIEvsupxlzsyRnXG2i0SEkM
jnxK4e6IJ86cmVjyj2wMk/rh0Epr2ck4lLaEgNdh1/iPS1j6n/YHcFSBSCPAH3Lov9oFiOd4rM/k
68S95CKjF6+u/b9A/MPJY7Shd4qUKSytxa3K9B4VTwNKGAqy1syX+o2+JEHii6f8+UxpIgrHjf8B
WZX/+pmE4XQpqzqUdQLBx0ii85VU6y4T0p+GGLnAgUPRqvyv/VgVp8EjJRn1udazyOKKzlje/AhT
btOFiTnZj+7KsJ0QwDlnk3pX9+MjAiPFLGdjC56cNcQuo8L8awLaNvhYQ/4RJPc651tDCN5H26ID
LwEmwF+mwcPr6S+NTuHb19pT2sJ79M8F4G/tZXhdPn2WpWTlL3WWc14HPnZMRA1HXTUuqFP1LXpI
42UfswztyDX/eouKp7VMCRkp66y2MSRzTeT+0qAF4mH+x+ZJew3AWALWj8iMoKFRMGxkH0X/r2z8
36mhXc83GZ7Dr6e8J0F1FMxv7r7ZoVKwPK4vHLfjVxqQy4cZWP1lSpuS2ew3ihqU2FuvRkWH/qfN
Box+k2O3etvkWCPpt/9RyerMStqAvDgKVnTmdsrC+fZTCdm3Iv+gdexmXF3SzFB3GKe8F1NlRaOW
+CQdeJ1qpjS72PmXLgaXH3qKVdYW5SvKVjjGYQjCBBj8Lsbq3W4hk3e0THJ7sWlD5J99KWaKG64N
IjtRQW/8Q1dKdfhmDsgWKI4r84D7OM/pFoCBf5Iy3+EQnJazni97kDINovhDQQ3DvDzsFM4Mj5R0
xMW0VUb3x+OsVfiPht8Mc5O131qg8E9qKltuGzv4wPolQl19hP8pcYgn6p07/d8BLTLgqgGD+HlE
EzoZV+VJPBXUTvcvTYttSvwmvHY5jqPet3XxLV3xEoZ2ZIJkz2DaAJ3xTSqj3G+Jodq6FSeDSK+a
t63tYuDIe8rkOEAj3N0y3F/Yh9r8AmKoFehxsdG8Jo9ZcphB4qrBGyewUGlANW1HhIVdth27RsZ7
y3Pl+vAfuAWhnD3b4hN6qlqJXN4CmfF8OQHnwjRYP2MtPgsP0hl/KlD0ZZrTPbKDxGBmVKSX5Dlk
8H8cUBrg5/buDSp20l98WYaBmH979qE3ag0ElWnu+5nkYnTTz71Y8JaqzyaRZfZq/GMdykn62OHH
doPvJdh7MtBxbM6byLXa+49Z83WsDsdysvtm6wZTOozJ73ou0A/CqTJZlnOOI8qfS65wZKaZs9ha
aqKDvvpy/4l/48GBPe3M9qshjfm7z8/C5081tG9zyh/cA7DQ+zHdN+9F04KAAFyW47rKTSnugxaq
5jVtm27ThqvDnupipQcrFTvh2T9wrrRmhBbQR4ZjPViYoRs/HTcnSvWYTVu/SovIwXntE+ly7Fwn
KVw0Gpw7170PmjvWhwXtCkuo6hqXJ5z463dD2HG3Cc9T27H216M45jpxhu+4vMcLVNt3uqUaHfIt
TM7kB7R6w0CfX0wfsRvnLSX6nhxBetiMH/vIVyb9zsJ5KEgC26/lx4jJGkN4Yoec8YtUFCqvyelm
67918127PyOkbheufLQgIeHDpWBiBh8xwKwn+X87H1wZ/I37hlqMrGxRid+C1FWowkr/iV+lENl9
BvOik2JMDK1BwQyRH3JifCKZZNGbbmKsIgg3vyyXA+LweOE0knhxY4VFb8ryn2Z2nZH+Pem6LEg5
hZ1iPISb1FY/kPy1jJchLlMK787Yzy4rjGawRcutMj6AHOsQisJOkjul1gmo9WjT6mvLxmE1ZXcF
LjwVHhMvO7NxG61AG+KlN8LSILlmx5Y+q2BJGBAQC1u2KeJ9RbDfVye5zRti2Yxg/vO/rupWgq5f
hysPJGpkqsOD8LNQPcOePuqjO8bHR3tfZlb8lRvwyMN/JOrnwKyuZHlxz6frU/C6S3Ehmw5lcTo7
jEBmKRWKe8CH4BlswcnIW2WgVscCRjKEGTMvYf3affn67aY3rJDGwe87kMAStZeVzBp0wa8q6o1H
bPFGQtvEkdJIdNvcIdAbKh+EXRlEaaZTlgQlTntS4tWckvl0mmV8x6TCu86WcxYk7ALMw9qTifyk
4yh3YykD4knqc40tl0XnIkstY0PwtIWmL186SAhAuyx4c8ibQHHyMEKFC/1psy8hM/XpHSV7XMin
brQHjfTRTKGxIAVkCfrQmJchjlp+GrgJJHKGK0EInNocxpRAFEv7TWI6zb0Y4J+oopyKqCRLt6GE
c0DFDKXP0IAydDnCjoXLT8kV/6InWnezC7PWako5fsqZ66qc9QbF4nqa49XxrGqalnhtFEeEND1C
nsqwG5pwXAxB3ayC+WvxBD4VG6n7q8SCSfNIk++WkzWZ9inxk+ou8Au1lckxjshblP4T1lM+ZwdH
2xEqcaNoYUpB2bhEjJ6gQtJv/tt5229Q5sN8Z4xQNSZeUxDUp7WzvOibPMaPXeUPSZ03szQX/Hy+
clwGWo0sg6frhznnI1IbNaYNq5K0pumMEFN5TteTqTBddGK/ACISUOZs34UMkKIMRJzGbJGLg6S0
+IBZPxP+/dps8V4nEJLtQxfBIWaSGSA6bl7PJoje7KFNjNgmrbx53eXdlF3OSYIqNTbtXL/RNKNq
d4Ck1PifhvF21GvVpdQTq4jGQvWUS8Aa27ExtFkFED5pu4KxAnx6Myihra6gQMt7sLZWUampjkg9
MvptKAJYihkseIPgPfJh8dkRfAK2VvcYT9pzQ+G5SSyAXrI293OTm2USnm7HnZzBRVPmfO6AEFUB
o+LbU/P3HfhzE0BHDJoNWw1Y6NLmE35ZN29Ej54e7/d60Lr7mbJj22wVtP6hQVx2p99XKDlsBnE8
tcCV8K4wSZMPN3IGDdlOTp4GNk7Q8QyVxzRELoWxM2BbLskUBefr90aprK0NlC3fqh6FxpxbEAHs
UqEL7Q7FIcQ2JV7Qao9Yx1mVl9xDGLUprC/c4BHdpd+eX11mRUFY4QbxjXfAJ7Op3Pkg0HIQQ40z
NEmL7Mwll6JDBg0Fh1DSGRVg/8/Rt+MRoI4zBSCeZl+3ei33wCIoRkBtbo47syNawvITJo4vwNWy
Jkc1TEcydS5VK7kU/NS/xXTWA6UykHeLm10UhylglwDOj0OiaLYcYWspPM1M+3qHhN0usWeE3a70
NLCjDPvXisbnc2bCltabsRX1rsQhqZWrERhVDNugIDNdesvG+PBdFwbQEEAUmWkehsWJjNJojHMy
Rl+XDj4QPYjkL4X7LPPCDHI6Y+H81ArJVSxG8FGZLmj9NOQzbhQFFwgjhluNb9e0Bplo03+AT1oG
3cjlXr+rKShUIZSxlu1mzKpbQlEge7cRQ4rllWlC+utYDdOaHR9cdvldURFzWH+v43eoN1YwlRzw
F3KCWV/RY/2VC0YSbB9nR94cUh4dw5SXTBP1X3cF4KBAzalyyeMQ+1Y7erreHdDjb1PNcNees59a
zKLiFW8JtKPU3EwAHMjlI7fQ8fe2g4I1NrdNfORa/zzFgr281bgMadXnlCaYzt1NTzr07CaNMJBa
sJTcm3SvEsNJ0lExRUBifI/UFSXwC0rAtnpqwPzFjBJ/hIL2rwYcrrEd+4+VlaX7J3cm9BUMtsQ+
NWnwE1tkN7wZZPfXMkQe5bZZqawnNQdI0kAVJPkcK6TBp3nw+tEdTzE8KfShO4/nn5gzHyDXyA65
BY5cLUfu6DPhOeFKk4Nz70ramjmtcJ39cILrwR9VGy6+V0tIewilJGYNZkOsc9n9DoJs1CglOpgX
+14h2DOil6WfJb51eknhP2qV/eGkg/bfkcF53WzLHtBiGHFIa+5DnRfUDArgpxoHEn8e+G5mtwcl
YOOiLl6iOsagwtA6L8C+DlRi3IujSXqQFd8nKMKaIrKeqm6rV3qVzFi1Uae1C5KLgJBx0yZ9eBlQ
720zSjhKYT/q5w2QvljYKC6vuI4LTVnEB5q2ssXM9xZ9so5cKvDMrR6YZJuSrDnQ3CqbZ8GkAYl1
qu3CC1227qkucK5iTAQ5cIqm17ShfR5rkPNpi8hY4yPVPZcMpfgMxltbs/aErcdFW0Q7j76vWB11
ZUYlldBQdsJOc+oM27iqlSPmYRUW64gLEAxwYvdB0pINKXOAosDOOdCwCBMVMegmfKAu9b4cV12N
j+m103NIzCloixnezwXr1Ul/7Ot3HBc3Kac+fXsoD+cE92zGJjfR+yj7fXt50g1v11+No5R4QOzW
7Jz0UY4MtJ9y00ZXtUwUxyrZBl5CpAGA23PbbvmDKMev+zoBX8cKRzRYpAlemE356bzxp2Jqq+5k
wQoLG4YLWY6QbYYEEfrNtXIeUchJi/hTQ50+EqajhMMzGcXX6DAPCsPf2kz/u1xJnpOok/FH2/qe
ILp/qhxvhsdCNcRHztVwwNYYT/WgEScp3o7YNP3LOPJa4vU1sA382BeW6I/iGm0W2+5UADuVqf8L
h4miSGz4a+ZzTOtZYVb2aVE6EIufmqzL9fB5+MGI3gJWhm/OXY4cAIdATdfYe+rd+8OxMQ3/k3YT
yxnhxuwH3Y8vFI6sTb52kPXR77Zqxk49FCsQfby5OfG16HtSZTK0i7D58jsz9zgVNYSmyL5JdNOF
POfxnua9xD+WQNcxkjI9NbHUIseM8cuvBPwFoIcxpkuSCY7LlSHjI7mWL+L8TMopIVSM3/oHDqY7
WHcdoZxu91HIZSWq2RcOquHhVjITqSIQRumMPi6ULuLoLwiRzXf/WIdE+Obms/oCDwdPaB+vUcNm
epaiUPEOxxiUi07KTNiwwvc+O5KLibkTBiWCJ3qZVh2FScT20LvQ0zGzv0QEensoV2tskq2mOXkQ
bKwSUJdik8cbG4V39/rcT97QNQsyEunfLjLBK8IsotvXDniu3DyBgSFRbwEk7fSpP6gaf0XDZXw8
fTvSsgF4aexb98sx6gm3iJhG7HeOzJdJrmuQaKmjAiVJWVYj1ecHnFoXddFWx0IaZlPzNrEwJtLH
6hRYlYMpQVQ9z707RAFraQq1nVeFIzQuGGSB0CkDr7ssCMFOzg95MKIrVeDcU6R9V8aeI9ncYRfF
dDdFL7prkORJOxjwOToNgSkrLNfdU04q8fJimGkyj155sVXTG4Q5lGwufus5nZ5rQfwuvNi6MPTF
ZK1QhDFNDuFeqjQ3fKPaWPcihpfyz3CAyrhrmtNXWZjD5NTUOCEjzUVkDN5FyCNT+fZUGtTcQouB
HARFMIZhnFddbxTCWQ2f2sQMzsD7jXdI1hO19Tdjf58xNDGZmdGQCp5eeslZ0jKHUPtegQaMim8d
LXT7wouMjXqeuYTnIkm9hJBEFGLWP/b6tYmzHcDGTO8lQVPH3CsHZwIzndEcmnAEtmH9Q8avAcqo
apl20QvKZ+ngFNCZPUnkZ7bnE/5K2hQkD22ZGomyXnUrT574rOAMIRm/16wcjn/UcCUC9V8jni7J
pdL8tEriPDmzsyhmj68LxEdwb5ok9wXBTnZrQWW8ZalPpuNcnN2bPcSQQkvixJWBshpe+SYJEfot
SLviPn4AyMHEQQIiwjwdUwQ2DFRlcUsqJQpXEtTx8C0gZdVV9m2ShWJz26cbMAaPcoSM2e2FuH3p
obsv+PcM+NwDQqRcwpXO8Yms62Y29SqEdFKqVo18QnFSMc7UjDafGYSqkT7LG578kB4h+/6vlKCo
IfvCo+2ctFgB0J/gjj25xygNfVYHoLPhf7pVQL9SOoI41gbhhQx6W4ifozBeiSX57YQzWrsY2sji
Z72BoJEd4CNYCd4g7/4WtH9yB04z3v7U2A3mjHKGmBVPaogK7azhSdj4LPhOTmUM4aOzVmF0pamZ
wu0sFO9swqwbru3gyWEzzHqpx6n7816hqkjPFvZ0PhkQWyPLuKyvUY3QD3IulX+IpXLTRA7CZ5H9
P8LyFZMo3fMlP97rM3YwDetRQuVDCswwXy1pumuDPv+h9REgFkD0vSIX3qKCCZofpQWZLdXYqG6X
e+Ze6DtDanOyAgU5p2ZFTo+qfvHm+JTyFDloNf5EM8nrddIlVbI8wEqJE3mMwHTBLQ5aSKoa4Qfy
dVJTblTN/DGWhChp8E2aEK12uJYITW/xZvxiwegoM2sCpnKU2PV4E46GODRvrpxsUDxdzexsZCOd
uzOjJm8sTAx/aOBlQjpcuki+lsgO3MLu/NG23Jbtnua1HuvzvAX//je/Zm2ojvJtguX58eB72Qbh
5aJRd7SenMkxktYcw8imqgJHso+g4QezFdK0xT0nf38HwXRYLJMbExGk1kI2k95Dr9oKiVW3gv91
X5NGvMCvKVnT/VsXaHQtQTDtCVJW/IvT5H6JcFQvMU+tq8ePGBE1OsGJeGuyzdxRI2jQyD7J03hc
Yfi2uJaC+nekm11l8jNF23Cb6u8Xv8CLcKMwPKmq6WMziOTUTIP8OLLxNOXpCTzRkxnrcaMcukd6
a/pkS2dEAq8Vsa6AF1q49eJ1p6x7k1pGob7tIE0+AqQjTMCO+7StBummPNQrC53RJZUOgu23XKvY
XY/Lqf+xSapUqJQL47Hn6r32IR646bEbE7lrq3zqdPumvCkWtGOu6I8NVgZ/Kk+2wIj6aR7AI7pX
+ZsVVRojyltMtK1Y3CO+3GblBM318JJSd/qpDV6pRJAfinw9xI5UBrIWd9Ix9ZGTLCOOOBPV7c2E
K+SJZj3o3YuPKmCE1KJlqkLuBmtCXYiHqhRu2U21EDUBBxNzRr2KWGV/eHHe2nUhEImF1GK4uxJu
YYD01aKi6gwFwUWThAhJRKCcn4fDMLOA/sgagXXd0SRFaScIBlrjTtBZIF5SDArhBTLpFTyDG8P4
Wsg89AK2/z6hpDL8qUuEsEpzfabpBrav64xoSsK6ELgy2yEXItMfqhJ6flU5HnNst/LZGjIHqcL2
4Fl7BFMtHI54gEw59qBi/sxLpTcHEaJktJRonMZfq5K14K87qWck3w74BGWhDiWl3UMDzFVnTJZO
rMF6k7V9aor05+SQbS42WISQmez9snsnWlEJgME+9id6t72YfzlCIM7nyGk0PxIFkAjQoEUCt3iZ
3vHcFNnFgHRIxZFVfjA+gLaqud9uvoxFiF1AObTvmlu0tlDwSLikixbNGmtig10puepkLeFjxxuw
BHU7/cXv/SrRj/Gre++cYQEAB0GCARosohiCmYWeEZh1cnu93jc41h+3za9iYUUwHZf+bjibtweP
VgK+7UT3wV4IMZr0ChNq+wwss2GBUtlyCZ3c4W4B0eQ1pjeRry5iCxe418GoZRPijEG73RGRoEYm
cOOqujKTSdGMSqEz2ZsAarDwS7fXHo+xWOAwODvVWABIwf/eVS8PVofOmT5dj2owYjw9AHKyUb5E
iF3EjNefCYZ01OsKZlUdsHkBUPH7iNXe4Nk4nCCq90nlgvw7w3x02PVjQGRj22CHxe49uN5DHPI2
tfQgBzl8aOKGqtREm6H0eGLwEn01hecSm0InPKEcfcDfXvQN3neT615rVz4VfDoeC8A7Bphhv+J/
w2tiJjRVeYIkubLhVgt4DN5lZpv1Ay7b60r1ClgZhRaroZ5lY2upp/k4mQIjQ+DLBM/Uwf3e03Vi
+lugpyJLIWVPqeLJrFDvHVnSpdcjmKk4m6SHzX2Dk6Bee0YCZDJDj81KGMK4QoTD97fy9EEEztS0
NMvMVzysKiOwM4gA/YXXY+arB2d79RxRo0iDmJtounkkD61+4s23SskdFbmfM/rX7i6JTW4AKtUu
Ei/yRWkOvOyl8ETX0DeiWRhVI8qOnzOJj7FlsftsEs75HQ4DesM0snMWX3s+VxjzBCZxtDIk3rpC
FSxbJTCuZUCM6Mp5MqH2/gpTfNRWQaKMq9C28BzqR2dhS7kbUWBOczzRtYUiccryZttowkC2W8wr
dXObPz++KWuMGjMv8Pa+0IYNjJtj5YFOLzh/C30/0685AMenUjbBaL3cwgQhLc1avlwhjX8dlKc4
82L74S30j81d75XKD8MszFXg7NyCrsbRsPe5Hi4yZX1iJqxadd4uav0E3cd72HJDKxFbtSgnLCqU
6dIWxmNX0wuHMAcOefw9rEhTFoRD/ppMA0353rTqHbnT9f+U9KmUh6k+aQees3w7hv5rjobzGXs0
ZKM2AN+fwCLrU/iECTGO7NxBhKPMCrRWvV1WtG1c8iTRMLRT4HknPnxFoME84hxn5Ru3qlcU5I+I
xboBfgddNsDFm/A6CiYACb8Wasj2lxhLo/ymWJl0zlAbSMRd3sZ9dQuz/pvRRc5mGtkenRj3zaZQ
Xt3dtpaX61c4NpER6f71venjUg0tDsVamsuwUMtuBpkXoLLmtSXRkw3aVb7zdWlljmO8A4IIKZ8V
u7jAgS9WthdD7FZxqWGk/1z6sS4YShE2+5UbB3xupb1T4ukGQEKTk7YqAh6PxTspO+3ytkjyF05E
Pb9IYiCDiinuoIhxG1oOW0RtwhWmx2C+T/ZPy9HyvvbtOIMZSIGQGwBdL29ClK5QwPZGrXjS3vak
3FCDTl+rEzrjbT6niN6p75Ealz5LwAPMWz4k0BRtyXYNtSASpYueHL1CkZLchHyGBHeF9mAvZVdY
gKlzfg/Z2hbfh0qUYUU0UXMN4/eUctR4qRl6yoC0RoLEivP+QGTKrjVCdPWYzq5v/aeEKleLin+W
yPYPdfjBPWibG65EQx2UcLrs09Xr7dSzXWuUgmdFo9kC9P1jOxMaV5lbp139F84LZox5zBA3KHfx
88aMNpb0kOvFKxrs9l8mvngvqn5sMm5/k0Qe5RX0JYatVHJYCGcPzP4IpS0/t+1NWkAFRY9y5Wne
9kad91bOlighdwe1l79BMnwKmVUoYGTBx5R24hhJ8hQzHJtMeaJn3FMRAip4MLfjNBJkS/+YIuQP
Wko9A2Qo/CYxrsLFWSJS6RmZaC5EG7UeWM2tTQSKYZVgMAxtJPs+HNub7dJOvclLxp2KaACeojQ8
LgrKkSDUPLusOXUCUIQY84yQdutwC3UJZiLPdSegdoJDpfKSHrw5kicCKR8KMOaWuRN5Lh+RwDAo
kUr1+HpXdT+n2NH3RnTCCmSXwhjY86wlJxinmFHmOHiiuswMH9oAott7xujYyxohDZWb0Kp139bv
oS/2/HsZiyNmYGwQzim9F7bFfWCHjAA/z97veyBSimaEuyoBnArJnig0O0kRZHNJ/o24sgpbQ1UL
alCp59L0Tn1XnhSRSJrc0R+BEkJNqsL5eyQulpfCGHtFCCwYO5ad+thgcETNPoPq2xuSNMKHY3RY
rKUzsViUi6xRSju4TvKE1TzIxseHbJIB96eHwbTPLnEBh47CJkyW/OhastzcK5eXe6ga0OIkE8VO
RNvGAUov2t5p3+euGbSjs2RNXDbZbzhyCvecZjbziIadjWYWZcLVeYri4rB2aIGZDN+c8R0r4TyO
rzd0O+VO3Jk39QAOaHfzJsQ7RKuuO+aeufIeN7KpimkDfBWrh/mq397Rw89lri3RBRVJgM4s73Vm
Rl7asnARHuIfkZ8E2VQpMLKGED1JyAqMmK4O6Ja7hq4TBseArjKlUJUB6NdIIrHxQjLjwW6OyVpq
NG0ZjhnwGnUcFKWxRqIk3fGlaXNqFlP+zfSmeC7qMm85Z9HdQFEyRsN9URnUweoK75+WJHveAIYe
DCSXLp7CHY9NmihtmqXKpuKVol1AyXni7YpnVwSe+N30PfQaA6BV7JoLRrRGfQDhBDpJx3gjYvbO
biIWCZQz9JHEmOBIOnpbTTKsz8f1q/13qxUBDKDt0o8QSJYLolh3qDlW/I0HfGuM8wr9ADzklS5Q
GDhlGVRgfiChSvveQfH/mfWB6cW3yAXzSgYmd0DJtEye+4b1O0G3gKvpGmS6Gs5Bwz2U0OVa1V/T
WEBVpINCEQ0PyEbxE9PEBT1uRFGTsARkha/eRPI1Tqv10J3hW7bIKdX0/vHvwowR280ThHn8xR9p
M0JSm4sW14XdmwrOaUnzZfdpUKVvNN9nuB+J79TJHB9uUxS6311kUfG1pB0GlkDwmu8RLXflljAj
sX2Vf/rtesnipbJkhhBlTDXXRyKD7oeQxRhuEN4mVL0yu+1uzo3p2wNpJJFjGWal95mX0Hn0nf3/
HuFNhsEOzsJR7ycuqN8LUcpS9GXPffl3qn4VfRXU+nra6EfGyk5L0YWYC32kydGgOzY5veTNGGDc
0H6d8/BA0OaPJ58P4lZ29Vcnx6nCA0vNoYURERPe0T8jXt3IekTKfowScD/fevcVDHQ1yFNPZ4z3
DD9xHfpGAgTCOFj4mT/a3O0WNZOipRXZFsZ/Rfl9/smIVcOtC8No2tIKavkppCyRvDOvHaqBJDsg
M56v6sGgD/u37Svx1qqPyNWge84G9zyQyYTLC3K4hdLeXH5gI3OXx1IGSXxcGxPGsiJ/z3vOcU/A
hO8Aaapb7z1LuaTDAIx03Vjlk2nrFwnuJg+oFJuyF6eCB+9vhG76q0mHXPlN733OiD6yxzd5vg1p
tgqfXO/mjU1CviJszuSSPjgkS5AmE9acDENGgb4byCpQiVRWg88P8wngthstydO5m63dBxS+jNUL
wgO+U36pT45nopjqfqnQsxbSxRCsOA3fosVZgQhGxQ9Yud714d8tsQO0nCV/zTG61mzyfTvjxS8c
/mHexaJwAngiEcmj6TZVB9XapThw+V84KQzPUMwX5bzXfoEM793GNdkSwHlYhrx/1dR5y8yA+7xW
Uwx5m/SD3eGtO/vw75edOSz/YwovTX4Rg15nXbeaeEkvG/Ub53oqku30jMAWpZIi5tON5iU58ipL
X5E1/S4F1wSLFSh2FJtP8aWu7noW/ODIk0iwSFgI8AOClNYL8JDjigcQ7wJqspoMpJptABMZp2Ms
aerEAOnHsPkrLwXvpZQE/6C6t6KUu+JHLWFKNl+6+ky87MnA5y3dN+spukA3WzNQ6mOT9P7fRxdK
As3oHksuzGxFhHYHmqA61v2RRyj3s086C9qA0nPaGRYbV30odY1qm74Ba58AG9HcLZO9W2c2CgXh
Zv0v+I12khOxm5A4WOFhInV9LmSCbUctLQN9M62EUwY4k3WWVOPjBfQL5dDgTfKf1u2mc4lbNY9q
UQeyfwukIWzmuWp2GSqsxBRicFXAY3FtH3w+74TKNIMgqKrGLtm3+C8zBYIxh1WoisI4qcrWW6KO
TgYmsLaSpHqHTcp14r3ENNZCn/iNMR3bX2+A+Y9lv/WocOb1ghwDukiqKxpneYOmKWyixuP89rtr
tXan9FaIcYGNAAQr6zU0ybMsYK+9HzmTX9WG5l8vUpW1MrtRfU/Od2OuskEbSgQ/32WSvgdO+hiM
1n+l9ceUUpMTSzU0jEZuTATw+VoUUd0RfG2GwHnW5ddUGssqdX0Tr06DHCQwqvYVfjJbV4CQbb73
cpUORoxu4d20GUCfiT3k+mU3Rmc707Aag/kN7VCrNiLNjPufYoqBzQQI3ISCOhTjlju9sndsrDSI
DW1Wlr+WqRqH95zj/xFBxXHTYAm3YUkvj/0nCA3TWSVNLEku40YoLd7xdNZR2g6kZ9yX1gjVAMUl
hozfHK4yOIqPiCAGd/HtCmY2REYL0fV4A1TDZmBf30qDaRZibOLaHeaoUM5uPzGGOUlaGMehuS7K
YyGEW3QX3MAPesJt9FWfYyLl/7xVMbk8cxVFlZPVvJdFD5FVwvIyty9kHr2eJsNT2rf7YNl9URUE
ZTGA3BrS3YswR8wjL69o3QRxAu2j2lo7R0L875ClG30Yo12dIxYyuWxnL6yVKnVF42KFsvaCmWhP
Ck5ptfbAQm/x10ACTCN/3l8vNCcjdi9d1hiCeNmSf+6MDiTbPNOGFVka1N8eDih9P06dRgQNZIQ0
Tyb/oK4yFsgQI2GfLBfqvBENPUcHLkVCUw+1nNz3K0ewjPeKmz+CKh7crddUG+/6d9v2/FsbAPKj
Ymtw/I3W3j4VYdrnh/0LHRlZTe6GnDoKvpUgW2ZHY2nQn9IXyMAb5MRQAvEacmvBAULlalicAUI3
9VcVYZp0mro1jomAPZqJ7eKpUIlzbvY9TZ3uP2rffHc1x0C08fO5lgni1Ea1qpASJwbb49TNceAK
8sdpehwZ72azCg8azdDz/ys1Ug17e3NSsGNFgA/q0Zoz1gOUbQvNcjFb1dIyecL1rmE/fQ/uOXqT
nx4zLA1ciCUNtGmT27BvLIKhm260j2EjSP+bD+09wZHQHgn8OVxBxfiE8YGqmh1XyqE/CalLDeAL
1llwvu64dZb9rFWBSXupu/Cp1cwz6Emio7UFSkNnvB3WkRJFRJvqTNbErJvrpaJZWeV3msfGmcCD
9a1GpYwbE2W6A7wGFJecu4Lt9mgszWlIabn1LUi3Td1FcimyNXWFrp8hq0nrKs+/HdVMkJJizntf
18PtpYX0il6lgLWp8ssiwzMB01jiNLVYqeCnpba1q0Gdr0u2Mcu0tD0YfAZw1GJSCZzdiB2lmbBZ
OYahdBz7aCYzfth7Cn2bl0zZJadB1iOQ6L4vxgv5Ejlpdljv7ghrnIXMTnWmurLLsNyb3sChQcSw
vpu3O1PiHgFfZZ3hbNdJCjnyJi67yUV75s0tF9UDYbr3BtLRiX/v/Agd5MiVFdP582e1QRpIqJtD
tTsQBPKVuZcdhk16OUYct0QWO4p3ak6jA4qsmkfi6jVnxAVqKbLTYowJGZ8aVvq4rcLzLfzAqQZ7
vmkUadDD6OobWVDTDPUPtn8PfLX/1JT++/vYvF9YyuAuYkdCDFETvfPMyDBrl4KCaCmzyWMrWY9L
lg12TNaKcSElBp4r3BiMeIACZ8rgMWXeSzypt8IKid/soLhXUDvQUzQmS1VtYEYP+rkDr7DQQmXI
86pkbbeMZiy5yQrDvw+s2KKCJ7Zq9A2QS6T8wvbNeTpE/YBl6rG5lfEDahZ+hBYceWHMD023cX8k
kr6armQL9mdpUwq2JXkgGBtzBiI4xbcdG4GjXTKyS4v6/z73G2QpVOwA1yejPvxDhAD8CLIMkjsD
ANhgLgHAiKP1FVszaLAbDgS82qvayR5MartMhks9AP/0N2HXYD30wC004cwCWOO/OGCnx87GwWUC
LgeoRdowdma6pPKlxv1GoEZ21ODDwf9x9WHj0xHe01bHbg5E4q/yG4yYraANdHvO0+TMWdpEOkx0
BXM1jSXbiqAoB6MsyZWsWW0iXMOvgOo3ScMo2JF39VLEF1zERjKVZHgz89fwcYu0/1zQHvFY8qTJ
47u6/AMZlhkXq/QN8S1RuY2F1eEai2GH8t912UcIbv9KriB4JUW426ZgrKOGo4Y+VHRijmO2Ry1u
DdXblwFGhHcDpucXCKZ7sPmM5Auoq/o1WyXpf2n9H+E/GQK3VgPPOzBsacb0NGHh4UiM9Qo3XCQ/
xyOoDwRRDCwYOwaa0PoOTyoP1SAQsUXbJGodFDDNhhkAeBGwY05V2e5D4P/3g0hh4I6CDO0E4MAQ
YnDcT+mjb0FKLeSJ5jikuD6EIuKfUq43Xr7IJMLB5F3CQc3KaLFAvmVFNd0VKU3Nann92pZiLsZY
Eqt5BD8x4bu2uuLdyRqSENFGOTmXSQfQObNgnsGW+8xXnDrnqoPN2jjlh/RwmNnRw/1Tmgxoh4wE
eYlvHi+pGjBd5Sjqs7EnnQiohv1ofi9As4mT5XGv5mvn0aNXgmQ0pZagghD8gtnfqzZ7bUDaPWd5
axYc94SyFflwitc4VsGC2/V+1mDe1AiUD+F0AInzVoyFuxfHaRLkqB1WnmRlQSBz3dA5FuJm95RL
QLB9iVN1JKRqMjWBWHv/XDaT77n+PpifESB1qs0Y1+pAJcoGJSN4ybJPyNxlp5AVoWiVJx2IDv41
Md3GG3x6Yu5BbKz/VXmMjFFdlLzI8wIwf34BWPgE5oERmsqRRQyPxYVr9HLrpx9NS8dSrchVofI7
swFo5mW/Q68F+9f/n6KQ/vv+bqvxXmLUj5A+rZONGFxKfIk/isZDufIW6hYs234K0J4ktFWFAV+J
UFZkb//1CKcYrsgpMTog2/Ct1gwrVWsRLYp75n2xrs4IJAOt4PgVva3ohbujNRiiAAS0nnblRDNT
TEbckBpfwY1jq77APMhKZR8gbwbBW6Sh3+WRZ6IprMmmp9oRw1rwBG/EEo5px5ZELF74UPwS3IXC
KsR9V1Re7Z26fO8CiMf9niG/n2lW5POcnJ2qUPQIE6upuWRdDJpArMdky0VcW3Do+wWzVu4e50Rs
gqf1RY0SqhsBSiqyrr0y8vTnwQuwYoYJyurPZKbWSwG5eep5xdEtel9I756CJ581SlU6semz5t6k
O53iQRulJGy4+M4ZTPg7nOcMwz2x3EKZvDVEvtkbe5G4RXPJ1b1C/crkalBJxtUJGbeF/S31e92s
dM+NKTpwn/zGyimvAHPTuAmItJzHSDqdlE2BbgTPydHMwMIYOBmP7iMYzHnoNCYoKF5A8TFeGJ3n
aZRhHiC93AZyEydhIx86Wlesmse4kJDMSQkTt8RbEVp//UmAiR764Ye3CotvgaS279ZhMWVxvO+x
1IWslFrmOhYx8LAKUvI75FwCcJaypVXM3f3WIvPf534DzvntX4mgynLdpYpx44loTFmaNWwOpwvh
qCxOSvbA7GuHnGKkNg/daNSnWZm58X0Eugqk7cj3nXylMWUx8D8bnsI8ovBsgghPnIIT9Vq/f2eN
t86c164MsrSzbBVGWN4Qu/HxAen8cPs6paRAlCqgdDpo1z6zIskgbP03lEgOgXoSjBf2jFxF+JDY
e0mCa489Z3JkPcMNIBFO/21AyWcgcVfqOy7PMWbAH+Ti15msgd9diyQpvYiYyU+GsgaKgGS8KvpM
Q0Uchw2gW3z9Lqq1Cxtjc7gOwd2JBlwZpxQyN/3kTGD3ZoF34Hm7zfOPUor5JTIEP05XSWps/yEa
nIm9WMLnNrS6bVgQBtOYLOIFJUUq5reoZMOoNJyz27ROqajlnAVWStKRiVTCLLNh5coDSYgFBjgh
hSQgmnSIAb07HNxbW9PxhrI2ljPf7wEGuaolUXsr2y9tza2WT0eWwERJsLu9r16Me70ZO88ADGe3
R7Dg+HSmjRyC5AMtmwip28S5LpRmWn5HeWqh2NBwtRnfyIiNmcWigHzt8HUq4lcoP6n5CnX/8o54
4vJFAOzjxs4VUMAKmaZQadcVHm0/BCU6IRz3ZMrC5o0Z5wddP3aZmVMwEslpZv3jr9ca8xYImZh4
xUdZxkBJJ5EoKkezbhxAs2XgELpMO6HqhueS9yJX30zpWdp/s8i2iXZanVE6v1/T0P+7fmywLQpf
fA9QTbbeBz6j52cftpmBbNzT4sy87zTKiuBWF0G/0KnwTbXwxnfMYzmkjD6vuUG4dIyt2f7wAxdM
ijingl10sgq/EPilMTAPB8Py65bPjCTqr9Etsyz6ZmvoRMMi2Pt+XohoX3WxcBEQc0OOtbnUTXgH
PG7EPcjybahs9KdARZgO9bfJcRSi72Qv00Ssyz8TgBLu7cmJzLZ5+PLU7zPHieyNDnAlfbQqo/oP
ELnaZ6QxVM0HlEkMky92EHwDOGgSbNcIlsFags6NfSMiagpxs0mNiI2y/XNpwBEPJ42dWF+LnVBA
P1BG25RqCrVwqH6+eU108aWInOvgeCmXavWmabadxlY4KSQkrrXzFml0PkwFAMwwV+YgjsLHvVZr
hG4uVLg8rVHD5df2QFB6gHVIgWdqmjCTWrd885PKd9pqccPSHTNxdKWdJtJd0rZUU0Et1nzJmlbe
0iP7TUuliVeOxDFGuNqUkdQd6P8DlxukKhYqgtbyCMUfg4YvnY619bq3Aod5PgEcDKyAMRKlNBwp
vSLfF1UbmONGRcUKFuR8lZybmncCtVmGa3gY29sE3TV1HZCCtlvfEJ3o09m32T+WqQGdD4le3VK6
Isl+7yK6a8u65xJ+baNmORqJBiRYR6Wz985ts0iwk4Kr/KWg7+T539qx2tmEiQHgAR5m/a2GoODF
qqDwkC8XCxq+ABbqqZ1Rg7+9IaZj8IEMAXwaMoo+chG5Y2Cj6KlkcL7Dc0nOmGTQhJ5lSgdDUUFt
Nbm885d6jluKqo3Ro7bhITvtgujo9MmvL8ryV6wiDX3RyMCxj9z7fNsPf0CH0uulMLsYLPhWOFH2
gIZLSNEh2doHBESMZg9UO+kiVUnK0mEOT42SgCJ40g4pV1EShjUI8K+MuTQOmJrLf0LvYRIDnm1Z
jKsPr5nzHZkjjeH41KuvTZNmTGqKzHDfGB/Du1rYBh2HDzI5IuCQl0G4C9lwmSCv6dpRWHsGFTgJ
GH15qy45J3LSs3jWa0XhB6N9UEYLMa29TrjGQpPuuAM4Q4koBn7uBNtnnMOym8FObGF3+tZYjliX
lY3bMSQkjonj4EU+iOHWB7IEBsYMIIpkPkNZpGqn2VhcrHIHmBNJ5lMagXSux5ruW/le7Ey8GsU5
jIDABx5Q763ehUgCet8aUJCfZkqFZxT7D1ac5rvwY/hWCaiWVx5Sr59hjpxQTSPSt3NG+gyDhof2
vYndJ0N9wdPIXe+LBClSqs/arEpfEOkdE/jemq9Kl7oRRh0tDmpW2soq0tFT18reHzcU+8YZoBdM
/KSyHoVWOT1wOq1SrKuamwfQs2YW39+GGxcu6BUn4yiEhftIXZRtQlbF0XpeE4Acth0VcyaQxwLr
E4GGwS2RpYwFzafkTOTQRMz0qtn0jo8r2JuYDuu20I0jJKpnDwsQYASd136mQiMXoYqm2qNccChB
baItf6z1ak1aq6IbctWETH1ZPp74hG5+u4BwNTAqQiHe8raE88+qpYt6arIJy85doKRnrkmuS0EQ
cktBrq62iZNh3kWxy1wYMTMchs8Eren1EE73hFzIs7lkwMM2TJHSDVWRdtnwPMaF9Ho5lCRyDUGU
t/sSLMnVoTmrEnxu1FGDWL9WAf0kheK3Xqh4aTVq3cJEHl9ZYlal24CWYD0IPjZ3WImIJ++VADDV
B+cy0egIR8SuCQ2XSz5vcNkBuEEyFIW3fal2NfD9VJIcDq3ZP7monGZG4vf5FlZFiAqY66xYBVrV
g8y4dAoaLYux+MbAOKk6gM8pagFJUOV0w6JQpd1vGHKjVAU3UbL237sVWwTaaRgVO1B6H7eds/zS
o8+5q74Y20YVAuW6wiTxNCli+rRZ1V6uM178AJV0Ueu9BS3glyeyx295tzKt+g4DjKfWCZjaWDdz
PaxAhAjH4HGrUWnbrmeCfND4W4v6nVBSA18aKqC0A3fO1ssCzGFzcIcINGHpXnFqe7X/XP79szx1
CGcMIVtHrg7DHQWr1bo8CQnn6yHndTM/IGPs3kfe//jCaRDuJSJkma4Envkrvhm2HpWeoOkcoHin
8R3PLyrQf3OGdOxYzAHCOMohsYTpjeKCtNh2wy+K6T8N20EmAy1AmGYRkFphoXiKDWWd87fKp8XJ
zxe2ARbFVKtTH8KJ2uvqFGFjKNORmeR5GQmzG5St4ADfEwURo/0uBLNDIg33uALv2LAjGY6AYZhV
5PKkMlm3ZdLY+0Gb50jAUBcOx1AQxTMl2X6gQlVuSjkKTpnmGnsOk+TMwvwKvFvjJgS805syJxsq
V+thnzC90fS5pc+dqtbBDAe+jqD85RfpaJhx5I6L3CgW2EmKPFDu/ePSzj9pG0aieEh1vn/Zlo1n
iYsiPpZXHSAWwOgbDjXMLquVmPBcX1eLuoeoYd/U8eN0hXdgNe3N/qvFClYoFjrI91Vct63sIVgi
ClQpiSz0SxSw/qyuJ6bUa6amG5GoEAwaGBJVDGGedUocwR84RwSiGQVtYB2DJr4zg75fLpXcAhQB
MJ/ZQMvAJKIQ8tMNMgwqaK4/kxJ3Iq1VinF8+G7ZCdxxl5Bq+5ZAvR9cqIzWxRU97Ds77IdouGqd
Y+yue11+EcxouG3PgzVVYWBt1UVcMwKPnoAHAOV2k/MghkQM7386YMAYdbT6jZe10LQ53qr22gOT
RRw3JmBwJvDnjwh4waVfrGz1SxXk3QtVfOpsvMafK0l8HLjamjgEVCvWrTf8uqbfNe6LN9ayxYu1
6kczj4RxRtGtpBL+uPE+SQnuEelh2sFbzMVqB/2iHVfBHEQRT6QQssumcGI5iQMR3TdpUA5Tepc6
h2rrW82pR2gyNKEUwnw5Hgxow3fj84RmdpYVzcVl9SgthiW1dz9tz27CUCCd+rL6YEZNWHiWvjOl
+a6sUebEsWLTAwbPaH+eqc3zTdFwwtwokYyYP8ZYrEedlA/HG8p7sDi9KU5ssQvORLJYSTlX3mTg
bXW90TCtbZ/L5MniFzG/aNtn7K2Aiw6p+qt28QVRbqqJuhfFoDJ94XGLoV24mjkOo/zHhN49X8Js
hCBmA9qaZ+t434tXtNqFSxHw3AKW5bSytju6XZz4TS7/fHuhwcnmdsDIY5/vBayyeqfvVNaj5CSL
mHgFTsB6TMgbBTjTubnfrE+4/r64aueuZSrGAwTRZIFcgKmdl1qjmbruIQnkFDnodKjhIHVo5ZuY
DuwGFq5+DeF790gulQswhsX++2UK6rwp7ahf3qRf6HZFlq1HKbGGIF1eAC8ECAHbmztj333on5+g
qe6UUUs69IdUfhlfGTV26J10zHM5LK66wMa4vvDGyVEbH6VHXSjexits0xQbEJ2edUM0k2e0ea0f
ewc4uhr/Izxm0qimtJCuWMy124D9L8ZKnk9BA9gu15MSlygOmtMxx6wjLc8HZgVNqmhm6RDmKFZa
XDktkfuSWYJzMBEGn4lVxRr52d3zZQBG6tpWryO5uzXRepnpqL+GJFZGeBx2++6tfgSYehG0xHug
OBAIrx4tPvJRBLYd4n78jauP/44us0fW2kS3GOCXtQkGowjLq0AhoQ5QjXT20zt3QpiJTNwW2WDE
3gNAIleoEgO8Dde7xuptSAaAuys8jz1UCdH63t+xc71QkisLBs2OXseZaEXhigisxWjdpIVbpZbZ
0aF8s2X3Y+UaOsFvSrI/CAJxG0hXfpcGeVUv5/mmY9l+75x212VZhNdK/TzH63I46pqmyLeBrsz9
+jdjjHtZ+JJ8uSqFXn92e433o41RosJxb8gULXFkxjAxyyRUeX/dtKcyD9ixFt19KrK4KkhduNnK
MCAv1A6VvbpSFP60sK0OK1ufD7YKdo3LN0zfCcnMyY6j2tSftjPqaGdFOeMIFdqyuNBBiDAtixhb
yGpOf9OitXLbBhboX+McNuZdJgrNsA6PCfXITI+Gx+oK6EuNhJNK4hoU2p1AYERaePR8hU3neGyu
rTQaU7SBmVZVtUr7PejooEGUS6hXuTSdf1dgxc6QN9J6QlgF4klhjSQF4lB1tXYoXsfi5oeOOKWb
bJeKQ8XaPW/hM1D0QzkqNCfmK+q1CXchp1VIeX870VVzsFwxj5yMEh2KfWZqBmYRRejRZALeTeRv
cv0B0XnFM/0NFURFTW478MI8CniWj7ChMXrT23qq0JBl0iiU30z5uMS88PC6XRBGD9JrNeyT1Vzv
uv8z5fcVMcbPCutuq9MuMotlOzQVJbsE2N4pEgPjMHcxwt+O3eChiDDaBRv99RHaGKwCV4+Vy+bd
t0Fcr1Zb2O18eFPBcZ4nmbR1IiHOVHwhJCxV1OS+h0QB+U7uefacXxkqAAW6NjBS1Ek5yTZIdLjZ
Qi1d5w5KNZ5PGLxg5agfHzcM6FZ1BW96dNPdyDG47dtgUFr/S2/kLsXGPWPLviei0lsksKc3qDJi
k0Gn/amIQEK/reZRj0L2X9qdIOt4ezTCMypKls5W5tCVuutFklnqHt3QWxz4OJB9AU5fhnaTrAqa
xVF1pW1l6+392Bha3JyUfY6NOkaTUHbMqoAM9q3uskPrCvDLhROczA3RnkGDNUKft/rAXkRU1JdQ
FQ0P60n6pw+TJE1+nBOpQUUqQAqiAN23jHopfrSdLqlIwLzLP2lbdo/fFj1tfWUu9TbtxKeMLuQC
LsK64g8AqkXza1dfaE+tBhAewyvAkQUnHT0LJPraieDRPCQYG6+kPJ8GUEeGTzFnMrIr3WEI32WS
7eh/BKW1QluedGsykW0WVSz+WZ4dQEwVghz0H8B50v9b51SK0MywlXmI9kVUIZHPdV7rIJpFkya5
3GqELaQaB0dzrNRTUzcgmHCBTMUSUpyRiXaZ4IZtREMr2K2AztgLLLtO2HRYyC1+cr337nxoiwAI
IrzKl0I+1LKA2rM0XGw9EbqzSxIP5xOXkkcJ4GaDfTcFunWVH+3R0lAKvPlgx0w0z5Yi6V1G23D8
TOwGbRnVu2QTFLgc7SHvSFeVOR8cnoVLDl9tfO9kmdmv4dQcvaEOjwIERcH4dnfr7qYoDBjMIQNw
5RVd8pdzBTmySKt1kmrRQoWb6N0cwVW37PdRUtGDdaCrGm+QFQf9yGJxxoIvzniJ6ER3wLDyhnxM
ttyC/SEOEagqXriuJG1THcuGYM5njAo+Fso3MPl6GroCylXpv4zWlMYRzsFNOb+tT2orNOzAitPh
loDP+0wbmS1BhAOJ/+iR1FaT71OI1K2EERXFnZY/59yYzgN06DJ0FIwf4xU+DwcDsVDAZDBs6ze8
o+tmXwhahpmdTmNLP8oFnOi80FeOOR/jPqBDcm/0HGBNAMGwenW99WfdQqC4V1o6MAE1pOAHb3Dw
f2YL4dZoLmiTPA52/DZ1WH0j220p2kvziaf+Cv5i5LtEXn3vRr+B51VS9pg7+zXYEWAOdCLkqPA+
e4GP77Jtk5mJVmNW90erjMZmmPkRw+PrlQcO9jFQw7wmI7B3QKJcQy0zhBcc6c1LKyDgrolWr8zJ
HsVTr6WrOnaDMQjJPbfdz9Kbhq9kI+j8tQ6/2ng/OChm0NnfKKFhkb7zcY84RtaCCUsUrY//vq0L
G8MSUzi3oNFpU5Ma11Dncbseh6KA+cQQfeO87e0yA0smByOYfzpYwPKJesEzmcfgDavInOeQml/j
Ty3uWeYOMaqvDkPxOsFYIgenaxyd3Kv1iqTYftcOSMFFI+T8PkMW8ofcccofwmv99xt3DLW8VAK7
d59g7mq6pCT63EmhiTKuQBFcq/bGY+ABcE0a45MNVAODMSqQ+BjAh/Akye39Sma7oAGeQ6t1Qa3H
DvRV8dCdoua+fnOCaScV/pfbd8iEflUi1pVuyVfpdJrd9Q1NJoA22dFIx5NVcM2w2LEaiTQ/dtHt
qanFPDJnPi657JQmI8ylVUI6IlekPClZmXQXcYye4GGSMbuy/29JHKfYFIzNCHi3nC8yK72YhU0f
W5J/ThkYENJ9cECNTVHx0o6X1a+vVECz/bLbFhtnXPIJ53RVqvr4jFXlKbNZEubRlpI26+QvGIXa
Hu18Ykq1L6WPDQ8koEk2sYgR9NRqQDuxVlVYX41MxEx68sQebK5pA0Avbn7UsREVYrtaWwvxmgEp
QATVfv+xssAZBONI1uaZ2tiOlmvyDXyOo9YHYNWM1AJmhGsWoQJwnjurZSTBqfMO2wXiUIXelVPr
4GLNlBssM5D8CCT5ciH+nSOoR8seICE/Gzeu35TinANIUPhVQU1tpEziugHE2Ov7/PsulychCKqy
o+oyRTRK1p9lPKLc1uf4oksQPzqsE5yKRBTbbwkVG+M7BD5NjQu1OK6KqbZjeDR7I+aFtuw6ZFXP
0d31N7SlH82hRS2xrKTsz1rkbK++f7HtmxECUcwcrkmiX2PPp+4bwPNLCn2IQQzoFM4a8UIZKIb4
4wHZ/WNeqdJNAAi/a7LzMt/0rlWx9elg9Y7EeBtcRfayRYnMS3phtv5UvGdeBC5qO7JRBxv+d3Lm
mwvJXQo7SgRYGVv3gm7csvAmiUtOLNQ86tkA2WN019MT00BRrUp4qvUMKQ/C8Gw3WlPYiIpT3tnc
wI22LSmRMlqjxNU6q5iS2lL6Z3+YFSP8nKZgBNsXmcrnRL2VZ3lrlunxCQ+gGH2Rw3BnlExatIOv
SFnd2YqecQcJxfwLddYBbeQwy9t3k+cIqOa/H/9iwiBTjKsY1GX8q0Ad7fcBKpLoKDYZRQzDVByE
GzbqAOJWCKiA5zGCwhN/rGSmeiKx7Shpbt/Z005NOaHO50wiX16gjGVbmzoCRQ3wCYrC54kGeoPn
8uB7o7GOqVppyikUgwyO/EQ9i1D9ZcW6XNZgZFj0dntwMu4ARTjuvA8VgQcTl71BlcP3sxPEUuQ4
qS/YzJEGeYdeKWNheP/l84NAj0PCbJBx+IyJi3Zwe7k8f2VzNCm2SKDdbGEOPRmUgAJWW3E2sCPx
JUJIj6i5BUwmjt4wVcLDO0KyPXzigLr+FI+3GEAeBILCdYYhDCcPsdVg+YKT0dR+iAr36ALETKt0
AqLEiZbJNIQnyEhy6cChhYzyXHAXZXza+pJf+a+dnJ+MinbQLh1N7dwYorLCIN7VA7xT4vQxtDid
W9vuQyFKn3zJagc75wy8uB3L7YisNDbClTzgISqpn2x6nWTAcEzPKP8pHrSF42Ba51A78hAiL97X
FaJ/jX9JhmRvV6kI23v7iN4uHgZANWd1RO9x/ZQ++yChr8GeEdrdzo5JJPD2f3tCcun+F0ZzF5qN
vvgCCOGLc1oHS2dB1TmnnBq6z0Z5WhPc/M/OPJ41QvcjbzKhqzw05IOtV7ogExEnqY89uk6+023C
slNko79MRKsCwmqK47TKtoz4HjakCV/qgeP8bWodAwLiL+NHNKUCMyO3titNEhEeJLIpQDeFsY8V
hbKhJ2NWDgSBvz5IC/svaWsBqXFBDcarLOfUOaDOajNjLjCEKQU3bvva4xN6NkZTL1/bvM3kc9m1
NAnPmGjl4QsCLY1bn444eqsSjTwzDex/bU92zX+/lbpVxxgJTfnigSTx2nbPAuRxxmiK+UYpjpp8
Kz2GUKvbnaSmslpuxhG/Rekp10I61aoIhXwv/dgBdZwayWlqu1rcEukO4hYynSGxwDPyMiYAJXSl
FqsyBI5W/atSKpl2rVu+7O8JAZhaYtj+iBs0BbLupsfm8jMVfsOzYbhgrpGQDfRBcOSsHVGQ7z7x
raLngRTzDwIASZQKPlzsYdNUxGqgQkJKO25cNhASsnM3YB6Lro2Ren+KsGiQyBIbx3AcxDnnLU3b
vEj5n7OumQyot77iwPAhBsUzUiOjfHxN6u7FGpwy4/r7yA7YfDSHeZQLK9qcGJY+HssQBpt9o1jK
SkV+DjeCqMbtf+wCc8m2WsWlwM05Vxkk/UBzY8BhMbt+OjDO5KaeNugFdDARby/EKSeis9e6xLHZ
KQsNXuw/ytu0916SPfx5q8wJaalgYw6shSPHAehhgauI+aDifldXHUi9gDP05zak6Ncfi8PYxqDX
rU+sTVqezY3k0tghZzkrSNRA8F32YBrJ2bAdIBwsDGDspfeohKmpx8PAe3JP+SkiVGBJnIddmKPT
zRpK/HCvVJ6F5njHJtt0hfcAX8SC2NVE2XXXkyZcn39NA9IorxCreXl0gztmMwEoRZbcvWZU5/iP
wD53Q67902XWSiQwv5LVBxaLdj9wq3UMqPbUKz+GkS15DnaiCQ6mC6yVgn2kIvKNHvo4DG7wrxsA
jLYcOtpe+rqCLbfTuQXpReREoqrEVNQIoyzL8KuAjePtWRmiOBQxG2aXl13sCHkzlcJm8ysCsBto
5fqORSQDtymYY52d2V6Fq67q6oGxI4+r1CAgAg/1nPBulUgLhS16fL3A0lvNhqHlGbUCON6J8rUE
HqjS+fJq29x3AwrgY8Z/iJA3ugIUZ61yoSweNZ8u43RmS8ZWFtrDgffsV/35BS0iGaQi0HVJKsr7
dZPNuATGd2BbX3K2gF4JZ3mZ1xiUyGh8Ejv6/xNYLK8RXNozo+ZBe7XwyKdNlTCZSO5uGtT1RDI5
PZb5Z2gJGV5hRkvo8p9naxK1DbyIN0tmAgdeNBnz1KYUXfGYQlOcyq2xjZvBaYc6j5rQ8bWRG1/m
ildVElTOWPviH4LMkpJordIGL8OD07O14xBSwvsdLFB1k0biqFBmqRQnIExuKjyKmxC9Hremh0kF
o3ttxaeKHD2fiFWEuRAPCSFeL6nQha9SAE3IHcWJMB11ovrJKkI9qM3gq26zpV7pxYhvPbTxACuW
ezy1yK7Ice7OAcao33Vc9DF01sTERKDTwbK+5lNeMgx6Cs3vKK7aB9wS1os1IMgO8Fz2ILPOMlbt
lITB1T79v9V35VsTOfWYGkBEhAEU6x2dxlxx5hMNNdpHD8eSIahkLBjxCoDF2sfjTECYLA0zrzW5
HzlFc9w/p3ksN/yDZQI+YsMGwfDR9RROpwpd+6ZSzHN8oLQFF/vnOD5ZOWCXQ+sDuxGr1iAoI0cN
72/gu4GcakVXqTsjgkmvq2hCpTEiVuWJA2ctLCZ5n3yrQ6noz0OlCgauYZbItlvF7i6zpNbhJrNG
tSK3vR8ND+22YsK7i73VBaQHly7wResc3C4XXzgtLuF31xzg//fmaiL35/aO5hbTZDYKj2g7efoG
iMnUtvmM5MMDBLkcK5mXPylHvfyS1rvT5FPixrDClRtSZcg1H5W1lsZFAaSkNbnPUd5lHwgyLbKQ
G2r78KW8Z2z9GBhaHWryn9I7pvqvZYHFl1ss8QH8noZZzN1Mi7i7PwxgPBalteZnz2XdPOAPfxxr
cWt0jjpfEkEewy76bf2Vq6n9xUcfy0gvft2vqtBugjaWBNW/UYTCBo4nj2/EWqcIcsgasuGZ+h4M
dCIB7qk+49FrhOVQqKw6stfyGo7LAI1Dc/LX0ljUcC44r74a79AKiuE0iB71+H4tVTg2oLagAGnv
6Cmpj3vmrye2qvSa0X91yIYNBuG7l4PynE85LC5oy24DSMJliXCNVtTy9WWnw5jwxd274U0Z0KLI
ryR4v3K0pFd9KfdnRoUejd6zStoBY9x/pBmG4xiSYMnj8HsjUFVAHnuW+KkIIWMUWNPvNzRl+Trg
bQvkM74SJDViL9TDWzWKGpguQj8mMNQ5B69gNhUWd+0/7cxSGzvO4uy/igAZT2SCzY4MGI/w6d1J
iSskTc7jH9dX8GwPw4V5t82yd6wr5u+3axutLIg0ue8BKlgSbEYcOY5W9/O38PukPRuqbLbAKQrs
zfYrHHCMCdBJ697AEFShCSPpy3Za0qXCYWC6PyoImWpvmrll7JbTURJRbTFZaxwN/8AZMuMJ6pGN
N0+ZSct1fcLyxBGhmR243D3/fp7fa9O6dV991iVuJEIR06X38VBqMgVNIFy3Nvlu5dsm90URHNOD
d+2qmNvb8F1lDyDjaVwqyMn1XI5z/CSkvglI1PPeleAFFTjtxXs1W3wKzk415y+H9D3T41xqoisB
IhNgvxkcBukvqcCfygDolRUzK0ZUZLIPgMRi6/yvaNpY7Tca3ycImdGc+odA925B1ZzVPCgBIlx1
C1l5y8HQwTGfVne8KqWQ+wvg17RUv9SmWmfm06GywYH/9taNsk1PAcZDPYTnP+ooVIZojVwT3c7K
H4Z4fJX+MvlJ31Wioro/PBgOU6kETLxKTNkwealUDT/wV+zHD84xELGWEeZGgq835y2JVTGJWuE+
9f9ZugefrIwGhNrhkEBy5jfVOKf7r63dmq2lFGdBb0w+6ghLq1b1so0DSXQPE1Xj6wlZFo6NWPg9
dP8rHWz39YonG+dBRSnggB3/gfCG6KMR5Tr2X49YgJ8B6/eHpx73TsMG+wX5ID1QalLqlVItxZgL
2VvAp7yX8V/ZVFFVC2le98csRvhyeyfTFnwLn6igl7+1uV8M0Fiw0Di0lOcZFsxS/9dpH2vvZ2wb
tA5RLrh+uBfxdcpUf4qIirAxunVa3iZY3M+IpzSfccePu2AljkZnjbqCPJmC+fUZxmhYgQtO7lNG
djEZh5y01ExMmRSTt8HF548LbOaLQpNUK5imj8hX5v6oPUjdH0BjBlJdQ3BbdY7GBaBJMhw2BmCe
EqXrwwyI8+DGH17RaHGUVIpL8V4mWM558Xs9Ku3g/2DYqXmcM+jeYfhyuyqlEqyCMHsWqCP6RDZq
ZTYCAroqwK4oOwbnd69cTQUotoZ15mlRppTDPT9WMNvIXQimNiq6nABMnA4s9QV/lFseGHyDWuQE
VXPdicYiQ+MGBeqnT4B/SkGMGd/nm+GryB9vtXGFOYT4rcoz8omh3WLWCkLXei0PtgS9P0Nw347A
LUvNZlBpKu7boBYfTQro+S/76tJfbyiQvvX2ueu8P8Squ+fJVycHE55wKT5ebzk9WvkPQYPB/ts3
SzWtDWRUyEU+lBOR1/WA8FeMtV7oPQSbE0EIiX6vNDm6o16u3DCX+zwVXyNLrGPEecZTqKVJ8vmr
kJYWh2v3ruIwFY0K1qmtiNCl2taRQdolrljvx+0bHJ1U6QL28JYpibJMCD3SikQUj+CgivCevAgM
MfVUdu6peUyljQCrQV+OM+t3CctiQ5OdPBh4XOadTGDCA3+dFkei1NzCV+cVfPIBxK3S0P9L/7o8
AOYoPXhsWug1REA4TMCu/KkWl0hI1UPwFLXhN1O4x06wd8QB84G6H1njhbzFSoOguHZrKJSx/dsS
MV4XyxCEZlMn5wpbkQxv2ndxHQhOQiZwEk2kq47OiiP1U8DJxI7SKQA0lOly1uDWuxqNcf3RANO8
cbip/xT4DLJhuTN7Qgazh2PCd0uawjATNpSy/h4EVtegdt89bgNd5uKRqgeJhfhEil+RE7GuxIlp
P8f/KNBSrfe0uJavzKfZQGtSD/cnSIvEvalnD7iM3FgaXzCFULfns2QaMGYDqdYfhvVQ6NyNrvaz
vj9EqsriBiMxVZoZbwNkS9XSSp+kRck6q9RK3lCiSVlbgWp8mb4JLNrbLH/wlfPNSMzBPf/J7ddo
HJN91awKPFcLAiE0poskW8bjRDIUP68B7ZtwUSzmUWP+XrcOCf+HNTzlw7x37L5GCGy3vpYVI5Hj
s7nN51RUINOFIktSWKWSjSqkB0wNcLkxE2foo0PcR+RPalGv4heqOnNaybiH4fKiQ0py/ASdX72Q
9VJy330zJVljDmafv4dST83si6TGu+sV+cnNADMBt8AhG24dA7HcvGhX95Q+LWqfWCwQcVwz1sDe
pAj9MkhwOAuPIUX0OsA3Fzq+gC181jz7f2miu7DnGqKCE6/PN43PoFBxuoXOnlDFqc4ijcIzaIO8
53hKY9lVOWnzUWFSz+td6phdvgEgApMNN2guzI2nzON4GDuYk5Opv1ing+EVDBEj1jKqOTnqkyDy
Olqj+aW15SL/B9NXR29EFwxhgkMqUlfSPUTNcIOKlc2JAHRyB4+8lXHfnVhJWQQccQXmbsvBWpee
iGbguDqmGJQberA2bFj2GTn+1ds0jNQ4LkxY7mVfc3/T/meHh+t++p7fq9HE9U4lz17BFZLGpsmE
Wb3bv6wZsQADxpHZrQv/atTt7X7d4LUrGDNgyod6BPQu7QiZTi2O0fWT06GrPmFXhO8lnZT/w3af
ZuRdyWTYxEauEHlKcfpkM2MhIMhWkCBMiU9rWQT8qkaOO8FgEvcLIucP2AmOtC/sD265uRf/YzSb
hHRcVCzDbugjNToo4RC8E/MDcfoQcPg8C294olmODRBnCla09Aw3hQc3wYpHeA5975oggIilpVzU
wbNoxOFaz1oNyey8UuMGvcgCGedi25AqaJGr/Y6klQDi7515a+/dE4Owpf/zWYI7YMDFHGlgHNsq
BC/RqcObv7pQHXoWWLSzH0SiSUkC5412nGsBV/4W4BKVe4Mp9m1KOmNjo2H/tKiaxlVG0BiR2X9x
KKr/WVCSJLO+4wd5s190YLVIwy7sEEs/7Wvp6yPnWqm79556aVSAVEEAt5EmKlrEiSDBck9yWPge
21fCigj4jI6vjM+EiEJBEZAUiHbnvwqwnaK0aw9IxS9gbH5hde/RylIMQh/ReZ1YLzPafMMuHZSo
+kFE0VsCj+Vu2LuqlPrgG6SikWv0HMPITQ8cfsfOqflCdEAiedmLb7oP0hy/T8L6NL3XQKF4hsOU
9/a/XANGCP3SPLbDl3Vnlk7dhmOjTKDsbrXssImUtzyJQsuN/JNJCfWN49AZ0ww3+9Sn6+/BYj/T
ZfIvzfsfgfXmmzuT6vJ8TNw4K02U3JSmJVxwUmfpBygHEYCThLdDJwpsAdGfO2bqpJFKj2C/YQjW
HRP4o8UHkFLtndcIQrz7oZfR1AqAGUJiKCj6lkLzO72S5xpNaJhDRD3QLFHFw2QvjGGoQSDRZpvI
+60/OsrBAOAig3XLwHPgAlwZdWtowpz0SNOT9ZRxJaLM2Sy5f0D9dfEHRu5rVM1NIUM2/LpoqhHt
IVtAVkuWb1Yx5F7DtypQMLmI48qqW0CSmtTJB8lbJdmYOSExQOjZRRVZVR5+6aefT1CX6IB0n4yn
FBVFCf4Rts2QlrFwP9pDJpBb6H0A2QvyXWQGZMvdkaAdMI2/1o/q6hMXwWAsAlYep1zXEKOn+yeV
AKrEW0htIJMvCcw1bM6TqDGB0T3P9ttKL5879ANVcDh5MKU0Yb1Afth90valnGswhosHmIItsL/O
1aBj/e/erKWq7MJ/DTw8V/CC+Moa23oIsZmAHw39vRwMJoslmW/xRT4ofNtfkZ4q2VOCALjXzPWh
Ct7ir37ZLDuiG9/1oAgq7ZyCJ0Yb8jg9m/XA6QnFZSz8oppMN5b/cv2ujyB7F9m6EJXIByh3xc3q
VqxgPOeR9R0gXF4ahVX/sMw5nGDIoqE6UBXhUOKuJmzR8Nm7HfVyEwM1bhme/D8dEurHEPiZtN++
t3je+fOVaLgoXVzaHxQeW8zrYl7CO7MCrcdRwnQZQsDHWt7fMnHTKXs4H07x5TjhkEXVt5RPtSyn
8kyQoKBHBWKjHKFW7RxNNz3a2WiPy/lIHgSaqa0zbrDTyK1ci6Gc4gNwNw9dVsJhN8J61Zug2um5
BEEjE8d7+ptj6t/qLvvXUQyfGerfntaSEoePTBfU9DEHIZKo/PAFk4AsFcDvEPO8nqWK/GtDlL0h
5R256lVx6riQ1+b7mjP9tA61P+LN5IRvjso5+/2aTK8SARN9Es0qcQh0f0E22JHstXEzewBD+wGE
Q0qNTI2ZccjkrHB3KJwgODZ79gtqOwNUeEzmTw9kPdkbXwhbJQy7F6gefgmtrgcAiAtJc7gf4EBM
2D8mGNL4MGrlPSQSN88BhQ6wYK2Dk4euSOkbqGlk9zHShAIJfOPSjyCDh6wlERaEHSwsg7mMcdXt
cl89EA3xMEoZYjHQNg0h6HyLBCOiz231Zb+47Y9cbaYzocqCFRhXmsWMcITH251sQaychzHZ+avC
OC1vQPjxoS4CD0SjQKh7QK/vVXBb5Bg/rlnGLEwM5qdOqNgM+YRoQXUk6fgQInDV180CPRcI0ojc
g+jnEm4xQRToQtyArMA93/0lGcOZfw/TorrEHr7p8oQoyO0csM8hEOH4kUE/9K4W8doH7ZyhlW0n
KIxXa+s8yTuSv7rd7nEELGFLm80lAp0u1FnPeYDTht4nRvXNfvnXtThf0BSvBphL0KA97pEDetJQ
imbhEdDXFDIxuCj6+w5zjZt1iXd6B8deOZD1XQMc3GYq/qYANdKmHHYt6FZ1Y+a4I3uAjWy4vYw4
g0XAFRSas8oSXL6boFI7bZp1bbH6UtCjWsuivE0gHGMRy6zi/xz4gXUlK6lpfl+eqgRIhEnW4eLW
oTLPbuSiE2UmmMrtnbNejqFNXTlHMkEtEzyrhH1KnFFzAW189crvl7XmXhSegbV9h05WeZID5pqi
kwafFBEs1+xkSExl7cXVydPUvr6W0TyzwSzjY0cee8aRzDsB6kOMtrAequ6OfWpNn0JYDaL9X0iC
8HpEsXWbaI6LyvyaUU9l8mhDHukk9seBB2l5Bu8dOOOLidpB4yV1DIbl9JgbdKrQOW9A4oegoH52
pWL6zkhhzBfJJkV8HI0JVfRUy8Qe6c1xxzoI3gHlY1f+4LrgruVE/pTFYNS8zozFo0S0nMm164Ug
cdZumJVFXpGE9v0utQ1hSvXf5yU41FlOq/L4myS1nbU2cHu8+jn23jfiMOePb2iejoAT1gVDUfNb
J6EvDt4CxQlTq0HqdffZPQITdCz8o+oAhD32evxBlzZHCHuKvDwTOHEoWiqfeHAXQUSDAdx8y3FC
AVk1NHN+01rlfra1aED3CRpjWjnPn6ktOuSCmhdHOeFBUfs6K43aBcliB+nHV8sjNYypLY+cdN6q
egb4jhkfWtEPIPfv6mQXfb4UG0eamyIww6im5ARXleQS4ZDXjK5bIiKZ8v6RcSO8XGm4iYKKOmbG
pwcji5wXKYObhLpe3XDSqCqUZ5HwMOP+d/L0AFA8d19/KrKR6dv9OzXNddv4CPxQY9lQscjJZXwc
KNANifEz3fv0b8PkIanpPTWI8emEJbjCAFnju3tM/FkUZtxPGaj9AjFujSZvhA6b9+VXb4iANtWz
2nnAhxyKNQa0MwzWxY/ovFGar62e1VjP8ehOEgO4AIFEfDVkog4zxu+WzKvt6DhjK9Fp+QQy80TN
54eGFPbTzSx9QKgJwuugopqxQGOV3iRA+ZUHlcFNt9A39MXg1ej5RaK+7p9zvhz1tqvwB5wU29+b
BPIiLw/aa8vspYfTVNHfPByFoAwpVsdG8pJG0eTYe7Co8rVT8Ix7CGbJUnXiViPxzy6OPNU6dN+k
Wu1np7fUoJPFOMZv7zcTndYtUz2PzfhGM4Oon//Cq8JUaBdsvabYqt2QxVVJ3lhJNUQ4agbIHsgY
vRiYGrdi4UIr4DkPdEpVzxpzkMhOfHjrUqK7i120jKcMF9FZaq31Zocx94I2zWOitbD67uLCPowB
ojKZDYraL/pq+1qDz5rQlQhJxDMI0VL5wk8cT6OB6XPOIuxmp2iWJyx/+mNxADKxAi7hVV1WyIWF
L60C0OW0Gfqf2sp55DHZygN0fr6mm+HVZ2xFn5AZVuhSGhO7v2jaqyMByT0h873hsEikytpwIpIQ
iAUcF1ur4fUbfR6KK3b3RFEz8+rzWv8t1V3QBLMOvBQDfJRuBuMphgxnVSOClYbGU9sSsVFKDmmC
Ivx0etJdOmCjqAyy/oqmpMN0Ue6LbYQPJ84Rn+MgMRYo0c8cNveobtgiqxjRRnJaHnZwVqk0G0LP
AOTUhq2JTVd9XAYv3qj1jLe3AVHGknPRN12B7g5Fzed9m3/XzLimOPUg5InfBIj2G3Kq1UXarXz0
THcErzIl8aDq9z1THB3ffWjw0FCTBySl9PeMxpPMXsHkW2QK3723DeeinRrXsUeJNMrs4FyYHkxM
/jxyYPNVijrfQ2n7xG5DNRcB00saPUSi5UC2J7TZozosx4kVJnlChFzwY65jTZUAmeDgfLGbt/0u
llcEOPY3Nwz3PlKG0UfEB88ErlEPRePUQAZ85m0Y5hSnWRxgeKv3dir0cPARFQFfXTNh/m7i0WVf
JNTV1ZckMVHs4+LCA0v7KlllTD/tB2TBV3VRXAa1EhaRj7lx/zcVxLxzcPziKLtpdrg99uKJA4wi
ye5NaE2tFQ6FSDYskOTDPKW26/4mEfAgdnX5OhtKNHvluYV0uvPDxmHmssA2RITq2gpXF1ECuLzN
WfYxWXjfmD6/1mtkkMAQDjYK7HCVyxthKGcx1VGVk6sQBSD5GCPJWQhRhMuPjtCW874iKpAUJamO
1ZjpL5FxavL+uRv3hNeiKc7J/4RUyAxF7/8qUjB30EShwnwxniz8EykkPwd2o6NUxSSucc5qv9tN
8w0+DREgxkV+RgW47y4Z11VAVDFzwo6el5sAHuV2s7ofqRoHlFWnXn1yrv80mlU/bFS7NUyZ7X6c
jZauH1PIbfhbQjmR4TNHuxS2pOpfb5Nbaq7n2e3oIXYaxb7RD9obyS06jY5ydOnzHVh7tLKkQj1y
Ay4TvzRZAXTn2hQkzTdAPTDUaLRAlLd0DKdateGEBPufbhZMbKBUK+doltiy357I+yf239tUH789
IWjPToor7RbFiCwUAOW2RD47NfalgIW+YmfOOaDyzdL57W6DqhO3lciEM0AAsxTOgeCHysloRs4Z
Rq2a8xGeEMpt74JpzhQMmqu/hwDOWDgDJAv9uKwKUvBfje1CBekhm66WX7Iie2mUM3OLVIohnQZt
4c5A2LYmMCjRRFq7VMl2kfe5C79CtXkU3RbV6vFdXMEwK0x9baIAKMswdKQnNL725FUBjMwI+iAA
0HfRgNcp7UlfiB3+ed5mCpqwTD+Cs/GCz7NfOg1TPxM05v9BYESrZ2UFiuesnwUMM4xZd6wnNI6x
Ptky1azz3AkBkd6oVNuERM6GEhEFPz0ml/IpKT8Fo1/CfDfJai0wPoYYidhHsT3K9r7z3xyOlSX1
0oIhJ2Yj9Z6FwW3llSlFZXVivXlPmTJk7ihG50vm/ON0LVp6UvDINeD92/0N6VKEuRLaouV4wjvE
PFdZQmDhFie8/Apmq2qQXfW8ERDUMR1WbkDRHQDVChX20BitzfDSaaD20pjY9c6CxQpv4pHziWb4
fP1EYhpABVtUKQl/mwKGifIwUDawqKcfXqxSP5KkM9Sf6iC6kc4SgHzHwv33+km0rmwNP3pyJCRy
o/B2GkirIe+L/sQk0EW+ymhReaBgJHBT7LmFZ1n369Ja53rwhfhd2q/YZiA5mTYw35By1ZsaCMPp
RFskwSUPyEgKDR5Lz3V8lyrgJL59ljGQIUY5+GChV245now0ykP2tvAUA4OWJYowKQHmO30PlQTh
WY+2pNVhWUT9pFeZj6Be4W8YU8W0fHZzK3MNTbD4G1oUCZU/Mc8zntLAqvnbBPrtkHnYttidbELN
WsAqL7lRPw1neo3DBVq7r42Zf/5pzcBGAZs4q3B3zN2KtACg4LPcDp0U2SEQahYm74nDyKkIrged
oZUZw1Y4+kfrDHiY4N1P+XHNw+za29b9/ISPxJIVLuNcM3KqBiSPqT4zlIixpBnraS1HA2li7BBC
FWBCEXGbavVnWRyQ5zQOPJfj/xWn4ADar2xE/Qyo2GhfLQ1XL44R41/L6lQ1SS8wNqbIigDBdraC
zzarz+QspQStYmPsB5CW22ohmu5T1uts52ZPdyA5jqXAud4tkFYmcgoTG82aA9v6RPiZRatX4YMu
HIgT6JeZHIxB9y0JVF1+kxxse4xKjB8woaVC6W1KR+W8OGv/QoUlxl9DozD9psZtlUAjsQ5oKxr3
dKOLy2ZrtVI2sgF8yPal4dy0g2VrfGXWBm09a5FhkAgDouuaDCyCpk1tgIBvrptDp2eF4zju/Mk/
2a29IZcVwx9A3sFjnkjzXk1CcVGc0AfrANCNHCvCjQGK7Woch0mRrxJyRTXFqObzwzF/f/sCTcsM
5i6UDQg0i6eXCSg9GBOUPXC0OVeFGe0IG+SEjPphYMl854z2G6lj4DV4n4mgjLDVK4Y4m0eZn5Xj
zFppzhwUGKEBkdUXKpeE7k3voZpLgO99f/ou3W1DIw8gjS/7iUepI/rpYl0/oLiOM4OAtxUPr4ro
YRkJmcR4hvyDVD4an2ziUSdF0Bi9INlKS7N/J0Kt8l9r6X9ruJL8zzkEFxqG/tIV7rpxhtcJ1Pd7
RO3d2AYP2PA6bLaxu9SCm+s7ywok2KRv1Fbe3/V5L3pM4Zy1xugk9llJy8wj+dVGoIUqdm/wVA3g
bxp7Q1zo+WKSueGisdlgfmULccX//FjSrOpbyws9OJdbCvT3egIQaueERproI7/+C6oI/Vj81Qt0
JzJTh2fZjvnNO7UQIPZ2smj5R1hHV9HgdZxYTwXUSB8Q2hmyg0aDRLxIQGhFPaplabm1gFCillqF
2Cx6iMZaKWo2qnUXy+SBOuooXfRaOetataYwm2CrnrfLUyRMgOhOQG9AlGIpv3tLu1dfBRhBwpc3
g5w+fZzpyHtKpqqk3z1e4l6Ilh/ZcLlGmMy6pUoMHQzM6SIqzUMxIC++qBy7Ni+DVHMeY1LmLHwx
WNdN0cWvaV+T3LLPCj+cD9F58uqxelhke+WRrumFk1mDxldp7UBcAvRF9lCRqFNdfHbUm6MYSRkl
ZpIpqtjJa8GBIDW3IUS0eOcDWjxLZE+vIFHbuJyV9sWbMIA8YXI3f94aQ5B5D3x3/BIOZOvkSPqj
+rGnGkgALkbCstELT+SfSnF6PBycRe09MFMfgW9PKXpwFx6vIt1KYaEqGttPt7ZOSoqUMkdPUqol
UPnLX7SbETx3Z7sLQqAJRBq+JApCcoKGlQEAOEzDOPKn04K7iTgSf+jsIZQOSRdQHz1ZUkND6dnA
wwAwMq1tdwPg0578WxUll9cei12TmPtEeFaRq0t/mqvXxyg2oJZQ7nMZc56HindTnw+ql+mu5BDT
MR3txnOQHYuCIB6UDKNaxD6jL8Zt6AXkbsfYIc0IKr8TPs0M5p4tZq+rSnwkU3u1bJXt7A2gnDv5
Kxd+jwLXAGIXm+OIr3RBSpeL3A4/TcLpPJndX4LymMphsiOafbB7leuqUZmuZMEJaZ/TYe2YMjZd
cenokTIAnMIMpwWtEt/ymDikaDFCa00lnN5KV4jtB/e/P1N2AXQYqNzdBoqJzuNNMdulxDHgAFPt
uaR6+Pfq/no501gwVQ6bAEIFHFFzBjKmZ31GofWtSdBN50NZMWjGlV4kEtFHEca9QBZ4WciPoG+8
sdRJt7djCuNG+DdrRe4Sh3lN7kr2L3uFp/3cQ1zNuon0c8fQuFiJXsPHKo6slOqUogiC7RKmnlOI
zVUXqh2p7sOFIQmVR+Iatal4xQJIcyreW5cl0Wf+WH9SMo18bCkJo3RDfg+9iIu0z4cvYblAsDfF
aKMUOHJeY5Ig4Xh/Hv1Gae1yWraJ4rYxxs+NlmyzpmP0LOCkOcDGuRjQQolERYXhEFnCaCEWsau2
pJx11jb84PozUQ1zpKFkCy6NW8hDobF8t90/3FFH1fQZibaA6Di2yJkxtzJC4Ek6HYRnnFtPm247
vNiOp2z85VgEnUdwID3VK8opv1NGGBHp0X4NwBEtJob+eC7f1kZJh4XmJTUpgaCPNcUPYbnOdOXq
9OqJv3I7SGCMGAkVh1kHYKgjzchXH5x08lv4QX5mYwbMvDjTYUy0cUKuHfGxs9m2h1RccEP//pEf
CtdvNDYVY1XRo+4w/AnLXmqHjaeBqH4BTBnh+zmSXH03o6oLuOdPzN80iGCL3DlGXXGk8c0t9q21
1yh4GWcJcKTxhShkySPDsLIKDiKRgWMbJx1p50v9hVx/3lu6UsiTdLo9vroVv/ivGPOHT2PX9oH3
V/Bqtr4oLrL9FK3jxGhqcaRC21jK+y/dm2WeQFKyS4Y7pgwaOgNJl3u/7s6ODHMJqzyFGPQ4zPHc
dRCKt4pyYwPEXSILDEdLoTMoxjHH40cju9lg15tJuDDkSGjqa11W6Y3FaWUTcONU2r5Hvphe4Lqp
mdwFfdNrbb8TXKgurI/ccbOAfsHoGSu6irxvEcpyDNgyhPIibXXFDCX7DpKDkhq/mpxnqG7WSAkb
1qO/VmaIg14EnuO8o3kHMxDGauOY04x324dwEhY7Rb9JyjoAQIfuh0nZolScX54Lkk/Fdp0yQEMV
ICHH7sB+O3sxJFiMMOBJXOUkAGzIG0NaHaFrbILxan7zp58ME4ONG8Ape9oeQbN9BoDpmDSoZchh
U9wnXQJ9GTCEcpLThPl2u3nOke5pbQZ9pRVPKNx7CfazFRNEKDYxO8eGtnyZnkrH84kd5lEGlDiq
O+ZGdQfEGXDeUh6djzi29YMVPQldTDUkDkqRt9CVcQqZ0lFQdhXpz7BTYWlPOh3vSyS0erFkeKFm
To8F7UrZ6am8mfguvuG/vlw1hFi7OAw9w5VluL7lk3p80NecfGSfN3MTFZp5JARoN/BcoPnHmcrn
IUzGfPrKgUdYMffCQagp0Dd2pKls4TYjYSmqk+2X3NiPV7dAdsEINyB2Hpx+8isAnLocD7TUWOKc
c1eaNZc4Cts5LA1uCwJGrrlo/r8qwojsqVLO70jkdqCqEtrKNcMRNYWBD6bZ0S2LjGExccL/fXzc
rCWTh+ufI7rQfgX1lnesJyV0vqBn4i0xLt9kjOGe/8kNzgceFQYkbSX0wLPbftc9KAzMj0xM33EV
sZsXCF5U3ehHyrejXwH8D7ORWjg2Te9Ybx34UT9u/d4w/T6EeQ0EGR2dk7P82NieRFZ5u4uNuH+F
vjAA/L61Eaee1KpgssIGt64tqa+5UC5qBrUxM85ZDEpxJF9dGQT0Bj3nOnxWSCJUlSPtJnekqu/v
MuNxJNqlBp3h6J79iVMNtdA35uaHSzp47wY4Ec3PwdjOM7RzavNJ/bsfjC7vzFT6m3SqHEd182d4
3a5TMJgJkSajuPSyejIErepNEqcSVFxQfoCIsbczgv/0SyQ7EbXgod63BaWx+TMomMRp/gZLOrDe
kZyDgc1ur9XlQh1AYvme/PpWXQq3xIkK8YJ3Oh8y+1hdx5iBREpZLBOLXIZCQ9wSCWgMkXR8hd7r
zC7CHh7CuITvnlzoSfeLSuiUonbGkvtQI3goaD2OyGBT7PoKc2bC0X4QIARGONjBXZeXUBOZ/KHx
er6zxiAK0BrM4/UOORNst6RNQUlFIZD8cUsNO7GLWj8JUYFfJnjnIZ4XChb979ScHDODUSBVlT4b
B0MQtWBHNXUiukosZWXY7WazcP9OFjLh/h7m6MpqqCbKqU2Ic/SZs7+YPPlVE8AWBDxfDJ6j27mz
lJEF1VLl2u8fDR8mdwO4RjqpW7MNVtGKc44QKJnMhEsuTqSi/yFyIhKnKAWHU0k9jOJ1RczjG/6A
FiAagyYBB7ct0QZb4WqF+I1qydUaaB4pRFoILuOaHcPTqd2lambIUMz3cLgJACIj8bj5I5Ys1+EK
N65gfHDAXEOceOEZ9vEBagjraLEO9IDi9aGAFDdd9cxmIAZI6nlFErxqAhUJI/Z/kTnJ/8YexH28
vxRHl6XRmKBSofDwZKxkJaUcmA37ik3t0dMNuMgI6zytU1VMFiezq6HY3euJlbvgKNtEreDLaSCa
7o7fU7qp8dbmvGbQSAAh05t+TuVb8VpWNEpiVOUA3s1EY5TKUgEe4+VQvcy4P87XL8Sf6oHC1/6a
bxk2DwMlQD+Gv+9udqMAbUKy8JsMXJ/X9b1dhMjZZkaCowGkIplW3+J1BMfE76L4c0sSxQecKZjP
CQFLrg0bN21qiNTx9r8fDIFj6BygvwzzFvfAsVzr5b/sCmmLWiwbr0ZYvv2pGCxmIsSGSbZcwLRB
MM4zwwGuNVUAs9tk+BTZ1o9UbXMuTFegD37R2LMBySTxQTkbzzRY5kqL3YKBKa2C0o5RhdWJ484/
6jvPBuCc7cqC+lWuepeJZq3mgPnzf9HrirBFuy08BLmYoZ3FV2k+Cjq0pppe0lY9a/1FNS7dPwrv
S9I5vA3fusU5g/JSp8B1pdpPonOHyHE3uOIuNWlessgrlFzxh9iPcq4O84TAQecnL9NJKnLo2a27
C1HKR4XMN7giyeYKAKRotZxqWGWb9s3WV9AsDe+3jzS+b+h75+SvUhv5upU83Pd7fRGvIiClZoML
g37GVj0GX9ZLT9MOck6GTFvIGadKMZha5LUrhiP9NOCJKaSY2NGpxFToyzMtK/MsIvF3l93pCQSm
n5Hf3wdlhaVYxoyVfjk4rKglQosY/vZBEwzSb+nr6xni/BYsfdX1u+IjQF7vKh81a1K3DNOx2bVc
Kz0KnUwZGax7QNen5eVYwZ9TyvaKN3ioTtX+V9W8kRcSBk6H8td4FjuwqqC2p7ETFcCXrrKYM2Xe
kCDt4mYkgZ4C1E4cyLH8nasGdDs6QpyJzmLIdskkeClYiUHiT8dBNXPNT/q0FwXJwAZyrgQ75B/T
5cFKTQYK1f3NNwlZNH7eSREbW2gNvC4yLWqRV02Dh94QQpnN/EaQEWEQEaNAEYHFcwy7PU0AmlUn
2edb4uIVmMHlZdcSPIDdqdqUVUtA3I3MG04O8vENQBsd+/2jkn/4GnhvKOOnpGdMhf4DpYfjkkrw
FYKwm3S+AOu5kVxso7+lztGbj+nXEmDY67PAx1gpQ94cAOqy/2QzYiEpINdZCoDkiFW1HRgIKUtY
Y8xohIDhqQyzHjsThpg2fhuXR0aijw1Y5Qx84ymw4z8er12BRWQ+9xHMU9NYiXYQM9s2fZaeI/2F
uLQfSn9t3t0HBf2Zgg9rF1UxxK6ErqBCPHI9R1hjxel8edSwP605syf/MVt+0r2xBs8J6AUL0mDo
6ANf37EbeapOhL3Ep9z+4pNCQpNussMjauvaVMAV8O+CuTtR8xozsNEV0z/OAUWsF7lcgH2SQdIE
uZ+MB84HDFeRR002fKp1qh2AhyB/ghFzeLXfxOBPi2zeHcFSuLeoEnyU0S54NR/hkSLk6bT2cWbR
CHosh1PzGe9jAY1qUt7q6tZPPlbaHbWV9P8RsMj06q3iUPDm9i9iC46nWIAm8MM6QDELubzrRXCR
+S/hhtMUqHIF5tHeWVpY/tdtg5KgP8ljXB7OwV+/wa79s0Vekn599t5GsVlI2RT+CYK7WgWHGlzH
i22WDqwmawJt/G5MQhtkiGlLuFz6RvC9BfjBe3ztua3GebDEicSbVp2803xkadUt9pegVyAB1y27
Wtk5bnFjAgZ4B8qjx4vK99dhoHkQvsXTfaFBDCexnTikr/zYtALpEbLU6jvC1akeM8vUzGrhLVrZ
5osn8ulxgqCIrVsN6R+j916MXKqGPWlnBT1+W713k8U13K4Y9QBBpcccIc8NhxTVbNgdSVHKP6Tr
CVwe1i+Cixc+FF0qD85sqkkHYrGAkqiDo4cCWvFSh45gyBmcgVCBJ8HZaOEca4flcaOY14E96Lnb
UbYPAiov3RGGWgC8ayHJhdIrk39zexwU/zJ3rxueavDAhBZWHCAFkm6qJQbTsZ3xtlRIRYxqrLIY
TxZe8w0hJlnqR5ibbX85oPfKPFuBU2LOMU2bSXeznGkXVBS+ZpLAxY20vSOlRbmkPYCRZnph4ldk
kjLKSmSQMan7GNYFQD4M1qI5Ea9d7do6qdUH2UbB8+XY5RlXsYU45duIOCI6L3BpcuLFzp9+iLik
3zc9jmR7xaTR4+ykqC6Y9XtT/U3qplk5cK0zENiCEhtSNDRZmySmtInZOjO9Aw9yPoralHABoyZL
6Ebjf44NFV3fMOckVReDkSe4ipjuLZCVwGTVHQLU0FMQgH3OFzTGJ2wmypSGVEjaqwk4EPX2XrxW
/AHSv0M+jog1WHkdROEpTCeawMuiM/cQY3MpHiHOFclLYlhtNnQD/VUFfxPlsIrGA+v5mFCEPdVS
/X0moBWwiuAEURU0ohbLfMLlflwZNx4LrXHL4vwyA6Epgccju/AQgUSAJSRLSm0coNZA/JThzLYd
PxS8uDa4xAPYSjL2KhLZKTchQwpwTj3NmMssJBWOX+U5CuvmXPRSncwiWTTKCw0EHvNNKMZcWjyB
Uh0BvE1zt8vY7k3Wva/krniyM79Y1mKsTetBUEGHI4qaf/kl797VRkBbRPvdi8sxpzX9s4K4K6PH
Gkb5LJr2qiJsURhVDKPnRpmIIRxwf2ElWSKbBT0UE6xe9nMApjqMVVJe4wklQPJ31ftIqzYvSegr
EzfrbIE8xF6lmZ0B9oxvuFwKn05BMomN3fXpzWBP9DnI1xCnrfBYJhHAa4scmcVSHpDdgCuaYP6i
QkVFC3ysuvLHaDYQFwckmMfb/kR4niB8t/qNEaaJs1KFj7yc7ld6QX3Cd8jHP7nuO+uRC2V9YPlr
l3of3EZYUUpW5INR/ScSx6rVidC70susaHyJNjnv7AeAGOZtB/20k+ZOQWAXY6W9B2G55OVmCvLX
1K+l6/TfHzv2WyADvILUUlIaFL9fdwSl9kVemZ+xvxDtXxojRm7Vgc6naIuFis4OcRWKB4Rnrqk7
6o23i2jKsdJJUc36AiIrv71e9dDLv7mReo0qlkyVyecqe8qTxtHdm4AwS8QLCVW8BiG7GPWCa6Ej
j5hBx/Kavirr0FcUADzwFYHnoCZoZEcY1WOYZVdkh2rptXij2Vvwd1GSPllpJ1jAMZiYYNJQmOLc
HsTPDQ8pFGxzmeWt7tAf02g6d5wSrqbbpBUSyFuH/NyK8HfQZDXU8p9t/uiMnWjlvjiSV1TK+e1H
HXEGO6PYrR/moyMEQSMBp6ftKyGYDVA/TowiMa+PTwy+6bcVOUMtRCs9vPeGZPbX7r6ueSvl30Y5
FPUJnYcEr1XU+qTo7Kg3qVJIl1BFZVB49YR7SED+OfGBAg27nh5IoXXoqf4yABJT8aRqVOp05397
g7on+NWSXTEBjnei9lFOQ2HyKU1/G7Cw/SfZX4QIVYb0QPCZwK2Igx4/D4eqwUSZpM5ge97wRVXC
Aa/CRpjZLxeHAXcs2Xl615SmYSpNZV2TU9W8P9Mi5MiYLw93LfXfYt6R9yv//8W1mEQN08ptjRa8
zQst5kxwhi+Hv4Hu5LBfHceF45x+jfkdUvTA8q++0rydg4a0SRsNSZiZoKTZtMV0vyVmhTjTAvw3
cn6JebfkSC6EBd5v/mbX+0ttS6TepLleW2LkFXsGdXMhIJ8s16juZmI7RVBOHnhIOHX5EHQoz1Hm
mzqvwKjq2Hk8XoKFfzH2Fq+K9TEqUn55FuNS/nUU6lwWa/SRohspBmFzYXybJK3zmErFXwIL/fqy
9x9beeMpKE8xQ8WWTCnl87910jiqxhqHgpLCapowBT9nGX3puD967eAZZGA0HGjwHjGzK0LPZl3x
w2ih8sqoiWiwHmtLisoA/BJDBF4kPrPvcZhgPiW9MN/nud5sC63d2pL/Dfl43UjUwGSTUeDHD4YD
o14EwXAGYaVvFk9VClxllHOkyBW4gfeE4qbVmFqUKHD1kJFF6YdbMNry5jL0hI7wjUXbJvUFxIoa
rqFW/f6t0c8W01dV869qH/jVndnOw5T9JkGj2JYER9AXi+VVg69kQ1i+FJMHwPX7qRYZx0/8Ia89
QQfl01m0umZ5tEBzVtNEF2KjlVy3n9xlmRoiC4JmmKQIVJgCJvEOgy18kZKAZxRaLJ5TOnf9UTAI
wUvtzqFxl8geoR7Cm8AY8rwZ9GyJYuhK+4rB/+lTWVy8wRUeF/YlT3aXZzkDD/RbiAeqxPn/v9fP
KLPYMxb5P+DpwJQGZ2S9le+p3GIyeISJb47fj96JzXBbZM7bmxF3EtTGbGA8n/eW9cJM92zmrdHE
mZcmp4uqpfBgIyHQhKgst0LrKB0XC2SQ7SexP78Kw+kgQMblbLHCeiFT02m1MifvQWaIa4CcnwCt
+vRMwt2MaP3ii1u/roltIasDRfAzmblvFyx5QPoMA+3vnicR74BLAmsjv5J6gSOpo1s+9tsSwmaD
3IvBujdlaKMtdnkXCkCXvTv8fTG1lxSwQAzAlGVMMnJ+a31HDYwLZLCb+NXPnPk2YdWtuhHSpMAl
y7eQ398S37x/NBoi0dGOa6kTwOtjkJYk4jdgC4n+GZDL65PGAbRYPELwW6Per5pQe+2vsSsXLibi
adSu4lZoEHGqZMIb7mQ3QrEZCIKTv7H1CErlPswvGVxrohcd/WvJieMhytyiyKELX8PXE5ZLbqFs
CGwO8cZMFdDa4qFL1qTPMVJi0zCzPtwliYqUfSrfdVTBEeIynfnJnKz9C1VFFOTPWgkbrnrtkEnx
ny4zQS0zigswFdt9kJO8xYDaILrEIlk9xhLk6BYEzmpgpwkhLfvtDkTjOUHFGbXxwPDVn9gSJhwQ
fA4EeKkAzPpoSeQBwBeUxFA+WEdIH/eMsJCFw8rm/+O/YG+RGcp1fvNSDdErftFWOKbYw3b9Wpfa
lz/PjMY5i8vT+7i+t3kPlDgsFIfKVhx1Si4OUTxJ7wJb569qgVzFhMefqVtEcl/705UOEzIJfOTb
MkBy5rgklgwxG1O3o/HI08BBaMcwUyH4nMHkeQp9dcbTAwz17NFBNXlTftkdcfH3CkPyVxqMp3sh
ycSlJR4FQHqxlVdeNaxV7i91GCtQxlkmxbSQHdD5zXm9+LiW7PkSZpWL9lKzL6hmHR0oz/TxHgmO
llbxMYuMZhw0x63YKFgxmDTrga/GzE2SAwUlw0sdZgrq53PJ0AmfXpAWfT71+cifWx4IpdVk2MzZ
jNHg1W3gkx8ac+mEZLEk3ro2Em4i7zF86pfuWN8yQTdhECAM+2T5oLyyoKdOGMIbZ4N/6Avyj7ae
Jep7eLjWhv9bBdaewp3ghh0Lif4FdtdRPvwGfeKKWYoarnilTBp3E0aJEY7iKIBj07MScnuhmqyk
ulgqOcIwQUtEQHUvaJwk4GZFpfKoRITAvr6KQ85XqHA04VDVJgPw4k+ycV/9N/odZkf6bXop9B4/
PzpDxqohD/gYzr6E+/VDzBehUlBlBChjUIMhYdtljEtjnVgrNCJH55yNw8bQusNSrAZyeDLgzN/l
h7oMFooJ4kcz7M1pA4Z/MH6qtQ/TllUS/0HvIjz3EKC/QqBXxXGcKj7MjgSMZZYlhLV/fJOddVsL
3UtKJd2nFSvyINdXWj4sIJYu/dKbk3AbHGLxyyXPC29l5boixtkR6yd6EHOu8qOpH/Yl+wKB0cN1
K/wfZJTHvd34zzrBPjasBOEkyxs3xPns+YyIRHeY7fnNF5ANRvPdjHxnii51R65oU7/8bnlzIPPY
vhUPjqjH2B9xn+k7Txga8pShytI9CupOBb1OWIWe8f28H3jatxJ9MzRKmuCIs36L/vfZHAWlddjN
zX7yJ6qdtufNM/uck6HkUqExlH9FXRzkYFqJnxnsRVGPBsWRwfS/Hy7iw2EK8+tK2DkZVbzh9hqG
M/p81cIgM054LA54OxLsn8khNex+xqJltwiERA0h2n7io3oYBBGBjeL0RuP8D6+KvaeWMPz7p5+o
EWx78oO8rj5u/LPLz7z9qrCuo34k+lUPNpwYicvjjPEggZ98foXJVYJnc5nflUDg0aG2n67WfW85
1bq7N2UUI04GOyRHTxlYFXC9I/hXjGeDqCebq/ZPPL6s3ENtGTJ97/YpJreTirkFty/xRADerSQj
FuMybqEY2RNZc07RDCLq1IZ8rupBPs3BYphdUHG0yMav37elaQpHx67/0CWGnxXYhoRQfP2wwMla
xuXrlpv4ynwTp3wujoZmhgXwDsJxMcaYPSXzoP5/OtIJP5t3k1YnlB0J/KlgWCqdEMYRHdsDWDjW
QJ3p7i9BUq3NPGXYBh6QR/z2p+mcrsaystivcQwBydluwd0JRpOFNczzaVLUXeMnKwLrFKB4/3yz
QkIrWjzdujsxjr1xHue9AzTPqHn6inKElm3PrBP+98CwCK5zbEWXtny6JpUOFUdnxzLF0BPrxyOs
VcTmAbAhGBEHm5a45ZYMHXMopN4BlK6A/JD1JD+EpKlUfgcwk71bC5yaVslKn8qXrXnSrOiecMwi
UcjduPr8jZhZLW9QdnvEkEFxbJtMkc4Cm923URe1MEj8SGjGu9ae6LNUFjXlZAh8+bFQN9eL5K8n
pjWp8xpJuN/OBQnR9GQcZ+oRXuqx3zX8WJgtmltVHVEDOTK0Or/J00zrh9/1FRgkPPjjjwxJKaKc
kioc7DfJ1gwoUKf3OqpUBISkAosjPp3TAvx8/v/ELIXy+8P786zLzycDNAiTwa2A2+sXfDp1G8Xh
uU8J9oGgoClO+ERJGg90ls/9+NZMGkT/RzcNf8lasqZKHKf39o8AqCkgLCjG8APVrnv1vJuWCmAx
/EEwrXohWzZ3iD7n944r3GFsppdUhNiwM8BruVUooR0fg5k5qDOfeo7568xlwTDnUl/wXdeupGjW
pUPFXbU6cL9QQpAPUyYGWvQe/EK1vCd5xblzumhY7vAN3HUeE2TVbpE7qP0m1/PJLteA7q52IndB
DzRe8qfEyQmGwMpAVALgs9oH01AvDsZnRPymFtIXLduhsX3PKqmYAcWWH5dWvrlZtYVow88Jt2EH
VrupSdJw6R5N4GBsyb54YgeVkVni4BpwiasoI6lf3kBx70gm1waNThWeEqN3Is939BNeZwNF7lzH
kVva8rPKO+gIrYogsKn0dR2YdhsvFGQNQiQsqXf9Jwx5IITA5Ae2qyxJzFCVkRR1lQcJcvq35z+D
Ao7wXZaY+gEr+un5yLoLxiGA9Kq6yvhuFOG08KKXaFhGcYpbnIChrflVo0OowpkWVefLf41O6Aqs
N46zIqpXJjIO3CbxtKSQTF4A2RPB5cXQura6F635GcK0q419LQcxG1fGpr9ZU0kMM7PU1692hhYC
uZ2gek7DLVHZRSjCjuSkZG2dtixYISrUt8920KIkmge9bMuY7H2M6lV+IB7A2QXExbWI0UrA5Cn/
YI8TRSol3JmpLK+yczXnR/JiZSrs6Nt5lKDmeGs/vGazStzH5nnFSZ9fBDEQrtpl9i2w5ESvrPbD
lBwj/bnpFg1WRtvV5duyv92NEpc+c4lQVydkSfGHeUIYjTYsAQMcjeD7AMT4Lq/Sfy062srlKadn
MMguinmSZnddCysraYOemM5/ajX+j3EVfwrSBw3RRmtt2Tp3uu23UHJUweHLwqVVE9tuYVJ1MEQT
PeQldORK0tacUCxBcXAKnmcJ/wHWFzqkI6Y2phc3qimNPEiWd+WSAidd1dBzv0TVP0hsnHv7Dabt
JVY8Oqq/ojMb1o56unWEIjeB+Vbp/ri+//yUQK9+6H/M0y0UIIWfYZzhsc976A4tO2TvnljXxgtC
wzl5PjiFLoasxnHV3CWt2MmQrsMDpx1RIGA4h5m0anRrhlf7kwi+ad4BpZ9ut8KZnChdt/0uFXjx
/2sgm+7vQGuxsCjtmekX7FZhxKv9NA9nYh7Mm2MruLNejein0c21dCez/pwrKu55NO1Z+vY3WEEh
T2e8ewO0oXz4tlPCNQUZ8BwN3DDI2dGulR9cQcTomYN4CTNP3LIUARPifs9QodvEKMncv9t/DWy3
LiLwIswaVshilAfjOT2R/lNvgIbee0Q1vzDl83pzQnI9Qh5ikYUR1CHeENyuppLIbhnqNnzmwX7b
t6SetoWURe85zlsaWyioQMYwrXUoVgGUNPFSpwAF2mVyX+EmiPqCENJ+t8zP2IlM8ugjAZ+X18V8
Ngicf/T+eIGzgsE+scpOSDO+4warzGdAwfvo4OItIZoZBLVjX94K/vqyB6BwePu7UGHrDwBUcCMJ
Ez8DL/g7kzaYUOcP2vkk81OsaniGvVDd4Pxbj7mYbv99jVJagCkComxKuKgYghbt2/0ENjIcYLuH
Nuk5+EBu5EcFmJYWwfK4xdTTJ3ayS8EyNE+YFnKeKFkrbZwAS20uhulUxUnPpFYeZNV+Jz8loCX9
TcMNiy/iE9Ttkl7dVXNr69vO/L0G80E2ddlxUmGRCG8eyIIlR2Ge8z335c48KdS/LnTw5rzvL5Xq
Jelzu0KP79801nVpnNTwChcHpjwILMfB3oCkX+3alFF3HzNE9p6JCaiD++DDXPREtP6bX9+u4/uG
C60FWb0nI4DZYgU5zOJVB918z6fxs0U9be1J6GD8KrE+tpmSqKrgqd5KymDQVGqq2Q3MFGlomKO5
J9HAX6KQpv53IyA5bPYpsLLhDH0lIQMhxARmj7/YrHm0I09xv1/QYa10WVySlDUm04N9709MOgSW
Wm1jsRzz0YGL8gPRd8vYky2/+mXZNzYExi25d2vO79DNz3EyzCmQT4jDpIlVM8ERXKhCQrrcQ81e
Vm+eOYRJvvDXuqoDZy2vv9Uy//WpB82t/gYjovsJtb6pEYfNXWzhevA8QK8tnkbDDQbSoCyyOiPg
iHkRYic/XiQDJBYV+xlyAjHpMVMuJohYuVuqRuz3PfVsqWL0BoDMc744Rg/TRuiAVHX/nns2LAni
USX4g3XaBI4eNybFoJ317emZVjNbYYK0zqXVqrkp/P0PDDh0B5SsmHnM+yvILe27+slAxoGPreap
V1D8xn9nQeEXQR7Ugz18PWmEi38A3rjQX9koYkvEBDSN6gGlIABUYfKCebwnRxXokqvn7YVKOZYu
YWwk42gHSn5FJ/qZ3aUnWw4JUnssqiVnGDUulyfcKyXBN3LUQ0QhF5VTfoVMKHWIByx7WjxncpaH
sxSJJMGuBfrLNAKngnwGa44D2zpajigHEYrP6cr6fvDAdd97cQPIBjoiHJdJz8Gs5J3lfog00ZqB
+BedpE3JZUK/pAp3TiLDipdMZJ6lTECjijc0B5HazBv7xWbbsmQYGihdn2Dfvh2g/Tr0ubTE5phD
d4pHZYnVFz0itXDbNvL2mOinpadG/zA0T0MHjJUKxRgfxx2PFlDHB/GopIl3QKoPN9Zl2NkQ+dgM
QNcAwz+uVdfAdX8+AaPsXYasEQnzdwxwNY0QuqeH3fVIuG6W5z6bzhOlzruvcZIrmwWHWmXVrLtB
lISSN5hdhRc526oi2FqYMReKo5lVH3hOi9J/jGYgFPgjTusuth+hzTIK3Dmdf6PtqOKVtKuyWOw6
KHtjXs+yoK4G1Eg1VZi/LuVt+TaijVs+t7Hot5znR945R2d8xBdPxm+7pOCu2NFkZKJB01lrcgiN
gMb961CiCi3xd9bRVm2jQezw81PyUzziPYcf+0gE/dffc6Vr/ul+Y1ZHGXtjnN8cdvinw3z+M5tl
uBcWI7ruXMSL345sE6HX06ovkaK6mT/9eMYBNwNvI3i4ub3To+M02tBqO8OU/ObfogVeFUq3ah/l
k5pQRh6AhLdBwRCyxeBzf4gZgdLbECa8dRGTR4JMeHBDLtgS/L1NR3LhCMv0oG06x867TLzWh81/
Q6gK7Bi3n4KeRsKn8Cbv2xmH2fUeQYM4EQZ2JZPSA4blyJyLD22uCS4PA/WY0ATQMnfDnRqgSf1R
KFm4mxWp5yMi7ga+ec2IrIzxDmfDeSNZcvTUXA77F3vM+/d+BWhOX0RM5tZxNxpRB3yW1vDFcNOg
5uurNn0Tx1VYNHm2OFImAHufHN/uIIAtyCEimt5SxaHHTIIDbF3vvhc9AssUpSrt0583voOTGzis
LLIPafrlDT/Zr0of61GKr7DclP8P65sUTZBaX9CovxMgBNXSvh3lrz7SMnjoFOIkKhEZqou736C5
RWpR8rGVRhTwZJfgkaqrUwAyt7comiYLf43gZvAw2NZjfoGmlXSGSbfttIRFAOWQiBEInrs8Jb6W
eHEKE34uLF5CNCW6AXiQeDQKlgFYDD2GAubUzwOMAokAcE9aSmQ1hOmEdyk8pv+27hvzt2sqxEaL
cTaoSRdngM/03onVE0P1C/1Nor6nu3IHt3KCWwGYGp+yjt+aDWvIfLNPGf7X4pk8SX/sxbHLddbn
GDMaCGk6nXcqjjxgdOzNC2SGF+PgctR4f5g40a5BLOd/aYsTY+UBjTlc6nqhOQ/QJCQFHQcSuWVc
e0YHz4VojfhC6NP88c95C1asB2AWMwu6mQwR4ozB2Mn85r06xpZCtAj8PwR5DAzO1FiQ8fBi1eZu
1Bgk3gLssyfyPnOWMVW45c5bSY8QjgFEpJuvzuc9fQ/RZQ+epawuU3hRqTSnlfwzaObCNF7ftzt8
rioV2KqLWCYzJ+HgLc+O5dNzDBc0b5rR0ov8TR7+L1U/dYMT7ON6RnLiQYXN5ZkUXGgDQOit+zc3
EMgV2jEhgINTC66dGGKlaFVwlEs3iJFCYv6WxlU/JtZsDRs89mHtih8KAfNBEzJxKJOFCiRQdU6x
dglOvxeGxx2mpMhdXACDkz4WybEBYrkakPOGkyOuhRCkqpVzFtR0XU/mdtfSw8pQAAGPpKpGdcJG
PeqWFTU17tW4ENDt9A68z6V0jpDDInyZyFnxK8O3sIqlHAdu+9o8+xnmahvJnkQwIqdugT9du9nc
6jYcwV33FG350F0W6l+NCsk9zZGkCTFQoGDmHPSZQs4FAr8yjf3TpI+ui6cwIdbo01egdciRAjLU
cytroIg9DdRAcYogxMvni9eFNH5mZuJ/GaAF2YZy97yd7nLc8e9CQhS60Mmxaj8xxhsn3mox6R/6
/6LSg4Pgnq8GnIJB34vrxkhX+sIjRRPtXWYh20ZpgMBw5e65QC2UTpvZnJthgzhgiIPeKj2WverO
451r7vLlx952Wz9nMB7mw8XhHWU2BV8Laxe9d5gk9x/GIGY+36UiolToepJj2DR7dxun7yEsuqx1
S/V20HXjKLH8kgoh+fNAklnYCyym8FXZyQk1FK4MH7JbH8rc5vfZnZrGCdEYvQenXcd+ejknARVO
nhhmNPj9lrJuabJUg4G6+EET8Wt+A1jBVt8B5h8nLyXtP7ftdDoPK+Tm5CpodgRo/oapzS/Lmx0d
vPoCBX6evdU+s5nNAd0qORVunKkRw+eHnDb5X6W3g1Y7X5lOTNT1yL80Y+pkCrxaoC5Aj/IQOChO
0eKrbLBQ9Caiu1TFVNQgmA8djC939hjxw/3JoTEXfPnyy01syRI2FuQMzcdSxAhYKzSPbgSwaeIj
XRPO87irSaQH5RjRdffR8LD+AHs7NkvY49+xFofCPE3Q2s411Qp0aTfTgGJybZWB1kQLJBmavTHk
+kd7ZWn/c/9Ki1dAi98BfB89+DetEjexefCBvnNHWYqaBnVTUFK0pX/Cy8c+MHbiB1Ybycrck4fU
C9Mv0AZyYiylMbBqvQY9L4kS5JHuVx4szjCEvu3PpQladgsEWaPGknff7tQABh4R8uDUXyBwACHE
t1N8trACA5C+p0U27/4yfQ5WishSw2Z9FM0D1FwEj5I2OlOJUecRFxaKP7ZWsqJax7oc+fIWwr9T
UvcFBNXASg/Wi3CbxO4aUpZQpQkPTT/377sWrRJe0BysADbQRMAQXI8TILTDqCo5cKw/jPaaTonx
bkGeMrhxEU6Oriv9MFA5hxDWVpMllzX7YOcnTzSQiNInTiNqPER/LSmtaNWmjT8IUNZwAT9IL/7H
QNrRZWBYJtpHe9fUFGgeiddE9DyrbCOCmPGqTJ/Yu7d0xW7/pVY6cel6u5sSpsdvx4U9FHOi65WL
09lnTd/F4+qPYgEFIrssbCywxsi+FLIZINAAUF3ZrR2usTOhp5n/tx75c+UO3GQf2HXKruMCTLO9
SAlq3WsCAqAiwRB2g/W/FmAWBqc+rgxCMQNbQ6w05FamZz8x1d5kqTKMNqA/8N7NLKQ+RHar9MGP
YscvgxlDhzr0dQaMzuMYylcpOhJ0kDKoGrAgKbqmkHHkxZzF1ZXN2+jbagSRsh9UOtRysytNoWKx
Nbzy5khj/NmI5c6wNby/bM/fPDe9JxlMEh3gXzpc1V3071eLqJLIYjQXCNOGGPe8hPFjpqFdjLCm
6VwEqddHhd5s6rcBFlRAFYvSfy1OvZtpUJuY7Z9O35wrmjgHRefzohJV0MYGWnHATfH/6GypQXAo
ycbwM5LUo/RRwpZ2jXfqSiW3t0xMN9H75SWypOLBA2a85Q3j6qDXCRdtlDUBGnFT2LwbpY/dFkP6
mvjkVAbkDJf0x9u9FW9s9ny1QY3zKcqI6HNf+6oJXiKtmYpKYd/NTwtU0yRwrQRmHNvJ3FDfdIX3
W4TZJGUJpmKbwjqq7k7TE+GNKU8mWXVXg6pX3nu87+KEVpSGmlqO4nHhtW9cWhUbeQ56wejdnGR1
mPg3hYg73dRnkfebHEvQSmo5aHV7w/jOc8FcPWlzg41052Vx4Ax0T1iwczbsrmU+VnHdJckY9RLn
Uf9kz9iHubU3crMVUP6KTTp8frlyoCG+KdOIZLetmGaHxKE1+c/HFqR71P3ujxEhw4Vef7wwVO4V
L1/JL3p+GEyYQTnzhycuoN5vqqiKj1px6fG1z6KvApl4HzUcO/jPUKCnaen6YoqbU20shoAzxWaz
R1ZOpOrdo9Im66OQoL70pd+tvJVmIrJiSZyRHnpgGx1mMrTtH6tIU56XakPEru3XmDCG6erEZ+8C
V36QBKawpCH8+uAZWQyBx/5scMZaxEoi1NuJXTSWHZuDp3gMBXER3ehEgngqEuf+2u7uJPkqZboY
gEq1bOz40EDJ+eX2Rcw9arW2q9pwrJZCdgjjTK/oW+ArKsULOMHyDzu/1skR/7p1saYGSk+CvMyF
SQeBhKaEdFpBIp4al4QgdOaukUrqzqBsL3Er1Ho5gMnLn/6jUMC16Wl0K8jxuGfNrtXZfEhTRHYv
a5kTr5X4aZNa3VtQvaiIa1t8YODTh4R61Llij3TI453IjCZHgUdO/ptkT9e9Fxp1Zl8m3xtv3KVV
GXZrKe6mQ2xWlMOs2LGz0kWQcBl0WI8ZtRT29H4htCpz4uos1INYrEHgkT3ebBUYaMeVLA19yeiO
rNZ1IDa23zzKc55MTL/b1XqKVP+aXxF1lI9l4Iqnpf03/4rB9QpFZRsze0IT9rOP4GOisA70UFta
r8grxB5Qm9SyS32kM7N1e/P1d5vgvfFJV4qD60/C/M+Chi7MoLpDD4TcaC8ldwJ+G6TWvBOaUmtc
IZaQKBn1y/kNjRr3ftHM8Wl2wMTY0Uc4He2y3jWFRIF+vvd9TmLfycRNnJkPFp/Qy6alLVfUGtB6
SkKiMY2TjY76kPcFXVmSFtRKP+mHJS+pN4sB4b3ptUK7hvp40mqKmjhlSKj86zoTaFzD/FkF911K
rzlgRHCryspiAS3Do6pn1nAwyqXPmaeHQHMhKXd92bE869yB07FN+4HboaEKaqyrNW8pF9Bzz8xa
oEFgr1mRR3h2OUGiaV+jqXbcgPPdpiPRtJ4OJNVsUcNwyU7uX+KmoUqUX/kqJjqpkJWEa/yUKEXc
n4+vwek0EJV78eMpBivMHY8EJwSKyCg2YQJi9VNBMaeRoyUp/IeGt1RleuIVJ7mztQmqnR95TC/r
rY2TJ5sjW49wzfyd9umOeBrlbRHHukYNk39e9eLGuYXJPh4t1sJsw0iWrEOAHWXqN1NZn8MrKcn6
k/xc5MVdBWMLPrjZ/zwg9oSNNu5IhuBI9grurglt1t0qDKLYA4zKOVU7SQPltuvJ8JYMDEzDHpPb
le0lVq3D2LNPh8Xak9G7NLmayNNlmZV8enyVps3/fKGwFgq5b1UY5fhE97brUs5wsAcX3yqrwziS
AFSZfYSZVFoLPsmma9aOktxpHNJC4eXHAJoFAUY5t8leACkou8mp8471AwKD2ozKEjyDUMiU5/A9
KsAr9DZS02oGzBOCqGatXuQUHUl+9OFLQmRsRwmxYuJj7FoMHChX9ScImxiGp5Npc+2UHADOuO/v
szFPhGB+a+fpd8ZNUQqQLX0S3HUPHbEtH8IwjiTA5CX/QL//O+PhVWhESMR8dxSbbS8pJNEdxGDV
4ZaZn4994jLgWv75qjtEOtSqQEasUS9cra328MrqvoGTngtuTmF83sdw1p+u20lW9u/XsddSpv4U
avvR0zKloos+Rtv1KPxGvfkUBAnHf8cf64NELmjru4Txgx2iY31lSt+5MDgfOWDRUymXBziOhMDW
J2XJCqyj7MSMTRFaxZpb0ESjTBrSyuL6yp8Rln/fsnYRXhq2yF7xMgRk1swNHpS0FFuO2jDE8n0J
ObY+xalfLDSiEbhpZvRs/1SkcStZbdsEpqNfPhA0UaUZmbt2Zt2hQ3Vh0DphZMQIax59kgoV0b8Z
55DOKpRnBxFIvHgJ57+/EZIR5ivGBQ0/OBfzr01oPWGhUza2EhJcqNblqwr9h3Np1LWjhp8hdajF
4N1tDeDe91AzExdrbs8M5l8zghf10hDF7jKgbyV84q+19iciB9wNyLHOooiHKbk6LFQgQumElJix
v75V5eqOQESmbuB2HUITVh0ogSwfCRLotJUe3nkspqBvOk0pUA7ynYo2WXREpLCNU9+suDW/AdPm
AzTBI9F4eagERlZrVRpEqNp82sqr7DPsQBWotENuGU9nk7OAmBGpmf+abnFnY3099LWVX4b1SoxO
wyM914a4bkSfePXo0BylHnGNSivP6EF/9IjKUd2fcEwJa+jWbfwRAkzDHNJ2fjZXkzOEPbq1qlkN
rQtheulRH14kVHmkwVA9SpDlbJlhMURjixXBt8VYKAIrtU5eAd+LDh/eTC8IXADo12WzT0Ev0s4w
vnvYVsAa1RMk4ufHJFMNeHEj5AFvxBi1QFzmY3qUC+JtJyP/whv4xH4ckAAOeg+25KJGZLGw+6vk
ylXEe6unawgA7k4Ne/oEr+A5MeMBAjK5EthNl5dc4C3YOb6F/Z3qbULdNe9ZIv8FinHY2NtvOuEe
t8nKpZyKrIJ1cZTPK0IPEVhrSOC+dMKrRFiHYNKoIki7YSlcuI/81vi6ae4cCWcdxTnL/Dc3hUgA
mSW/VMSa4epU7BbROv98pLeTEeR7Ffe7PEUaFVE2HdEvIbGqnUzyo/PV9t5P5BuQ0Gnz/E/mp4lp
3k2qPv7YUbS3YKWWIPzBZ6ApKxfzb37IDGA05Yj9wmPfSRjr7ydR4wt6I+BR8oVC25qGYEZv9xY6
n9LzxR/JrRRb+by2P+3zcbttQXgvZlNvduR1k5cWV8eJ2yWgip964Srv1frk+9xmQ2N0u6E/v3pu
3OTymU2AkfR8dLLZOM/ycgFiPJQy6dQY+XSXja3A5FW1W+w7S8RRQirnJR7H52COcS0/5fq2fTHb
VloPZ39yphxMCXUVHGaATdAklk4c8Sm7ObVUPgZ6CRRbEHx2Jtg5XVGQAdUHFo1p+nqGGolu3YJe
pdzG249KMs6fxUbfXwL0l8R9T3heJdiujsy36o8tw6hNpfNV/FTbY/MEWMhsjDV2G27sVzmKeRmL
Hw2vpxru7NvBQ4e/qebMsOcVMt2YiBs6/lyj31Mqa5jkvwBbmN8GjorJRT5Mm+80j9lZIsvE7xgy
rC9nC5jcDuEmyuaXUc4mSYoYTxu3ycBwz29Lkl2C/0sE05HeBwHMsT3/lxM6788rJIpPNnmDfjca
HJKYViLukWKCkNCXFgyOe1FCfBpIRqi7Q0tW079tIJ/5YThhGcrNhZyDJ+oSVOA8WKgUGVIMTmob
LgGbTAJlINs7e5bH5iFqtkmvYGmjq106DZDUvcp7ZDZpMVjv5kWucrIYAuetyEXduSFMxYoxmVzx
CZgf5sHdGKv8A/06pk0J0mYfqD23zk7Wl7pujvLWugXIRt1gKOJFuIsdJs27dY+eMcmAcqB3KqoE
gK8tKoK+mTxhjLiBA6VvEiOe5awn47+mlrdNzxfO5A33HbcSF9czmJ4o8RlRCXpEMeQ8dnz77C7r
vdWxZEzFETuttyZU+yEei7//Sb5DEJe6BjtRocXgnNKUpVcMUIehYrZkLWSGjZR5SojH2fnZzoRh
bZAtaw0ncnA8Ceaa5J5mHu4QIs3b/FKyZYqKkrAYggcO5I8wxS2Z7lFmzQpJZmdzKqF+kTu5eCUc
amYUA0NTSigiUismnEgAMadycCqg6nx1JKitPbFE9ODIXWORQookKXkMP175AvxY+YX/RIOTgPDh
sISn52uBOi/XJWV9hcy+O660HEBjK6tnaZYkR0r3KntLytluqBwdkE798khGln4UHV/IXBzOyQHm
5LPrYvBe8S8IfBukGV/j21lLMUCm6pkd1ObkoMgKHmpBUHRv7o0Ywz6k75oaUxt8KinyzlRsID+N
OSGm8xXvptAwkSaISUpnRTVxoNCPd62Civujvwvzd3SNjphwdAF7UEEgjCSDFVuVZB3U1mCLX1Fy
2/APY5wMkzw0hlaZvG8syc7ysxP6nVWtP4Ggi7x0qoe2Tudsnp6KoVy+3YSBR/VNIrVsEKSFSCwK
PhSWQbW03tTJ2PtLbFSJhuotfmfNu0wlXvhky+gFqHgWrmrVHsVJUfRO57EFInuV/talxcQYJOYD
g/weLykGEqcjibrM1j7VMHYnpQY57FdsAOwsv4SXLT0DhePpMAQbTvjKncDkfKaBFuG79TfQ7fHZ
vibDFPYligD0gt6ZWGHh36GAfC7Ajw/2HM9ZhL7JKIv3YVX1hoOYYePVLRRRDSGNUV4tNyfZ/+wf
dD+YqD8HvDUfRmqZ4lhYFP9ZfVhy3vf5ZkqD0v8yrYQoS9Gh5fewUB6YnIa0hdcTpJC1poZ1kOzs
geNU6F9ou3mon3pt6nxeW4wLn1NagaZQTpw32vHEJS6bjx/tWlmIVM/IXtis8ax4XjAq4mmf4V8Z
ppNGFfOfzug3n+t25q2Qi0ngh9IjxSptvy4az3JqVQgR5MIEtASFSF3RxCntJ4RVeKumv0dpzKPk
CeVDIQJ2I7KbF79RsROWg84rm0zbCRTklPfhdN3JmRBdaERaBtd0jU/BjpJZzfTHzP/lJOy/hx8d
ieC7xMACDKJjdvsffiBXTLVrzUibKIApK+VEbbIEpEKfplJnj+ym3vwuMI500kSLHcxniSGR52i4
4CJr5nlgzHkCpdpvG0doWrn8kE5Fp0SvuNWsJ6YOvuPghRLKVJ3nxLnYBk6ISYx8GQ8XwnBZr0qv
OvquGJLmtNjmBSX7fSFTovpZqEyEXst5W9T5J0yGMEgOn6pSf8y02QXpRzPq1EwrX1pLsAAu1Y88
hPif/IN8WLyrnUY4WikUe1uOr6td2/5v2E1cZDi8gebSP0BZs4bPnt/n+Wr7PiTc+QwnSW5KGZOA
0W+4uVTKNxAdK6L3Wkpx1KQSYXSzQjBP0SCxTVydm6Mc/+dsAoTrjuRMWuChBZYJZbHkFu66CETW
ktjpPhWTAdmpw60cYD+uM4rsBtg4e+F9QNLY31R0s2Zohv/rRfp/obHLPw/aZ7Zp6e5nFOLjvstg
rHzowiFHE8T9yL13fQSWFB8tugELovMJXXs6t5WWqOuvswmJf+d3epB18tp7V+IYZnI4ng7X7rxC
PoLEAKz53x6rl1wO/DyW8RS9rzloCYfds0/goau5lzC3qoxfdLV6nb0OQIzZoPYnYIavmy3O2iUB
3PPPlI+prrR8Qd++CrddA97iFLDUuYqZi/wfih/2oJH4MmcET2/K6yFO4+BZO0KXXQkpelOvwiG4
BLvGUSjYimxALTiH/dNwTgG3Zn9a6XjfZi2yl0WPS0CQ9EX2+c1opOotcB5+VaUDdG/CUJ65ei6Y
6yzh7bPVWrTACduFdXtjVe31Xs3E5BLIDsYbHJsaHnIWqp+dlGm6ayEYrlQXbnlutYAmT6+4pzkH
ncQQlLCBFlyoFRm9Fz3p2BIqKTk64JOjbuoHWwxUCBxNmvzoJf/GxcxChRH+x8s7AT/oyIDrrJ87
DI7Jdxusy7cgGSHUu7nWyq1G10YqYFDJUG+AV5TZrXXikVJM80swQUtoHdDXAi16yMgthPua3E5N
+KrPP15D8zzqfLn28Nmvgoxn63VWgd4bKYxORuGpMSOoZDX9obMnfL5mknb3A3pRaKnE5w+dXXCF
OYBSh90IHJ1zajVMC9Otz9ZG1jhjE3rnjC0QJz7fUIFKeE7OJXhOy+kOay5JDP2xrMStjaeMKtyU
9CDdfy0WkFig2R58c0k4s2st+bC1u2ErvOtPgt6BvaBvq1izo62ssojX+sSs0a2A/BVQ24imkwPv
UNPXnw3VCfrM1K0ZhB/2qa2/PXkpTmwnBBsQn56BdRptkPw5P95AQBP34Na96NMtkteOWUIP8j7F
BtVbw2DL5F/anzzQUNRojo/BxX5lbFz+j4STdhdgx3sbfDbvNlBcaumyrTCCWyslZlHB92YoZwFu
4XwgW/K4nwcqcyVw1I7pp9EmBARf4plYdIpuHUZCwE1KsBcYxKV/9/YBBZZViI/k8FUJLaF77vQU
O/LbJg06e/FcO3lxLcY1+Os2PFCKjQ5b6lEah2Cs4aH/EDlI1HYSVFwHPX/n1CFttEVX950Sdm+Q
a9pEr1Tat/uh6gTXjsHJH4msMvR0PhfuHKGbCD+sfvBmuxYmV8h5kUsZ3yFRV950jgsCB+9lPU9P
rlCErBV3sS7qu/PYUdF2wDYJe01IV4Ly8l39OdT7DQrRhxz1DWRoato9n68+HaQXQ9hzgowt78TS
qzXzUhuNAZxkvgAhVzAklSf3IU/BmcUbm7YlEm+RRBkxdaV24L2gO+9uPei07x4I8jHdOf3IvI2n
yInmyEgI0f7cu+Fcv4+n0aIzSloP0rGMODImGrguYK7eWHZc51KCcfuyfcOES+oRTfOOld14eQhK
iQ+Q1YsSRfYgevOhz+EK01IrKixDixXrqBdKTaVf+lViN/2MQdU6v3PDI2vtRpVOLgD/AKO0Pln2
8Y1DG9ShZ2MvuLQ3PGsmwL711gY+6T47PEUzq7uk7q2KK0N7nnXEusSSbcLc/Ow5dMdpyzqy4mZQ
QzQ/3q03mor8Bfzo7WjfKpYm/Is5M8vEOjVg9vpmGmj74yLL8jEfdQsGgBua/vaIegTfHbdetK1Z
h1DW7+1dOaVzkdYjWw/lxGUJRrrWFj8BDBLj1QWzYn28k0NWyJ5Fl4Qn3gumWLJcKueIaWXlITFp
mBXeSdDABfgHUCGibVcW1BeyP6daDbJvgYIIfWOR/aHek6dhHU1BbGV2kn7ZKUBAQuuSE4hktwW1
vdsrt6FM1DRHyMbyMtVs06VaICZCtQjcFz4HOUgjMcX0QQz8MxzPVCPO7bppH1nnt6dIrTHNXucp
e0mkNHAdj7YTd0KvLKTUuW1qfb4XnGc1F+dwhReD9dMP+MVehmi/dUmUjN8oFO0pR1lHAYVdyZES
8MhKocuws/FY4nfxEJQDKe+vqGLlxOaJNN6d2ECtr7Sq2qYupc2QbWdi1cKcX1it+6zdewmP+FzC
AXBFj/TCFxV/EsW0zDRjo4k/4fQlS4uVSay2RO30ev6h/zwBlCjuP9l6yBQ5lmpYFni4+L8SdTvN
WNN3VZA9YKSbmV1XY0a8uSksHLNPH5NfRqbmNRKGJf6Gd0mTp0l8pRZeV4dnrQbXuJo5Y/phx/xQ
02w/mhinvtB79+JLfGb1HjtLiN4lTt6yWB64rURZtqlMleGnsRTzq0BZuJ7k00OTDOVM7jjZt9bP
IdbZWzx+QSJYcFCqowX0r1nf9wrZ0uTAeA3Wc9uLs6KB3fjQOvwehGPbG2+Mnz9yRiwOGR/HlVd7
KlGo1IKVxmjHeAen92CldyO0YxcAoPk6LmD1l4JLNgoh+6GDcrZBCE1QLqoI3NjRECHVmEqE2e+o
vYxxQdppQ8NMy+y64A6ss+0Ap6Cg38j/PbrG9wlqZAD/wpbCGYbd6XoEYDIhMRxT6m1Qoz/TgjfK
AoUmPGbiBuAPcG+a82lTULxPzva/sZj8syj0IzCoB1o37sCbf0Zhrm08bCs8qc80Q+p/Yj6BjLQt
AYHlMKZ0Tq1etVZXZkvqi1LbgoiuXLEtNLdA5cMvmyYAVxnc0Vg219yRrvig9raw7TMb04E+T3+j
5wRn6kVkc5TIr4eX0nemzV+1SEmTbmEw74u3tvnzMo2GDTB1fF4a/PuQ/L0ybHWUAqhP8nHi7Ywc
wUIOU3vsdnbTzsZUDQKa5+dYs8ItqgNttBfQVYSBoLRSR26uijibuplf5oGx1uDQUD2w2E6Nqqn/
kU9AMbz8unj6ctSbKNmW2yRU75xafCQGiESCOfGZirzrpsFWvxqmLxaEY8H3aHKS7P2t5ew6I6ev
mvwsXfXQvIzfeDle+kBQjTOWELQAFt6jp5zXKhZaHseaJkL6AAFU+gkcVLzt4tqC9EMfW+RAEQX0
oVOl1vJ1xsCebqFhcA+9GJAWAag0Ca+GgtXfVK7r6fsJPliPO/GYB1rPa6uA28INR7qRVm02sTD8
d6JPG90falLmRfylfkM8wLq0Iux+xb0o43JFNYM14KFoZvwgzbWQkcdZ4HevNqy2m7HA/Xf9b+Gv
j9NXXPNlJ1vpr5bsjd8dx4xiycCd7xBhoDteAeZ4+7mBPbGimAePQjDquNOgB7pTv0Kg83QwCIBz
UR0vMatO128psehzVLl3PUtjCD5BlMVM5E34zPmn6jbvIVG17dzJtVVQgTE8R/L4p7ZY0iyGoQSZ
+rYkIWXnwkxmPwqw8CHKHUN8nZJ7e1upcjfwYp+NtKdJBpt5lg4Cb1sTMvycoQhpBDB6Gdpzs6W3
z/XbUTqMJW4usrAoWbedT8xbEIsAPQB7239f72BkParI8xSHU1L+vH7EvSy6Jg5Gn5PuqECB1tfQ
8I94QGDvb4v2FH7+6BKqjxsJzXdF64vHTF1N7/+dgpmzkOlmeRY06glXF8Hg3IefJPdGu300uKcp
syywVS/s/PMHCFVj2EaWJpexH6VTs0Mr5jJd3jD8t9M6NDcfPNEuLlf/Kh1KAU6X6UsDmxVbiWFR
tfL+FY8M4ixfWgJ23iWnOsxJKdkn3IHw+nIlsqt9I83sYCwdSgrQ4gGxVd97ogswcCMSBlboBzFw
tjcJBGFXSc5MfLBniJ+YTmwD/kT8NjNnZno9ekHbeM48CqR2qcKTdqUuH9o6h5sF0W2u2Q9BCWyX
MdYW9oibpg2AyQBpNertwCXFyhIZMRbi8SgoqQwVtqS+kcD7QqB5sn98aYpl+dqAQY5wDZe30EQ2
UJpmpnhw+ezzkjgdsjhS1ExTPkDCgojB/h1wDCxwwhuox8TPkVXXuqQQvUuN10MgcA7PKIIlnwEK
SIEp50p4Ceoi8kDNyChNi6coB9yldMbMhawfhSd/widc6PR4P+fV0YZCOTEmfMeBIKudTkJ8UxXe
51rDHEQmoACOsh1QYtejGX17dY15HMGHBbmoXpyhKT7atcOjOLxdZoKpP7i5a9JudRsd0KUdVmXV
AglgY3KJ8zBxrQmkPvdW8GL9fmjKeEkD5TYxPnlFr9wal9Ph/c8iqWMpr3kSAjkfL2QyWs8LQF84
8kPboYIQDa1DHIR9h6YH39gsfYdQv0S5FcLfLTSkNGEF2U2qbY2v7ix00i1UJMYZdeGJGb4Z0ayD
kSed1eFWara2eVjooDUGGG0SaagfpZklwPU36YHhpm5b9Pi1emQO9K+uHW2nDmINDQX//2eiuUL9
nqB9hCw/WuwcUH/qcPIDZ/rnM9/yMKi+c7t7qX7um13SviF46wAZFBc0Ly2GVUO7SkLJCwMGXt7c
EVdCek1Q5GXSy+XyqprZH7xK+Xb7lZXaB61YDcvn5/k+LwiTFO8MiCptwFFNkUn3yCNsfHcEsSIX
v9P/gUxn/dmkTPrzGGz9v628I+wjZpyiEtUk84DyVAfev4/ySWEdy1vfnRDBbN/wvinN+P01uBss
CFO8q1wNR5zqU19VIjUtHWh2Y7fIwVMP9SHxGJjKozc0CPAfYH0Xg+mXY/Ma6N3hCuR+62R4Ou6v
vdec11H+nCgWN9J+o1P/7sX1SQLaPPi6zIAH2g5QvU7GWKgOcsp0Nl4+vDZbPtMUeKUjL9XdRqMp
TkYS0XbenX68fgfe047nwxOelXEb5ESlqYifY9NLfjyzZq/A9riiL6IiGdAZt5qMPQ1QRLjJux6c
M0OkMcv9bAxBg3SN0EhHgiSPk/xz79/PPxe0OIuJw+5v+ujbIcD5EpfVjLSQnwIkT7NBo2Dt9Voc
ZhJpJbWZ5KWP+AkISQHVZoUs5gY6O1tRykgrmxqlsOkfQC1CLUl6IybqXas6p18xmAjwL7VlNEZf
9yXIyBslkNSWZUcQEzQJFXcGF7FLI4nLrCripsHcAsi4cPSFqh1u4DJt/tJthe2HvUMRd5HpQKT5
WYZGTA9IdPGNLQYS70SA95WKAMwYiWiNvMe+ZVzj5kZ/ilQ/C60/yrH94aZqNn/3ut7E3EpyxEGz
ET/ilwYhx4creKneeThwOjl4lWkDeBixLziK/Vf2akeEFD6f93fcxqwSiEuBYPVWL6WUYf+tVi6a
1l6S5ZvyEGaePbL9/ygQKZzDET8+M1ieQrmw6rWWtey3sb1RgZGjCjLCfE8VUSkCTW3ZVOOlU4Ue
23zVGAnvzToDo/MnJ2zfVJB+/dZbp9jZMEAFtQJsiAf7NmOfYXAcQyetfIXRTQ337G4L/IwKffyx
J+FUw1pcUE5S2XCy6nC4fSdoDksuioHb6XQkLj4APIcEtEcDk2Sq1kdZQ5SV/roi6uWIj0bY7s98
B7m+NwbP+K/fNEjZ+LeFkT+qeH9EGmak28BAb5trwKaljdOB3ay4sq5PYx+q30ICLN1au4Rp+Cim
OxdTh799cAqTtcdebf18RaibCZ+NV3FPMYApA4AvBOWAeV905/pOyZQrXdc4lyDBo65vpHAH9oGi
PFv5gv/NFjI8W23YR6cAtvFyNmnjI681nGtJr+m/JtEdhWVJTKumfu6WnTxy6CW9YSvnNZauhkBF
KZrcGBCFCU8uoPCtax6Y3qAMHGTza57pHyOvHeyL7T6JVCAfdKdrFfwi8adLbxqyAS4Hx9IB/k3T
qXE8bKwuOfLEN61P/aM6XlBGro8xoodJMzW8FtdYwrmBefYDRoLazRjzAYLDwCPAotV0Zzj5NiSx
/3GQqCKxf54LkJ1B50rp/1FuI5rxCOAhKtqGred36HIJ/V8qlcatKNl7uPLtQ2KUQUNDqxUuB0l2
hXB6CStM1o39XYR0u3jvCQV2UpVLlurw43cuRE0QfnzAvfadaR8lKnUrS1Jwg4DRrzhVvxDu3zjk
O6kJNRLwSYUTOMpHAFxro4uKE6cJ2uStT/jZsP714sIi1x0JstvtbgWCnehzFLQmjIqBLnQCcxz0
PsfEgy1rfV/6jbYp52khce6LjDW5Hyj9Ae7ElUsDRbiycBTPoD8KZig2cqTrqVXbceYikl0wuP3R
vogJJBWEaEgg816ZbhBKtw2ah5xoUtvrNWtvJ828sNc2CgOfmN8hAakSKDAtGeItmFT8m6+bQEcl
D4H6U4O+C6rj1cbCWtCinwgnf7G1QWZE2mXB61QJnQUU7awqbeXAnkdU6wC/wpMPN6/T1Yq67of/
utM6+MAfYBeuBOCDaTcKJRgpevwLPMl2GZ7IqgtlsPPaZ7wyoVgMRMvY99xZ1wd7GbcS8okSo1Pn
t/+3sEWHYok1INJCkUp/Bfe0ZHnExsF2JiPGXE5mtgoTGcT7NlvU9gyY40tXoa9q5FTNEvOr30ag
JZqxnvyaS5JUdbnd9/EACjmYiidIsEKdfDOJ+FmIomRXfp/Fz3ko8cXErkoVRcYmvN8VgJZTt8qC
RBHunTCmjKEM6H+c8sy+DMzrFM4OjxXEgW1OrS0t0aZGEdH+711MrUzR97mBRqLtt60HzLhtMq5N
WUvbXW+zq8By2epaoyhhhVPAnMehIWDK8pS9fhZoITW/MnnfSNFAl2FavGgmqtxxk7IiE+OVN/NV
Z19uT6qoXm+x3GCoBp0qztOcPCJ2zc0fgvVb9e1AKImVxDAfyuRbO3Y57rBnad9gKu3oI2L+gCWB
/BrTO5T00XppGw2wm88x9QwA5YauMn9vwOmdVZ0lycnUbKElzJBtqpOVJHViFJd8ZvjE1C4xwsJP
bXgbVeB6N1sAHG0aRjGwkvhbl+0uHcDma3FrYJiykoSkPJaPOFbApOPFNim0y7S/zrvaotrBMY74
ObZW1lj338hzNjjXqrVgzZwfK2cOixjHJZwZHdd7cxrGYOhthoxtWWKQsZWCLhIubLDRRE9opzpY
l8xFurpCPJb8I66PiHHZZKbAubO8scCmNYwU5QGTbeIWFBkHPMnvB6BMiD24IFT+gVb5Ddyp6it2
/3KPiSQiQkujAIJxGryRa31By3KERJvvsNg0jz0+F1gunZEHqAShTeITWCC6dPUsclIUFQyYS7ZO
txNwj7es6wfIN9gFXXiCEbw5crT2CxBYJEoOFVIe0CQMc64gg2tlTB6V2tQ2gLzhnfqliLBfXJUr
6O65SXFKzUOfh9xQ06ayURdTKbnTQ8eBbnCIzzTHTtZ1/DRdH8Q2zjtEZXV9CzBFIWWEpkOJ7AjQ
/eD2eSrdF5pSSHIvIP34vWJmb5tOfQrgif/8nLxuMBtG5flUhZ49iby3ByzNMfX2wL72rPHmWrUc
asHw5QY5CAl7+t4fzmXD075uodvHbACbhOiRvxtXetdBj3DBbHSD7fJRyLTpoIjSy4vJmDvIawAk
FrU5Kf04XYd7VMHNopgVj5SHaA1G9yzxGY8T9bRJWlLp6Yahv+oxrPOlGnYwJ47XAYK0SHVpYdMR
3X9xAeezKQcGZy1YuiIlVMBjCHHciNKyowbut8Nk3tiHZKXnBREgNp/VvU7j2jS4Nq/9lgM/1kzK
oeiBdnxRg4HkXR9K/+GzMVQaoAD0Nw90kANbGt3fBwMLdbSutrqQ2t4JqfF9LIlh25MIJUD5YpIe
gdFGx4WmQJzFE0EQ4SgHR0UtulcE+T5U5rjHMAnTboRXDdiKRyxt3RSIc2QjO7+FRPlDwV4OGlP+
woHlmLSBZL2lPaZ76ogylERDChd7Z7oKngaJOgQoulJ3MjBcAwH1YYdX5XJWGDBV9vU7/2eYggaB
MQwbvp7ASvK0jjncc8s2zn0GcBWUwdBoW6gb1xQl+2OAYOW1wI6kD2cOsVvsH1tMNST2Xis/uTW7
8aWdg+nnF9e5ttR1frB27BJdTs/5uhZqM/cjRUQYQ29hP6UkJBcINJXlgL7AYoRl/lXeAh7KKge8
eqO1yrwydheZiW9XjWfBsNSYDkORNc3MZiY83kkz50kYbjjCs8teosEAVXWYvLag9/YsW7+yn/oS
pbl4lQvID9bK/4+n1NgNAWAqS4HnQktHBPXMlX9EFSuVEfY1lIkLOPy+kid7LObeQfIlP1OspgDb
dbwb/fmqF07IZeuUb2KWgbjJF5Z4dY9erH+DK3FgXWtXBE0c2NDlmkdt8DpAHBMbXRuMwo75docR
csxEoHvyzB4xWOWlWnLbP2fknLo5yb1VbfM04l73JoN6DaWRmWSDBTe9puRInr2ipF+T8XcpY4PU
g9yaHEb1BT9LA5k8cSIG9sBe9SOLxDTHEjGc/Ol9RAH4eZcJpSKPS7dZrg5wMkV7Pey9/hOoVGV1
F5ID7zH62Lf3nw/yOVb4xdk5L+J1ttV6OWqhUSWHHc7gy7g5A//bw9o+9gUWVfdilheYCdhkZowM
333wmhb+xpjkdcRiRwBuKAitBojd5NkUgvlMkN/6Rs1jcm07Emw4xZE32SyOAK3iZ/drcvHWg/az
MqNSgFFesMWIfL3+1PN5zJRyVdTeJQYp1Qh7aXCNapGrfuD1Zu0BmWp/I2ERKhh+ajGWcguFg/sS
gbn3Pc6nuEsRgjqT8XvD7NZh3fx+ZEK7tHheM1yOAMJFuMzbXOS6P/ldn0/VhtcrKeHbQpUVm4fM
dfhFlimvj1yJ0hwbs7QPSvDmu0GFs7E+4HLw3M3OsqaSmSIVJPUiD+wVuhZKaIgmJBNJiSRmnBA0
dvUP4TH+HMCfkjQ9vFUZB7iXi9aYmq9xg7i4+fZoLjYsmMGQazsY9ByH3X5PYf1e0tYVfl1HSiEX
T/qjP9loMC1GEzRIFRTNdUhUnIRNdGf0kNwcUdCJxPeeV3XHUrMbIvnlh/6Rx7p6yrMD6cBvLbMQ
fGizwSnd2oTv2KG3BYES03NvG3k+oW/whsD7bBqt5oFCPbXnfH47Aqdgjr79qEVhrfe0QZT0c8Sr
/LmWgTrgABs1tI3i3D65Unr4mP5l6WzQGU4sXa1hUTd1PxhVYCr80WxLcs006YLYx9D8F4NFVyhN
TW00n15rj4CwqPaSycMBy9fO3UBjoCWFr3xEwLAmhgBB5S78puQC+gA/ZYpuSQCyrOxqyvphqWKH
IRFf1cFvVUUt8rysLJTPT8HfKwhEDFj4UsMsopPMay3wqE9/RigdtepwCX7xrwQhC79YIWWelB35
n3k90fsAy8jBOZpmk9dbn0PhZJdOZcZ4QN7t5mFvfxgbEzrhgF0BlsODYAXV+/8muCMJa8dkaPY6
ZP8yFG0GiMMARKcq/X+sX2x0qKw6kCK87sArfZWFUc1wJonjpOV0fF3rlAnSUVBeft+AwiybwUqL
osNna6A8LR8BhmsiJ1BQs/lEbeEwPJEbTOshqmtbOT7tPIjIZD7Y2UeQJgdiastYgyN3qUQhpzTd
FU2ij702hoCAaagMtUgVyKSYUpQ4eMiE55xgbDUsin05TgHghyeXtkg504BFTMAeEgrfD4CmAo3b
drZse78tk+pPug7MvCCogYYWzKG6uxC/ipw44o6fX6JdiLzUnFQiKujhrvZNO1fw2vvynXiG0vCO
Pc7FWlvC2gzzRwKd4BqooTiiWKLrchU/pHbzMxV12ty+Mx0GTYiAn8oATT+9sPv+28JpACZEacRH
7fyvb0a2gLkdK02lLzgelQ4Qg9sVvvmqBvDmJ3YDGIJL58fGmOj44mMXBcMPZfINvgAj3zo1qGC1
w97b1aq4H3VBjkpIzzCGdJxlkYG/Vx0B66ITHZKbcR59xH2dagF0aVxzSoMKzLzxd3j6XfdYNZq/
Jw4Nmoju+DGmqYXB629pm9nrJ1UgRUgQeP0dwKADGVYh7lKA8gAxCgvYDC/hB8ErwApJBPHa46iB
7tQZcFP2Wr4SPC1t0YZNHZnKqANtjYOHszMn+Nk7YO52vwmFCvpXfgw25kflRq7NpGY46tcrkeu5
cqqo36a0xhzMo5ipUXELE02W/qLvZH01xVxrbKoJwLJK9TDxDYFSsLAU6TMXV2d82WsI2tCIh1Lv
TManyFlnHZ6zuzxrf0osu9Ki7NXpwruGdFc7j22pGbY9b5Oq7Zc47iSAfoB8rNa/TOi+LYqA/33V
+hliGgcuaobtACw9Duij0OUJXZygwP/MwXwEySZudt9LCAOcRfHzaOe36nO6m/XQlCMcVwdhTXEm
4HzYmml9rDYW3o5kYgsEnxoooKhhBW41ZGkBf2p447SVXRdFIKMf0SM7eyvo+voMfgtElm0TBz3m
BhNuBrb1h9R54eyhc9iA7sZz6zpi+OnxhncxoWUamSApVkScMxHP4zYoktt8sRcfKSf0Gytc4Rhi
OYz2Nbf+o71Cyufg5VcUX5dBk8o2ajEq1AtoDbFPJVAWJ1edwGDUvWQbelTfy41Nvn7odkN6gPfh
69ZAem/Fb5oWv7WTSGPM5Nt7sbyPeb/0DMnaZ88Pw4XXWdq/DC19o8WfKV8ucNB+VRMtl0JEXNBE
x/8fnl8643LwrKbvKvPdafwCqE7qCocsnwgT8HS9cEshHt5MqCeaTXK5RZgpoiBDkf2j2Pv+JjkO
U/42+WTyuHU0ZWqxozBdoJGJRr5ADWupxobuT3pKoLEVN6Y/qxvA9mefOvw1x9PVeLeykJkKSDx/
wX/e0qnHj9a1StTOY/yzNVJZEw7Mgx9PIYk/5LSIUtB1bwKZgM1Vu0+jI7C82ekS3fCj2CoO05Wo
tPe3FLxpu15CxSya0NQEgYbFSv0Q8HDjhT9cNxqtgXqMmcaqZfS1xyA8lJO/TRqNFsntq0S+B9X1
6kVs3nL55+5Sb45frbH5guZ90kM52m3W4PedW1r+CxHnblxHLY/Q23LUqCFl/10/f00uHOCh3oVS
oMlgw8zPPOAfuYflOkcJtTW8r/A5IjYJaEhVMdMQTCjVN7f5gGMdtaizv6RiEEm9GMUMeRcEaqDe
ETQ8VqB01Cy5mYUFcAdEsn5K54hzm36TYydiPSwHKMUPiLo6Po3le2REkLC4/zfuJECSBHw9fi3Q
gmLrjCt03PWh7Hog6tjPbPCe3Trqe6aNfdiPAus538zhPasaqsiOQzgnVx8hS2oG27y2G5yr/WOv
+RqCeQvCkGGBaz2ibs+PQYmAnBEXNK+WwNtRyv/92Kq6nCbQfVNjvKvBDctfWV7j5wzC8fhobXaK
U2E5DiPSfFM/I5BB3j1WPSgIn7Uguuy5mU81fO9uxcoovsAh6kFE+E6BAGgDuvW5Q/+XOsVHx/vi
aJ8jfnoWF7Ng7nsamVXALKZmM0GkJLjp3enkpYfPvuv1nePxYs7VOUe/0V1ymhSlW5rkLKeMc9e4
DKdjHW+UOg44gqNM3tkmvdya7Da4VvcmXfIMGsX/LRi/SyRSwoEhbmCuwEO+DF1tW/z8Ga6eeq24
h1m4EvNS9IlGnYLHrcehhgjL1qAxWsBXAkxh+hKAaNv1NMOKR0lQkpgZAsAsZC5KV9hy1sKWPNye
JW8hN9sfvTONsQER5nMq09ffBRhnXTi2G7pAgm5eef9u5XsSYF6QbD3PJCxSb3FGD7mNGMNz94KK
n4hVs5YgUsI2g1AXLYXm/xoJhaJ2E1+FtkqhpfzFSujaud2EP4MF5So3YokvUOH8mf08dBX1iyPJ
1LQzmEMq3KL1izf8TI0CSfKT3YMiVEWX/Iw3ULn75fLCLUltn9yx7aVcyim5egzFT5rpqnM3hPvu
ay4VlL62tGVn987SPs15o38EIBEmRyffyQp1zvZpE5tCFyOy8eljSYNOgKKMTZPuoQaVwUCDLUv6
+gu63W9VYX1BeIJhaugEny4Ge7rZ1wsUBd4bKJT3YbsTsNRxnVeMcJgDnAeGxCH6lSny4TOx/Ds1
cQl85s5QQMLFDVsgjSaeZ+MQcwL7qunOpUtslObr4vgOLCzK4CNKYJaE52sKwyQuOZL/gIizr8s5
nL/qN3YRdDa5vdmgUU8MMYokaAg9kJ1bvEJeWBWnrPAORX1YrDrJnkE8l1zDU1NKPIozmFNVVVAr
kJRIJ2mZVCaj4YVC+NgGUtqoF2e9OAEoVVnlXUbRlLxMhoP18bIrbXVFYpXJfegG5qbokDVa25Pq
HN95StXbbGXiFVX9ZShijDDgHmtY1elnVPAzaswIIfWyS5SSdMa/sAAC3YTVqcxAgwfnmX27fZBQ
01CzVhqN6AJV2omimtbQv6UHK2dwyIDzFJMRn8f+uTGx0CMWc+PoaZCiWykg/YzyCHZlSZtm11I/
s79UJgoNOjsAyNIPx9jrzCEF+kmZ+HrwGzXV1k37y3HLda5e+MX2XXmE4Zv/UOeUTgXC3oGkZudy
k2qEQCBCxH+HADYVM/8G48yvaWiCr+bJlkeda3049uJXtnSm1v3OWeDJs/ILpw8ZLo3/LQjHTsCB
27VizZa6IvqydIOxCUm/465DNXNejUqT4qR8BnHnS/uwF5YZpO8kq+HDfpx7V/4BRjPw/hh4QgCH
bIyKE6ZhPbCOXHG7XOd7sYXoicuAb2JkFdeP1WSmOHkO0xnXdS6GEYtRoZnueZnl6voxuxMkqH+y
J09xIm5V9I0ByHeVuSLak4pNtckLTIR1ya4jx3EfX6ZtJpKLUoM9txsGvrhFbqq/i3qb/jrkcHyz
3C0fyn9JqTDu8KNYROIwKmX4pKtiVkypiqpyXTtyqmMVBm18XhABV+FKtfxzpkOJOtgzmG0aOJI7
lnESSXgMElt5CDevru0yT2xat7f+d6K/k2tWehhbTRaoB8hV0zHKE7D/I64JDWoSZxQ1kbuxZG/3
BDtjdn0mtjnyarriFZZIpxrbuYT2llL4/rCwU0olj+78wWBWrkroeG4mDAuX5B+g+2y1V5aIckdo
LljJELFDIV0c2LaXqRIwDhgol9PyOK/I7ZZmpcjtWHWCaCllRQuNwAPEiQN91UHus+Ki4heTwC6i
dud785/AOMxUlQQ88lSGHLptOmMj9bnzloo5ssUjFDnINvFKN14Zhw9F1F6rs5zAy3tRgG2flV/h
0+nGDLOzSvN4njGxn4I6wONXNNcJmuK8ShSTmAPVmFlXyEwjnsODVNL+by8A9v+aSwehgAhO19o6
VADfGkpK35pOO7uG5griHanBBN26OLqE4A1gEQypSxP2fIei9Gp+XRXEJudhZ9Cku3BuLTHSJCMy
5GNXwweAlKx1qLdZCHIRGlGRaWka8tqnjGw5s8Ll8628+LtSJqiJ1hpP2M6G3ebxJDY5eTwbO6WD
Df1zDOgsnqkLvqVzKHG7EcQ4DXKBsSmf+JzazaVjprQKKj4vezckaOC40z0ibH/Yt4KqbUu6VoU/
7kERmbldjxBrqsbOWcsYlE5EgCteLvA0C3F8qxuhOYR0BVBd/uEIRafDg+NRN6axBdQxanfHRw5J
jnOWbg2YZPRLaavQY7rflfb4IMCsGz9+7XhTv4YJjOH2J2+F9Xiwwq4XZMRjAbvh1dkiWK2MmB36
zMl8bilyPWuMU1LD949vpLrun1KV7h/DpuMPMlwP2dw5fWap00l9LCtwHx3g3L1qAWkNGfuGUr7t
ld6MQAsBf7eh1xbXLqRAokBMLNprIFfMPv6gZD4sHtX+2N1e3L15rfd12bbOLaLrOjJ4BAOEbVOR
nzXlBZHDXHJgeD7oPJkAkOiF6p10NoyhG2Tdz79v5k0XRsFcj6oGdd15oDUq5A8p87ej/qNE4GrF
aBN+TrLR9beVoRGgeX0htrqKyjCbvxrLFFCc2qTKaeWjsnUh1DyRK9vUf/TDp9u5zn1Q98Ey86Dj
4Cku7SLMLMdI0eOD71WPlguGMuueT5NNjtLizL1yeGzaUN/n0tD5H2ZfFk6iNiJJZw54sURR4evU
5uczH1cOzxEC6vXSuV7emexolHWfuz8nKW023j10mVxT8s3F9loypbWNUxxao+rm6mLlfKRU+mTm
6PyL5aoRhFVWwbJUWI9l6KbPI56jlcw9ghIFDbjgGFROYtTkzaBTCJgQMDMbC6GpYGp2AIfZObIn
cyEIDi6V5mWmPRlqs/l9g/hPR2svIgdTTv+R3iDncXCdvntqrLaPxytMUYM6HXPxY5wzcAnt+cE2
o8seEHOHyzYOppXGPSCy/LueluL9wM/p6rnYnRt/fBztsi9Bn5yhLmRx8Wpp6OMHrdoJjzZgyeRq
6OhAErFRUNNcGt3cwncbFSxtmN6zHeF0tvxP+RYAXBZbr8KHpo84PWBVDf65lEM+48Iz+SnbOku5
kbHQ4t5xNUksvBb4I1jmi31LrFwXSXCA0ZaaBe+pJtvdqbShtt4cynvX6uBB5aniN6ojZafWivS1
50vD/Ymk9+QQHxCMppzSBuSEQAvIVo5t36TNK8VkYzAeBu08zqqEqkb+9EdMRBl0QUEaViUQwVXD
X3yiBgFT7q/rN+9fInEuvNdOEzOmY2D4TxydBI8LoPJlFEQgNR8L2UTBi+kUENIvXF/7hxr9McGh
8owygGHCrPVKMkQVgmH3mPpHfNfYND1dFFJLEnzOXc106AyXLC5q+FkpGjspfQuInoyQTS35yDlr
uXZaMTo9FECU9Kdx25kaBNNf/KZTAm5lJjxEusfvukWcen10ttAENrfygL8Qk/aG5ISehNVPKY6X
wTfKBksvwGeFQCWjGKWj7ojU7gQdzOdkNWltNSdZOH2VXa+21fS7oZwUPw0pr+2oMH/SPvHNDrdB
brvjREA+MWCT+tzwgRKfTMu4w0Le4P8jB6F+jCPfZTiQNJZOJuHnUix3M7z4cTSj0eGEGveter+A
3t2hUQvaqto3XGD0D9WpX5M0Lp7fcNCr8a/FkGEXNL36CNBfYx/i/n8v7WCCJ03+CigzgodduYjn
QS1lnGVKRL9oBA3+ZE+D/s0pQKShLBzkv/wX/CSIzl2bxgMiFbd062lzeT6NroiwRv8t6h6Gst9S
UdLY4XaD4ZZApRzT1wkNsQlXNIQ6pkWqInZ23FNaU5zHLYXvLMg/Fdbm+zE8MKeRsLsd95fsMoSv
sAUubQEz8lHEKCJcIVsz2jmt+Db6A+kVow/cslXWkvuZ6/KiQcmEPmHNv3qGKvxGw5HFQe7G6Cnl
9q1Q7dcQryLeOW8ouK8lZF91D72/RM46IpqWn6WYQMltcqwFVwJ0ETok6Lc5g2zlI1x1w4KDTA0c
T1tRSkM9ouM03SC2ueKCP3JYAd7WJnyYLD2U+h3S+/LkVeKHzPlo8wyqtey1PmP+8z8zPqbfMySv
ntg2JIZMs7qx+heAURnVRD7iPRNNm4VGWw3j78JekIlHoI3qjya69QCCU8mt2o+As2WRsBgi0hob
JTZfPTK5Gmo+AGvm2MHVdClp8f+g5vvPNRcNzocA9ov968kkAVLLdY1TpB/AZb8fzlRCaYaSGlqg
va474PYAcSUhw5h/OUA1ZqUPBOSkFEjenpDYsaFJAMMdk30jHpucrRVEyEbCJUTXaSMmOcWIxuPY
KlMobxjnmAiSk2cXSii+2iTI6h5mu1BW8AX2WA56X30jT3NUhVVhLVKNb4KSfsdHRI6YfBQvZD3+
xr8kPRKsdMsmqNQDCm1aBFGAu96t6c2c8MAwoOQKFeilbcOlUU9h2w25BJ+fGwu91uKw/isaQDNO
GOLw7/+vhcHPxR0sFw2JXv88XnaRJv6xYEoRg8GBjTAREC0RJHlS0ExUrRUpecInE2oPgweiqeNl
S17b2RNN2+mjAjSE4UY19blyk0P3BIJIjYIMgCmWUX88cam+N/VweELyrYfiekNl4cAa4e9tbKix
sdH/BhcON6PYwiavCnFCWMN9adPbmL+BZm40fiwvZ5aaZVA+qlOPgYbTQMswNV6X83tsjVOR5hjL
JEh98A3If1nCv4BNtIdfGLa8ZF75jvQdm2KsVMx4Mrjkt61Z9RTn3Dbhhgjtm++elrOAq/DZONHz
K2SMF9WqyOBPdTeOGsPqwlx+m8xKj0yDpYrHeTFSDbaHgIWgkL8nhuvFKFrxYUwIZlkqrD1/aKS/
NMQbXeMSY0IODErpWFRLOoRXdaA35BupHgi+6/3dtBNqzBiXDuCaeYHirFVKqKRy9l/GESV/pcHe
YWoCwAVbkSLFsBpx//c6X52hv4WfcYCw+YWej7eMSABb8JaEhydDh0Dm26nRZkb9Z3rNg+566nv1
tzu2Jsl7UsPXwEfUoXaRDk+3nAH/Oo2rF/oNY9dr7171Hfxv6mYZl8t4ykbmpkDyhNxLn2YW9tpR
vxezAmvWndYPjI3JghmICR/djbPTC0iOFgD7HvYTu9xo8g1rZY+tD0h4vXYf8r5mRgva5RLr0N3V
r3TJCXZUv2H5Opcwhhv2Fy6ogbZeBXG+AdqoyI2UrWHpyj6CCR5UdBRzQzmimo8+QjMNzhZy5qEv
W8iyg4a3pjplp0lSklmcKDN7wRdDzaRiN4iM5rWAKStKxAr8WhdoW5y2W497TwaZxT+mj5rG6Lm4
bu3dpkgfwDGt2m8zq8ZAf6agsGPn7LPIhXXkxhM5ZKOsiA2BXYFD9bhoqzo056eh1F/XLEVErE1U
pscZIGmESuQdsBxPeqtnTy9nVtR5xPtrnIVXg10jqFAy7sDukEZcTtB+TUS+6uqO8j75tk8+yL73
2ThmAmPNrek+alR97oWfpA6W2ak0090fu3IPfNpRZEcXq3gafoipScqPVvh721Dl0r3Mh4im0wBx
xv5b44niIa7DilQHHV7uYBAF3pnt5oKBv2YMrIjA5aU0RThPUA41crK65udKeQlsiTLGKQn3v4QU
yQDTh3sl1+BYhNPPJhidVHpFkUXEA5Sas89px6EIFOXtil6Ryfj8EPY7gCA3DcsTomdVrK8cICCb
Dn3PQAIwKm1UVfKemrTIIBv4YD4/76szfnZcesQfNV+ro3jtOZOI6EF35BREcxQOV1ZeHO8WWHpP
PjP1N6A2C49PZ2dn0NUtiJSbfm9w1xHmqj1VnBsdtAC2zyU20IWgWcgfMWheR3A0quTpl3a6aaIv
dpUOP4Ik2RbVT/zGVEDgHXmbsItFGmFjtXkkGQJYnlVDbGzEmXSdPqND05sMdY076V+JOt+vI1mF
azGKAnUewK9DNzz+AugDYDJVJ4Jyvq81tIZPG0PypU/VPSksIR3mEZB2XI9vmTehHhbBzgslPRin
sZheM/4zzPCgcDpiE16ON9N9b8SJmLUxjVT22AF3UGb8D88oHbop94ToUJ5pwwZajFhPYNWoOOzD
6X8zg3oh8klRMuv2bXIlN4Oi4tbOOibOCzOnVeXqV5DNCn6QTPkBSjHRtMieeClN8RMgy7MVeWH1
0CcxpSpJXlih8KGA1kqAUiFo9/LFeI2iM298z7XiUwwadLXK4Nj6YurkY/L4eW7n+4mBRPf96VF2
dY0TxIvsGPBZbaRJsSLZzEqNAFjM/a1gcXomWsbVh8k7Bwts7LNRbGz1VE76zjEZJ0RrWflt6h2w
RRswzT5DT00pCMnyc77i7n2gtudUU3tNPbS1szZA0Vklqv66rwezmEHtLeK8mwqJ4rvRxwzGWygP
4iekHp9sDp0YD/AQ3lEH2g37lkzmlwvgNz8VbAGs6y64MJp70tP+vGS6RC0oBJj1uIno4EIygd5t
0ltDtVnzhJKgIULcNAdlOdXUYlW50ZU4SnEs62Dl54IGZxgHR/AmZwHk6G3CsHJ3y4OfVVBt6YsP
dOz/sJnyByVzgJ141XOpfoMX5gwoSDRBQBzCD+BwjacpcxHHmC4zwQOu7ozs+4Y3Pwq3FpvNzPMi
XfVFmIWRrFlc+1IjcxiJQHhvbQ1JUhqMYPaFiG+2ZjmSfETH//KOly4xHwwD04F5quctaxLt0pm7
GdJrU9nD+wlYi5UyZcbLOpcjnGUwVE4VsfxEbp3HDVOZLX17pvQKIGZj9Rgw0Pr+9ccehE3kJ+YQ
WDJNUP+uwZ1oVLXvcY0kTuCP0ZLWlj0KuFCe5eUreW9SKAfWI8nV6AkTqqgMfx7p06jWydImHYL/
0dqOBiO4VVmiyjCXWT7I8cqOZ5auG//9Zd+agcVVm1WnkbP5ZYGRDkOzr/pqS6HEZFUtg0+r9D1f
ofy/FNYrtgo99/hlsa4Zjh7QIzSwXUYQPBMDOxUQ08pSuVbAT6cIG8jKluYv4yr/utJWK2oaUnPU
z0gIym4AZxYLOP9nAQr65oNdMW6ivB/90AGIMyAR1YX9Vkz4C29PDPGPeu2JIiz/1N5ZcG00F/10
IvTNYgeAnFbjjeZ0wzm7xYVr16ND4VUBzM3sLslDM7sAEAamaEQQfPQTeWhlfBzMc3BBnzR13b3j
tvVdY1lBu6qDAi90fY0VSGC125ibbNerup5MTXPdxC04pKL+hnZkimt1t6+dIzNUX6V9y/aQWQ/v
YHw12g8RbpvCKNJjtDumIl4HIiRMpVxQ0LUcEvb9DuZhA61xgnMuwMO8/pQWGxNHn5wrLoFn6CL/
BZQYISXbFoVpHxPNeqXHtxEIxKRZwoZwCc9CfdZQJcogIpapSerd4Krh62EbFModYROY+WnN/Xn4
G015ZSobNOG19Bcx8p1BsZtwewSPjAYdNFw++sZ4RVXYYcBVSeU7pxcvKFO6pKZBICFVJZBqQd9F
5ckwl+Xbb7w6bM8jhT1r0VuWZwaN7zGcPJyA7ag0hBIVCyq/oh07nDaL6AWD/BQ8ODzJByQAMXN2
4hLnF4RV4zwfKNE2JfURKGJLHhtw4RvQnTKCkbLj2TULvFeVr4Pq4HG3VEN1Unhq+LAM2OUGgTO7
M+qeETmIko9pH+mo5rmNS88U8ak+AcxlKPJIem12JVjo8XPgnJg6p+2LMmkA/aub8y15Dnwg5TXi
3dELKRitz6QoaQZL0Mb2icLGu2pUearjs5QoZ0AIXjS4cm9NqYtJtljJv891aGVV1H5uquVO1UCa
/HzPUKYJzO1E8wdJsaYzDAd4EphxyAHc2XMeX6VPy45Asgob+2tpSC9x8WMnLG8jh2a6q6La3eEk
BW4sJyee76n5RNYph4ZddrmWuMUd/DW3G2CRLd60YZ0skfJEqBDb3hwR9s2S6UHGTFj9n/UFFWY8
duFav6j35TCSA0/TB+T4Lj0q1dBiiQuTpq3SWMPHKVdPzZidomTlqf3iIM01QWVAt8SuuoZO2NHg
cKA5o24qhghWgTwvDJRoInLUZNoMKx7zcRCZ5JW+x9rVHgU6u1CwAbQB780FxLRCR1C0FqlAtS9w
7xWYNN6/c9a5m8YLpTStTU4wAToafa+biiXg4ua5gESZxmHXFBFk+oRYmynyzmqAEEHH8EgDfZWo
doocPpMnskAfosnh3KV3frieS83ZOkjFXErMRzyObJkou1HJRQf73IRVm/Nn7YSdDXFTxmbppGa8
EDq9f6x+SroGRkfpnRZJ1tvmlLl5+W1bCFRE+MO09j3Q5z6lc9INACgdzNIMFZgmUTcY/h0jGHZz
fJJT1zy/+3Dmk/qlOiivKz6updephsx4ZQfF8MJXsx09NQKZRL4h7Zgqq2hwcjOWuJ3yIA8tZ5Q8
w+yt155Gh/WaLLmNAhCk1Kn4Mq6dqlSpGM26PYq24jzfCr0mo3DX+zxDZaBKGrnHDQsUpL2/GFCa
O0deavlDVeox2j9/CWReOEbz9tVDuGAzPlvHfj8UUnfmaV7YbpMbF7hufkEICwnOGCeux/oFpwT+
VaLXzrE3YrPT289u75yfeb4uqbjLbUEA+qL4yJWE3S5PVEIR/H0JuXhiaEW5aKDzW9aSla7n0gJu
97g1fuEli27CoPsGRkRUJY2/EwH37w4DqpZDdzXFT3P0TYa7fjPiQjsyWkBz+HPIqhwmv1Hr4x7a
CVFB2nDJdOPNVRupkwrZtGYOV6B9QyZPJmPKC4qQ2rcdosHmQjDP82RQaF4uf/lXGikTHgUJ0LO1
mT3x93443scIqLJFOzEoubhhUBATymobMt2EQw3mmHtYGfc/wAsOpO17TbyaenSJfOEIfF2t5ozh
UXyRQwVICyAbihLQPuhAbn3ykwEVmrC9eErzZZTk6FSuGPuDCOZk8XjvSxBGwRYpY8lyRF+E8ofV
IPy+sabVCVXdI4ptvO8oSVaCpmJ9+9ytVinb7hPLanOmHCiD3M+nJ7h+P2oZo75aKDbwwSWzp3pS
HPjz4X0/oPwZr8ufLW5xtYUJkZPhmWIMJ/PIoYngtxTMZ728TSGejxApPZ6cVF/XR2qhbd6bFtuT
wFoSLF8Ik9ZLos/oJ1ILY31/JrTL7vWGKhbFMORQUuE7do+NF0iaOFtyozZ1NQlbTdksaHarQwIf
ORcKVNrX8HmPdiwr0aL+vuGLSmJDlTA9hhDTwrrJbhQPvi7Ya/FIZNdfst9qcaUMO1UxhHqi/G0V
J9fdPeAYHcPpResNvdIkM90lOhPO8EuwwMyGM4kF48GZr+SGJsEaGX/PideLGcXIj5/c/8BO9Ee5
GuZDDJAIYzm2wkEcXbflAchKmBmgYjZtAkclnZJzbdJ2BBrFGeUNM0pKczX60z9yoMUhNs7PRKqD
hjq3tOVLdyxz7xPExAqje2Gp18b1sGo2Ov8lFmelN8+sqJDOLEfSimuIB5XKJBUfov84fPwVWNRi
rkszgvMaA6bGdhi4ClTHWrmli7loSY4CkfH5cV2+VwDBEWgZGe4jDe9R7Y2RAbyXiuSWsTsmRZa8
tB0QhF2Rako2+77GPuPHot0MPywPNVo2pQm4Q8lvW0yKXaYN+0Y9XSDNxVl5cKq01LctokZIxQUC
0lJo76nNdgqPO7NtMRb9fLFSl4QtOy+azLrMzcBqGkR4QB+uYK5kE+LsM1/lMdgIIlEGoowunVoM
aMf0pkq/E378FN/zo2c4rVZ55yFyUN3CfnA6LK58RErbbfOH7G7Cba3hm0bMc6NJaWfcxGt+bRON
D7aJcIdUgm2rbjl+YYXvT3O6E8Zou+C6FWNcpNuNCt5UnXXpjBCzKcHA6hW74a8r5TcZGmSvaV4D
zHGxssbFARWCd0xMoWFdQdnn2+4zw33P4uT0a7H5igKGGNHE6J8CPnKtZu3YMootC86rxr4WBkc1
jUMpYpFdHOF0I4Z5Hfcjfpxyod3LJKzvHPXTUVRqx4mfpkqjnWDRf/s4+u5StotF6FQSquGlrVul
P2VbkWwkbntcDvt8XhYCEK+btG6aidexvqKKYSGvGonP2xA3poqRgcdkkCiR/kka2d5GdmbWAGbk
+Bthmvz0yKukZ3/y7nlSkIUjK9mmCkg794lTx3xmXXyz2nmO096hnOCBYAdYWt5sIYCv76oEpL52
5yXWnIPIo/sIDVj+zzJgI7SiRrnvK+74j0ML/XHJrsdxAIEIYgjcRc7dtOORtnqHtuGI1gvh9U2G
xscELmW/oA+QbVTPudZilIm8X3BM7Xs+wio2OxoP0qwPmOv/JsmNczUS1+/JX1Y5U+qGVAhZhWKP
rPybMtpjhDhJ+QbzoaarbIHNXbHDUl7ggiZkeM5G4nmrhnxsqNlo3sLzuR08IcZop/FWWfnUCNKY
aYAY1dyiOGzJhJCcx1xYU7WlDqx8fWRSD2R29up097t/yBWW5kdFZMFvvpOS/qQEJXAqx1jn+DUx
IcLrhll8H7uK6LT70s5cUHwbDgjDsdhBgMisXI5nrhW0gKeqj51OMKm7XsMClhDAaUqPQ6OV5/l6
XpgsmHYMAqpDjGiB8oeXAvjkEZX5Zyca5NLPOKhhPoIdEkGI8IpkkjXCXPwJSoX+XqDMf2VPw2TG
nkSivawqXO6gnAkjqp+YUOiaIwm23saPKSItmVdsFa+InaO9K8zBwB2CmQqYpqjNIItO9VqhxUfY
V/9EwcKl7Srawlr7M/x0hXn4IqAUHE9soUzp4YXbN5HSeyF73NpO3zAiRsBv0rqhKgpr/z+F9fRg
q6gYBp3duf7MUL2j4xGCEN21E6gRKSIM4qKRcQp3/HBB7pI1H9iaJTRxj8P1ZX5p5LI8f1EmUjUc
7iFAq8NB7HkD6VVEKWswHqj39DNTfxOPjvR1IB61Nz/KrZ/frOS/f/vi+5UkDwxuccPYkuOKqlHM
flZkuhUvAG4r/FNnW3jxh85bphZic8TmN758BLuduzjRLC2W0E2ZxSKAi7nbvrnE+PjmRKz8E9xd
PpRHAPdTW9bAf/Nq3A91xnmxiWTy1ZD383B/kwkTY8mVDr5D95CJvFL/sUhqwZj2s3mu+yfIe0/R
qHc4za0eoYutJGzKF26tx8ahN+aRo/9zTUHkz6DQtcQFct5TIOSkooNVMgurWPp29UymaZ3HMab1
EvwK2g4mt2f7HM+245VdTIxQkBZneHcW5VTjRm7QVghbQ4ZBY3amuEvr5UrbHFSfg+FqC+W8y/um
T2uEXzt1o39+CSRSvTmqW74YzQZd/5tVYMWOCT26+z6tAaRQzXTKgVC08K03fUYoxkPAaLtf5jHx
6DffoQROcYr1JzE1WOBQb5hPlem3Ezi3gWIS1Y7vOrU697pc1M7FfOIAxMLyC1zsJRmNicR84LpK
9aZkQ1OfIwnzHjZKvXDXKDPQOK3+oMYqzaa4FLiJnZpzTlb89JqvEwI3o164g+QttAJSyI+vCPNQ
kdieJ1S067xIiMREEN/UN/nK8rHIgVXB+ujSfaqTNDZ/4e7v5wRHySGiH+CvKlFDBLKLoVLifrY6
VRhukqfj8Q7Ugi+i3eqOdTkOfkKu1xUZsk3FEvtBMDmxht6YJXjndaFPDBzj5RcnYjHufcNbYPDK
Jn0j+pSJrlIyEKbWfgkw9PElQav8/WjfH0/I5Cpx0kOvg7Hybr1T68eZA0E0RPWaPrL6yrV8kmaf
ftbwsPjIgh0MjgA8ZGKcPwiqtv3iez9N/D+MCQuZaVcW6XNVjDHUArrJYXnZbg2Dg+LoIFbCsOlU
Q94AX4WjztrfUfSQXEcqd/US/CkbnDJLbeWz7wm7GYlJWV0DjCF7J8mvbqfnE/9fWmhYeUVMH53z
3hzHgQE0f430xAn9tyqLWr1Y3hK5T5QgTFgOit4Ladxx0j2Q0W6lONRHKaqbIdR8SR+mbsbRnLEQ
G/eCUaDjTZNe8ZE9iDmMB3Vcii+9cKv5CK58bd6erfr4RLaWLLAvpqbmHgCDpWb4+bsowowQ0zPS
Wfm/CTay8ckqMWgZzKnnS8mONCpoQd0JUSPOyJWrZ/542dU17tNd45aHSPqcoTjPhNYq5LU2gLmC
k41pU5TikJieycONqjJ7oXaWwqNmcyLbOVgbDHfLL4KH+Vogtyc/5R6td1YX5HR+4PmK6mVuNSB8
K+sejffXuEAzU0pTWEqjaLaQAqlAaFNWrZal5TDvY8NjRBnZlYUG0q4ozYWg0/LTBlnyezh7s26Q
81Yx/fSsTLNcKFZO0sGiDaCn5tK5cUmuJ7ewvvsN6QelnO0KMxKcy8iUuAZ3rHZ548SFsyVCP5nS
pUIuDUUimoAki4Scj7JVWbDO9Uh2mBhIPltUh/5fdfJHF1/6k8NHcPEdFYlBwRFxcThJ+vU34PN0
Ez1iMxuL3eXEz5h/XFdIqIYKvc11OY1gMieeBytAgnUpJrEFDg0afgBbeLZ8uQwJVZ+HPymwjX4B
S2ipVYJWlTXzhqZW3cN20P6bRUkH6+dPZfni09UppotEqzK8XM4RGSeEYatdw3JZ+y3btiIO+hir
mTphHPAry5NEIQUAwlIAoaAQH9u9KqPujyw+pBqaZR6Lm2k7ATCjPAzjgle/upWdOJELqhsKYsqg
N0LWSm3Hps4823bFfTpEBGY8qBeEjhpkDAqg2npwwCIYrClabXqZFTYmxhvKBMfK8CDkOOSc/EFn
BJgLnJauZZuR9qFCkgFzRLEPIICoXPdNsiNyDTz+x8kyRu6+x0fLy7LAwKSxD5GXk7ES3Lijn7Hh
Ixj3mc1g5XusW2zpOoiQKbjeyG7VzlxtTLReJ+ORmHeKE+eUNhM93lv8nk68IZmUVxNFbdeUWu1T
4/Y27nb5gsi5+ozP99U6Pnewp7lH0lF7XeuWzNY7nzQpqvEA68PENTdYW1GJFeRR+eSE1tEa1gDk
WntbslAni/VlnIn+l0JlBNRJHk6M185Jac55AMMZY0BTKHJRIdyc0CUb3l5uqAGPzE2wntwDqOwa
0ztoE4nFKsoXHDBRb3zktUu+/4kAvDHE00BJdUHzT3959WHO82D4/CqO2pHa40aEF1jFNf3YlTXy
oAxCeAGnZeijpJptqcNAiBCpbbQeMnodCGJDIVgbox/MM87bQKJOcpYJZszb52IFAG0NAxNJ60ZI
LVRmYJGmbj+F1Fovi6poNetYU3pLb/3bIH4EtLhYQybiwXKd69QI+j+YJpCvFAaq6B4rBk2SwbuW
OE8nu+ZsQtADbCATsOPdZIaHFFWeXlQ34IgszS6Gm0yNUZg4eM5HvKnyK+8clmSMDFMAbwj5dNBk
b5ArvDT3a0vvyI28nABIXiyeaezP5KXiH3rBK/0hSLJK8+I6gvi0OERJOcsTZ6on8o50Dy38iiCw
B1Oear0zF46nuxvQsq5/L8EP7/kgI794QMB0ELjObDA5Zm1qXQ99zBtf3FeE9GEz2fCDA2AOG2Ui
VxchgO2YcgtxS4m2Z+MsAi2rbDJ5gvMxEq+5AUiDoisSpNoSpRYlBvOAWEIyLhwQElDrG+5qHku3
kqMM67dYMnh5pX3Yji738le8dvOZOm1J/CEpSoGmyfVJxr/77nG9Gv4mJGp9NMODpxfHojpSnUd2
4YMzgF4xE2v5pAqnYo2Oo8FwJ4CWd2N+V9F2itQBoKuNnkpaz0HAiwxh7wBjGjjP6Nwve3XSQLaD
l9uIPqJKLSdKDjqI3XGpoNRuX5SGrkwz8F8ipL8eQDnNNuQz6siSkuOo6Vp4EMlxWJuwNstORvpk
oxXmXNBYFosCoYEJWIqWhlRobCMStL8ijvBnfNB/oA3Lmk46Njr46eek5JvGklh0Eoyd0C1eFIjs
SMBkDYlFaD0TscqCoB0K3LApVQem5S7mqJK8fwwH9MYVW2Nebkg/tt+f0oTvFIcRfeLx0BhOM2eB
GFwtCPzQvCx75zglmcZ6wq1KjJmqKQpem2UJftFbQ284tP1mtvzh2NOcR7Hz23tLzutqZobK3gk9
1EKrFXsldIXSBR1G7ZVwVBY4tGllar64bnMYoLFXzxiQgSZCA3nByR3d1aJKPawEmHptAligXYDl
ajl2cHU6diXZy8BS3GYoaekQbwAz/9WQ59YHGwaiWYtPIufwNh9Dnvdm+79jkYOEoZh6tcfJRjqm
aEqn3EOGoLi/HJv08KeQyhT83FHvXzLC5YamoFbHLmdKRdX0R9kx2YFgxjEVQ08582elY3t2VWd7
74/2N9R5FLtQBptiGatLNEpLm/MXbcoy800wreB4ThV9RdQpjjwVrUXW5y0BZYjXcF2U8v2ldOo7
T60+jWH+wo1UPm1bFgVoTvT7tzKxcDyKytq9Lu5+lQ+FqM51SG+ftEC9iyJTqtHq1frTf96IIrrQ
bB+TR/CqQKaPBqG7/odJytn2XrOscu4geNzGMcg+rjd+YKic8VAXhSlmg1mV6/bvjVC7XPqnDmB+
3GiZCd8XpBffZJwXg4LO9fXxZWkbaZCJ3ceNYtcm3xaQugGOkMU9mfE8Tgyk24eHgdKBL5vAphke
3Q8Y5ixEIOfHPSPNWRI9+zQSigvFChm6wNqBp6ih40mYtqDaE0IhtOyYJKqo3DSJzmQcJmeOB4XS
+5oK0TeH8dQfls938Nqpmn19P3KVhul4wMF9N2wAZcnnvPLcL/MSyKiwhiVeSUXdW5ZRExEIZ5/R
du7FAst7ZxbS2VVjfIoA12m+M/dH465DPT0O+c63mjTBd9oYQefuyNoQdioUSsKDHX8ZUsNB+Y0+
4ZW94rDCH1hBHalrCGy5qRM55RnVZ8jV/2PJtiazgWO78dMm9MpLcUc7wUqObQ6sDG+G601K4Emj
ZVhFf/uuzHv3Tax4bko7A0pmqbzw4s2W4FmRrglTTUbQTv5e+G4XktVEVY3f9kFnhtBdztX+A/oR
z6K69/e7WUgnv3Om2jDG3u+eWCFDA51rr2Qov0FP5TBAonPaIgTQZBp8tXeZkSIUOhLXTlVznsr5
HxA0G7+oBNGfTDTZcVIUn56l6ixep4I0/PS7gbMSUzGp0Aa1JZbFN0EZWQdE4EJhCUrVOVwjXvDt
E8m1doa0dpd2DaCbf7AlZw/NxODvMnIiFS7RCTNVjJvEpPskJmIJFTLsa1HLsLbduT+4+wCBJj33
EHrQSyRVAQoMkpATjMKNvEjhHf8ITPFhvtVM/QsmxNNKf+T/m5GIKjEF/raPPAHhf7Gxl2Az5Axy
ljr+TJehSVFVMDMekWYdK1xALsr5358x5x2JPaHBG3evBkYIz0vPFYrorqbUMaDno624+6eTgtZW
S4GY7T99G0mqv6M1Q+OLV6tItGA051aYuKhcRqVdBR/Qw8y3tstQtImiYqqTMDpl8tkmo5gBl4np
xEmy+soeeaFgwH12mm93YDxChDT69BRpA+7aRM8q/qn0enDSOjr5sEjsWIGBnInSXgStN28xWPWa
LCEIeJDfFuTj3wDzz5PPqkKkQG3hSeQPZhHaP5MyHq6GE9w0qXRejFOz6ka7TEQLgZeEhrFfTwak
AuBdp07XjDIsVF7GpH5pC2dTYoVXheQdEKpCaT6rmGGcFC5fKEsXmp3TSnfGP6ll6TkVX+3hzwYh
bGaaz0mqINROgyVzE5fIRzznGPA5rPezF09QNkoNwB3MjqSXENM4R6xNfLuKXtO32rfiOdf5yyB/
MtfEdL83lmVWhsTC4YB8rYqxKFZsUuqjvjl8Y+VT4iUZfNalTdyzyj/Lwm0O2doc39XKEAiKIv2R
PJ/Jua5YxF2B/SvSQdEJJ0ogHUyP2H3x3fqCKYaV6SRFVbfKBVqHxFYXByxMmXo+jJ9B0brOWHXh
xZmpEAOHQttH1RnMetRslQM/38NKuPNYlSrfBEsBW5bQrzv7MbrYKCndzBy1NKNSKlSKYsgQ+YRF
jYb+MeLyWyF/KqMRb85jHoek6xS4FqGdRmhxyuYBRItmGXz5oFzwS7dm2Vp1oQaepqh9EtypYP3G
LfrTkGfuE2WuJ2W/4/wJQRywLcApebd4Bw+/d0VXISnCEqecCW+/o818VeLZFXg2u2IGh56wPxVS
iwtKqUh2489ANSYPuaf60Tq2FvjASqhBpIZ2WZPJsEJdGjBWUpF+MWokjJPnRpVPJ/wkiVhj5Vts
51iea9rpT8T7dyvNQHEZVWsI8yN5DJKD/xY44w9N93V82v2XO6o5yxbzHSY9d93y234cHVYhmJ53
ABUNS7lcj6MAhlXhjSO8OhDXtVWbFC4hYuBF4Cy4GlTyDz13NmeAT6GIezAcpVTJgDVHjvn6ISRh
gEC4Qef0sCD7fptvojHAcf08v+DoUhdysuZRoNt+knFSq70i+Ge6nh9MYlKwb0BjnLH/OY43vfmc
xWsjdLF3HNJplt2MW2v5KnsW+krkpKGgRBPhr8FtlDI1VSfwsgDdylLciSLNttj+10fN1kKQXLhF
MWB9osMVW3B6O5SN8eSZSUSc5YpzON5Ydgt8soCjKu7ySrEt4iJSqkoKW7pMqP9crNba5OlooReR
AV2QRvnW+z4t9iUKWtjjvmw4YQK/ei3nLXaa62CCUdRTBRRXkelld5mP9S5qlu6bXsTrTyHj5v0W
2MWW7vKvhz7i+HI380xzeikndyTE1R4UOFKbXw90DQ0hxkXDNam8r9kP8Lj5TH/ATWhjQz+wIjqW
WUXoM8sjhJpMnSHIAfJ68ybnSUnaeIG+JdXkoW4ECL3iGpH35KxJGqZB6rnjyJAe/Z1iK+2FQAe8
zGU+8ZiTosIH8n+llTVtnMwOdGLOXbu3ii7aClndcbc1khDMXs+vSTcxopFwUVtp6HP2/BdKj5b0
2FyktIesr47mx+5XNJrs2vpAbTOLzjVIGblq8MHS3VfOd9/vI03uTzvj6l+D4gDiE1jRQ5nH6UDB
ZxBfm0jGStxc9kSrqXIninKKbGnWL107LRgGqHYkH5QGeXXrheYoEQKF9iKOspiB30F9IMif33mC
yMJDLyOAZ/sc93HiGIwNpigG72eFwfCGb4rSvW9zwVrpGOD+u2q2dGW2Ihh9tyLFQRKvJxK41YWJ
0jEOgTutbUxXS7Bicr/ZqnhP6+Ka1FLnhsyBIWe5sttx5kNZqrKtREZmzSumtF5Zle45rzUf2xNE
xS8PygTUGe1umONRhxc5T3qTj2t5gUDjx9j3nb+oEo99qNjqklMBp55eFbcNr7T9TBpqmHkIgp1C
ct46jmTfcsf3pmkBalY0HDsrns53rb9fSf48ggy/RUQKk0kDncI/ZZexzEb5KYe0WKlj8pV5bisx
BFH4BxKTfGiY8JfJgOBcly0eT2Pa2JZGibqspRvKNNUP9bsXGTXn15YhDgTEWWBwCWbvWXnQPfQ5
UmZmsk4qjtOSa4AQdzuJBPS93Q6KJaBwk1Ra+LnVz3BeZ8HNckt4C9sW2IYVM3W7DIpxRTSA3kJx
WSIYMdzbViaudvFx+ZpQ44hCqYtnYnIuKRcR8uWqN8R9Yfb+4NGHa4j8vGnqLVUOQxbC3ftBXswp
ovLtzsccD1aP6F5kW4T9pvegQidBw1zefADJ4Z7CXFjhVjHy84BeFhQSxFy2uyy2BXzzqMg7aF08
F2+54w4k+THTY+ncqPPZsypqA/m2WVgAbImwKWgC1sVkIOJeQxilOT/57Rd0H4QAmWTJlNn5x0o/
hOrRZy8qkBi/BoDmQuGFBFYKzHH694qkQAGe+dt2Ur96o2voNRDNPLWyKb3DN4RIXMR8Svw4Vy0I
IeGA5+PMrZ0bHSdfNONpZVNPZg8V4hcVI64GjCCJBBu1maixGCQCabPZXEruzd6CQnetoC+5XadP
BA58rSAl8Vf80owBDbJxmvyBhavuqRwxT8cGvI+to2JkmdBtCYsQSagND8bNes3FmFNGVroTxB2K
e0s1e0rLIN4ZPl22dpdvbPevW/B2ARPRl+Y1Su4GE79w329CZp86vZloqa2bIiF1tpkm8c2an+La
6FjSHcH3KDaurLn444xpN1hz4/VF1NJHfQsttOAZYsYG+5yf9nV1i7biUxUvPZTOAqy8jT1yzfnP
9ox54CEsL+87Y7a1DhJYCAGQHF3BMAzlrj1Q68s+pLEebXgRiLfyQGI/K/8mk2RJBQcOjafVAgHn
8VA/y0gFPCGCAqL2M53txI+/+QYNyJmy3XNzzlrJRqLdHzOXIz/wj6dxF+xncHsgNps0aLi9YKxM
7fpgfFKBlh3zS21R3cNPnPCY3NnC9rYS3OEvL+laJ/6tM9C5FTB9bdayJnlIeS9AWWF39xMzlJLV
/Q6vLYFfyrUvXZM9u4p/VbKl+HcV+jRKpeipzw88jxxMLkTWsEhr3uVmmKWDkCHsL/uGlficp4sb
hZY230foeywSwcktPZMicDHRux5995Q/qGQNvWis827lij6qOSesa1XoqicXBSRQDtAxiKfGMUPo
RYdCM8h8jzExprs1ruMCRpyVtmwxs1Icv1u22y/Da0mINNjG5y7Iih3FT3SRlKcZLllRcwiC+vuQ
twd9JKUCFIBen+PF4CDUG7l/GwHK3CCWwtY66W12/FdlujbugqBRKauusiQzzOe7PsVVrtutjMmd
omS3JoEHEKgq3PY4CIwUkgvsLS+SJzROAtMcZ4uTV5v6Mjb9D2EzZ0/pj8oKIREHCyLshiY0AX4D
ZiCNSlAAwb6xRLz/+F2e9y+41JzzLkgD20/FLUPe5yLwaovbtJP8oSkZ9lsqOWzuMy3O6qZt7ByS
w5WW85hUqTEM+oFk1m3L1xuuSwTesOIsRInVdgqSHLercVM8nkwIl5aPDBO+eujaH+txJXr6TxIr
Q7EnVxEz79GH1RjXWaD4YVViAOa+CKAmgzyiwcCXw/Q8BSLvoyvgr/oU4RyRWnjJWxJF3tWefJN7
7qyAgTVOBWsz3t/XE8n1HSe4BxxC4gYWGN3aXIIN55ww/S7I0TNDQpxpoej/ob0LYcFr2/qvV9q6
2X3gF56Fai4UlNPt11IMyl09jZdgMgk2VjKY9gksu+NN/xnRs4wuGKS2NNBCXvHy5PiEtf39Fsk+
4Wpit5hJ0Xe9VeNTHUnq0hxeHvzdFypeyekYgBPAEk85xlFVLLa+Zw7lNUjborGMPwtahJcZTIZb
T0EKGTJfmM/ztgJZr/lrECiqUX8PGB3OldOwIBYFUfQ8aR04Qj982f5+YPBgRcbSZT0IawQOAjjU
9s9gTUNfed0DqP07CFeONqG9xB1H98OGjd3kD9aXoO1OX0l2CJmOZS2zB5w7z2fvojLPQ16snOZ0
Tu/ZcxJBI3SjnBvbpn3qhC4m/i2yUvlgWcs9Epu77IHrRFs1GJhKmfyjSKvBEXYaBLRkXgxct1iK
vGFMqEjYHMNEa+nkAh2ToPqF8H5itLmXzlTIvwO2psIAVrm1uTl3dw+JB/mCtE87XU6Ss6tlXZep
roT5T7HO2nIMBxUrZo+9jc9pH2T4egeOzucZMXpBL56mKn7ytYG1iKXM41NCh/M/I6L9QSLtMRNn
8FfWkcwy8K3xLUMP40/lq2dEe8TF8N3KWgC4g+9WZRW03ZxcvlsfNM+i3afD0GQ5p/GkGE6PrqxO
E6RqUNy9qRyTfFbbY9bG+/gJGJm/XJxuiS8M9B/C2LY34CGirIMh0IuzEj/QZARIgMIg1OVp9gmh
Mchhd62YlkIcJGf6x9OxB7Z1FLe5pJndogLDeCnEQWL/15lEjEJKPSMmAs6DM3u8YCBLyn7nr0fp
fNzJ7RGr0qt1tdm2DB4rPFgL/SLwL2UTgqQOliKV2kHew7+AnxVjNfTQR48hvBR1gUmeqOEbVglR
n3M1+MrA8W/pgZ2z/latthXZtX2nUumBL74RCM7JvImVVvryecj4eXqNMVfUlqRSr972pdEXfcXy
+jsy8UAjzat+UdqlBrf60jtNzHQC31O6ix7nRaaYTvC3Cq3QwGkK97aICpPCAlMroyS0fpeNb6ba
/r4MqIxkFgfmSj82ksq2uCvZA9z3BdVcaos2yqm5SJHssvGDLGcXKDg1HIV3dSmx4tn0K7/UK/mJ
l6CcotiJbXjAggPUX7Pjpe+ryANvTlYWwQxP4SAGzxGxSZWUJQXkyGEAPIo59wCBRJu0Iy+vgqmL
6m1gluZAFqXt/GAclP+sk7I6CCD84FANVdp5sgyQrCr3E5upqaT9r9FHIKPfTJXvztmlEIYrgXD9
GMZWeeJ+ji7OfqFkh+ruqIoHKYDGFW5TK0W2QNK3tZ0YwLf0nKhxIvpfe2rDaRK9Zua6+B1KRkmx
y01FhJX+HS7lkx7UQ9pamhBL606Zd95AjJOGi3QbpanJI53wyNMyzNYJM5T4KYhJ1OAP0ZofJLBQ
DK9qQ9XwYaK3xGc6sNrCrLIff6W5k6OsCEL6tcMJxJL3Wyq2lo5p6UisQq/7BKpz5oJa7UtWXapJ
QAzCJDzwXsCP1eN+9zPaelbl+pawKRLXF95BsNwVQMMLCd3qA9z0zM+FvDmnOcCjNsIySya7G3YY
NbpcUlzxpUIiPhlOibZgaNPOid1/W9FWTG2LIjMSWUUdDd3k9H8XmZ9Wz4e/U0SGIuAYY756mrHl
M6wNaDf6bBgGJJsf/8bK+2MVUTBiV7V5ZqeB8BsAUk5HNSSfWY9J+J6YcfukbK8gWOPvXgSSgbRZ
lugmHgpH3Mbor49tUzI2bJPmylKCUqabiSrHlM4oxbbFprDhkeoFNq2+uRLZzbgO70//useDD+jw
8SLZ2ZSckf2pqRqFXhyAjtWsYUF8FyOOJw6Hv75ZrGgiARYo6B0w7ZViHGB0VvZCO3zEmZ2CGl08
l4RUcYYb3QNU1QXO6ulXv9gZYHf9axpDn7W/6QpwEummSKv1j4/wGoupfm/u2uxR3rRlLk9nxLw4
nAUDXv8Fz+zYqmdNTCpCPW5IOr06SL+3smfU6DmSvXRT3mX+FiOiHQXyx7rn4L+Qruedjy4UIOPh
X8LH4OhL6Ds3vhrOc6xchDn45RJRS470uRNuvQTPUXk0HVNPtfW36Z7YQ2preRtK27zDvdGngGQL
A1RIQjWd4cOnhppEHtxjOCC9TOrusdTeh02hvj/dGAGF93OxbwMs6XGiaypZIPZii/EprpuSelCu
JSD+TfdyZxSSauNo3II35uXtBjrCNSNP4QHlMu5PRafRbzsxlD1H8y4yRTEuwPRI9yWpG+iK0kVY
Z7UxxlsfK6JW6w8zL6EvLsCv9THJZ60AGUQl1ndcCuCqjNYdmT5XWnySDd2WSs8K1KNTe1cPyZdS
Kxt+6B9QFK0hufSUdDcpvnoQ2hEAWKA9EKVLtw0gQl0IFfmkD5wvHMjlYZ/QwXoV+J/HoEKQLIcb
yAPWJkTUG78W3UrrAXkJhRLDAXYElWYthwIo56hFhZSz4CAyf0RiOWga/F/CaEzBK7m6dWMk/zJm
UBNU1HC41CwY47+rXj+h9/QWcpBSkbyQdleZE3RINfFv7H7LcK0NG3awqgG1DgcAfznBLeA1pDJ+
lTxzVL0DGpD5qFw332x9zgNo0SYSXBd3jd7Wxi0egmIgyCCebLWz0eJKbe4w7OHR9B8MxKaVswPk
tgBx6spUiWVCD9cl+TVBSIY/3SQTM5tMqoXJ24FVFKYOxqIiiyz6UxGHmNs8sAyPVkbOxoxBMLEB
0S7BmUPL7Q+GC6fxOLkPge6pfmYJPEKmeoVNS5tHdBoWSYi17okcm/lllsjV7virPT4Y2rmdds/P
a8mlxr8k2x2ATtZ42epj/eq0kD0CCG6Hw3qSfGqIr9aVSToIUl7yQCZ0shtRlaL3dZLOjKrM9Vhs
oTrKNSBIxMIbCk5UuLVJrAf16WDVA4Kt9ECPXZ9zLyHiT/2fjjcmnXMbYrvewx/dRtGpYxZ+w3iQ
mojIdXJyqOaB2NfspXmP9i31b2N1GMZGPNY4Ku6ZDPcI7Ha8zl1pBQPNCdb0D/+WANLA1R0PEUgN
slTakQ2/hOMnu8y2sbEgqnhLQ0WN8e/xczaPtzIcf5J1X9ERYDNIAtprbdCkCRf9tqFm9Lng69dJ
HiwO+39QDEsh6bVEuGeRQr7GOt9PvX914dx/XjVumQoL6oUwD9XoDNL69eQYzZtOYi06FAcAuDYh
kPYAYUfw8CbLO5cZt4K3TdUtmW4wCUm8TFg/fBFMCZ2ZeEiesN8avMVHMed/JbNiuZsBzO3WEkPr
O/LbvEocHHtRKEZOUYIM+tnDx7UiIJyvc+YOMjDsn9FprtM9CTu6Vjh59w3p74JDXPAHxSkHM+wk
af8iu1VW+gd1ocsQWO/FL9sZo/5v9ZwDsle/7CJtavI4nwN8hyuEr6E4Rql/Eo05iAZ7no9u8aiS
XPcmj88CG/EsVWlat4gBncNCBITsOXgsCWjjycoqt8cFRvhJKd5zvGscS8Ij38Sfuc/fT1Bn7Q66
mMAUAOEpKcZcYLwVHdzZnU87BVdEbUh1h3bwI6aXfl2/0gBVVJRwQrSkpYT2uGkW9zWxAEF6XHS3
j4MyJUJDmfQz9P/L46EIswcsPAbGe1EgoyISbf3IPLgFH05Qfz4ZboRYGlyk4oIOJGAGNVa/tfxz
N2fsiwamIwXZ+nMBArDRiHmOj+PRKyAckqqVy5g+wZ9Z5WvgNivRP6cXg/0omN8pSdGUhi1/T2Ub
CKVTuqrsqnGNhhHfJn8ax0CbCTTYAKivm/bsX++V/XsMSVxz7iihq33wdlgYFHi+8ZnjElw5WE8J
BFkGDfGxUv/iCnccE3x96KvV3ZS/xxBOEcsd6a/5zBVrKuJ1XN9P9+cCtsucJ1PIaztcbX1h2th1
pNKLHwCxXzczWw3QiQIJNTQKKRMiUYfpdCFdi+pWJr2VwTlOUIqPYOgcTQzY4XyQZT7FAczFcSwW
+ca4xdPPgT3upbH7xpu2H9XQ7ubE+HuFLVUdDqc7x4JVRlRIWFlRlOmQgM2Ikn9+zfwZANHg/u5D
xjOsjXgI5WzOr9RHYCKXD3wEUzlO2TRarhseApvTO8QDng0dAy7Qs5VE4FfYFFq8stPW2IgDsjqf
NZJpP7tQicFWoAKC1ZmM58XLgQfRIl8gk6PsUryNWVbBYtIj6AGjl+TNrQ/M0lDcFGApbzAu9zeQ
slLBEVnNmdF0Zp4hHTpqupDJaPC+RHi6k8oVK1bVEHxB/z4zXRyAaPCDDiwIux2bEQWSWpzUlxle
IQkdCdbWdOwFjC+tM/UH9lKviSHP4JPiMVt9ykJEekmFGisjggYuF5K7lEutQ9355R4bvF/edphc
p6rN183Q4rHE0tg2N7oJT04QgAvtchMEsvbZiIKW1Fkx2OcXPXENgnBhvSlOYgjP4fKhS4QmTVpF
sNv0EBkLmK0Cu6rbWu5YlP4z6OIQPyIJG889vR6vwzqz98YmYB1ySoJZR0wYabiIpBrpPTuMAL4p
JGRUoibL+wj1Ns4WoCTihiSMqS9JsZsDUAj5YR00hBZok30FvSY8wsbmJuGKki3r9L7gJV86gIYR
fNkJRtt1ss5cWgs0pZQKSSTWGlE7Yt4/3sK4D3+4fl41BO0t17fhTu59LsZB23SvSPHoIVnLtbjc
2KY7eCuk9oW83y4Ron2AOJ921ddqmvwcqa77nAvSLJm1S/VgS5grgDoEAatcUmh8LO8S04I5oc75
uV3HQdxJSTM2VNGwjQwkfADX80C1SJPpavXpLVNwMW0qxtMKiJhFPGllQxr52x38EcszNH1OmsBn
A/vstJZqx2eNrJHhXDyZeDj/4Yscg79K2Aj4HlK/d8cwJDzaC5ZzGKqKQyh+UElHbcmhMHakLJFb
JFTFolahol/4KE7l1eQMbyZBR5tRWYtZrxE3ysVtx7OpYiMI5nJIGgrKNC3oTLR0dU7z/AZZ58pq
YtFIBTEUo/Qk2q5GHwf37B4fqb8AocADJ9bd8hkHDIzdEi2S3f5yFWw7oOIaAe1t6OxfkDH0K7dK
iJMAyPRYUDHh4xL9FyiFEQrMfxnt5XWbbZdnGHGkVrE0+e+Df8szFGSQ4a7l3FGKA0uFFQdGF7ZU
rtilT8gZ+3PUY1edYuSvZZ241BH0MVntJcLePwG8J4TYZlWdW/+o04dcu0qynFQLJ/BQ+MCAWJOY
jXu7Jm/54jQOHi9YHDK/2QRbGMk8B87WO2FgGvOrvPJVw7t/1Ruq0sGe8W2gAMmSmV994Wfo6ZHT
u7gNm1YSFE81C4voEELFcop1FPHQkjfgDXGb1BoH5gM7RtnmrFUAqN0l6vvDvmftYJZkBwbrDXO7
LCDXTCZDkqvGHZGp1dccS5sLCc4ejRKJDTfqHrPsFdxcdSJJTQQ4zKQO/fCaU16mEoWftAYKfdj8
rGyaaDU25ncmli2ngLzz4M8eef+cbhm79Dr5n+RklI1QboTxfj5rqfUQpY1tDJV4x52Q9FzRhnH0
cueGuHMellRUnypGVp67G7GTvPJqU98bUVPqT9tgUt++dnrl/ohvzTpNa5pLCwogbNZb0IMsw7V/
cOf8x5HGFzKAxl7U4c8X0uBESoXQeChnQ+EFw1P0pgrxnKH6jLS/MLqVwsgGcvtSSv8qE4ihruGH
AoCutZyIs63T+JBHZxCNBG9J0qKJ8pvn8ecicT0lCrgor7BSmejc/HIAukcOaFLiN72NNBeuIBdu
vVPb0Wj112oMlXKSjnzBnMVxnvwTjcsjp34O3KOS+tUJYt0XmV2nB9dlfVzSi4ob03Gi03BO0k6f
vEectXWW7uAHXy/IxR7fkTIqDIUBx46VTiREGvvMp7A7oiJ/S6I/1qqPTrs7qbFC3juAgxLcJgpl
u4FA559zK0UNWMcsepSvWjJLBofII8aXE4a+5pCdpf6OmAT4rZL7WmWkoLamQA0UPA70M5lFYvhu
aBm8o4vmKf49bIREIk6GpOCr+yQWDmaST6UR+stWSfcXQQTWiZHDxP7S8nXa2KkKJLrjBs00E72P
gYm3/uQKQiEhcr0sbW4rqCqWjGPBX1MA/UcOD3oYIqdffng1lMnYVfkRHxjU/oJ6rcxq0WJJowxP
wG7ekrF/4Dk291sTvAQlUElSdLpCJN3n5lWQz/rKtBj3HcVAkbGkgiHzbAKNlFlkPz2mLyF13qf7
PxsSTi/MsyZ19ocJUQANA1Rz7Cqu9b6Wh0ksSSbX1E7bz6RD2hiKVBhQCP+KRv9/IRfbFaZ2WQ0B
IuLZDLqe9orMeiwcQCCrePcLJe0iq9XngK/w1SD8TalzkPbhInC5f1plrUwdf3TGoTelg++ajo1J
zgxS0ZQ9doBhuYVzF4uN5srykUgNVBnWxdMXbIQe0RUJunOOyxjjNP/K3H9O+OXYf5nhLkMmfk9+
4GqwS/njL8xkgZ3uVOXCGU/4np2KHbQN17tUk71kpOIz+QhW8q1CrsM+Ylk4sdzXMhF07hhUhwAI
9gkALQsxYpXRVAoeXBDoLtQo63VZRuIVEi0s7a2YnYH+UTSfn9gzU2ChcNwoLdvuxcBPdPej07vD
EVhuBlb7gUwOg4N8r8rjLFvvKT66sNAI+3+e5Z4rKMT7+GLMQ4+eGnldC7pak4CBKh6t8t4crb1G
XIPE8NSva/DiILPN0OMSpeRenBpU4FGoH43cj/cTbubW62+1lfbDT+Zuk/0hbUYwRG3eipFDBuSq
7od/6/Ne8OEpQzCVnW54H7hokt7E2Rp0F8r1lU+F/RW2S7HqSyVNjjl+ojLFpse7kqf3gD2WI3Sx
cSEOJd8HJnJ0qbVF3WRCg8jmkGqlHCVw5aSWbTMMnMDp29qKd3HwHdlRLJ5s6UUfc8/lHMBv0nwa
kl//ykaRfalwhDu4HZlTPnezeW7RpRfDoT0uB9mljXfkrHRDSmkBde/3ecr+I2h2RKNCg0OVacs8
VCWBDVuMuzYnHOULAYSuxX8rpCSQC0ZumPIUhmRcf7rOnVMP5fzA7ivJUtuKtiV+GVkjENgW4O77
776s4E1mfODxzacJWDfTQ/P3fOomjRgQkacPOd34GYu3n1nCVlBca4cDd+hKqrC+4gkBF/NzWBst
pWKcgEt+U1G9CLsZ1xZMPtlQDCinzJPOi5l6yGrHTBIu+JsdGDLAoYFx03jbL88OcDgmgL/UbbpI
SJgWL8dY5iSLSIgByo6xCca0dRcIKa5zvToQrc+EoM2WqwqVa9kQa7/u0chS4o97pR4zH9gbFocN
QvKDVPssb9c5x/e9WDspC6CDz8Fb2FA7FcIUPNFr1x47ivD+XX1Vcse6W2O4Aeg8JckhUyOwMJCl
W8Zkun1w/8g+veKgK9UKbjrNLOLMPUzMiZ2vhrLQNchePS4rLtLTUFt6PvgpWYbHwpZkamBj+Kvw
j4Y4zTaNbI5YD0PrdFRVfscNTNUTJ7fD42ej0LHGHsiSrKsr7jRQoKMeNH70U7ihPUM/9PskwsuC
I7DuaHwDjgDAw8bzj3TUDhRhX+Ce9h4gwAxmrpQGrFw1HHUPjDk7KA9YNOl8gxCP7MTxThb49mr0
nGlTALmMo5wv1KX/U6Fo0CmHF9guFPuJJlVjLHq8RnQ/s3ALDcSaP7s9P4SuakVeYovURlHZWfwT
5v+4kXrDmxlB8Usk83op+F31dQrNQdgnrRmXMvu+oefjQHVhPUHzBSdUkmjrNyO6g2XkU0HdRGdG
g6K+H47wmfxsg7iq8MIz0/zodu+yiVxZ7duJshRbDIs0PMWfmwDGwCRfS49aHx5lc4IqyB99ZqTb
5sPxJgevSX+7tiWgxI2LbUM9P9u6lPZONaeRXQaM3Xt9SvdrUe2epZVS2dA4F+PuD1tZvOospJHi
+d8rLTBKyre/DyZ/0YUqkPF88m5iy8xQXECl3Mtr82cP0NQFqQ0t57RZ2ew+9lhttxq3MPXaJYet
wWGFa5KvDhFpQmb0fcDmzmjGaZeomyMnbqyovV/HiJNkWvQb/R3L1OXYpnYd1POms3bLobXdd8J/
V9vYSFCAb3dGI8wpQOR7mxV4tIUUBFnEtWg0Lmbb+db0u2KZDeMEsm4cB70YHf3FFlT6ZTxLHAua
UcxT3Z1p5t129SWv3jlx1MTAXXRYjMDwmaIcVjLTlJaIo0fdU/t3nYh4ROyPOQNaDzULDnuOm81O
d+Voj1KULsfEKNyDl46TqzRZQUjCSObp/y6dBjBFk/zACfTBmtFOvNyL5dwdfH6/o2NetviKuWqY
u+Zo9uEjewSP31FugAmjq8xE5VMN3qx+s0ou+W9082U0he8lUdV9D1l4erpncgbaD4J2WD3QrhA1
hs0KfnnKY1O+ILJRR0G6Ev5VQlBoPGJ6BMtKRnWAryVfR1qOVCz9T9NSSvqL6XgqOvrZQvi+peij
O++EXW+o2u3Kdl48U0+HghzL5CrOmj0DELhuYEOhSfcS6lorvpvuWGJlu+aI3tSJRM0bpozd2OEm
gUUyzAX5zGb4mJnRDXSboUE1CexeNlZdlApST4hfnLLWFT0avrMVwWU1cNOYoDcd/7vFC84NnzAo
cXs+ImX0nVzBSaaJiKqtA9ZST4qFTdALoScLf5+Co2aixd6lVJf6PfERhGXpdB1nJf8Ilbc670YS
3aWoZDKWmk8HJe0kGRKRuCcXeGCDkPVwmBINW6+ItzNoGMnX/c1rNXR5TVx1+eQXtFxJH7geuZ7s
5BFIbkT9sh3ydlrAGIWB9KZgOkTwTPawsTKLKv2pCl/3xYtiimTIB2M7BcP6I5gDlDGGEc4lk4En
eGvbKZh+d+GGFUJ6b3XkReaKU7LeEvURiiNf2kUzZi5LMnrIoZBkMHgJgtAmD631lOsfAjoNhYfP
Mrvy8jj3KzgiLjilnwYWoIW2mTLCW86qy+LiN5zmc48YomOzkLuZK7c2kHlegB7nQvFZBqAyLpRf
XSmts3exOlo1kVrRU1zBrtWyKks8ezPsXjOS3ll4mfZ/mmuvVrXqROtyBK2zfkQrQB4tIAC2QWQZ
Gr0L+ZIPPYMr1ptvsaDBQ4SpJ2IrslKqEwq7cYs9qAdWbF50U6hUMhhxmR8kLd5c5Hm3TTxwMLB3
wp3GtR669LYPeDJDUiBKi2BipcdCWDFmhe2UFxqTIAWPlGXkljh+LZeR2TDIf+ee4bpSBbveQpIp
hoGUS1El3AFvKPZMihRGsSUBJ7slD1RkKavvbrWvvJDDJi2S4HLmaVOsuQhnfTE6LbxlGKKO/MWI
o8Hy00Dxp2iE6nE4Jl4iLrbQaBNGyJAQEUYMF9R5ts7N0uefFf1zePNInMII6pKRtEH+14VsBqgq
XIsYpOBxsfp5q+TXjqmKVqivO7XXYYUjsrbm/l6hkY4IqV0dieSAQLNg7th4DEr7zRO4d3WZTVAt
seiItInH6VQ/TpazODjhmqsHYr9tHt6qWRIPZ+508UA5DoGdljyl3hh5SsXlEcJzb/ApvKM0w/K8
MsMhpgozkwvggsYPvAKeG/BIdKErWIU5nUMvZWOS5c6NgaEnJ5qhrEAocOSeeGguSX8gi1EOwvXE
1q+UZQJJyc5dxh2LkrsC2vGpUwf4QUodJMmRR5HhOdm31SNeJ1kB52RRhzCT0NJ1VjPi07mMiRsV
HGnJEiIxRyi8QRGfu3KgX4/Us6oH7xVGlKKSUmRqGcnWx9Dvy6LKq0/BzvClllV/kiPlZPzgIoXW
y20m+JMVHlosu69GZvLPVGVUs/XW/2wdOCEJEC/S7mq/3aoMyz0Ge6Y2NJ3SOMArXO3frN+5VYsZ
YXZgbrAz1L0CtDsLvDzrc3BsCQLkEIFVWqdv52/ITHpq2aSqyW+awYzGk88/QGiNVDTYYM5j5L9o
FBmsey4VF/34tIqRkZZxCL+k1NgwQOyENxoHnccbY8f1BBxpS9+eVfX+2rUhYK/OfpFOusLwskQm
4H3QZq84dXpfWTA1f7rZIPuOcB+87CgBn8Bg56KYLcEmNYeE6+o2/J4rUz26Uxe7LxIKWzyddr9A
Rdb4E0YcJ5bhovVB0VGoJ+QsIuEDND4f2zljrZS9sYVoK60pCFbiI479Gd9krlQcNf30g7UV3Mtf
Lzxvgckzjd8FY1QUKQ+ZvC0ccSyS4A/8rnHyL8dkX7G+KPtD35vClXeWiafiIm0OgBs9FbV3j1AZ
B50v77mecCbg87Ku/sVDEq9Tfc/zKZR7XOJcTCa/IAO4ftq+b0kUD+z8YTs6GUYF7+Tzc4Oa/h0+
X7GQfhSJhNfLD27v3fPhcyAZ+TnwxWj2svKLZ7at8l/Hmn8j1dGnhFqLPGZkme59zb7piom6mIIt
pzaWpXv2Vtzfdk7UtkPulz2xiParqLNXhc5Mp9Pmxed5upLaJbPXRmHLFCDC7/yNO6qqVFLCFaJb
tmdCLneTm176M7umnfIT+8lUQAiYkIsLAU26XasqWvNVKGNeKhTOxY2CXQgVOT/VuA8OoEH2hH/i
CIVwY6RBwvbaLOsCGJ+2SnLQc8uhiFjZr6ncD0XZR7z90dSIRyBZp0bMovKtcQQe5V2B74AKPlXD
4aC85VBzB7RBJZ51JDiSnRNBEb3gEhzsPc2B7sRDVIrU6YEOPxZSfGuXB7+xXgkgcGIR5nYEmeyb
6n1hOyGJv5P7J/oC8zmRmCDw9LJYp3jOf4dkSt23DBNUMMoZakh4yKFfh5iWKbReFrLBxVkTJBHU
dWhGG7YZzY47lQkehkNAE0bpkpqgDwZ5GzmikVWz/ZYLFWgndfkFuQTdma6ciQYR9aQBoFup0Iaj
JhK4WkHF2JZy2iPLQRhXCtKtdYodGyf0OuwXXZDRV1g/bDusJ/Ys9GZzthMUVuzalAFYw7yoM+k/
n+kZi55F+9/dWch6dKI7Ebb1W2WNWEmgUEOKr/GcDkK29OS5iUURNySgxyyS+eKJ+LMt7PiBbeOo
4/pzwdhKmIfgAJ/miRlkLT4+Himozzah3OIJMpQ/vz21HlyKFPEsKBWpHUPGy07o1TcjNp9YLcWU
W+E80EDPCcb7CLyqq+mII3Li9DBYYachk26RBwEZoDi39TKf7/nHoXk7yFL5hSuq4VseYXxI9NYB
x8vZ/befusP8DXTEqPrWkpiVC+LIeVkS3E6JULyMcFW7dYy74B6FVbcE4eT0BaeL+xeH2Js9PopM
eH5PqtGX4xIM12jtQIjLR8VNLDYKU7FBSeQmB4wm8Oy9k/G9MNqOMWxWvBQEnRu5aU+wpbUAKNeW
4HB7eG8A3me6/Iibv7p1Ylz+ewClGEqD4AyEhMConvroCA6ds/pBRhWZmYkVxYZjGTmYxR4HfONg
l77tfb40wet7XEoHzlhSLag0bp5EBpjjDAA7A5FmotERklEz1N4CmokOFZGip94Wi8npldts4Xay
WDIpRCZ/kTi3jrqqiwiUIndWhKiUXFn1dsgNvSt2b8DhEUbCKM//BP8dRosFKE7Cayd2InIU/BMt
VBNCKefXtOo78VA0oxVdgzbfkGJrldYFErLaeW6D+dJMIW599Hm7ZXvsGfhQhOVi3biLw7pZZ+/6
D70vwLJBUn59sDIINhY6dgZai55CQIajT5GRZlibqRRbrKYPrYZQp3yBwoWmE8xr2uoVmN0lN536
SPIgciq7R3zPW03YWB/HaK+GcMoZ1/qZJXyZtso4qotkiw7CZmbz8HkhvE47jTCl5xgyAp07PwFy
ghCFjAFpXS44aI1v8v35/V66HBHMLOASWLspf9e1+0t9ZZ1NShsk4BhOSvoQWO4/z16xU6hdAXQc
AohKAcxtqIeotnlN9vtED3XLCzTyvanRj3YVtyJjCjdnX4DQXA2wwdCxcGa0tE9iM6rCRCzhTJHF
T+dhB4sfV14KndtSfvulbzUXKnsbNy6hTPyt1AnXp6KhB26PfCR9LE1h+rwNy3D2jYG7ag18b47J
FLs2/ZXJ2kI+yHUNLu8iNQVF7yb6Sxd7yq18e13tfwCu8cyuHKqaFQ4FdzW38OJapSa6jkWZHAVU
lbyZycaHAlf63TKE75oTeoGdnOBVtD2tf2QK8liGRN5Snuls74Hspd07KPA8cf5IcaypvjgSibTd
xpB+loTJzBsFLrvP36YA+FO861W9YbPyEqQAzxU19MmtjBj0L7BF6n/7mUpOcgMNZUFRBc8DrscG
5eE9nDnxtIo5fTxihhlAMc/9XEfioXc4lV9cdIyCQjXcL5ZlrtotiewktWRCICXeZ0PK4U3Gxlrg
pQRAexokYSzwWOp1DnoTfIE5Q7khX7IiEkGcDFyV4UiAp848gh8acOku2f++LnA0wld0Zi3kYgcT
gUmz4IZ6PIYkiYy/4XUgoKJsXMcFVC9oIRH4LcFuuLjbpNjs9iKV2MddAjPqE2q8uL+Id4hlOwYI
elwM/9E4KI6Znp5tjUuemJGvOwj+iIxBl7RX7XBVPYyC+pDN7jrbPGg+v0NMqynLS7DV646dxsX1
8uX5n3KxDt1HO7XfIHpcnAWph0gCALY1UFadg4LjdaPYwgVPTxxd3V8L/deUHeNyrKlp59ZAnwzb
ge7l/nZN0K8BCUeVPgbIVHDRLeFDLCzF2BZRJsbybN6HPgGXNxTB7jUtkLb6GvesM6j595Luxfcy
MePov6+AXIT6bFlHTqGZrhJrnQOH50Uzwblr6DDYpBU02NTy0xxAzdBEgs2fgCqS3lpesaNC1IIK
9CeaHW89tx7Sb85mqNJeLJlddfatv+tjQDDe1/WZYTgKAklL1AA/zgvBx9JKx3hssiugQi4r2Eqj
5dL6tL4oAZFkkJm1WzbMXZmnXKFFJhvO8LnzcV/FYBTvfxidkU5fNcKRBd7SSACMXkak/V5KiEnR
lH3GW0GSRWguxwwg3GoWU3lnU8rx8GKp5oFJ0cr6mb6G2Lkn4sa0TSq+6KZ1VefmhEiehIbbncdQ
tEgADOOmcTT48/WoCUxt/b5dQlsCmWTBsweS8PNOu+M1MZixQLzQI/uPPq9hJNHtgFvdxKQ01ju5
BzLkpA0+Bfkc2H1Jakf+fIsdi+qWO4AcDWCm0L27AhxxbKl7pkUU0VAirJrWrFExpfzkO2hbAf44
Mm5C4qfhef1iMQz7wWAvOBuVX48OWIq6WF7yixlZpG2h51sv4iNrmhyJ9QSD4NAPrsMg2MHKhJ6K
f/uCNt7wvcp2faWk+fop60VdrjC/kyL4r9muccjsEvdZbjtzUbYUXjKQl3KUnqBUpbkNpOajI7q+
4HmCqJNX79v+0Uhjcg/C9Sr+mkM+zF4dOqqkRZlO/y9rH7G8+0faSiqGzpKD+KI3y5EKfz0G9alq
yOrohsbuoyQazl6kdUH0sdLsQ1sGPrn6MdCEo64lvSKZPllcfvPbBbVVsop2zt38KSQvULBCMKr7
qKVHi+YYJYqU+lVQNMitC2V4w+mwX2TUQ8AOjjtG/4p+apMPN/2mMW4IjHqOAjoLboNssWF7wpeZ
36qVki/aeOlPd2MdRzmSgYtYg1Nh81vFVk1Swd3+xtYgN4gH6arnUq7/lOSkQvAe4lLPjc9dtAV/
tS0zJONghIKt2w0TScc4oMHY/rwLeFP1Vw6CSza/okelicewEk94WOq6nH2i12enc+fnf1nLNbzP
fYmLNpGBY3MM8s/wOM393sNX2STDaSdhvYp/lEfVZ5ggTrWYvaqdXFVhlhpVJaCRopGbLvKm0Y10
o39xMezsfjF+YGQCQ4+BHPdpFpQBilrrPHyJ86RmwAjs6y1Bly2+T1tJd8MjhpY10bPPqjdUkHpZ
BBHmZMpJX0vPrURyaVhkmDLcQzxKDyf7XY/stRoj3SwlAfwDJV08Xs6GebB7ZmZcog45/GU12OTV
4C/QjA/LzStT7KxIfR10p/yl4bFs7wnBIPuOkK5kKpDtINO6sauKXdDt8ZQWHE4yEvGPzYkSA4hT
Of29OYDYGi1b0efb4Bc8l4GNS24Ag7GRxBnQdj1n8fiW2dhM8z4O8kZN3A/aXzvb/meF5s4uRcEH
oAs4XC9+u0BsXaStYnY1AO2Wb9oVOs9Zm8Q2TEHj58aNb1ueL1rw/7RGH+5CECNQlFVXZL3SbpGy
9654hOUzeRS62B0CIKA+1qUnknmh3dtD0kRB+0J7n0/DqCTgCoea6C43IFj4XWGs3Cu1wNRBtyEr
6YOuhYIcBB+4qKZ1S/T12M75yu+UK4kgHfOghODhG4A6zsDB0BtYu466XA5OQnvpSzTvSQNStHlS
cx/d/ThjFP/mqNeLrKvLq7WwoTrn+ZK0o0AZr3NbVqEK0wNLA+96XTR9ADNvcLJyyhDP96tEbkuK
XYZWdg9ElgK6HLm92V7TVufJXcHd53wvtYUTYaPABXQsRMh52YqtIifUMy0d+lfQUtFonigv/YaA
7rU44/RtHqliEVlOB3hkqHH65pvWamJOf+vfjL+bJiQXQZA1CmH3e5lbmn3hBk2mtNoboOOUxTAg
J2R+jE6yAuhWgLjTEYGahaDjMty3ia6d6cfUnwHjNC4SagqiobSwTynWJfl4+fweJB5USgg5CdWb
1rVEWyTNfPYQNEFD6Em1RlBhy+9kGfIo7oiEFDB9HNAkt2OI2JZe0/rOmSCESAMn/q9P5zAoow25
SYiQehiSKs2kX9dkTuaLG6gH1tmgvColYcvPcZWUUhnz5YEaue7SJ7JkBzDnqcObYkn3JuAI/Af9
XnR1y6ZEX/egR/i70RX8aLQpu+h3331l0ybBrTb8gLetdu1j5zmdpLQ4oizH7tH+Fvdjt31CfolU
cx+BCUh4wQHzwgQIx2eg5lvg57NkHRpiTMKB5wt+A8jNUqRaOD0tI4G+ssMclr0WW8q5h6FiZVij
ebBoMoYsm4rkhGZJVcrZGFseYZgK7mw5nuUltYBcfLBEyB1WTnY8imcwzuswzhcM83Gy0BlAMZbv
Z3wXgxFtIVWO6CHprt08wZ5ClKBwQYWH6x8boN3iueyGgCRSSueSZG89uLl0/fTSO2jrlxs418nS
gcISVuvovmNDg++BJKaqaqTyv//icqOmZTl0qZbfFKyyeWXfm6vPwcMk6ooEc8bhxHSpuCWzsMRU
YcNctjbu+slubhI+zNYgn98HhXhOEoF54AhUV3sV9Bd338HH1M0Hm45yLOovHKaLhUBblVptJZha
0mnbq3s3XFKYDbd9XjIYo8dT/DMCBITh7g4T6gE1QBr4gtP/RMgDQ5b0Zrqggj2kFsRGe0FQzSfg
DptCSaP3qg520WvdfiB4UHC3YKGLJ73Y8euLS14brySiPXYnOl+BR4irwZAOs8PERh5E0NZjdg5G
8PxwJ14NZSOWZTi/BfQSvwsezu7RLBa/HK+IOyAvrIRpo8bbuqsqrdNWob9fwkFwz0TwFjs6BDD0
uJ4I32Zr14bv0znpAHuFZFuBCneVt/XeluTPzQIV47vN1oqvmIrZ3VFRm5OUyw9DwuMwCFdDko1G
2fpyzDU/7rVf9S0FfS/8Iz73spIDKinU1g9n6yPTgSfX6z/voAOW6rqx0I+YYV+5N8WbEsnQB4Y9
aTD/bKOUOd3uldu/CoGetE3oj888mffyYxgpyXiUc1MGUjqS3ugZDEgAQ6IlFWwXGTamimXWiXLO
5PCOe1Ud0HqtVbd6WMqdO9C2PnFHL8OJzS1JklSoOFqbpTHdywV/03NZRz7onlgPIFRszu+Exwfx
9tz4tdQuWiCUiWCrfooTJqZBr0vyzjk0MIVem0xAtxmYm0MQlKgTxNvXqCi/IFVgcdCbhDPRrDua
bzGFg10l+CySnYwUWayiWb/UZlZeumafBYKa4w4CBx2ephotpYO/1Mzi2dcaBYGR7PklCyXiRonZ
mkgIhRCUaUXbqGPDla+SvQ2t//Gfvk8S+BkFWKKjdE7Eiljrn/J1GC8NKvygJaAdn4GCMNFhSN4K
nTIw1niQqq9wW4cAJcA9Qwym4Z8oPi7Je6u+QnZU7qyQEFS53R358RKiTJ/i5zciVK/375fp5P3f
efSuEk0vqDlzUBJLl3lICGEV6dJ1e/yS+z2yWWrM0/h/6IyE4XcDd4lT3bAYcHBy04nGn8A49t+J
XLmfKfRkL3zBl+TJ7Dy/hTcDi3lQx1ascPEOayAdrLPRFRvmJfvqK9UnrYznzJeyunsSBepVLOOf
26yDhsedX7SJWGJhPquFJAiTETkodGe2IgKw3NibDUUuidEzQBwgBEF7C+cFSBpxyPOE0WSMfzY2
l0gn5CGVj0LwUMTMQfabWqYyStL1Rt+GzqSkVjmYEAKtxPaPv1XgMFoKlT3qSvVQcIJ99CiqZmQF
dIL6tTGHVjCxlAQLnBKwNNSAZNZlVC9xihiypUjZ9Lb8/U3NuOqR7YDBgERbWk+E1Vj3eFvL38K0
vT16/B2nyhFCwODsC/2CvtMXg99gqweVdURzoshGU2PjQ+9A0+yEBowYJ5Af/hZ8PcKrfy9Wvq2T
nH9mNEa0s6b4yM5MDN7vYeNEbgn9Cm/FwnrLZLJWUTOCXlngMeY6Ii8udNSwKfhJcJWOqEJFLkEh
+Y8e6tz4aWKgvAAEdzAy+8rE/M9neCikIYLu/AF/LeC/GlTLDx5rwteizRo4AlNF4dl5r0Ny8cum
poFI1Ws4OgYc/O7Fa0rYv/Z+KFFu/YXBh1Vud3FHiRCPh0PD17/iWEGm++KH2BZ5E0pcX+Ep/Pq3
4sWof8VXXapfEJfEoHLkSAXUtnoff/Tjibi41k4AlJiTo2DnIEwGIbeIomKi893yfjiyzlrIBPVP
f5+lHW3ZMFD/hzGCIzUzQbcHBN5fpv7ZyE2ebcf5vsLShSRupiIVbMPJrlIrKFvCDjcS5qWOIwxZ
JNmwIEar0DU0FYY2sAxS+eu91AIDqEa3rkJ7o5nSVuVHxkYXG5Z4uCtAWd7hsyd2Gq+qh0Lp4zW+
Rw/hmiJewOBdhCFib75WkXuKe+T+YvTsCtCvWjIqefs5ys5oV0b8e5jIRabU6sZh1KXBg3H6kLO8
r4pP+lv+1t5jDPf1tWDm1yhbrT77VKt/A4v3J5H/vO/UShwgVzB4Psu13Vp0EpTAfyGXCV8t19Si
VAqHotvUTyOoEioFxdRqGfJUNpDMwlbjEHeHnv+2GelSs6i3UT5vwfF+9flmstCJHV0t1WDJ1zR2
T+M8OggF14DsEzbo2c0gV/lWIrhvcsh+chN7R33sswxtjw7REvD6Aol0k176QWmNvbGHnyZzKhUJ
vMh6e+GtUilwDiAYeSWcTF57IGkNl2rpPz+LCGFQOBegY2lNN7oGCdNgkqdTDyqoaBPjOCPzkcTU
js6qDvCsGTrfb5kH6Ju5ymIZFPJ//JbRo9cAmUYNQQ9azvATsQoodPiaRBu8JPOhrT4FS4sPFG10
7htmNvZA7Cq5UWsUx5HxJjMSpy0TXNfu9BwdQ1O3pi3BT+MOzLXrQsYxpWydnxXiOtpZ/hP3J0dH
ZSF6LJnTfLSKR6wWaCQJl/T+8s4HheooNg1D9vYFzpNThRZDHMEtFrZE14PE3NIBBWtV1jdbNwlW
4k+nu62FfzQcTzDX+MPcWwB1ooBKNk+cJT2K2AJ9uAdrYeBIikTlXgICjKiAhnZy8rv+jS9LN828
IAQ1C4HADVZMeileAoEGKMadN7QUOOWNmKIK1x1OwNI0VvQoWpBz/RsCZu3eRWIrTPqUwsQ+u9ap
QzxA8Ku1Xu90NPI7nWAyOMcZ6Xp4hNVABV4PJEtK8PM7ix3iRauuOdfEn3SDs/GUWW7M1+I7hfRo
1DHk3ev+lzYfUNPVyLOKUwXTeJQvrtcCWUAvnr19tEpmgu+9zvywVmKMO30wMnmjeoUTKlSzPQ1n
RArbDryMAkY/hv/34KPvCI6PmjNX0tHn2EY21mojyrYRh03KGRM+5eE77whQtY184h+95orlVqOp
vpKbVnnIFDnlmH76jzqXTuKw7gGZ1ejlgRUt2DDV36gaEZ2V55nKrKM9Hr8hzn2bgSvko9sQ+13V
k2oZqwf1XhaDTiuQurbnb6OpokKWwx6BDMQvmZDKB+jq6lSTs1PgNTMZN9SZUTq83wiSNwxr8u5Y
DzN5W1L040V2VdaIvRGmu5cL8M1j//SiWN1P612hKtfwjJ6kVwbOsZGOPV1lk9Gff2zToE6erkpQ
g8dw0vk3lP0Q74+fTwxVvA+Gt0oBpWqTTJHmW1HZsEphoJ9zpr8fWTc68rILKVaA44186XDRBXnN
17FmeBtlwXOyBi6T04lHvoYVIbrUxwLS9XDomJQVmofIpTJY1QHrwjmDroBpIb1OZFc4ZIRzHeU8
z5LY8lULFGNvgJYgPAENJpqL/l8W7M6e7LIOEm//4AOTJWhKveVs9SQWiN34YhwT02ghLyW1dYf4
AIE9rdm0NMXDjLPiyKkx13Eiql2g3/JxigKYW3YqFl0tkX1DaOJht/xIQ2Wip3MfKOBIamYjLl1c
owYDuHSqPiYu6aAm2Kd4IiUw0jZp64HO4XXDz9YvSBl9S+MU4VjSUeE3DtWVDxF6ZtCDCLRxuEg9
CYXpoh6IuvLsutfwRA+laAvcp7t1oj/ZH+688KfD1+RcbBLDkCdANCs6Q3rKyf8uGn7WLT5b1Dvy
Mxu52ioHodbveTnjg1uBAn3tRFvvDEVJJBjlEC6aI0SZkpUhyiKCckjIoYrFWhyeCfYqnLZIVoyM
fVMcVBl/K+mpJa0vpZGtDhr/jc40fLZWlO3fUKh6datMbwl5TjNzm3n5OvBBXSVSklDOsazm6/DR
mciRrCC3Mdkdc+7+fAnsFWVTlQeowHlVypsLKm0hcJ1sU02aaTG9h2hgNBzw3hML1Whx8yRZnzTI
3xoD6MSUfTouSIuzYCbwqch8SQsQC4jhn5/4vvuZBnCTxJ55gRtd3K9BTTasGYlUu3NwgLeT6pl3
GTZepW+LrN6BpN07fFvAxmD/ENyS3ybJQwuEwb9YtOWC39vJzGWPWy+w8AvUaOwv4QKJnl/qMjyQ
WdTKLTaZRUm4DY3xD3krhDALIDKsbMlU58ebJejM7rZlnKQpSQdLursmwusSApWDUsMC+g+bGq0K
R9Oi9sqOcIpKsG3+phW6o8zVgbEZyDcC5Lk00MZTak46dpAD10e6aM69tP984mhTnxSnx5SMbVqC
zF84pfFgDaRVouC7LjMslZHLAlGxAn1P+BXG3Bvsp9kgCoydCAyavsoam8GPTEslfcWGLa66JY3G
jyDP4Fnzci23quD+WAELUNNF6kTm+U1cDYD0pViyUURTmXZH69htwvNFsWCrFhVMI3wzg87B80/d
E1PX+4r33q2G/oJ7oXZZHbgl8DwjL5V3sodCusMawpwPuUO1/x+nUPcmmCetgADLy55BG9RMCKGJ
B0mCBvAD0i+Y7Aop57F4viYDv20uu+hCp8JK+056sAuhavT1pY3rQ+pYmFRzXPyxHIX01RNROTBK
+nAK6FuXmQjO4Fl5tfBwTqxNsYnv3ZGs9aVgWiMUu8aDGriPGpvF0ArKXZZoZXIq0UuV+/WNiq4E
OhIoepomUffgB0Gcjc7X4/IBJkCHGqIF1Ql9O3MhN7FgqkZa4g29B94r68+pStqMyulT0hqhTptj
kPKvTcy2VeYsOUFVgR3gKEo0xE+dQRyfry5lO9ifCLeYYqIlNdxUc61hMhujnpnfQH08LItoi0lH
YQBS5+ieGZJVX2q4+4BWcAwgqJDTDzrOnedNN710twJm8THsGrC91+4hi9KbWOMmL6dl7wpXMUwm
TEjZjfyTBoqECDXB/sevj6+6Atc9XE1XwnhR5V3ziO7WkqHpud+9GIs66hu1IOBM9r6wtT+Mbx+P
w/ASt5p+k9HvBncFN8NJObPtGMOCoiGg8yHYh83zlv8LcpjdgYQ8c4FV+B06jyZqzWd/C6GXyFqA
jDbSxg6i+fZqFZewlt0daevPXpj0ODKNhuX5jJsRpMd8iuk/S85ESk5KEpLyVVW3AcsHoxgEFUKF
F8nzY9Km1sG/aux+73nFobwg5rTd1sqA6psemlDkKjBLBIGBysxvXnXWBEKFoJK7nOzio3yjIsn4
NmHxdGU+VC/ydkCy/KYHqEztvC4GD2eJxdj+YTG8tEnT18e9EM436rpX3XAJdje2PYZHSDTjTDdO
r2VfYycvxMvwXj0sN8srEuUrmM84dCmf/i8amY73iOxUikNEgSVvtUETQFwFRWtPriQI8c36RuX8
FTS72gOvZ5ZUbtQeKFf6/6YHM5RhxN/ijJurttn5zLzxTWIJImA+zD4Tjs+up1ECIKvwZFGM+Zye
vKGtzUlzeWOk3McuOMoY6oyIomYp0rYhTo4GyDyw60FUBFl8TOJ2OLZ49dbEnztQ76vdG7y+oJqb
Yi2JJkjyshzlmVQtBWF9MG9aYxpnwTlENd0Wt03U8RyDUYk/j4wuFo06v5lLgNPszNHjIG9NyERU
76ZyK+Qh3F3THKui++1jCEZz8/37z3DgB3nY50jr2AMPzo+qUyq84uHOO2yreNJb2MNRXsduFTPo
qChHKbinkcLiKePbpDQ3aHnen21Azwibc/8Z3FE3XfkCG05jxpCikuiB5ISLCoY2VZKKOLFTJ75R
922jF1K0eRdHTWBnCd7tFXItPxw19YNuLRqW33yfCbtwQhU0A8HtyMdBMn7KGMr/RG9zo5YC3Xdx
0eT2Lw1eb8D9S9+GER7GQl/OJR3CjYeF/dyB+2pkEOjpz5QfhUyZfWCHCGsT5PHIk8zRwSq4jyiQ
G/sz8RzxKoUUK26ybvrdEGQB85K47UknnouUIvZq7uUM8VnZO1yq7vqE/VRkFY36SFL711vV8UHZ
6QQ9/ZqNmXqZpIK/EkFkPuQ5fzUd8FKqaK/TlRozd7k9l0KnFpotMZq8wcbamiaINqrPpxW2xLC8
v1zqfcRG7/IGR0HexVJk0Muqv9A1cDVxE+G3VlSdcVeTCIDb8qrrUk3ElVGOYwxA1sZFNDYAOadH
GTG6stlcWgu1kVE638KHN0oWvrMZ2q/Job9Q7j1H33dwJiue6eI1F3FvLRan4MoHsdQRF5KRUnvH
oZm4Wf2DDeQEYsqLJpPClqMxlCD8yP/XbStdOUwMOSS9zwThjGpkpVyh5gHH5A5cTjoSwsm4Irb9
8pzKSCTjwN7CzNcU/b89f7cNkYvyJkXxG/MQzvjkDwFCTOwdX+bfWRU4s6e3yULvB1xAR0sdA+XE
19d/AOP4huV+2EYPgGqoGU9plu6+Nxfxgkj1rA9bNt5miXVu9w6FVmlhwncOVmwMa+XVriy2mIrS
gVw/VUVUjKtGwXCQeeNP/HqGBWiTPQwsVwxfr58OgCB01UIGs2C0Irqva17jJ6+CP30RI56B69kl
dF+ISM5BZiEFNA33af96FRk+Rs7CFyhtUasQczi3NG5SmR2+OJfKCg5TpouUc+kau5+QGKmQq4oi
UJcUGcjV2/djqFuNJ1EyOw7yKD1UzwpTtilo/iRCTKEnZySpKKzpqmFYIJqr1tTTJ/Zpu+0ixxRb
Zz/WcBqtksZkw+nxeFIV4ZtL/pWghTHp8j/mc+6drlF2L235QJ3d0auGQ/iRPZVpCtMNtUdUqAoN
+Q6KTFTZ9Jzg1ZoAjxWifDnUOYdoP0duQVZfaDBgZqTW0C7DbhLnA8LSerY2f6iFdZpqNnyctKv9
sy6mE70+AHSShdn4xacWOOal3gMrLTVmrwkRQqrR31GAt6cesyteaBrBR04WAaPMKp8UmdTMS2iE
ZtgXEYHw56AiCFWhTlEb/Q452URvwussTsUfKXQr5frQ0M3XAatSVIDxA+KtJuEDryvrdzC1yMgA
gEnQAkJuRxNRGVAR5NxcVFTEMqk3bhKtXqNgqcQmbIK9XDyXN8z/lb3uh+lXbBQXUhz2dMgckEWm
zq5QiKqrRjlAIXdlJbTdIMNavlVNAv8Ir5qhxei4begsyqpGsbFeIakAPIfyFE0HXtuIr4SDv94l
5YCoXq7IgMVCzMvyFC+8RK+bNJS7Lw34fCB4CZxMh0umFVu43y6+oPKHC2JnjtNoFV/S5s1ST0sc
B0Wx/tDPFgqtdrIGGe+kDtDOoVzKOcooESPeYAd7WGEz1qbkbKBGxzWZioJBhtwqm7B2aiM3c4Tr
kJrRi79k8PYKt04bO+FnYQ62CIbma+smy5DYKWeQcJtHYgLMdrMu0tNq3oC3XFrE+MIvmfCYDbtf
O8W9mWQqJlkizsscdlbTXPq/zira6soc99hTqBCXVWVSkiLkWazIMQvaB2+86UE4YoVg3g3c6k9S
FfYO6Zm78bFnmfsGbwC/LjFdUnIPE2sxjRiGUlwvvmU8K8aQj6Bs4kbkrC/aP5ErWxf54fm3tioQ
IiyaugLvpF5sPQj0wwZJE0gQhmOjaqaGm2z+otn8QhdLZtRcvbfM/WK0GfmuhCYCz84NzQ+xhRcv
Ki2MwQe/7FN1zy7Y6Hr+MMsgV3eqXeDjrENCly8r7K4Uhxb3EQSk027qTrdQzeaGVCZrbcwEnTlB
F4fphGEXwgOj9WGd9YNpaKhpozjG8TpSRnkB4FLFONfAROa4dbpjtLApWasCzOzqfq7K56SamI8u
+07lC87mLkglU3M81Y1ZDBF6o+6DFqrCNbxUqQLyFwev6j9xNW6aezDEoE1bnfCPr5y+SyGxQT8u
5/ObrB+nxRNmaLtaSRPNdSfTW4TiRlfvYnZNrfMq1CUr9pcL5xkAnFZe8OzIYBl1icWMWOBdZaMc
ge3VlKhaVSXpZHwdS15H+pzsIJXEVeGQ18+rMfLIdHYDC0VZoSkTF47bNFN6Uq38dXjqfXuh44a0
bPbD9ZmWiCLu5GMqOPBXfT4Cu6t5wg13PCLb5hNWh9JRecxkb7GIIKTb5c3qeXaEoBiYReX+78f3
FQ5ZCW2L6bJ/3my/XdmoHQYT/qu25IhCHEq2OsnAm7hxItX/RI6J0rwQDUA4OfFB6kdveXQ5LCUl
lFfdWxoG9s1x9fqp+VJFnvtwY4nOwFkSVKDJrwxOIGe6x0LmmnM2hUSYz3/gx5UGWzsSXFURD3mm
XSzNS9vsz/xH/b2DQ94p5AZGvP81Yd35c9qYWiBdrINAGAacd1Xp9Z3cJ+Kw5psPuL5lLUgndSqG
a4SnmChO091h3UTakOd4Qb25cx4NR2vtIRYlxmuG0VQLPNSZjfbtlwZszT/1z8oI6es1fiANs3XC
9OJx6UA9IvytbfxdaDyLFcUjvErl1yE1nSU0SRFz97nsjphPJlBa5Gd5SN40qgNEnDfyzvl8f1qZ
U1Ty4PiBBZ16UeVs0LQjHrfAEwWLv9Il2ibDF6WY/9KSb2pINwqInC/Pe4fIJjCokNclQ00EC9qu
/DK0KF4uSei6hEy2vcgNHLgZvlDbNE2zjLWAM+duqyrVVuI/lEyxBg6ej4mxxkm9707RQcuiIBpG
fwselpKR4Ks874au+2a8uGMQkeS/qypEXuDQLz9/coTqQ0Phvnyy14R3UXskNFgoQ9mYkWldVEXH
GzL+TP96pBSbGKqYj5bKnkVgpPEzRqZ3A/lTRq77+6OxmOifd0SiNRuwaKFEo5uqT5Z1YT2Op8Ko
CK4tQ5IYTtSfB121FXk5NnXY110z7xL3WXdlrgX355g3fJMGt5A1kkOxVYQvqM3hit6+6kXXaQHd
jnlsal4+kU8xeJCc9uJ5aBWjpsGrhBS5kSIe+u56CD1tM+qYO8qutV85K5GI8Yc4RyLEJyY6kY+a
5Ll4yXC+DGcWEjmy28Krcv5bRDUfk8GfpU4Suq+OBZDeOV3XBzyOxKyZEBnY0PHLtxBCRBUkmXsS
gpAHfFFBPTcjXHcfS65lIhvGw7+r/X9WV8O3I7fN3y4piruTG28VDNt7ot99TPzzHNHhywVs+B+f
wsNySRiqT8c/Jvsp0NdQuqGJafdEw7HohdL7gPVYzunQm7YwONeDBNofwLjXqdqMu8fu/WzOOnXl
ypCSTUvRHJhBSX+zyFKL7XKadgBZXEwHxV8NDEpVWM2dLnNrJtRGUEVXe1MAAcyPgHTcjbSxmm6p
8leyF8Y4+BRlqNex0vsP/qJZBsRrhkegQHOrW9ZXHZUS45Uhn6Lp0p3oPptYzY74H40V5O9UD43c
NtdluwyLyhPWMHZlwHHfDeBHVHARXYjlzhdQy2qLuCECnEy/p5YoNm/RGSc8TwYQxVuYclcj/PFD
oFQnrvESie3gksr3lvLgyMdvTZQrhaK5/h92TsEecbkgvwhPzWhXYgYSjU5sHRHtb4KOC1Y1PHPb
QXpaQK5kURpvS9WzgJjG/FUMbLjSsn9IKMI/ftfy0jVq+VaA2aBvGM+pJLJpVH0NhNRm6xZfbuOS
O0h2Y3FUtYbdPHT9mjUQeo6l5eclqYxpgs6WaISBlSfL33mkNkAdvzG2BPFvtCA1lvyR1YN/k04x
Z16mWlSomM4pVMSZzqmq7d7ZK2+TqESFIZUKxO1JZBnsRF7QFT9LYPr33WMOzjyd49ZnLP7gE5Fs
+1GJdXSYz2fRHSPwtzalDO5hYxyfygQik14pFx7BXyc3LFnDLzglKFYg5cUoEzT970jKKooesp68
sm+54gJWTFzvJSY/BGoMVH6/p3H9Dz3zdwOqcv0mssgtaU9PVyGcOZgmGeOASSLL9BGT1tOMSddu
BdlWPn+8sj7pYanXKzan8x/HKYEzJ0nPmYn3u5jlkWttPdSZ/gALP6x64HqcJtf9ai3sQ/hwmiK5
hd5IS3zamI1x/r+tYBR1P9qqUpU2/gfzzBkdnSvzJkG8jtS4tLiX5eCARN7a51gKaUvcnSm/mOZ/
BTwdOjGcB4UTpcgrr+jlQKVdKJZ7LjpZYvUdx6CddyDnDMHWMfuAn6TgwMJV5zow1Ik7QBXaqiu5
33i/4lfva5s4nQcTeeq86Bx/lQh0osbaD9euWKbRrENF5VFQkFDw+GQe8xsGBQtQndceyobzH77p
7W0BqCROfgAFX6b8TpwphEDCHd2xFQYLETETIbWgCWkpYmGMAQuuozq9U7Yxjy4QNpLWXUl6kCQj
NbpW1JBSMXKsZAF4GgmaKleQ11EyJRKdLpFR5MI/+rk4N3t4Pc2JxhIC6Xi3XgN16TH+B2OOKYom
mFRM+gprQBTcZ2EOGzZqUIj5Ai8UV/FmEqGBhLbt1F7Q81hX8uJUvjcQNiCfIFN6mvVZg9npD8gz
Y3BxAeXRf3e3ZDLQrgTH94MeZFuxU2Qeyxqo5Kpvg85TqZay7/Oc5LU+XB3Bv/oLXgYa3OB9BG2E
cT0QjnUutnqq3bD0TdNK2T9rVOQyJY5lp4p+Y1+Kgm5dwNCNAKup+E9ckzHc1tOkQPcZZbISh5I4
tqBmF1IqnDjEB0mkPgGGeh29IJKYIVywwYIJ4+Q2gDQic0Prjpumk7h4sydZoSYXXZbo8WpMt58D
e6eHijvVQqbmtwJ1Zi0/+SkUkuoYWGVhMtR94PysDUyt5sHWqFDAnWjlxfCpvYte4BF4HqpBiAOo
sp9ZY3pgwGQk/wMNbITbXwbpfdK5FBfNnRd0nhqtcX1JTP2iFyycCrjXbBK7cbVdxmgFTQ7vdLbT
M7xrBewJ/nRdi0kx3EfZD5M4VE5YA7VMXrzE059qqYup7Eo3BcwFIde5amzyNte0D1vDSn1L4fG7
0DJgmY5IwPDFR8QPMTvT+c/QXXdaKLcOYtkTPnUcM4o20qZmpRUe4C+gJq3S6odkaw6vvleiT79N
JloZKIG0u9gkDvbm9d2wLnPJPaLXpY/hzUyUAPt8gjF2OHTYbZOwwjnVg5bo9MTY4rkl7gUpETvN
GvMx631HsNYUQ5ffAU6q58BV/65HxP4DUbuFC6rPhBQun8FK8SpGhwxy5MBPHnobXVDaIVEzbn72
t5BKf7vrRpT3mmHyrS0vp8LdYcK2NECD+tKVg0+23KTQpaeVegmWXF8s07uPavAVoXHwNHjrXFym
Ci6g9+0OSjwXS+1lN5r9o5KOay8T+FgtukkRHX2ja4M4T+1sZLkmXmeYR7ICwDqTz6YqVPz3N4bp
TXMrHSE5fjKhwiy/h87HO0WSxYou3ljZDPOSqkAqi++2ZlSk3vryhxpxgV29g9O0zeR2INKsNMT2
hWKp89EmgGkmRqDi0sH8+n1MVKi63KocCFUmGQNUntAUAY7c/GmyZU6hnlNWxMixIurorDprE/6i
1+ecnrV9dNeSEUEDHWlvZRRsa3UW+uQkVMTXmP9hsANsc5jde938bWHiDFILmj4+8mtWPtVm0Z1l
4c+a2A4OiSga6GtmvDjUk93ko0dFIFP0f51VGlFds3fWSYhjYqay5nzM6CxXqlEDL3HIziito5mV
kAWRqV8C3+LbDqSTgclfjkBxuCK+lKgOfsyFzx2jHeMd/Ljuba7iMGaPI6YxvzdcB5eieCkE4Ejd
L9Zwyn6x/CN7Xq0HbJHDBdtNXpJnSW6asrsniR2MZGka45GIetuPB63c07phYNSaLwCuD1Oe6hys
nWLsyjMDu7sooyz9lrLeGM+LrfD6XK8Bg8ACXMBIypDxVPXM547zbmSanCQV+BvzjJrgg3MCx0UX
tEKXd9BqKRIW414jwSNKrLoRRfDSfTd1jkSkUlrZUJ1CIVirnmth4kYUmxhAb+kHGiE3fLVb7uL7
FSb/8//5rcbqgQOxET7a5cngmhEn0CAQinE9DPwAVTB81qOqNlO98DPLmVziuNqgPv5mAjJxeOXL
G7xxvH9LZoNwvFYZ9NQJkdSEqtHBKSr8PUzDY7kYh8fkvZ0hdR/wk2w9nkCrD59Gf4CC9DdYqSXR
qUXjRI1qgIQPdY48khxyooj3fOPkRco16Tw6ydv31A5nggWEWUBrdZt/jRMrd+PtiAR9nDwKfUIb
cXYtvbnQzkb0WqHqgM2wJS+5I1ldDdB7h0w6pYV8KNsxkuoXA4qXlHeRLntigr0HAZk/Jkybac7n
A7I1zQFES4sQ2PN2PJeAwWFDEW8FVRsLkoRHGflukHToxWE3djC+zs8KENcrbv6mAbX/QsbjzD+H
dMuxi/kFcHU51QZUkGqlXno4qbHw10xmxtcTULpXS7ZDqnI7BK6cbHfA9F2zioYoRDuUnMz5dKVF
YXhe6SMP+W73VomomH/xeZpy/FeEV7hocYjVGLpPG9pMHpw0YuwM62WB+p2Y6VdlmxV4MHiV+cB0
QYL3ksgha9O6E7hJBUNJYfk8TQBlGBGLgsbpekE1qfA0LDv/WCl4vgc3pUpcB/eZ9d0aPRPbpAmj
OGcXXjxZbsKZL6lloUwqjmAjsa2SaeAxB3PM9YZbC1Ww+3n2XgzHdbQqnaZxQlEkygdoWzxUtYjP
5bjQLMow+hsYp6U3UFMwNWs10k+u2MAVHPsV6jYfY4DspORpfI8wfwM6yGimFin+2miKDNPXwsmH
04susVUMjGqvqQa1LOfAXIlHB1CMD1kOP+n+wHLKyObTLvjn0rVImL7SK5OgIfJYlYVQx1ehWxev
eos2yZBBE0Hm/gZW0h2tAswJmCWNLUXKxbolfVorbOC8IhOSvzMcDKmpbQirmwueOD9an6w0qNsF
e4se3VPwPUy3f/x1DhadbWB1JUAoXlAposZ0/RIjfiQggihTOQYjA3TJF0M99QeCOuU/ti1cZEq8
pueoiSElfHgapspnk7qjwSjyLtdr9lswVyvoCYISM1ILhZw2NakZScXtCZlYjlzeUaqjY1O3FgIW
KX4HWL5LLyEh15Pki5jNdID1mHyWGIKTqMmi1V+eH0ehjQT30e2mSzkurwKCjyn/PnkrgrlItoLe
fvNe+qOpCmpj8GSX8WERhI0Qe1BgRJvSjJvIbX/AHmm/80Fz2NgpLW3eMLv0w8aPI0d/SDS/abk2
TCYjew6Kl3vG3xD2v13fkFodEs1KEgqcRS+Fv5yA60CIQhXIdvuwvomebvzJkXAXpojmRzRXV+Wy
EeL20HBe2sfOOmmGj8wTi6lmEOvsk8yB4pNdwbsf6XWDKf8f4yu3JDiz6MVWp+vC/MYb4XPmcqVC
iZHxx+hl0YHN5a3xeHmrEJgFq/g941vv2ZR6cLRHMglhTDIBXtvQZeoqhAX16DeazvlD91fSkijC
vkNtsjiBU5nplebkx9nQCHC9p6x9VSszz23xKO3LjwUict2m7EU8a0GZ5qs1QebYnW57FHoj3dPL
sW96M2d920zrNZU87SsWcYYpyWzZuapZK003ez+dm6ewNHagNg9IAZH+KiycRLSeA+7h8eMlGY6T
+ylXFbg0rHlA6ovMSbZJtRQJHJbSSvyUP1ajenBDZ6VNSMsWhgnyLjjWt37eazaVRLjLG6543g1o
4LxhPAf+OVsCv+yxhAeaPcNj/CdxOX3bouvt6wFrJSG5ZOqXTLs+HM43u+B2SxtlbPWm5XNjYuBJ
AwsgTglm0/KVK9X+g8ioihRPVGRQP7AlCFbYEBBXxSgY6jVv7uKZ8LktA1wCiHZ5PConoaYEJ8w7
gY0FRv+0kiFLaO7AL3PxC4jEASu6zeZ1bTEVYGoizUO5yFcOFIXbjDdaOykeovej3jPsLo5EIh66
ymswWV4wLdmhjh1C0Zua/CXuov42aTU/s5DFgKit7m6umrR8GtFkVl/ueiFBJxPKKEUYFMyq/rhQ
CHMe+YqWtkkU5zDdGIfYjOlRKiOz6ERWffRGrO0SlHTNWpQQ1fCeoOsoqkiBZgiZKXU1TuEwI5fx
2OsxWX3W0k/NtTDXUeSbRyo6gApVrSx5V4jYC4PdI/2W1pZlG5TLiooO1OJW4uhi8FryBNw03d3F
JQ928B5LNXBtBM72PJw3Hm0plpjkvJ3yuYuS2tnRPpU/FPpIPO7zKfrDegseXtGbAVSrG6hFBG+n
C6Gh3vJ1Ek6gRF/yg34wjkwdBteZY9cHHgjKJRN42pt/keuKUsX1hwGfLyCA0zmdT0ZgmEKGgbDD
WYV2TAsEQBYrRtvH27gnHKhTgEWmm+Enr6T4bf/SjE/qasGX7CM6/Ht5UuZVcTr7rWsKgW4i4tLo
AYRqJ3aqDp2D7jc4AorDX3odi6PqiTVSCt5oc+7ptzKkUpCCj6WAQY6e7E/beyQrJ/25ayJqs/an
N3AXuR0ttE5jl5hmogeUfOmdB8N4FYqHYXYJ9lXSjRQhHCoTWJl7ZiogzvUyxGCub097VVzjZvVB
Y388pa/bXcd+PObEhNO2tAMhJnb2ksUAkJz9ohdD4eQ0WQJRvlo0rjCoSKznRSuzm5fBw2xnZXhc
4lIBi38qZvOQHkXHJ0/puvzlHZq3vUH91kXynZaqb3EiJjM08Oxe/M+sj/Z02iqciclHWt8k2Dbw
sPlqPcEKonqF8pcJ6vzo+4CM9w8Vfuz6rhuYAltDl7RD2J0YK/7pD7Dw3gaNP5rnfyywMgDx1xoJ
QU8jiQjkMC41ht5aKYPwZjoEL1XfrZHfLlrbrZx5np9eYUleyaSl7ZB3GfXQNScSfrjC0KKkqtD2
0LcZdN2iNRinCTjgLZ1NzxVKCLveH8pJGYLY/BWfICo67TCP4pUuuBkOI/X0rwvCeIJoTv17uWdf
9PipbWp6vhs91lYQsld+1AixYaWIdc1tG/4maP8JNQlq/dMN1StMpZ36PhmZKVGrK3z0x/4vuIDs
vD+wsjbIHH0wFMA0CQ77wGmodKxBfeES9a5qRcw8TE3iEDgWwDDMxVXbGowEo8plvhhrhRgdVgtP
IPUI0u9S4K+NUDnqjZDJg+ZvVF4SyhT0BQgPwIu/QfbRn96KUj5wWvfczvbe1ZsMVqw76jJViTqv
YnIzwTrjubjE8pJ5dTTTfrue7J9/rk21dp6i5SW7L9a3H0pnNzdsVsgt7H6YXpX18QsovSuCkihm
ZlWqynpNX+GQW8ZhM+u10TguTo7lyPnS9cLFOefV9kf4pxAXvESlD7vcD+Gl0BIwkBmNjq7S0p+v
rhNHzo9ItkQ3ZCVmOfW8jqQg73yRa28zv1SiCd2NJN2JxtDxf7Cv6bDS9vCTbCR7skxsi64N49VK
UCL3dDitmD18/p6Xkg1POaHmf0H5jAXveZKlkgewS1Hcnf0JkELsZrP0Z9drBTNikGzTHyr+gkJx
TfzY4sIi6nb9H5xdTELfO8c9oW39GDrwb/3nVUqCQT5PGh/Jq5fI2sMp9rZofwEI14BWknpndkkb
DZQ40D+nwlzB0M7iy0TnFuVbPASzP6BR3bdTQ4MsYPcElodcYLhaAeyCjvgSnpKiglz//yYflO+J
uRzynoq+hE8X9h8mqq8lLNLtFHwIa2IRCMARqvfK73ckWkeF7dlQz+uMyXTz0rU1XaDWpeFkxdBJ
l1CU6rPgUtaj+VAx9pqkv1oD/iIiJYZiEvdODbf4cF3oq2GKv4LSGb+Xe9m/xwuSNGrLSGHH87Gv
w6bY/6L4+MZH96NK3wOhgEXl3e+q6wLgJNYGMb4KUUjXHYdHKudXeNZ3N5yZgoqAHNlUmyCCsXJd
Sv5Ol3Tl3ycLdCNQYiT2Xx3YFHFWTSnenk3fD41JTjBNXwh5rY0k6Vn5TH7CdifyDgq7dXgJ3avh
tL0OfIP1UPEclDNkP8HQC8ogrkpO5WW3PEbXi2rFlchosHwwCCEHO4m91PDYTNv7eIdqPufPD8KS
f8+YdfBs/fHD/uDGVXB0uz9BhAHV/p+bFvHIP51Bd9owujgxj7ED8MLlQzLlXR9GKHofsHzTWuvn
Rl1ecMe34YJglHrmLTixhC7tbiRLS5u/51MElB66d0Uw3Hp0E7iE9LROkJ/zOuLSDz6Jg74IVdyA
1qSlMncvLolvUnKnV/SS6qC429HJkJe43Y7I/Uxg0T2oa3x08uxLYI1ME9rBCTByqzwzFk9d48d/
L+3frQf1b1nRdA9nCBIWuGYIAF1zcOIzy10SJ2FFtlqZ6nmw2PbX2SIOwU9p2SSgkpwvbFBZ/pGU
fEmED/5r+1/9kLmcSJRlDuJ7qXGlW+zjc6CGjT4oTQqrRTDzqBIHHPmZakJgrt/0aQGe/dceU4Bl
8gAhmY9rL9Wy9gUxeRDtUBWkOk8zKldCpf4e8gx52TB67k56SqqDuo0xsBD5mABWTGBGgrFs+wnA
PipSdSgZIHbbEaDCcSTXtkdE49cs6Rg3ENy2qn+DdWAMiIXElTq86+6V6m9PCaBYzI8uCuWrHxoJ
jQEX89jjIMP8vylCIheZLLVXHOZq5UJhfe0Nb3KhLgOx4v7apDBOnWDSucRXCxR2aYH07Q2eWAUC
1JUt/YX2Z53uJvo4qPXOaqrjjRURxijebjgBPZf7rLSrtHlznom50JxCHhH+ZjrRGFBjkRU3e9LG
lyJInf7Ael61x2FpZb880trP8Udsk+geDwbz1GVlf6RfJkJeBKgcUyXfIpEshDsmDut3NV9+vW7p
8qEGAiGbez9qcS0Ot7a8pjGd1XPX+vQQtLxdQYlr4P/f3DARnRlYmE2FvvhJQ1n8lklA0tfJfFQy
cfu4A8rAdvyFvUOXvXfBWprCk8XPdQbn/lIoM4avHi/cpkBLJaKO7m4S7XvrR8V3txd9nEI6e1F8
x94JKlxPv8236IHxqLRoGUOvf7fz+Zqn6xzeGr9cU1MycUnaOhzocnpY+iUVXLV/xat+RbLhR2mH
RF78+4Wov0A8le8btNyKbfulkoXGs+du2soCy1JOUbVCY2YR7PmcpRfjbC/qfK+wTk8yLQoJ2ygR
Ts1nvDxm2pILjbC6UI38ZZ5VxhZxVC6E4XwOUGJgDhJx+FbqLvNd2Up7qSOAq8mBASFHt8EhxQar
YJmOwiwr1B4zoIXSt1XU8bS54FCmUl+YxUjpOBbZ4BuNjG67GDuhW0V8hUcs9/Y79RptnCrbwgyU
e7NX4XeqfrR7Ol2QYn0W9FdUgURL2ne1ZJtm2tTfQ3nrZUeG9TLb/z3vYNI/0iIGq6hb56ZVqCqR
6pmUhLhgwmZPel7OVYymEPdssPZU24dVDSkzkqAAXMdkifzWjDczC7D5IwfjpcymcERfJbGL0A7R
yMzIRXX9lLbRudiNtnEVbKhJSG+4s6nq/Y+QsbUXKhQIvuoLUENbFdEORLvLvG5vOMKDrXM7nYux
HoYczNUf0RDWgxzAjcnSb5SpZI4k+fyqBK6zkgqsQeIfGKk7u80Ol70wOsXECVK7oMhGUgLjb6qM
Q5slLkh+MWWj95ldggCE1rVSTulGv7a96Un3VAjJUxEbn01ONKYjc89szevI7+s6wSPPgUFmF8ZV
UlcK9YEvY/YngJS2xAQvKCv3c6UhdEhKWxWdhfDSk6rD5u2MqfN2xmdg8Sbf5mN7Hp6pSQ4Q694F
ZfDGpge9m3avCMKlEydxqeH194K6Ug8ZIbCHY/FSbLGru1Da+c9lxyor3GsJExqrRQNZaAGpbFrM
E9gXJMqUBOAwp/qW85Ymd5WI6Gz4f5SELXb7ntcEQ5oW+myPHYxsTaY68YjybMXygpzuN0NxMFK3
0VNbtFP9fffUutZKRSPBy7N0d/hObLgJM9My5A3uJ3PudM9tOxUlEFW60By75CdefIjyEtVo7bi5
wi8OYNKdBS8ULG9WqG61ehPyBekSMNmwQexFdQItYrCgdCokAqhI8ET2zQzsevCsGHkNkyun3Ysj
DWLJ3M2LHtYvPns/nR82UWqpBVn4svoi6XxfDQetxv8V93iq9J3z0SHKN+zPRVGV8h6cO5fn9qMY
Qmksmce1JWDkXKMAYPYDfb6HVCZflpKHiN3OCFPxATQatzVvFTemTnTCUY/GxSnXNG+ctzAwo96X
PFNjqpnqntQA/e2M8mk/6EeUIjz2VpqFu6XLKNa9n3cAuns7i8bLLK9HHu+uGhNCOt6WppYLx1UJ
uvoApZgqR83KtEwCBxUm4hhC3Q0HJEdED01LbFUK/mbnPf1/iIObKaEVsl3pnoaq1IfkskQxSUbF
lGK231RBVR80icM6qdOg3ixU+57cLGhDW6Y+GzgdirLCKU8O/nEYRLgF0QDri6pl/byNlEJc/7i5
x9PRjwkkBGPeOHpz5OC1k9nlaah+0z6gtWuOwIn1D3MUw5ejSmG4LJ6wTIr+EUQCm8LJHHkJE58H
amquDRq/AI86L6mrkDt/AEcYh+E9XUo6/FOE5rilabaMVsX/GoX8pUGVBa0UnJAo/WZCi0dslGF/
Gdmn/nNZDkyzsJ7HXeynLwWmsw6XfEotlWMNC5PeEKS4hWGZ73MROl4d8hTqtiXwPMWY6ejVyVzS
RSKYXt81JMQJJIRHQAq/2m6RzmenKF8+Z1CQD6T2pXaR1ytRwZUMnKxec9l+vPMkNdCEQhCgAYYX
v2gYC2f1i/GIsTjtPGnNvcRRwKxxoVtNueaWEba2nC6iMA1/vq595gqNUl/323YgqUfXhAp1c4h9
K8HOcJyY2GqtdxGT9+B+QWXAFXzvov9ZNxtFMJBqR4qXkRdm3CfJNQzfRFyenZIRj9aWu5gLUv4c
9Cml0Vy74bDArTIXlQrtB5XwXx9uRX34+iKVRSXbkPfj6e7B+r5XSHsZSCI6m8jfvPb9ITViCKDG
nyH5vfN+8DuzknzWzty69Sux/7CYnJUMp/PoSRlp7pU0OvGC61UL9XELYQNPRT4ZPtRvPtiQf+9m
73GALF3c1UU4p2WL0pW7i+lAgmCpugvfpEqM7Fd1Cq9LR9xpoU83RB8G1LbwAD1aqu5jXYBo8Xrx
CKnUeu0Qfll8Mpy1f2hGXHMGkw4Bj1z24WJ8VGoQrtb+IgFM79za36dWiUKGijD5RCRvU9qILhkk
3a11f1/qpIzK+QCYSJxG3Z6TcmgBw6EnCxQknx3x5KOW0mEqC/Ts0ynipnQZVNXjI60HVxKVd2o6
c+lZ9yVKD9e4uRcY1Ccax1tAkEpYcyg+eiWEDNlhwUC8ZuGt0zDbTFN0LBsLuTU2T7YYJIzIawHg
f275oW3m7gENu2IzBRvEx/nWcnWpJLiI3RkNTRqybWUK9OzXlvOCObqjJ1jBwElyAg1FBzXHaaio
wPzQ7jDkC9qw59RyGgTK5inIuwEPSLLCuMUXXA5kwZWsCmmOHLo+YbuIgHtWuVNTjyJKHCQYnYLx
YmrRV27nWsR5r5D2hGMO2vEULQUCk3VjDCvtuksaxr12nU8E+5QHAwFfvL3fIfcqN016C6eoNjs+
fivHaUm5U8LMXezIvFZrVj4ly+GbayEVJtM6h+VKgL7yfi9ck42EAWt7hZigei4teb52s3klOSoe
FecpnX4PV1lbT0cMtphemyehD4TGcLoTDj7cNcPd3gTJ/JbTz6UZPPlby02U069LFhaa3E6jovES
MAK3D3EXlSjIRspFXPCk4yMaUJJs3WM7yuGTCiuEY/oBRDt6fqKq8/CzoOspS+vq6xCE+LiHYoNF
Vq2dNdkxV6aL9/LrNRFmSYCDxP3u92LXBKDaWS5tYdTOAsQPtEbDXALPw+mwt0IBCsbol9a/lWJI
0GdZQHzWejTI311GhRWd5r0oyD9ED/HrrU6H8o7sC0a1edSw4uI+GzqPg2x3BQC6OZFVZR0EAs65
aKpft8ULAJdYmdz8jcMCEwfBfltbMpZpsFWeh9qG/+CV8eJBxhkNppM4+b7AlkN/01Mw8Zx9mgUh
w0jYsp3NK6dN+esuzhmuKEUUky64JxQaPhFzfTyzMGW3OqFr6OMXj3DXA2Sf+CQLVZM4e+1xpMpH
DgVslLF9hReuD7NNEQXCWqGbeSUNZmHMhN90A+3sfLKiob6AAz0x2EN1JOeOhaHS9cwWk1nNg6is
WoQbXVOTJDEahn7DYSYubE18XOodqgjfj2YSVMvv7hYRBSQ9VCy3GT/zaX1C+calP6beq8SWzQee
9H1pzol5XZzqoMuvkG0x16gAMFQ27GEKilmRVczaIANVuK5gfJ0G/juXIBUg0OjhMpElCGyKbFaP
WgASPoQu/SCcc0P1weVlYKlVP0WTaTz11wHd/ffXRpUZo/IpYjNaFBKXF6FgnEWzXSYDz1CcjkP1
OcAklMq69sSHM7so9YhpNzcowVuFo8Ba/jO7B3I6SmP9eumW4cLykTrA6dRQwlC8bp0XiOHNeGuq
TWhKybtqdMZTBb6q3UPult81fhxWDEr0K4IGg21aq3TmVBCFDbJ2d6kxNjbD+b1q2PecwEA07vFR
EqpC16xmltdd/XBQtbBkDvovndSuxnxGpi2rbX0ID43EioyZZq+LMFIjs87Y0pL7M3XgUupyl0Py
RTgtYsAgk64S5k46Lc01vGXE51wmO6IrpTH2w3aLWKGTGH+OKjpLmb63Kc8EO6B1bF8F2GeqWjmX
VVnaXT50lgb3WBstHlzeJZKNfX9xwDrvWC4t7+jGp47jwyLY6YJtaWlZSsliwb6R64GFcWxFcoQh
sX4IbJlHRvBYbN0+2W6ayCkybqKxtG1A42itZ8fumH4crMYWWCmpTLK/qdnpfPbpW7cg6LxoriON
/3jlUKLohzPsKIs28ub6S9MeBeyf9x1+HZvp2l+p4j0HGm7zh4Q8fO3ffbb6GQoWKewB2o2Z/oqK
8HMt78aslfcS2UtN6kQl2RjYCeFidIHfdqOuwn8a99Np8Zvza7zYQCt41aePtcB2QeRJXx7W4zej
ncTVnToat6M6PYFjqxr0nSfvMaGmPvHUf/0xJLkhU0FN0qvJpizDW+3kqTe8aMc5uhMTy+CGCf/J
pHzX6vEtDeKu/dKq83o2vGX55QCO9lSZigWiN19TCUKeCbRXNiBmoTbUetTPwI1s/sFTgrzCerhR
KZY5zIV7NbBPUqRoq15ozkVPGH6FRVh9PfuJChr7gqvDIAKn/w3qiKXL0P2w9UnT0ZcaWslu1zNQ
8qSrj8vMHvqssK52LpY8NAGu14juYG9XOtzLIWT1ug4jBVi1dsFXm8Qi3NXdJIGfDyKy356+UnIV
h8C+YH8soDrcMbhp2BOguGrOobjropNnaIO5mhmQZsHGat9glG9bKHwuuPQEZgKbBTVmZ4YyyS5x
eFvxtUVKrY9RF90ckaDPWcGR1iwQjBTOvxgVPX/J8GmOpKAnDmI6pzNp9TjHwWkEZpNW4ACzZMhW
5Jo1U8KgeM4BSu2f5Y1zVaXqp97cetZEWpgCjmhaX8e7caXdpq21fbOsCpAuHAOnV1g2QLNa6FJq
+LUpfF1tFYFbH3p+ZzstW9xshVGdtwwjJBNLa/CLMav0Oc9OK1QC3a5uKpvH4SP2UAcqABQjNwSO
ky5G9hTMc7AVYtpgXz1U6gU6P/SK9JqM2i/4Cdfg28iVZXfY7DHGnzG2rd2kQYIeJ7BD91NxX/Ld
7QBHCVsuD2RpM7zdlxYDpqUV1OhVaCX+eVBdBfboo1jBVxt0/v5dPLj9hoKP2vaSCiEqqK1mQPpz
0R8rbfnk+DQjTfeACwYEya7RztcuBtYhqxW7FxQxKe8PawMZtNxR9jWUfasyOI+k9CeVaVPjZStP
VN8JzYD96Sl15UCTB7Bus8Yf2/NS998qm1xUHMNS5o3+2I7rMG84K32tICSdBHJxG5GsOlIOJS4y
XvhW73ep5cjD5TuFBxrp8+OHV6tmYKw/+wVQZOLqT6dvXD+O/eGuhbpyxgpmipqSpsC2eLcXxPlM
69Et0XdQ3pr/4kjsSTHyq4TZDTLv7ZZQK/mG/u9ddy1mvwdUBq52Hu0sgf/U7J4AmMeqjs3H8edL
r4PxHNr1sAMUNV39KeWMAKhXvNR6ZoUindWGRIpn6ei+TESmRImKa8NTTyE6fLD3UBLqo4ggseyX
jeRGLOj427oBR2hQ2qfLBRe5VaNIDnBOldRnrrlk9+1X21tIPyQKkpNbV5SZbpFQuprww0R8mxfP
2FjR5uu62fHMdZBklt1eB5kivpHZkbSzk/JkLEZ/Oqffw6X0bXZRkO8wcZZKl6SDbzLMgSxvzVv1
xl8F7Z5lpYFw9zYRetIq/ziOk61/iWBO71nKMfDvJQUvF8zFwUkJuK5vGcYA7rg8s3xm1gq+Fhp8
9dUyUbGHgaQ34cN9qBzVKQFg/lbJ10WuVutatWmC86/qF9oHBLcHkAcje7T7bRyb+qHx3L+pLUt+
Tk8j6zjnMp3XeBGrgUQ3O/ez0BaKMEjriq00kUAgCC5MJi/AMJHs52bzBT0YbZ1kPaXQOuWgj821
J4hDUcR894bKhvR1CI1tWcWVqnI6n9L843wYZkAIG7fOas6EgXj9Ie7HnSlAMDnwaHwnlKOFNYLF
2wnu8P38LABBeh4oe5NnUW5X0VHhc3EocNs24F/5wdQ+0wkqAK25Th3vhgj9OvTp+9BTDfC/vGA6
y5u7BcFRohMi4d3V72WoIPka6i8Sd8N/8IWM9WUjpCjuxgUWgoPq16fooEnTNdBVJlfb/jLD0brg
KNW7t9P01fy/8Bq/u3PRoxR2QkrOObw3RN0ypJFMjLC9AqBDPNh5h7UZOY3oOWQ+F24V+Gv8yKxJ
R86eID+CUe97uEnIa7AJyeog9kF0a6PcTYby4RS5CDpBxCCniA7vlnsGJQWmZK+Zl68G6Z2akMg5
N9bi8F3+XhapfzDLIgGx0MU8BLK466RWsJGMD/ne7Oyb2r19HmMpxMSOC91P0q77s5/X5LR6rwNg
h6BMJKvw+4zw94bihNPEeyGzdyKBAfPWaRZJjpo1h2etrEhM0nQv2YGRBeVYhkOCwFfrmfKxSCBg
Jr+veMQJk1NkgaoCXGoN4lodHTf2ezsG1i/OGr1ySNpiuSSfJKUUQ+ovlwn/kHrFeJbCS9bjfZV0
rRByKjkxB7hNxFxPyQVO8ViqkKJmCrPC7qhRC6zSvoQlGwCPVYteqnPI2I8RjHueIUFkCqB752z2
pRAgkScQ4A6TrenJ7HwfoVHSkS6XmmtqXoXEaRXF9Qfnz5ijHOVVilLOqfDhaTAstjhU9rSeQr+u
AzqBaFP6QGlnZK9GptTdS1NexHAcmpUrUoYfREv6WqXd9C1+0wnl/zi3BPal/x1AJr7NYKDTFe3R
q8vW1pxL55DWKyKBJ6kZNcrBDBTx7Xnt0pDtF1ACnfy0kc90PFLuJkMZQAuEOIQAMDaM/LesUMfu
y4YYzRXQ5KBgOsnFai65EFQjmoU+mbXUE+n0RM8Dkbv7JFVCuain67qZXZwI3Xr6WAKvNmVb1oLM
OLq1DNa1fU9ixpKHmlrV5iu5Ne95Dia1Ap2To+R2KuwRG3nYcH2VlzT9O4TnbUPjpe0brK6Ef1Is
vjUSLkbIZFA476GjPiqFQqewNkIPTbz+oPoPF9YHtV1lstiom+yuiOFaxBFLK3mvBa7ubOt9fMwy
jBwdHakuD91ULbPy9R6Uxz1w5U6h65ROgqHl2Cq5Mnz8OFZhOOp3E0ynxpo1hlmuXKijFaexSOow
A8WFiLcuTwdbmLiYzQQFqRKtYDmhmkYsYeF91eiC9cXqF189wZBL3FvI/a1mdqZRDkvr7KS6dbJG
eUudfxZky7SIwscOrzAEKhgK5v900F4BUFslt/yg2JMi3dkjYhHGEGNenupwUSvoerLkdgk+fbXm
Jqv2iXRo+MUUZD+PkGT+hJanvINKnn2ZsBZ/LjicyNr2xbYei4+nQS4L/HhAOwnrG6B9ETnppxLW
6L5KZdY0XyfGwsJN8vLFPsoeO3P5ZE0ngDSYj8aQv5E4eKGPKbLCaDQ5ZtnU282v5CZYg3jrWejK
2xbYIdApOc53RWkMs9GD5ZMVCvk5PScawW3Sw8dfusxtSNwSUfIXQ/LrDX1DBUqijbub4ce8HCni
p+GVZ3rH1FsGtzRbM+01A0+2VaMYmoxPPCmbsadI9VPRn+MgZubj9VrPTb2S/IQwe3rVXMFjvRXp
BeaepSmXDXNk361sCQvDgpZaXDkXH5ngvLJQVUvRRsjmwrbW5h1/ZxJg/DhfZdJESeytGEndsgN+
4PuNKbI5mPek+AsVnkpRTsTNygFazujXz42nNsANoMOHoHohr4NCJ5ymsb2dRYcvXPE5/0/mmLVQ
+eixg5B+Q7e/APWUug9KgTK6eZ/qC4wD2Qqpicu3BtWMrCZbuWiiA7EyKTN7cwms6dqjnDlBs00i
Yg8jPdVBZ3nPc/QhUPGcNvj30c5vGxY9Yc2mVZBRsGCF8BIlLk7QkjHeIKEKyf1M6eDAJ858urwz
3aVB4zlYD6YXsbRkKQau2hCcLyA1+15Wu5BH8D8HgKAKJ74N+oRgCjTBnA9dKeafUkTBJnlpTNXB
2S1LXaSXlF/8Hb8x2jZeuUERMxLEm9OUxKKiUtaJqUByNCv/sKjIQY3b0EWImBXnmpqxpSlxLUfT
/AByaK9h4ORxfFPbJEubYPrpUdO3DHY+OwhYcqVQS6/tSYCXz6Y4KC7NwGSOEtm7OPrP6Splx651
vz0QPanGmYSN9Mwzs46AUAQRSQmB95sSgXN1yL7MM+CU48hPIJsFAXvfEPu6TKVHyS0F1mLDDpy0
BBTdUhBFb2Xgb4NOdZfb75Jqn8yBW9ajkWLxZbTZxCN4nNMW2ikOWBuqFU4tVX0CWwkBRbzW7mkE
xAZSMsRVxYbifan5dx/kdRonsvYllkoN2qb5paDSXetHBf6lWAEDMUst+wwFqK++eIYftjSXnpa7
N+ubJaryPEgz4dUE9/SHh09KNO1jPgDsxCI9r07AiDNUShwiqt8+lIK3nMTjbwIVJmgWJONCHITB
6DPHvjAyc2ELjKsEHe2NmqTTQbpbGt8SAtmD2z0mjyI0Z2W+Lx4nMV3gEaY2tnH6+R93TVT/izIk
Tnw/AIgy7pX6UP2OaCscB+nSI9lvdaSENqGyu0RH7shw9XZiw7YMbrVu/A5N0abzky6v/Hq4c9BO
gaMzPP1UvkBX77/Y5kVOCkkUPwzi8qEVvKEShR19xc7roPimvRgya438+PPsFy2kUtHWsKYk7SJs
vU0WmnQ4GmLk7aPadDZxObgpNrNNely4XDSklO8mEx8cz7lgzUMC7KRtOT7fKLmxOQFFe5dXY24m
NyeVUJtV+TsqijbKCmUHPLb3T3A4HNYpy/T0ItkS1iawxwQPVs28pvIYo1uHgIzjwkSGwniEM31L
69ZWjtYxGnn0eiya4DGckcf+bOcs82ZL/NBzOM5QlBHLit/dWqc3b7ibYs+dGvHDvDC8j1SEMA6S
NcLXQOJ4V5LnXbt0i3NfiBPpPoxnAENCuC1BsHsAutpmwTB3zK7dnaMu2pR8kvHxooBsVAEcpMfG
DzBISJ9ywU1QjTBIvW0sgF5FGo3ziNLrxp3A3PjXDGka7vP4IGuFmh2cRLi8kHRdrOWVYxBUHlf0
1hyjUfUL/Kep1+qIqPF1PFFGvrcho4XLA/BIOZ3iObBJ81E1ABY7VswVD4J4sDTpycLeUN6quucC
lHEKZVhcmSMnb3yvABE9uwVFHWrG79y6Le2CE3cyPcVzrx1LVzKWVZOpeFJ/8P4Gsdb/hEdCbbJN
h1qsOkiegxUkd2DECSadKm3OVFoMiAJUN2VnAtxozTtbBbBceN2OuPu3aPCh8nCUvDiu/Fuf3d/4
lIQ2wL0hfEziLVonkm63coZvUx8VP0mOSu1TxGCUMuU6v48RySKrPb4oBomq3L9Qv7hyvtclwVEe
5PAmcOlg7BhIHbQWz5636oAoGnCz383/NbcYaHsUGzkvSzDBXOGWA4ZqALPMn62vFak8T0ImxunX
Lq1gDq1g1N24XpH1hsc3yLcUEyLRBNhXM9/+0wfUdZUvxXfv2iDDW4ilpVjPHgQ2Da2hGxAWNIS4
Ck76fVYGB5kJjoFBsYG6cgJiZw5EPTRD+dSL6c2xEpSBvelVG3ex87ag+HkseMddGTWkqTH9SnYB
qCskDBwcneytTXr6Jo/WjG2E/EB+66wakI8PXGBc12M+D1K1agTsmMDCHWdGe6XBCagAI/1E2UlR
K8WJe980bH4qVtELdQ7MKaQ4uB1CUL7YMhTY7KHF6KLo5snzEu9N4KKu8L74Vli8FAkoLmaib689
j43+IJvs7trjNt4CjVNSyvxMhBIZ6xBbpteOM+jeGcFW6TQPyuvilDaS04kziL6nS9HhllBAV5Az
fStvhW75UHHmoHzvGtscyx30+sLVjvsQJNdL9433je3fVpbipWD0uvmhXKi/OO5aou/pruEnBgyY
06FZcapKpd/UxC1Ij7HqnB38b6XcA4hYdX9XysNYeXKsOgtpcihUYRmDf2YWv5DViF1Dy1LJb8z1
6QlfmC35B6kgyLksnPm8eEtecQyfS8Egmg2/3D5Ke9q0jhr+cL+gteoCorObDiPjGrjpxY23Volr
axHjKkWW4hgufZFKyiCytpmST+BL1oEA/VL+p8VcqaaiaCQcnWsgBnyE23MNGgvtXEiyAC6tDyPa
ow391zmcYvra5RAwOtplGed9vi3a1HKSUpKHLLbcXUFHpDC2WnV4GCKdOAcziI3yqIAjqM+1zvfJ
jRsvpO2HzvPYi1itKicQ3Bf6Vzy+zYupAyJpF3Ka00nca4ZPcobrmhUC7QcYB5BEkyu8whZnIlz8
8rdN1zWWZ1VQLZzjtvfD3uAuZ6joPc8nRwswql2ZnjgsoqiqGsh/JI0Asjvu34a4oFkAS9+nzLqo
c6pMRCvw7cXoSjgQKBG3FRuTBTE4AN3ssJoT/EZ5P+JTaugjO2vZUx5h7t14rRbsNeBPvDFkGKSN
1v8dSNmX2BX7CHs8Y6x01BQz/ubrQ/bGVpEEcZix+foejHSbpEeXwJvgEJBcTZTsWLyTUy2mzh/4
5jSfSotxAu6STMkIVXUO+UC9oA+cN/AYulNobfwvmSnYhUgX9XGx7HDsCGyeVJGKaY0BIF7PMrVb
ZlwO6iTk/AMn0vrdfEDDIuuTSELzqJ1bgJAeSuOOnf6CRkVexzCSv/DfGuQFyxpL8+dccGM7I6TV
yIDqwBy58HjAMeMb624Qb9qyevC+fWZni1iDtxCMx6qmctfQ1Iu6Ep1Kke1K03ZOUJuhYXlYFoJk
7Lgwl9SJWl1XwD651G3T6Z/APAv6gOp8ZvjuwbSkIm31ZxI0p/DGazmRRDBYsunAYzd5AQTg6M/o
4O4Qr0NZzQkZnPAZA7Uw02s4NAhtb8iKe2uTzIzOWb1wvrU6TwA8Y2ax4MQOGtWQcX1vCzJkBobf
hYJWmy4uS9zda2LusOTyWF2BDyG8xuuv8QOjRtydFMxJqx3N5hX3WMyf84St7TXh6rhrZrwdRM+h
rgD7MlNmhTd25pgiVS5HLlDXBjdz4130LgKcw0Mu0+7LDH20wejziE8XdOU01I6vWqVak7tuTuxz
9KtNRWPggLQONAT/KZ/85zejAL2o3ZFctHmrRHozZALvvowB0ldypLHJg9gMcEX5/pQzma+pY2/6
tyU0VHCDvHFC+tZ8W42sNwn2leSuLDH35UYz7zlNpzfpfQTGEUpDnJhk9WK0wFEGM7TerSnr27oT
C8JitEYCtLYKHjYb9UeaPvEgHNljHDkA8zxPxAu3RFi9txpVW1bpiVU687Y1fSjHtPXFMtbApmZr
m1I4kd5WAhDvwuSXxxdKHD3ceJKDojWsoUhUuS2Sdf2jZr5ra2t+LO/jeWKNb9YtmdjZ32WCRSUZ
j5EBKKkMmZB9VEQR/OIXCaXyPJaRSys925N5Rw7wnCOhNPRbMQMcQDJlukOK7yrqf6eX+1/1vRpn
bMZYE1I+CqxT8oBa27NWmbemA6SkUmWMA97nSzHucKzSjq2Cuz8xKymyMoESP5V/eRGETQSyvwla
mG6Yo/Jm6j3bG31QaFsCMoqxU3JZNOOwrHvRXRJhKlDrOQ3sN6p1CaxXMUdq2SUe7H/uxLkPCxVp
3QbMK9ezfB8071gSkXk60xRxrfqI/9lxUlGuzXrC+SP9BK6qGLCm+glbHvKQFIqxqDE6v02ZiAXj
XfngtBojF54KLCQ7gxUYlTJKR4gwH2RMiBp0VHSLZQsg8gVRG99GFOYm1aqfU8eNrG15csNsIXl6
5LWh6eeJ88kigdmI/c8N5viulK0LxQeW099qR9ogqo4KQEE5ZYq4HTo3WkteUSYE45hFTchyK40/
KDvHaGpjMpnVkaMlRyqFpA5KPaRHZZe7Ir01J7FSv6+5eR+6zw2cYn5Pvv1e0ltMN6Na1E2svDof
1pZ5+cYQCkMy5ZV3PCHuJ0OKAJlQg6NtMwHyevgF06bEf8xXS7DoxvbrKtvLyZjYBH0YyxrAcjnK
xkx6kN4Ya30keju38rH1sIinK0+JOGqoa/uxchWRspwSMNRhcgz1h9v98Hzt9KH6WvV2C7oIFocu
nfTILkfK0pj7H2MVliMX1BnwIPr2+Ap//ZrEgA6/2fnLh1EHKIvrNgdlPQKPMAKk1m4uPiutGYQA
dFn9dbltu5o6S+djQXQ43ZGsr4HM3Z5JpVcV2EXyH0BrtfvcGZ6V4R3h85RhOPZCsY7ps+Lfz0no
r1tDaorl5Oa3Gop+HEMhEjrsVkuYeTTaB5eJL/ABXcM9Lme1YvWMPRbQJuuv9w4vF74rI7N/xeOB
DushlctX1VTX1Pqliqk8SHwr4ZMn8ySzWqQNO77+Hm6bVvY8710+ESsVjn4F0embAQx+XaY8/Xmv
sHiDTGUCWD3GIYOMH8QP+BpgmTP4MjQmAHRBPQ6PjXf2ApXuqjczB07OUxOAAVBjKxSAqastNUbO
tuz8aGlnZp8GhNGgKvUKH5YhS1gpVZ30OLiTybw9Zw/cqrL1slMa71nTOb86rrQtSsPx/woHV4Ip
mkDQaDqvGAJNLnXp3Pgq0tpFyOp65xx3CQPRYOpr3IE7RtieESf0jRTsCOIl2ZgNi+a/Nh5pqY6L
haHGq5qH5DiAnOiIfGc0zmeCThO4a4EL5Wj6f0pWlh7Pn94U0itI4HDLCPLWca6LDW9yJ2Cv9goE
TEqKIhAChKrajCJAsllaWnXAfDPAcXgU5/tc4lUBiLZBPParSWoMGTl1edYVOY8029EL5WvMWIor
n02po7zJKEPJEgAn/eaKQYsFMknht1iHQbSyqX+T2IMX7NujUS4XoEoTs7sf/jwsz4J9/vCvtERM
WRiZljMATOJpN9ZUZLyV9Fyl6NuC7tFmBhwoAwL9tnMMppRH2Nkgx2Uyef4qn1IMticUKCcdYcJT
SCYeG9tnWvMOMAJ9l2hn21faBCZQYFf5UFaynV4+qYgsiaR+kgz/sY+wJa7B9gROx/4Y4ZvW6bVt
ncP7nk6fT2CP+w7Ya9c8sUgIoOFimWpqr3+0zcoxyqERUNq8f+qxcmwRshAy9CssBW9U+PQQA3Py
7dQAyrAjyQqm5oVpJ13//685lSu/Qjd2qulvsjJiss9+qTYHSjgw3o+MD20YiEHz6vhiSjsCt4Jb
lOccsOAU9MfSJ6jquDrt4davz0ef/A95FbqeJ0hq707ADGmyWwt1p77h5xVVq6YAevLC//mxmfgA
rOyK47xY8VNlqnDTyNwd8+fFhuQgIDbE6NqPNTbV61dCthGGD75a88YD9mM9/jRaqnIDUf8q2iK1
2vU+zrMVTh6GLM2CSCltpPw1aVV0mhi3HCzT/JPwIGUM4G9vp8fEGyfiQlpjunWKYiiJauA8cA49
4xMFuzdd1g9FNJ/5wm4PKUVtZpCbEG6eBWFNPwVABsqq2U+qyjO0TXorts3HggCcgqtwJ36/9jSV
sy3xt/VtSSngGdnoiIEStKcIVnVc44XHqRU2RU3eC1NSVs29UMtDew0rrRDO+136oA//ov0Kg1X0
nt0pMnz+Utb1tmjiPTAKuwAp3l8Q6zzEEg+zbrNz7E0X850aQ/rR0JslBYheQDUTRNVpTvawjSCp
jGmZrpTY5Uf5HlYAzgsScVJ6Ju2fzYi2OrI8opwIhKLLykJu9z7r0eqhOxswVekmoVCB3uRq+aIA
bgvd1mMZmauigHn3Ce/Kg+DcbP4e5issSuZrUnIE21JkRCJzxaBwIs7a5URzzq+qDI5RsoCfpXz7
T2C4dO++X2dZd8MSgVVA4Bdt30HzY4udEb5SwWrXA0tJP77MICHdi5ejHe7NWHUGdvhKU/hRuJL9
HPz8SITmfTvvb/RR4QyBwuMkUoeQCxJ+aE6JLe47rsUnZ/uRp45lIMwFW4/i1zKhlEOwFrpz9llX
TMCyg3mwYveT7YHuZ9NJKpxS1ykGepJCj/eU8WCAogjwu3JFc/P5HnhInWkwI0/ja8crJIWrPY4i
ueQWsbwYOQtMOhLlZafCo4cqKQOB3cluKmQuxM8fQGvXL4tfDjrZOt9ddny3vtlwwtVp8Qn5S6PP
NYH2HWAiK79IMlsmD0V6X8IbkogttD51Z/KK9FExXspBEIHYpihmYXPIEqboxVBF4QnQuIl9FUVo
FCV3j9tu6mQYPfUSEm5EzUij1NtvvcAbHXRkZj4THyOE5IYEfQydt9Kh/vJP9iccelWAb0l60eJ9
l74zCbLUz8Au83M5I+gAVrTOjzb+kuNRHFkIO1DUn1G8aGiBqKP0eDjTqywqQ3Cm+MJdzhg4exdS
5yLXeMTiOvFvXxuF0yc22C9kmaPybt41HEhlnZT0sKWVlTEhUO2r13yjPL2bf/kNFw3XDhfy5gaE
urjUktcQ2aI/3g0gKlCIOyOnA60E3rIVlVXZiM4Vz5+ZEK8CzTRjhTs5MrKIv7d7odqyyLbCEnDs
hoRjd3QE5psBYxODLGW68zCB70+Tpl3lJNKiyZxrWJjjRrLuW7Cv7E1UtdW4tZ4OeX4nSvJGpmoN
LlgWTF3QzhRS35gKggeUXPIz0JNFFQbxgSQJdT5LQPV44csHm3TyXGJ/SOnBzlA5JuqzZ14WTNpa
/3MwgAA/cd2salwbh7y9woJsxWNgq57tRsSDDXMf11d62Do39IsxciiukRRRiFZLThLaLA0LKj6l
1u1ZX8d6SadhqseY7rDi/4o0dIMMC6/hW0H3ZHlHWCtolCzOJk5U5WyHrCtu6RXy+deDxax5AaSq
5Jdth9DxhkYNniKy54mlJ0d3m17DHCFT0gf06czS1/Q36F3d7JZLCqc0wOST+f0oH44rh8hPzHLX
rzAtlgrLE8h32yp8Gu0aY9toa2a7e8nDdYoHw2V1ADV4fqyfw70JA8uoqRXWHRYSdx79mhZyYor+
x/7mq8DHn3W0f+Ef6uNmfdtxz3wJY9C8bn57r9i0ymMDsJhAnerz9Xs1zKdMNpsbi6S1ivpDYfE/
OFZBKTUwonyN1m3JKNw++Ek6HEKx1SJ3yXg4PMYls5mNw4g94JA3Xk9/kv2oQZUfpOobifT4JC/W
YXD+Op8QIgb0CGEWqxr7DWr8jNUc6AKUGE8hx0GQzNoBp4FYWHj9iQU3ihmvb4l5K0olvWKW9L9d
EGJN+TzBIqXhS2wz9FPxSUydkyJ5Xrc08MMWh98ahCIs6WfWKMM80opvWgRIF85Q2sULBGGKVvqv
pnp4m9B9ExM1/DdrpLmuUoQHdnJzUGQ7285SUkfDNXoRpkeJ77VIk9bBXYtsl5G9MTRD8EK1eMmu
+7CEcpLibWCIUXsRoqhvaacffc4+TTP2I6l6E5/KhTPnmyTgER+MwoV45DXZeXWVEVRRuvCfzI9B
TDo25GlJWdM/Vj5qlxAb+Y2laMJ1oltD4tJeTrMTqCzvDde40Vksgvzh0PuuOQyYe52uXpO/2xTU
lWyUFdwAOafS4ewqvk9bg2wgkevsu6ol7SxnG+nMGudwjdVPSJtDyZphFdHxW7wiH3jwj9zW3aim
SaJIiOPWwy7IuO6Fk31ex3JEHQjhlgG4tQXfanii89KZAGNTdVyHjn/cdL1WCC+DpqXT6ih8vlQy
Yt+yLJYXXvlT/Kq3X/6ONbUxJ3Q/nmbLmzKZwNq5KA9E7bI1tSEvEefuAUSoxoy5m0LHVmhngB90
WEWFecNDx1nx+tEI+oZQUPPp5CTujnB6u+ySu0SEDRUgiAJFBo6V7QNI89UZSmT/rgJolnrMn9p/
EzWPhgmL39iYgHX1aqcxCLhpu1FX8DRLQ3uQwdqZNTXgYn0vMNHFaGwzAv5LTnUzXt+bZ8Y95z3i
zlOU6zvTPzAPOr9bEGeFVQGGLLF/VoEjO2L1yzGDlJoi8YYbmLwFqiYU/+zVmX/wwBAWYbKeWxvB
aq0SuopMYKsgd2nkk7Tjd6r4aC3exABprDIlOZfEX98btiB4FDvffpfDdyhTzrI2uXQBsdjDP1PI
NpKNP/j9RMH7b1e2XMUE05F9VK6Q4pfLvwyUZVv3u7S1+KoLXa/9lekqUeri6Qnmv1nAWn6rzxCK
2xx4igjaAhpK1kJSvy2L2vBXH+E+k9VGnWcUnqbtbkIJAXSCfPgv+BG7MFYMHtI+TrL5vftqYpUv
Qt5P4c1nEwCTVzyQ8NT+WVg5iocnZ+Bq2RGnBfOrYG9yNu0/wS+8erIiG41j1Va+SM7U1MzZcPss
TM+cEXuVsBfunOOIpJQuGGsUqlh8+yFZsWnvPfSoRW7B6giKdyDPd25q1s+TTR1jIcIsMcFB/WQm
DhHH3qQTZ36N6Todt/uuDf8vsQUi3AMSgZyeZQTmxffD00fO4FXqJEQNWbJeFpuMANaXzV7IXxOv
A55G4pqI0PbNpxXWHOu+VkGycMJhiapxQwQf8z9dk8doFZjf6EIvCvgIJg6sciJNLO3V3x4g5m8/
G0ubdcieqydclnvBiWjjXjvJToHTlOs2TL/jaQKfe5bOko5SVxjhxPqS8+c04d/Of4xHGAYyGIfz
wxF4yGU9EZERzLMAba90qJJTGnIK+GALioNZPAfPGrlXhEccUWuclUMROiayM9TQLIQFaQ+pAxfJ
uX5qReXrJ4Y4XdKcYsnoEAi9OCKmgTDgLrLNp93jrK34aK9tnCC4F2XH/pQ6PjCkdRNRI2NIYHG5
iBYmrnfjq3yvpV/LvaRhdHUlSEUZbUYrqGnx9A2TKDn87SAm6sXQZ70kFd+tv2Cg/t1BQU8h9pZR
iErleSxkZ3jLDjlwDofiJccms1XqdComgppHgvtXg6ClVlm7ByFef+7h/HwZvIeQt3pogbn48Xwi
xkE3CsuzkBX61l4plMXGTdhuh4dlOaPjaSNh+H1JfWCG7udppY4QQcJpK1hCqBniUC/83G2JIl6y
FrfA+aWzA+OvhPXuN6Cl5qast2Pw+SjpKPMedrTy62r+fmMFq7Gocs2ILoxinTGdYtMZRr/ql6jI
3oOterQsg4dBcKnLbYD+zB+0rK4ycq+gvzvmzRaZ5JeCW0goZwFzGbaQB45h93mI8d4Pp6RYWf1D
mFqBmBwkbgAxRzhWlP2vQZFJk6j233hrPfMve7FNOFA9UlL9ne6pMpuO1bCXag7IzN+KImcIGVkt
4hcI5PSAScgusK/st3klGjGBUb4i8eRMTcYoxhdcCu54YEDOsxBp31nwyXwqucQRSbhdQMqF+y//
EYlAWVjm32fO/T6hSNsbZEr8KcrmugnlgkP896gxWvCFAdixZq1Qppedd2Jn9An2yvqGEhazpSWl
5UPIGnCQnWq1GvfL9ovBz3KTRjF9GLt/q1JxbLSAMbuAU9iMNxljkIH9SYZNnnDqwXUeoh7xhqP/
QgtHxNkqVVNSKbwKM7clo63IzJ71wtNA3+tZKYQR2KNbOPWmSaVmNJBE6X68qrrjtOo7WuodU2dV
46UlAp2UlZPZU59edaHOeR7a/sIGVZswH3mm6E9tGficXp/6xq/hs6v9zQVpQpda/8Zr0T8AxFj8
MDIDBemRKfQhyzTmul6K/DIV6ffKrOHmVQ8XUnjk95TQ9F/2Zonx6TvuK0+I5OmbRvvNzuLjkN/p
PvISS0rZQQEms9/x8t7wx9JeKVfLctize2zKZ3IqQ3zehK3iWwIK5Y9GJxXlQwLxQAXpfodkOZ9e
46+JjQdo2Q7Pt9PkECAhosbH8nmygadY6qyKhZUsRJmrugS8ya1hUc883frRT9wUQvoKa3GESmPi
z1dZQ2acRNaKf8YVesAc94yzv8EPSfujbEDx4dk0CFbRDj+PVbXPxbDwadVPQXQomU8Uv8PJL7Xm
cq1tfCTuViH8fbjnaEQtg9FkEqW1Ptve2KTedejO9aXm1PAp+ETsfNc5mpmB44kFyi6zirMQB9tt
DCIELJl9bq3a1be5uNM8PF3poJO2zNwtCuDjxPpJpljf9eSav7VrP19MXtaFnQdox40jugVfEpj3
Ho5cQjv87OJ1swQKU41ZDLliActdJwdojRRL3Oh8XD2ZoY327sLn9G6zJhQTtxwXXsiPHqepsP/5
hEqavB1TxLHFTJLkg7md0PEjlvXY9Qu9ks0WSUXrID4l7iB/l5+CQ8B5D0x401mXpC1dASfuc4q4
8RNwKoUXUOiSr2BkB0mP2XfkxESPcO2qHSR0LCtmyp2wEQdszUEYV8tCef4cyLjpVFulllGWaLrZ
hwscwqUVeP5kbekOm2Lw+YynjmvFNlnXp4AIhULZj6B6kTRtn+8rbcptfHeAuQ2b5ob/iNuJ3VwF
A5x+oRONvI8WdhrmWB/5eqj81SQeye2aEYJixrSIVSuBYd2SHmJVnpqwzC+mLMJCTCLrVJQqbXa1
tew1opdoQteQyc5sSVGdGIhpsPGYzX0uB7EHilxRCiIFjbKgmAgJW+OtiWu9kINVnUAt8cHN3Cgb
e4sO936kG8SZRJ+MxSzLkBIl9WicIvXkh03wiOpI8pbOx1JbMiDVPL2R2NWPNyJs3hPTKtZekqFl
gIRzBgCrbVCht4Aa8gLzdGMudKs9kpShp4jLNjMvDAuTFE7aETfSvyFqBFnoQhB3pNZwnSIPKvT1
RQ+EpEgSfBtchl9PWg+/FSz+NLT6w3EFFJgD2WOMFpKQhuK5J4wJYXmpTVV8wt3InX5YZ6ZN7PPL
UuV3LS2Zlhhx+3KN902W2z+OF2RWx90yEvx84Xg1yaZaF3tLXUzUjr7b6mxNic+rGztlDFKZelI9
LvRhyYRel0T+0dnnNUIHdxed65swwwJPKJ4SlKiApQk2XgwQ3sxz65uUsaCny3gjTb+0Us0xKYYo
zk0N+sJ2MnxDBMsO+RGU06M6zvze7csBZk1hO+06GgR3pmHyRYtOMX4Lfbo+TQH7azM5j1P300Op
2W5NL7fsNZiWA+xGb0smf2FWFEUnGZFcb9pNb0JenP0/JM+MGZAwIXqpg5TRT7uvbu80AWrTrmXl
p79BfDnktzlmSAaTkAvsOOQcWY85OGdCRcg5EU5Tz/jY1a0gedHsNS+PSCtmkI9ztW63n2DOhveU
54rKgEj7tQkb7M1fHEs99wb+Q7Elz5lISG7Fh+UfbdbZ2civJmR3lP9R0nnTUv7KsnOWVpcf5o58
gZyB3eANZ9txY2sTf4Kkz66x86LCS3xphKt9nX6DRTsxN17JhKVbhDQhMnMGYTD6RcaSoVoCV+qL
cBsC8XHhkMXx6/FsFHMAOBn9iwF+36PLD+OUcAeoX4cHpoPadm2HMJ1kHHRF8WVZDxE8E7jXe++r
iciK567X6GKrvSi7fGBs7RZNW+2KMsHnTkCJWFRegIGGdDS7My4KVU4vGlbB74il+FC6/wS3jW7+
KtRNDJsZkyeGLyru/a3WR66YovfRHbEnuZQPj5CkaotE6l7Z2+w9KtlcOflfTx6zJjLOHDtg7FkJ
0fEdk5MuLrdgSkW74Tyqd80XM+hTZyIn7RkuGGdwiwRlzUAHZ9zjuLPUyXhciH7HskMIRyOaq+Pc
Db3q4IMT0guZiROUxI9l2MdDVGjmS/J1wKy/2+DfsHhZ/owy6WL36jnOBIckvdLbE+FWR545F7sn
0RDL+b75aySnNvMob6rzys+y/79aSS/4Cdhq4s5p++Q3YjALGADcq54hRt68vLzHW/PEBlJqjsYW
Yf0uw1HeAzQZs4Bi1ncxbagPL8gQJXOyDGGi5dnZVZlVdqclbmsXswqGbMhHxujnVBi1IimOJzYA
u8tSXo5xMZHAHr+3jEN1TX5GpPcGg20bzUAKx5xAkyFkpx5uYOwF2+vIQ2cDsBR1UsbuCYIL0R8s
/t4oFLYnjQOESB4KRLmfkMxgA9Sz4VPTcoSDEXqH8FK3A3LHuvfd9D2PW+LVlKb+e1hw3Dky79xX
YOFCxK4gCqwU5OKgMI3jNwF5ri/mFfypE5srmaIyE/Yqv0lJvQJs4kyANpDmauuM34x6ycRuzff8
bsULt/VYFj1jsIrHEWKYShFmGob4J6YDSSe0CV6ee9VljDaXFj6/b4YE1O8KfdHMP20283LALw2d
2TSPfLF8nyZhT/fNFEG5wGJKbt4PlcQQnG0TlpM187pnWyYhVZYKuXtCTd/0KgebWcpDZMTWMa4B
rAydxbGTEcxU9jISHEc1EV7OdYsIes+ldvhxhfwZosX6GA3W7DeioWS4N6FMexLH6ousLZ3Gt8JN
SgmTs3zTSBJbTf+mJjcyTIR93uKjHSCp2bnAlAikAlXyqDGF5lkyt1UJ+Z9eGyye1N6G9pNaG8UY
GJD3OBqao3RjRKkipWt+RUKqFCnwsKTEygZQq7i4BsSnTbOE/rKrekgvDu+ZEr8ygOL7T7bVXyc6
yn5JQfBqM7Wwnotx9jj9CKIT1tVMELn9KhGSNYEej2Ws3A0iXSDOdISzcCcMTr/ixzW77SsST0TE
Hekqu/SRV4B16jVOteqCu9n4GbD6zqmlFiH/JPPok+1v9NVHWgiibowHeTQI3hXDUzcnlREh4j25
nbZbJX4q2MRb3JG5qQyymawp8DB9IN7thXU+RFfZ0GnFCU716i4NwN16neidAEvXDrIfrU7wBk2a
FFKdN4U5Y8A2tLBEf8ibVo5oK3AgRWQ24p8t+/h7pBkS2d9ecz4JtK4ZkEZaQQ8yGnQ/u69S+YKo
eiozmOGHt+MqIe+UFTt9jnM6Er1VPbvQz6WOXho2jqc0q74PO3fs49/ycjJhc3ZyySwjD6X/INSE
rySm4r1N/TvqIS91EbTGP9wcJY9VXTV0s8HVFN+wqXEcMc9QzrKBYqqPRxNkD1R7OsMG6AKaGJp5
B+MguVP8D+qe56kRs7VMVmSg+SS3V/NjtTUdlLwPDs/JXlu4U6iy1DLetzH5kjre4p/uG0HrDNyw
0gD+M3hmu7f0oEcberxojregEpXwBIzCniTxv6wIqt/AmmaNNqTsQAufBRFuTXjkIuRBWNVrHvjA
KcBvMkBzdUf3ovkhrJ8PsuEiOUwJEvJJBYKcwMr+W6H9o9S/Md45IsrBZsU9LtkQjprpxO6JFKgg
2s6r3+EHiRaZL+W9HW72GtQGu9jHC5GDJK4gnKSAVMEbHSx29/5ikqTxDZx0Eoe9Ci54HL9x8wPi
P0pr8TFO0AcQX14MscZJq5N3+JtLJBbTWN0pRy49nsaIBNPpUY0ewDcCnCmnIletgoaRy6zAxWOD
lJq5gO/rIX9kVrSdTg5RI5jQPHMSiLl4hIDgWBIjg3zhr+hYqBQisvkFzRu+bBq/qWDFzeJh2pK2
8/ZOk6T/AQXhdIJRIezIfawY5ROqXoP+kxdjFk3IPNsSwBPHNPifM8Dj661+qaAyuTEilvRMxxz4
+yTzCfOn4iw1c/gvYJphOGOnluwCIVaM+6zHj5LaRrm9E8h8PK7QPmD6Dgk3Paf9sz2G8USxrP7i
xuNRa9nh+p6glFuWl1yAqcX+++JWYlJy1x62+94SGhuDaEE933KCptPMFp73bFjd24Suj+qHoSFw
eKqw9r3/OsDDtL/cjYR75ZVHNwTk0x73lqDXSrHnpjDkFjPKY8j0gvVFrWRXroa1fsLT1FIki2K6
hUsZKfpw/0J+IDZvoM1yYthHYA+K+f8dkb/JG2d8uElbTzG047Z6/ssY48mHg/zY5wMJnmKvWI3N
1WF9ETqYhRneTYwHD3C5Bgd6A6Y/k3tA6+sLlHEvjaRIkonFj1v8LEs0K2a+bYpBEHfDAFhMv1rK
IqEWQR0H1EeEuuUXeK30y2/xTq2dZTMAoFGn/XuNnktlcqCHEelMqyCrb0hrPXH9PG8N8mBZXo89
vi/RZmDeogI1L43lYnA9WmM+X7aCaE+wQdpsh5Z9Nc+/Jre5lr1Y5bnCfp4VQhqitXCeyLIcJrpA
PQoqStOHxSF2UXXPvNaG2LdI6UrqXlYST681bpwsRe+50Ehc2gLWI3m3HZQ86E0BZcj0iEJpNfcU
OQqVa0mxGiHmAaCZjPEWRK25BEx19wYEz/j8vtQhOso7spSjq4/qeB+3gZz1L2yHabon2xa7s4eY
Qnhao+smwB8qtPITmcS93nytKOpICrLWVPpnxELLtLCzSBjcybT4gS64uLS5YLhD/gOPPXw1P5ic
iozqzaMXEdIlGMMc0+X6Pb3FhPFPpZY9CpG26czXp08eTB0PieQLPCWFf4sT4ylL5Q9/m2Hk4MC4
nQbR7oe50X7C+fK7lSTCZlCAPE3BIkp2Wb5dt4YxwUzs2f6ondrnUa3CZQIrsh+t8Zc1gUv6SJdB
DK0Ae4Oc2ddnEH4R5a+g5kwdxjBlepHnudIzYCSNCRBU4xZeQy3NQhT0T3h746wWXyCmEmFvo2t8
4pSe5LIWyYaslMxxOBYpry3gag9zJCbw3fmye5FEmHPD+YNTFOYGc8zUyPRJ9BqVDs15bspf3Kxs
z/7ZgMTQEAuzaaBrwGUq/ODPItCa7fFgqnL7TVbqkm3anckigRPdrlGgYAeO7vnwNgMvVl+Zr9Pn
QWGTkiE5QGNX+fS1VNpRKcx4ZMkkljxa0RsA3IUkf0xAjF7TBQ3vdkT2xvi5+ZgBrzyyYNAvctyA
2vxCA2k9oti+Rjux0w4bVCQ4+p8NdAZz06XvIhzmMVfbIbnmqMO/jcLbKtuAoVm0DCZ5+jXlqfqj
RG2RMQNXMiJNCC5OdxWTdl4iCXNx10UJDUM13fKLOpqQbHK8iTo5jEAYsvbBDKw4wxFAHj30Qei1
92PQ7xB1S+62ebIHWe454XffJggyKQRzle7uf3WvqODusyJYXWFEM/1D+QJp3egPkxptArpHsMHa
zVsWd7FDxWgTjqHqGYu/A5GI9iPko+Jx3x0DbAAKL1Etda+RrvhPuQeMYXPrqbcn4S3npjfBMgjK
MhgibYpvDXhwrPFb/z5d+R9sLJBwmSQjJaI9qg2BJQDKZjnGjxLlSgEoG1XxURbHotS1ry0N80f8
MVTZd3Yrhpe2qtyVzI/VSVH8JH9lGLKgN+yfLyYE9iMd66LHKJbwimXWHI517NAv1MdAI3nkUYZu
5o/1jfKLSPUQH6gn75revwqB2XQ7yr1Fn3JvOEFEN+c3BOg8KLRGJ78/tk80ab7Z9sTz+WiRQ4Vc
001LPy+eJ+7jP4EP3Z6h6pOjAbh71OYl0NDWAiAi+9JKCbMrJxskD20503lkR3wyFenXSYEgg6nD
YOil++S/uw6aX0hlg3QY249Qzv3p+inEOSXHSXyyrvr8LT6fVmugUrqG+LMLkBquLzfZWJMd1Ujn
M9434ZfkceIiEu47A4lH3/CoyI21T5VgocusdxcKgoHCgs9xJvIy4hZmJPnJuYDc3D+2JO5L1kO9
qrux6/4apDLkXURiprK5NBzR89m9Yvcmnu0/c/04IwBWmW0BDcxSTyQWtiyvmR0FTsdFyCJptwJ8
+zRz57s08txYTJscqa1GsSsQBzETJ8/YvY7meT8hCRkQVhmFqk8DUVaNQqc6m2p2TixzeXxLXSBK
tcu06Vb+6Bq4OBrbJpVTh3RRAdxBXo/xfBhFkhQY3q34j/PzOizp9gTS+N18oy3eXPFw/FInfvmY
58hfwfSMRu7U6MCMz61KBtx3rtREMRT7qa9pQNynyr9LIVqPbLRl+XTueNLTQTV9pPsI4ZEdt3+D
LAtihHC1V9rFT8kxhM5/xYNcrezRsapbr3BE8wNhwjAoYVFJfXPpSOEbJQtzCVzQJ6kVTAYI+JCd
p31z6Khby1CkYzyktK/PlRNf3uwpT9W5cc+Cf00oVYBX+kOCJjZwqHXRP5VXf8qzdUDV3n9YMqS2
PehKhDJ6HvC1EzPCg+40ieEr1SFXcBRKG8iEVTUyind7YilznOs/9ti6VS1UDfK/hTw5AFUz3RVE
RKQbg0cBu2svBbWPMsMhwNS4PkP/KKs9AqVXXYQ3RiLBEUKzKKtXxXPCKZswC1fZesaFu3lXsIa4
9YtskN+rM3lTUonOH/kHD7XbAH3RdubZ0VLt99SZ8qDuX+xJqXm9HFWVvXc3sk+muusQAg7rq2EI
0oFxeT6VlcZ+qRPLI9G4VqKqkE85NiNJWs+T1cgwcrC13uTqd37+S3oGL0u8Cq/8i+PGrxVl8xh6
qRLBq4WgaS0ssJiXSxg9MMgDVJHGYCvbyKzguGIRmO8KLO8172rbiXbHwWb/odoiRxeqjX/K1gea
wPcoYtBUw9w3iuYF5LqkNe7bWEop3A1DLBpHc8+IQtN85rKsV9QEl82yFJTVtE6JYMYqlA8Cieu6
S2of0Vd2CY/C1DPGi0OUAs1V468uywyZLs4llLiwdbq76iww+FYTw9pPqQDgZt32gIbmEAxigbmQ
nJ1djRf7yKJScrrHiWY2pMBPvzILY+w+KhD2C2T85L6MJQS5vRExuZ9DxQ/EqfD7fqlwokrWUZI1
khNdJdyTtwmfehtnTHbCH89KfJIqfjX05WFdp+W5b/wYF4kbjyp3oZgp8gV8LkhzNHSWIHwX/th4
hZkcdK9henpfB4zo0LePYPcc7yGglWYeyqAmZ/kZQ6UTK4fuhedgzec+2I6MFjet+I8QVf/77aEI
LBU+x7k0alv7Q4/UJo38vBwc/BZby811YOnR0XFWGShPpWoLGypNRIksqhz+GhiEfgphgjlRmY00
yUaCouLrJtFsIEgHM5rYrFmtCh/MxI3MkbPYa6ptqKSAT/h26bu0qhXKfSHSgJzWToozlitRBIEj
2pBAc1OaDlU62kCvLTZNS2xwZqKODVTHvDh6qPCT/cWCLM2L3M0U4tNCsvqBzgSs6Twrq1rXhDwQ
RqfhZFDGzLlahZxfgNxXkRhTd1m4wpntQ9oVxandojJMfRM6PpeiC6Ca4VZ7CR/s437r6NEdb7DA
/f7Y+njOXu2DtjiKwiyaf+k2y1ycpqJwuZuD27PVXmdfZWHwX5hgUkpZSK0fyyRZ8uzDFt551Lj8
QUclEuKjJq6Nut3Pw3DDSzM2obLNqtyrEwCmZsrrw+vsbjHJYbQzCJuNFBucIOrdvKn5l6uiIx0k
j9SC/gDn0RUjBUYfnVd1CZ28DKaTgo1XFyZz2DWDUHaWsFtfw1oxxG9JTsTXvs07gAo6cA91+8D1
UxTK77LQ8OgZ0NWPNsIe81lhLZo75kqYRaABQ/TaK3DI0lIPZhKZ2/XIpCR4g6yus617YhuLMUYS
kxaM1ZMnNKl3trNEJApJtV4ShecuVXqkhM/W9BVquAJm0ETRJ4ZDOf5W9PTC0S/5Yk15WzGnksIZ
HiDhoe8sGBoQ+4yNObp7gfUuJX3OGQzsksiSjM7qutdVUlpVZioHVZTFRb68EyzSxFiI2W4J6jW8
gdC42SXiX4JjHatSBPudRtZITvNceXtxsM9rnbRowm245+26K849UDybRyWjf8mT5h9RpR0l96tP
3KiGy4o0OYmKycSmbV+b/Wd7YaDg2oCdHTuLBbmbHKC9wKNMrwOmoVGVG99XBNm4r0c1dAeM7njX
f7zd2MWvS7o2xQ/h/3DkyNB8EulyPwVxuZYLx2/2OlqJnX7VxhKCRIGKhbdvjpUxm+0jCKyB7qRs
llETAMF6WsjRT0/1Qa3ocBvPTTUTUUilinplVyR0hib0OhH2+efq8ay0NJi3FkyT76Ey0Yk3RumI
SQlxDf4qYGTz4LGN4u6HcZ+Zb+5DciHJWYzWpKmih0b0lKsIULBiovyzgW4tix3+vhN7/dhUxB1G
IPhsq13jiMlOmo5mspz47n5SEe2ioomyB6TTBWWdz4nLYYGS4OwV1sUyr+rcMqqKXCpXfLpcNU3e
w0ID095d8kAdfzF0tfMRAvbKZwGyywQrM8I/rtLwHOuOPVIzZd6KwGszQila1QDhGkuSnhGQTUCw
LenhI74hAMXrL7sox2aFM5Z0uFDhNJh+NanQvHYNb4tf+c+O75YCUPRXTkHhX88xJHnDG8OqfLHz
Gb18hT2L17u2kTKggxZLSlCEVso2/reBvIdfwQUFy6rjWZkt8FmZXZvebTiprE+F8sqd2r+EdL8R
FUuLYzqOFlsbXJkqFd2ONlZvFeOIZpeYmkVqMwUuy3H45BcFsOTueom/oywsXKdm7xtoX8c6nWGF
hNi9+JVmxhGa5kbRVQf6BWIgRUjD3/j4m0FRF1gq2n1dE8cK4VnNaIxnod3h0G6OPv4ib3rlkGUT
5CLDGd72Ior3XhEV96jF3dDur7ehxURnXWitBh/jFWGtXk7kf5lYfcDf6DcgTsg3pcaS7IoMSVa7
UvRYBvg9NGGsexuIj6+yrvGRE1Nna35zElb46JmF+VQ7418lxAfxmy2HhVG9l+j48Pziui9uNZu1
+J3BfGQl4/HByNMBVgn/LtpQcQ45LxVwsOxKh91RcSbyW+dBdU5y3junQcAQiCyGyvwVXI0EiCg1
UGoh1otdVaxXlmGJTpX4QcRRux7v9RZV4vNaODtf/gpSHRlAT1y40iVkyg8Xcchp1jkK5YjWcdNp
D7ofWfwq5RNMoyv+Aze09f7S3t1Xwf5dGz1PeGik4V+wIfD0N/+icDCznoiTRo7mnz+IocW+V5p8
zLM2biruIyfdIy2TbG0WTMZ1g463aVvnTUSOcMFsQhXQpo72aHuLJQQ+T7B7gpGR4/vltO2jjIoI
pmbl9hPegBfVoZMPoxq/PDiar6sP4CVjDr0PwtJCcocNS7EFPFfhK2NRObg+FW6+goLijUMAgs81
FClNbsd1sJT8qzRSKD4kSniJ0nYciavhk58qq+1lkkbmcePUr+lEw7/v0qt+e/4BMN+xBoLMkBJH
wHyyfSduBEjiJAi7ok99gJ4Jy7LvCUKiGumWuKi8WBjZasFaQW5VWqjYzjq1RkHD0KPYq/iVcSl/
yLwuXV00P8v0bz5VepylnUVyhWXvYylj5crwD7vDEid5L8ssNidi2x4Q/Ra/KGqc0Q+yGQTBHRKv
obyHOWT2speUAbBIDXiemM31IU8VfZNY5nxWerpnCDXthw8kTZZT9aTmAxXCpsO8q4q5WcTu3WZb
CzHhI0mFmVnddfCHZksc1W1Ew0uYjeEECLnEfgXnpZLQME0r5cJfqrFyl3yVz2FHcrdxZiz5wwm8
9vL5jwwwcrMqNQYdYg7aFbgmR47LdROBnyU9cWW8HV45ZikApOMwfYMMs8sh7kYsUpDHeSwLOwk4
K+5iG+qRjXHdI8MMGAmAxyeOu45azlcrPLfHBYz6yo03GfY456ylkwIkM/27aPjOWXEg37q5VyBr
sM47iqvRXX3yLfWml1m00n37aSXGPA7icoWoSN6VMnPZ4+if6WCq6THtsze/JHSyB3LHkafgFs+9
SDhtf6VtbI9uSv0BkLZOCETErzgqLYuPMHk/T+Zp2EWx+nwPP7g69jGrbTKf5GXqr/Bj/L4fRvUJ
V0ytN1jOcUEzmDSLLGeEFQAP65wSzxWtz3kD/Seyr/jPj9iNx/n7Ilkn6KoLtHrVbK5MnSyZswZH
YehNV+/E9Sq0LXN4om1cXA0XcXhM4GkqGepxpxyrL0cq8RTfi4kX6wwaBPDaLU4vll9Zzy1qF8d/
5QhBCGVmmuOZAwnZy/VIWGxvCgEaGhc6ecdEN1hma3cDXx+XesmTxH5FLPFo6Ykd3upKM1j5RMLi
2Qp7Y0UnRDAs11k1Dr4AwA/VPEqO67ThvjOSvIEJYDfqOK+AeXKyJQPIZLafK19iAUbrt6F9emVK
STcBIjqR7k2ejVF4J6rYURQQStvCKBe9lcnykFptmQBtA+t7FuqCuhg0WtQq+BvILYVg72t04UW9
OklxJOjypZ7jjcQVi9GZAxa6Y9CVdfl1c9wdB6/Z1pXzFLyjn262zIisBjrRRDo4ixFN2s/6WoBO
Onba3M3GlkrJ+dPMu9/tRoxBG98sirCigHfQbPXHlUx7SaMyn01atRghdpcAIV+qah9KYaKVZ/IR
Cw2kiVh+c/rt7o+pnctF0aEa+ZmHPeHMRsu8sj2oB+YQdmaEj9KuJYRx9/5vqrf9zOGSjk181U1U
ZjC2jw1l3PsbiJcppSYFfSsq5oNiO4zTPkDQbfQpi4D+bvwSRVUfLcjgHmKip9gqkczKL7zczMLV
DMe9xHZIhIaUdMk20OnzIbXb+3oLKAbW02KTdXXUmRujx2IyFWeoNSUnsE21VrpBygfN9Zcs9Zqq
Ce6HvE8FZZ4Qn6ylBSquAQf9GnCA0lPQtKY/P4yMgaIKXF5Vt6enf9P0F3/AO+MiSzgevQfZbuZf
1pK/W01BBctvx5r3/mIkvLrcJMCKy/FLs3oMqh0uomwHLBmBiDzbCld38viuNlLnG9Mq5X2rMzaB
j3Z4Ek3rGdQUshUzcUCc9DE4fBfPsrad30SomOePKwL2vLe0r/xaOIupqk3iYCBEHCw1XfRgs97B
1325vp/cSHiiIr+Ge+DAyS8agdTyzulQEv0hIjvwwjV4pgjoMIJppNFrf+jCG7AZIs2Sqsv0N/m1
eUr8VDd19cEiz4wha+s5Pgu8pE8aO+AjbH9MuJutThIThjUjWpykWgCGmWsT+ceg3cei74uWyKE1
rLAdbzmixbNCAkhFixD0QYgfBqqbkaIcOhCrkUbMeGDsKA7dt7Mc8z3zlexkQgzA+h5Z/nxX6PrR
pG7cIwbuLjLvr4jvof5T0uuUdvqrqmzG9yvLRa0oqxeWawNI3Biym+BDLFgwMcaLos9h1BZQyyzB
RlIK8wawh9LXJ5W9s65NOq29dvatZZACplToJFFeeND/0j5EZPz1BA7IkpTD1XvpiswCQzbpzRMr
DbMKNNMGDQPP/PyaDDMrc8yAenndrFb8dW9qBlnco36A0HGjhEmCpFcNWoyNz+W88DNHm130/P0S
bH9LkggyuYeTYc6EIbdT81q5JkuyQzTfopLJC41KeUPYHHsHOBu8bpDnjHuZidZwqf36tqlPwTq5
jLE0c6NmDazVHdpIjjgcQzQyEno9eRwXTn4rkvIg4oIoHU/VdDlEIhPe4c6905oJsGGmn3+vqM+N
l61LIm/eSmhBdpstLOHXCv3KYMS7qUPR92KO62yjX+C+R02epD6Gtq9UM60bodVGAStGnZ75AeqL
GXoscn1+gigs+qtmrO/tP/Q8LLXFfZ7RadLw0w/k/TQz9/i3pbkmGbzJZBm5t4RJ7OkAu/rsjuIq
7Qoy5lJetMMFki466jLR/XoTni4oTshuxHuyneMYaXa1pGL9N2wWReR1pVTy9saeArlt5y9/Z2HG
zdPQCvVKEfrHlm1lBqlKoBXWRleaIaZAcWLeXyTISk2dUGQD4QzpR4ffXBuVEGy2DisOpGT4Rx1T
+B8VIhJliFLLbeviToT7pJNVYdW731MOOpngJlUhbSQgTaJZQM6fRfbRaO77/w+Xpwa03tHukFMc
s5z7DoqP+6D/+4S4aFbzxj2NItVrUWpuclAj6Ss+z2egPB0n5gYK9boW6+I6FcltsjO1RXgHk7fI
G/DRFVhUfbzSNK7y5LY3zhlCzBUH6jt7FEhZ1GSVL4DNMbW//aagPBxxB+R2uWWhRZWOiM1DjE8X
3/OVhFh2CT73d8o+49YU5guqSq5eVmbdN/U+UlKF1e9ahWzpy2XLJfz3ijbubdVS/tcHHrhAPEY6
s6jr44/oYSPIR1Kv1/+HuUo+LxooVwORt4ikP5WYi/Zf6Y3gNAx0kHZ//k3N05CM8jt6HiYFAjHT
9xfJjsD3kwYmG9kX3N2FLq4UaVgpZd4VAHOp4Ku5tsj8SYCrsRzvnt4iWLs24TWhkazbVZTkfMRg
4PanlqrjIoOKSpp5nvOQurFZAgQrfjRSsufIk59kYKA1TgP6uH8nYdL+Y0f4kVph27LtbHNlMN4w
V7XWoS8WumdnguHlRghJS9HZB2uqrMWTXCzM2wDu8kXAxKLM+gDdWU9CKubo70a8AJGVeoj6Dsnp
ZsFLJwG2jQ2ryxTfbwDRUJumbUtBjxHtR3gkG1zFwqfgdNNCE5cfkA7/FfDq4kJ8P0gDvPCkt6Dw
0DADR1EmSrsEsZX2H4hZqLSl6qJfPs4SYQ3Q+Z8QBjT+5AyHozKGUpQ4s00vUQhM5a0r7jvIMyQF
VcuCHV/BsUPao/spVSwnHPUmEm3gs8FFLhZTfJUk30TUYrdaLpBAIGBypAEDGeVeCa7D314E8yYm
wTj69IxTlHctl2Wl63twuoB61d89NnBLDwqG3K7t5Kc2EuBbSofRqL8hqBitJHxo50UvEw/8GU4D
jtZlqyWpGD67hej2eMCDWooBDWnbjRsZPngPGmq3FIfF+n72L+TJaQyp1plnn276FIKs2ceuwsK7
dWexh8OIpsb0ekytvGzD4vFU3Nx0dG8cM9UGpGRRFJ/yjH28jY4+NkIRYk1tboiNc7x0BCGXiaI5
WvMupn/zwfxSE9w6XSnN9haGDL7dLOZN+bMuoAXXNEHMESTmQJ5UeYfY6mDzDFF4deVJDqS0OwNx
B8zozpgpQw5vD5/hxkGnTj1iOaEiq4N6syl3vKij5iK4UGeQzm01RuHRKfhwYVoPvYOkLPPHsrJT
fDHc7a//nLrvb0jPZI7pS+8paQHYQ3yF4dlTvamWqp7rp0rsq70TqkDns5OLbTBLzYkGKAbaSlCd
NjyyGWoiD+NV4NY7BPoZaq/jdRdpH4ayyzsdhwjKLCu72ju8Oc8Y3UQ7HAdRB9AsLb31THveeV50
MznXQNF8wvCXlDR2tVYny25jVBma4UcT/cBZagHU80VpHe2hOi7gVLsTw0AQEIFMc78L2DqFdOLH
8MADLXCypcr7anBUe6AghB51ZyrY7rX8nsHbJehuHqT5i3Qeopf6daUjMbNjTlRtHe3y5zP6SrGR
8yUfnNoy5/JqwG8XSgSbPBKncuyWujJUamUmeGr7ted39u5tj1rhjAWaKAOC9yi7ckVXMccAV1ZJ
TlNprjJildSKggoA24xQM22WYRZFMO5XVgk6f5Sv1SzyiBNiUp+kJvypnkpU0Sf+fC+AvV97agXi
4azhs67qxssUHYWO9Ot6M2QreJC15DWg2ygRB2pLfVKtCRpXCAFmFuFlWRFR9MBweTdLk4zswDo8
Fr70VS9m6BbtHMdYHVb3KqxsCEbZPKInqA34/O5MNKfnUdW+KDduvpB/rwszdxgibF2K8Irs3MZU
tGMjCgXQgJSqPE6hKilH45yEPSRJMM0taEEnlppa1Zmbadq1kd95DJJAn3B03N/E0vwTyC8crVys
t4Cp/affolxkbOtffQt1nNa3eNBfHcQWnIx/VZg971p1EYJthA12U35kgD2bDICY0/vSATBBX5bi
EhDWPcgSzjR237qoLh4R/PgnfGGJ6KB3Pmbvdvd2swe2rreMkQwb5A7oD/+t4i8eddo094al7Cc3
7dSOASRpFs6hP9SI6TtDrV2QsjRNhflPxx1L0WZ2pliXkOFMB7+IFuHZTFoz4y1MI0IbZIr8jGhk
n2Aq+VOAd7csFPsK2IhyOm5M2+pigYSU9q8aRO1WSQOG1hQL7BlZHpJsCrdrebEBee3gCmFjLCC0
P5QK+VvUpr8+Nik31ERlo6ijvDq+tbpLFG+if0mCtYikjRUsUwtGbYd7bSZPGHOoDiM7Fk/pSKqx
Yq4FYaNVmIEOdMik0BV9X3dimU7hfZUj35PD2734CGlCa8/rh1H1qHGoZzS44pqCIoeHEey4vUtD
dsVKVdkuxdE8ohCS1FFKP3XQ9lz//IOAahgiiQzB5gZaABS51yY1uwG3gJdLZflX6sfasFYSt/qk
vnBzgKen17BLxJ4ufVi0DWFlBb4Q1NwG9sPH3kiU/mwnfftVmRRVmyt0k/Tc1MbwUDO0deKhIqne
ZOeKx9OSPftTZX47qC/0xXpi2LR8/xEC4XlQg9xuqHqJzx3pALpIFUnc0kpPkrhVWKnqvgjzJsW1
DMvVYNSpdgCqqDHLZf3+1OyCcsOjHRs9fYsJqHmY+ZIQSCpBIoUHhKwzHMBrlKbJvsaC0r/QahxD
eXLb7lbaOijJXBkutJTTveJ6sq/Ix2wPRjRXUAbKGf4TwNwfqGChELzyc+K8oBJjsGE0PJhNdI8t
3D5+dWC25qzfQe1/8NpXYOzdaq42RdOU5A/M9AjLpHAmoR4yto5McvBwxO28SveVR7FlStWx1S0N
zJHTYuew6whItLW6LYqqAi+l5IuamTelxtINTCPaEgmWlDRor2jy2qAr0hOzZrvA2HKJ6SUj8aXV
Rg8PBujPRbJ3Oc3FIKPiBVLjS9nu6cJ2nXIqOTrDTaVikWxn5J1jpVA6p8ykd1OuKZm9PNvfxnaD
FG6J51/vFtft9kqcVD5Kan8n4yW2IhKXSSFnyEz69jRTxyl6RR4INsby18wwUi8Ep11NLKilHJVC
8c8CQtaX3ZNDHR4dyjZ9vlhsexNRX1E81rJSaUKlIEUXaqwCPdsjFG6JWwlXrBxMVtaLcHPliOru
kneA5m91fL/qKTL0ePdOAyRMH0iDhM7xFIj3YugOLrS+JNtXJ3DerDZQPJZTn6TcCXPS+R3jveai
BLdnghGFnAR82XlG9vb2sAOUZ0F4qcPRKbZRTRAavgv/kA9quppFYBfpf8ZAxZFdXpvHmo+3ov+p
wXng+yfv+9pHoLQ2FXo84sAGJkigK+5/d94IwX51t4tZuUuBd7zOPN5SFIA5RLooSAHDi+vS8txG
8E7GO3dAOZWcN8uAfbsh2v92Bn5PL2HnFN/LeKPfm2bxOg4DRTKTNcWOQgprsErQrVBZTwnj/rV2
/iZ2ddmXCZYn0yRWeQoLmw/6i0wWXtSo4TRiWHYXjYyrWWrYuApRghXOQzS7djcwusIkIHbd5NOP
8o29KQrIBQDG3BEsPTPZZUk2Wc6T3RlDDYjzRz0IJbOjntH7VWbLVwGpi50jbhOLi3Jo6/VzUOpR
48iBENSsDa8t0w97a59H6tY9mEB5uB9+Zs9VuaVOteT7r/XGemH7dQMb9c73z2prQtu4SOtkSAj3
F/SVKGEcjXsqkvmXtTeisMJRCmVkeJU4WuATg508bPEajvEupZv3ISeTU3OSBArIyVSzRHw0dhFw
WOVjE+bjhHdFVndGlb7jrgwtYbKnROcBd6AYOfDZMoMGLe959yg0pWVwVvv50psF9W74lR8JJCUm
3bsSrvLLzrZx5hY5C6gFhIYCkhbZEOpKVx5svfAuTopx8yJPJwRlVGnjWHjYCFtUPpgqs9Of788l
uTM4EKlMtsKUcDlx4Bb7bqO5ekmQ6oejn1GM7iYvnpC2FNfD1NgJWLVIZ8/lAjpqVOARNR5ZIBf2
ZhV3aw0oPLz3qF3HhFwziEtAs9uI0/ZzavEk/entlDCgbZhajjPo99EL90Q0udNNBJ2P9RyUFU3Y
Vl1aTWP0OpJctAE8f+1XBnnOKw7UO6i12ga8jJWFvBhQjvn3j42E1s3L61JGg9DPPTjGhjKFx8a4
azieBATiLjPnUW+586OKRxMOQ879SuLYoldd1OwVTr1657jAQPBJ9aQPX5wuEjzCUzaPEcvfb08D
/8g7xdoWjd26/9TZlpL6ikzG60aIF1SQYUrug/ltz5sZnXbFb4MCSQ7+CMsLoFLbYpPRZ483ZeQW
DupmiKICREiFxg2Ua5EtudfliGi7UhVOXtdnKnjvXI+76gdZv9Qa6AaLqoPaVN5xUoxQ/SSkv+7/
1YZWWd5OG/CuPochZvu0IRxqQyYUR9GPSI8j97ENwav7Yq4lUlmcT0pAxUC1rf0zl5/bC9NTc2fA
zMHhynHs8kXMEsmfXv+CgAwV3Cs+jxqn/ZtEPDeTdSQeRbMzsYUHKB92wqROnkH4MPCHs9GXKilq
aZoZrApD/MeWz7Gdj43WtAKDgPr/GQ49em2P8LQX9azzwzH1a11daKjV5GDQLghHAu8IucAXDd3c
ZcVb3fneoC1rNvMMKLWlZ9od4jW/msJZWZNG+h1YDNvPSC9YND6+2cx/IfAyF05Nu73EOJ0vVPUg
YtQBYPO20XoN2TPmPY9KXJfMglvO6eBEt/1CvmFZN9/QRYJg9i7b6jxQtCGfwHsPDcS0Tliux+fE
P3qiEK/UjTxbUnlXPrhEJ0zwRIMMPKTt896qPHG/N5LuLn2um2KEF/xfNt/z9P2r1YvTgQLUc+VO
0J4SGKcNqwjdD8EaoU3GiCfT8LKoRFRvKRohOoALuVbD4kmBkSqzE7qA5eto05qytz0mOObqzP2T
fhhfDCzqITX968a3EVIYflswQfY8lwsXElgSX7o6lcB3g/SoM3TLwvW7YNCSqPpuQ6psBSXCnSF+
4ZUQfmja/Tc22ntiRcnMwcF2IlZZ0R+UTBTMNlno9HwKuOZUUoLRoiT8qDY69Juqj+4qNA53EaKy
HcLg/3sceZr4hz3kv4KpMV8jXTUFHuhMXeuTDcX3Ry3elguvIzSuyX/Fvd8ODxW8UdZMNOgWe3gb
XJACPu8azR5ny9sZAJijmlwfdd4pzegfKSR8ftZNYmkDp9MzTc2hfviElxqnWDkSOIZyg4G7Kv2E
113uVjQTc6OKjEmiMWo1/k0RoNENd6LeDxpU3SWnJRkczhth9d2Ee7Vx0CjDl1XK0Gro1ihyNgWn
tGkOIrWlVBKirsujQqThgk+r8HyDg/vmLRc091khzcXg8O8smz8LBYfBGP27K9TO2yauO2ZQF3kw
LfvmedH+rCyqoYC00I43lh3NsZlHjoYc5yzYWpoEUmAZmjmnutNw9Nawfmv9fWsJwR5QyJ6oXvsq
Vwbgpf0v8CBy3nOnPa4GHxPbw3wNUUWBn+MT+3YxtPt7GfgpbyGnQ61mJlF25ysso5b7VNY1wFGI
WgCBLuC0I9mHkgQB8xIJJX3TKrGr652qZd7bi+8MY0hGqlOzfEC9vfpUf48uMjwjkBhE63HVPJ8y
+/3aViGTuPK9eo8XRTjTw03PDFlLacQBdWHtOowTsdwWQUht8ELtAVEpPiQzhTk7OErnMAZF+pgS
zmxJp4PIxw8M/PFxiDGKIj9sYWyVg1xh3/gUbggMmGVTt+fuvlelFo36Gblay+v0J3W3W+RI4JbO
xwctLIdxjiQE/Ev2fsuouThHve7xRN2/a88OV1JnVLoYTt7ZnJPzq9kDohkxH8MAOKVbrsVU10fa
HmDMGuaPzPLOgR70TyXMQbL1i5Mir5APC/2q63rxbpXzghcw7gYMA8EvOBj8G0fgRUkG2udthGIh
pc40b05jAZgxRpOgMF3eSj8dRotfN8EJPLnXZQwAUuvJuTFN3lhNF3HwtjaNHdNcD9/1QRazkt8P
OFHilPTLF2KA3VWnJjf47VVDKy097PbWarGa199LIvRrpL8jQApNhvaqZ286NNLsAKSqidmNsUiH
TXj9z/ccHbGA8lgCBkCtS+JFsqkgl9qyWEohWmSkisqepY/47gOt5frLrveCjmrbGkvhnvYV1x6e
wXEPmMb5bvrABDHq7+MvpejEfKQurXHVn5DD37N3WnKhqfhQSkWzjrP6l6HpgTlT2SYQrk9xnptp
W3aqZgXuUXWgOiYY7DtOkjSMvDPKS1XsEhywVjIcxK8vbW/Wr+K+nyP/sorai2AisGvf/9y/ccO0
lBcyDXc/2WSdsUeYBmfoe7OOHq9yfZKDWQJM2ziirFiKbDOlPZ0jtzyjeWWEE2+A7QRuDmGIHV3C
lR8lB+FkT/vSD+CWf0G/dhhafuazvnalU6WdEFHmDdTUPNCiiAlMkVZvtL1+DeandDT88bv9Sfqc
hLXqMR+lNEkHaVkEBVwvgQagwrASurzftz4sJkmBquBAOvDv0deIfeoi7lVfUs64AHn2+Ct+p0vL
XZ4Crj4kOxTL5vJ2RcntxxcpITwMq0DlYPWDPwZWiakzCGH5SPvfMcHE8T9UltiKWVXwdHtBsrSh
r/727RJov08Bv98mvNeNRMzVw1RE/cqokavUfMxFbvSNeUrqYbI4UamRiLV2qopwVPfczydtOtQ3
Bu/YJimSzpC5Wlh5iadmxtsOrNA5Uc5JOHJ9zShZnkE9nS/pnOgYQsWtJsOxssCvXk3BEkXhZVfv
ghOEhx2inbpePvgXAaQ01KsBzWKSAGwcnNdFgjhSYc5U6aiYoqHMCgzDeKBssCK8j0o9uM6cWyah
E/JG4+9UbXqXngXTVRoynyV4TRQ5Rws8Uz+CpqSRvvijL1vVqebCYpautfforxvlXj+BDuY4D8O6
8CYYmr0EdhzMn+SFpCBFU4U1nX8EuYQaduSKuPYsQNA83qJCTMkDGqcnu0x9u2emd/mdp3dcxI/3
6GoSMw1Im5YTfsdmIssDHaWRAeM4Yw1UyIrs7TdLto3CJNZRvFaeMVxQqt+JFgu6Xt/O0sr4u+Lt
ZGCoB85mzbBWPbnc7ya+QuBtlNlTqoGn4tW4ed2NwPavxwTqc2jJSoRvas0ac4zrlXTUTQPy0i1u
QfRYXR6gDRSVA+8bwliU8aJY4wTVlzNAjK/HmGX0/6s74bxZ9OoFQ8CQfLkJ3QJz5EDlakTfQWlD
Kcko86+TkP3XbQS3PUzf33+lMQcmbZDhKmmX9SysllU58queU4VdwoeFIVSuKG+XBxapUwJ5KKIQ
QRrAgZarrnCOPPn8Gx0815nuiWOpAO+vqvSX6sk/3yOi0Xu02b6FnzolzY1Igw7xur31RiGjSsud
jLq1XWJRNBEl48NilK+gUTuVzApRImTOERkksUxhKInJ7q7ohEPUJTAHwXhQalcX92ILkusRrYzS
Ka0gH7JMUO5PY3glCOzk2URX/ICoRrxbmhnqRuXJFC6sAYZ0mxnkJ7a0qmhFwtT1Mw4RSGYhQVTh
URasaXNBm6bnG0iGqPfEh4/3XLxUTDD3ym9O5fpTQV9QVFJLe67mWdLugwbqmwC48kjRmKHDs4bW
m1YbAM0rjClxjo+rfEfYepGVCxuK3DjzJcLXfk1pRMhy8Qid8KMXe1xUuH0BehzME5iuv0f4Fvmg
UUrEuq8B+1NbFSsCBEfFjMKRg2G6wXapO0U1woT0uX7M8xrKLkYtBs0guBlSK/6Ut2mCFgabuOAp
Uba2EPbZz+GT//GEVPWknea1/ZmB7NSzGcb1vh7VhXUHeUv1t22xK2JbbB5pnS8+LyN0bFpcvXCF
AqQ3yimbIvTBYOB+UI8lU3ZdlbXNjqO0ReA3X2L/loTDsUvErRpEb09VDXOJNp+9ZFR9TQEu45D8
9D1A/e/f6Dnq0PVcUGftl74LkfWqbBOXXAihFKGJT4aGcDSZOyIR0YDx0GQVCT56pEKEevFgkJR9
eptRxVEDJZoxwlFLtLbjfeOqXABUSPznfpVFJyHQv6cGszwIJOs0RpqniX4Eg+YoexcUslIUs2LW
5FxVkRgqcYXtWgAjPtyqbA7l23ZHV4eY5NRw7wYS6SMafPu3q9BnBVN0QKOyP9AoSseoIBAwNgvw
stipgW+CBvo80Ysybuo/SHwsz2hIoPtFQl7as1ODvBoeCfW0jkYymMglHBiqga2rjV3VM5oPIMDQ
CoOLSDmCLn7Q8QWb5kZTPZcRpL0j5JRhpWP1q1RZJMyXDy3iv+M9T31wIKFRrjRHOuTY3GXnmdEV
Rmt5kULpvD7YqoYcdb0/FTozAKMA0+BKQAVKd1ZmuW+p7g9lQCk+t2Qwy26poA8zloYni1xQfrrW
QgtTG3gI4IHn/4gqg7A5lt+lJOe9Mi2ESoWHP6QEXKcpYUXOZzuca4eH2WaIJ7PBGajbI1SCkGVp
k5ZR5sCId5mmoPF4BYCA4z3n35cxTHVv7LLhfsYQrQayoe/Z/ZV8KY7xEN1qFYi9MRVvi5/a/jGM
+AJs9nA6Ts4V/5mbmHVaufvu6R2euHfLhcdgibYL44X9HPV7XvmwHxfXLXhOA/o1zawWmCZ+9Fi/
pQ/qTDQJK15Fmty5DmeLu4fT/5YSEGsMJMnlqiuiwerFN2TidbneQagjHWcvpogcrfnQzusipB5g
iyLesL/7eOuFxz8yjphJGDD9eFHNXDQrfBls228Sk4L0+R8KVFrZs3nshFZR98mIJEkGV04P3khv
81IbPIcDhu3o5Mf+W65lj0hct6Ywd1wWCR+bEyGnmyKdfOdXsUzDIAs+6eK1h18cotdPLf28GUZD
StSjxmSgS7M3BcS2UzSim4tU0HyU76QP76fDLsIUXdEQEiIXzG4Ncs3AUxTlkI1C2oTWsc5v+608
b3dkELTM7qkhn7Hy504RETXhHtJ7KmQTQeOaHaVjeyIKEeQd6tS1L5XjlouAjz6Hux0wYBlggXA1
i+w+YoNyBsKXlXZIxH/kY6sG/UdW25xXtw7ZTuvueGj22B2BUFbf/JvuWK9V+RkN67r8s08ED10N
BT0Ar40XkbLviIur+D5a8F6zO+UTgs2FCgLgiP0a7AyuuCAsIzrYaWrnMH278Xej5DcAbrkHPq+j
4psngkWRuvq/b52LGAmwEpSGSDIogGWxmQw85m4T2m6lHP9cYXSaXXPyTvEfUQ1icGpqG0jAcskL
UIvGkD39blnE6yhGobLeLa2jqqSXn/UaQ5q674bvuPRax2/BYze7lEZvhoxf7faNxqPgQ4W5gQtV
G+DDSPF745CUhvvCvMyvdF9Y/K4edFs8n4jwfr/MuH9AfNSDD4fs5KX8VN2O7L6LZl191d/X6MuY
aLD3qIK9k3pfkfE6m/e+32fOU+67cXZzEGJSBMiKsqkW+Dvfp8ve+kxvfvsyFZJZvJiScvOltYSv
c5qdPYd6Sw7dKktp/wEKmako82sMls8/+SquNwe6H+91LNjRmaC/PM+Pg6EY9TxEjwKKjXhK7Uob
no4ORhnEgeTVAptoGEbi8joDABsuQ+iMxEH7kgIB5kdukDzbvgkXwKgx3F6Yrri3TJ2rpYhayRyh
uvs8HMr8KZMku5Wcp6gMbUBllce4NGvTXgNrQ4ySa0YReJ3QRJCPqzBxquMBqEo3Wg4kDUV1xwEj
9qFMHyP/P2rCEbUE7qBSL1m+SHr/0ThKxraVQ7JjyabkbQWVll+xol9Mz4J8njUMZzdRX5olUhfQ
RHJiCVYw5mLDBv6qLxQJQ3u3EksWwW4Eza3nbBctWOJ12RJnQOGF4xPXc7svO2f+4lj46bi0wBJ1
vnM7qSWdoZW4Yt07+fNxvEk+KM4mdh3RntOrhv5sJtEJ+kGRgYzP/851zeZ9RH6TnsR57kQ3bUw2
clRTI/4HWNwqqe07lIpB4Hk46d7QNEM5AROoyZPDPlX3ajs0R0v6T+xJ0en9Y4/6aObHFzM9XoJW
PvVDFmd0GsQF0XvUZ5C7v0hkj1PUlnP9quXKvCmpTjqHC5WBNsUuK2SFYVQ6zSVq7gOqCX56JW/g
fcUe1jRTo+fhI/OH7eRimx4XTWsSAS4D5OM1a1VSZEcEH31Bh47iEQH2GtHty5hZnEyAsBmcKF3K
Qk7pW85GNt5cqCWNg7QBNIETEMDHF1u+boMsWuogY4JUSD5ueHhzbljB5JtZsEG/ZVh/B15H7fXn
ba7+8xH+53BesomnuIYaeCx5nlfl2E0iUOhbNp4qoyCZMw6UefOWxUwANRI7doM9SYYD6/1r2FRf
V5idb5fB8dA4uBvPJC+TJ+ckLoFbPN9nLhEftkgjBtBBJYRWERQEbiM8Jcnw10qpJBDkddd+zqCP
HukXAFLSmv89XHsfig1Ml+4tuK+bNsPzk4TBWvFS+fcwVk4qD+QJlFKaHjzHF0UnY1XtsZxbqfsf
HTob1roYehA54eMrToFo+8ypPYYdNAbdrR6kGvUdMpAXWAUcs8VesHd+x2AzDTLBxKoTVt0vxqLc
B+QVhMwZ5Dh6XLLVDH2Vvxr6BG+3Ru2zstsd4Sj1XchWmL+xWOTRNAMKbLGN/LzGw9I6ijkVxHTy
TbLEdObEk6v1BOgf6Mbtzot16a4DX6zjTNxuHpu1H1yEIpbO8QqxS0CR/5k7PTY4i+1Rsve6vC4W
azYFK8rwkKSQBjqKUNInzwUdIz9BsbfHhbLoFYhzoRNAYSAbwOIJ8g2Ae459dqi9x+y4jdfQiKpl
ggLyPqGHyWiupG17Sx9+Rw3elE+FWwmNE9Ip7cpGG5t1vbKU/qlENMO3nJxRSdq0F09zQEIZAPBo
ypJEvRmvQbcTrqg9LsvLelHFBwiun46WTQ9rnVm7ed8nTN8SwX2cKat1DxsznscC4fqzftaOOhx7
nSQNsxCnp1TsysRvoJ46T/AqaHtZampmM7AAa5ah53SnZdGRqJIingH+l7MrueEz3svND18ooHlt
raGk9TxtmMM50iolJNP7ip3feRm4wITjt3rpxgpM5jZLvDpnJCbvOXYLLjrV9juMB0VmiYErQ2yP
b+IBDiHkXx7P8GAHA0q8e3hf2YuSNA/MrrLPhpiuK7rqcqlnpduzl2RikhnoLGyNWlv8blPGfGLZ
mP8qoCKTWGWwoXP8odrcs+TTgrxQES2EDzoG0zmuJjpNtjKSjYBkEfg7Mv2mrlC0gRvfxqIQE4rd
C8+5nfN3PIkpEmST/7LyEOHaN1aAcsjE16w++GfzdycUHga0G2RA1j+IGynrKVGtdQZaYQv7VRni
evqG1Im/C7GouANQJ1hCS/BsF0QowBr/+SXYobUoYOTXcNl61TX09SAw9q06FIwFtXLqGphU8Dgc
79I58NkFIsTXwrgqczlx11W3xsvyHdS2qbYqmF+LcKtanXOSH+OXt/g0sPHjpyFOMktO1Vc/3Lm+
Kq+UJ9EeEVWJEimIL+KTk+6ZZyqwQncfZVrCy0XAzOw7UXPIrAmiAco8h7dvbNvfbAdOHyl3A8E+
MBl2K10gyCZGqRgfoLocAoQASGeYP82HiYmlIEZs6czwXWtL8Thc1NlykJJ6sf/sEJ5n5sTIDwxn
Ba9hoeFgz0lFzEEkmKq8bWTIdbfOF4dDspzHg+gI05YPmie6ZNkWBNXuRGp2UEZfqaWXvULXX+wr
QXueVP+wFr2VC+DGfVCDgngFWwuIR5a9bZLOx5rhxNoFMIpx9jN0HnmY5SEDCcTWHLRzhAjVJ3vR
es6SHRS9Rb7Q8b1JDAQKEwSTKzlsroygKzhR09tCxzZhl4OrjAsrUrkmb4RFWF5/607E03yxrq8b
u+rLdL/x6dC3Dwddxc0Ffzpj7ApEboBD1JYqrM4E9M2aAZbN56CXo/JpdDzwZzHQdLrSnlVIs4yC
iLD1aHAk/EGiDXouBH3IRDWBv3/DeQyF4nmPqd7NUkMqN1YSc+AIoc1dUWrCzU9YTYRL6qZ28JXn
fmJs9G7oJurjisZ5UBWQWcFJwbbt2oUR4gUEBnBpiMUmDqBvl7dyyjOGDY4hEV75ERzJ0PocIS+v
RknbsM9gOun55U4mO4EyusMvPj/oa0iYjEq4VWhp8kovbV5/BgVZk57Xh0tGGJQFs5rnTmXTSjrO
BKFfP+DJ3pChWcI9kuiyoxNey/VmHtOeuz9milXdGgcUclJcpJVchAQJ/agEa6lU0/ayBRXmupn1
BOF1CiEC97t6ylAh9uRQ5959OxEZCdvmn4kKK9YHMoCqwsLlwQ86EQpxs+sJQEBudeA9O1eFFNQJ
P3kVb++EZDMVEJRJoI9W0pUlgEpvVI4Z43gKzp1We4+vNGtagyGPn9tjLDZC1C8RITr1+Fs1zrkM
kqtErPav8rSmJcBS8MGafkBHwn2irT2NcIdhgJ2MRn6lKc1FHC9jsPq3bvQnrGBy4QqHjcttUhhb
OeqZyn8Vc9cWq7R8YUb2V1se8tpb6OodsuDKlySoHFuHiDy1hWJgx8i8n55F9w6InTulimMC1u1p
n26+bWOvAUixl5/BHHeIWRuA2bS/4XmFavGWu16v+uP7jHFgqTSoBTodHAJehwyK2P4RUbHnFNHE
3OUZGbVvw5W3eyYWU5c5KMY9pMRAjr+0H3dVDjjIvWGYGyDLY/1U2/G1XUo++J/asgZj5J4DHz7h
Pn9hjioKIKyxq+iqzvsz5orrTs2STjKYCznPCup/t21McQVGFsFw5UTw2s+OEI+wfgUA6Uds+o7c
IrUuKtSc1dgy8MobMsdZVapOzXWAyi8uJI80bTjyBuL9NeEPfZ+B2PJzTY3mFxRNw4qCgyq+20Bk
xc6k92lK6kI8fmYgDI1DTPTcZjSFp8D5yFOBX5Wmy4PBBzfcHdjRI4nbmggyZ9TFOUXdb57kHVeA
mr8qFK82+bzoZI1BKoZqWCqzbCU7GLECOKj2mNvO5+AknNaN7Ugt6SHz4o1kFdeeBuOuleNaM004
6H8Pq+DszilzZAKo6LZFgJt89gTWkbGUYvDavslic4AIO4/btjn8MDrThe0ThpbtKeyxt9GGUGCZ
83HfLWJdOf8fp1DnSRwTWwVLHmZWaX4H7aI/LglR9T1cWyETPlj8BJ0vWvEXNgICoGR7jS0XfL4l
2Ii1tENO9iYvHaSRv5Qv0orJ/aLQzC4PaqYODd8Sd9DSl7kIIp9wHjnq46HosMUzcGOl5w5wwm9L
AnG/ODHRHfyTZ2N1xN3s2hNloFYsW6lt1GYRouFLW1xXAQ0bOUThGaZ+UJ3R4aFYsTkes45i5QAl
bMKYl4UNjwJKvtqDB74xyJ33II44gw8YPfV7eUN0Cu5UfY7o4KqPkObeLEaA8rW9zhyNmkHAolVP
l6d+wt1df0oQiuw2JzHH22jDLlmM/ziR2Npg1OWVpjBp+X1leXn08MvDRBlB+I1IzwuG8BL/ebZJ
XoSd36tX2KtC03wMfLNCtx/o822ykEnsknrTVBxWWwzOoH0cgOvZ/nPMb9HDncYFwUVjP5p1hpdu
4wIMBiqcZ0TDseka+TNu24tx+ebQMEevSmtPY2FZVUHVciSA1tqcI62Rbw7hiQ0PkCmNlmFmYOFQ
RSUSkBnvJwQxKup9ETBcsifu/we1ZnQIdAfJvjhEq9fjBkBoLS5AMsNJWxEVItpnbArc/IJbtq47
nSTEUerpERUC4jPcwOkP0SR1t+Mj8kmpcG2MYpeHVV4t/NxeEbPwmpV7HS6b048t408LHzeV1Hfn
JVfLuJ39AeuV2jqxvrQjiGUUEad6l2+Y6/XZqvojmQNrUe2mX6wibRqw2lfS3uZPiuFlq/Ac60DK
yg0oCTVAh8toPNHn9keZOmJ6yj+NJm4ueohYoAfW0YEHLcwkwFuWAwRu2TjqIuENY9zksSdhfMlB
+c6uayxTuLymC90p1eOuDfL+Rs1NnNuGOraFOGtwQJsoml/rf3c3UTKBx+x8KHXo//X+/5ReHuVV
CTG4QrK3ixyDEf9jiipksNdTfLQff2ujxwy+ZkjB+MGUrII2q4vjn3/YH++xFTP5+l1pFO+Il44A
Cid6p9+oYWfGj/KE+l4q3N8GHs4GAk+KyHpDIRrhV3V4BLgKOGwINuIn8U72e7B7oZCRkbHS40U+
NNUG+ZaA2EliMKS8lYPyj/VO4Mn7Ztynx+nK3skgFsZaI4lweU4aJT8C853JqpcOjwtFuWt/dG5C
l5zyQwjah6S4RAIzV79yNrYJAoEdMcuKIsjcvRLzVwY7GVwRVdqZOc6xJU90ju78tpwAPpKGpgMv
stgNxeYpNd+YxLgSacAbuCcjszqfqB3adNNTNxz9FhEOUeqOM7J0quWEw6AWWxPyx0aZDrrKygCA
eV6XvymkruRRmpyqtEpiXb0QPQRKCUYW/1wJ+OK3mat8dyXIqbEOBi+AJWtzsWIFXDKm09jxAPxB
mrPFeJRfR1VPSpnv/CqtAunYF+SgJ5dwZaBV0zBQoHZ2sIkb9oXYSfbT0nSUIpbgIlVSm/WWt9ps
t3ftW02Q5BM3znlcAfuB5eYEhJw/azaCoGedRBiDYzSJEnLOEN4GW/Z3oPE+Yq44SEbsx8lXCEoc
e+kEbDHrjyIYe3Yi2TMr9aGjGRktt5oKp0ol/q8aVgmuZr0B3MTsFTeJvPyq4Fo9aXFHD4aHhHwU
RSgTtLyUCfoY12AuxEAH6smvo2CbTjvRQUtFoVTjCPtD9ywcve4IxALo6j9jiWnvrys0Mi0V6mo/
cH1d6Q8YzDd6x4/fKOW1G+F3ZBwkFFcaDoAcvtviy3M4HdxrHxquLEzlGedIDSR1gj3Xe1JFUUEH
NsUeJ/GvuomlrrsEq4NQWnnFIYclIWj3AuyVwcrkaRgEeKF99PTnkppKF4+svYM7t0FCuKtSWUwq
dEmepOMBgc8uuYOLLj/+Hki84z6f1XROoUGtG4Z4UfM0knIeLKbuG418MiomMhfdFF0t2zBgZsIi
ch1H3R7AFN7H+O4wAoyDs9J6BiBMh/wjlFCu4cFNQkZOHH9nW2q4mr37NvOkOT2r40dcyCUDUIYI
aIAU6QBDDE7faK0w7TOOsJPe9jMPWWSbED6dXaVr8evy/m26tHVmoTLzscPylXMAMY++VYnZaFah
MZXlX+daeaJRlVI+xOJCGfRNGtQZqGAEnys4hGZk6Eh9N3tsjBwLc1wfoEoBV9fAL6trOnMxJr0J
R41b19ATH47GMukcX5e9d7dl43BpFZUkeTMKmAwfdSQ65GMfJp7N0Z71WM9kgUIqFywtBX5APgZh
znQBE3hjVBmMPxbOck4fbjqsj6DY6G4JFQC2ZcpigXyIRiE2yRvHKDk+YPcKQ0ocNBDQevxqg8tr
m1hgmZRrBe1qwhRe5gaWQd2NhzPuq9r5npx7j6l97G54mp72+RyYnGonb8UFsBxxH4Zn3MJyon58
+EjVhGCIKtb+LkRiWcvDWq+idl9NPtgg6kbJV3GXYRlIx/Lw1XrqlUvO3ldh5cZXztO5X8aKcAtk
af0wFyKXM5PTMgFuKXC43u1Lae9yZMGEipgn8gyGBucrornP5HsJJYwiZaRODnsVgKdX2ZIn72TJ
2TgM+Nr7F9ikObofbMGtKA2hgmjVFLwYR+56q+xTK01ETsBZiLaEu+b4l1UErGdtx1QZG/sKw5Un
VmK1coQ3zm5IJFcNKzmMnAS2+h3OE5rrkVeVBkjEx1CTsMHiiAKqI4Eot+ad5s7H86pgMiGpcEFU
ThgwpKdFQQzUVvsjNO9705CwycvoCmN78wxDwdE9cv9FBScQWS+IJGyBLgKeUD7/J23qbN6n/SIB
nJUu8pGIhrPHdNrDKCoQn4Sc/GMUNEUxbMz2xiICM445COhy9dLBH13u1pc93fc8b1bo2EInyS7y
jE7ePkIHWz7w82SFAgjHH99OFmSyIYA+1GvWB6LotHkRn6jrj2oi6sbqrWs2hrJ//34ncFM559OL
NO7/LUT5RhLBM0VyytHVOVkk1OioOdFCBxyBxFjq0q5bHiMMwWgS5aXDFq7e+49Fntk5fTcRgyJk
E2EaxKS2cBFYFqfKx4H1DHaSEzYYg1W29euqTIsVb14TqpvGPcf414a7nxEpCf95C3DrZukk/LEA
mN/5WZtb8gwhZDDrHHU/6FrlZvOjkgKHXqJPFCifuNFDplFaAioFWBCE+GKoxTIco3g0BnKTqWDV
t9RNlPpvKESYWe+H8pw9FSWoU6d+OUBd0O3fjB4MbeUR0Xty7OoLkQq+RVaWfwEFMyKWA8h32Fyp
3QV3cpVLJYoH9I/mHoLb2Cutz/u3Tr9GCWOR7lPkwynEFNVlTh4y/9xuD//V7twb06uJgjJNE9E0
KZzAXREJ7ioY+xFpT95/G+iNZlTnJQs6XmHLe5I6vk5FwRXm78CzuW8Jx3JHyZsqk2BybyqhKCYi
dIm/qxOpU+pzr2v6rrE4uPYw7+Fj1Ciy2oq8+eGBdxKUySCBKjrgNIMnI+NjZsyGy8ZjqRKd/+IH
x+kib1vNm8o3tX+fF0taIe0ECBkK+ti73hL+E2du4e3fPLQSwI2uydK/dMtMm2Bl/vmhi+vr95l5
Z+FWe6moNfKMiUI4xMU1r9EL6g4H9wA9yV96Tmv8YIRo06MjiqcTylUu9+boZgCaSDq+72G9xsNm
CMVNHyLiYuZTGoQowb6/mtTT3TrrBG79ASGj4YqEqo12XVfNIZNAnbv8PfioidsUeUHT4EwpRxU+
L34ixGyk2bIqJym3NAfmsqc7YSKvzrUNDFb70hmz0h5VKRzii4nc3K7ftX3BdmNagA5Q1tlMW6s6
3B8xtsmFXib6WF/RjKiukLpU9JIEXGo/vy/1R9GpaYeAsoGOrb+p854mMTf1tbSJpLc73w7sJJ0z
vfG/3T78RvllaoYI20NHK2jlhCls2XMsO9dmiXh5Ej67LnWQ5szWFJAn9DLUxGag0CbkzzNCZ9aj
IWEgmxV875rkcy5a+dWCjNiwoVaCdHI7soYsox9yQ0OmhSdMeXIM5sXKC+8hVlbMTzpen33KtPQS
5gZOj0JBB2kEwOsCZ8j4/hupgC0Eoo4psAF3fQUBvMUHAkupBcmvqMS0+CVJV5yDPmOhcSCmP7j+
JUZBUrpMnYfW3PFe+ACrHbgFaW5Qc6EVkxc1hU6vaEAwXnU+KsM6QefAtXtOQ4bhpJl1+OSVFa6V
m0iAeeS5M3Zau9CeQZo3D9WVOivneNZdLsPD/YHbHOOFgSW7raZZ0PasL5GsBnPWupZoovMCl1/9
jEk2mqxqqWOHqr8rRrJa1YCaTWyYATBjHy11+QMNk8OoZ4QWHBh1mvtpEcFm8sYuad7FMeFUtVVd
FfXic1JhHHESRDnAEdh0V8l/53usFfdoCYL4cQLxX5PZEjbg6oZeFQ0yByreRu3QRs27dwRtgNbc
KyWmAlH2pA4wchsgaAdmYPAOD/NRB6gHTiGbMoa5/x6ZKgXZV+exkC0E9BlfTHfNs6CIlWtCQPEy
OH2T3QW5I+HSSSj28CrfWTOiQ1CwREhiOc1iAMImIAV1jnH+E5dn0Mh8avXY5ct5rhXULd+ZxPFS
9d9aaacxCr+5lR5w1vvpFGK14JeoyAD/gmRiGQ+X/2hcXzFO7Ssw4npXivg9fRW3g+YyjJ8FfkXI
eMK6cXTCddstG5W7YIEr2Wi109H47VxL+Keu8M5CAHwA8i044cMwHqn8aLTAKUT8GwQvvkYhx+UK
tRKxpfvc5q07hbssTiIYDNRQEcgEcvBpj8I97gvDoYEbSKsIhNqGXTZ1rD8J7W244Snc2XuSNWen
UVwJFIb2UD8nDO1Cx120gJvdly+hSPeIpDORfHJPCNl+p4Ilw3Zol8PQrauj0oq/f1HH3XYnMn+v
oE/v1LK2lPwo8TCdrrPbSK2IF9fdLs6v0RkwuiWXTqG/R4GydBiPoT+7U9iMKVFURBPl+cYTJZxr
YvIH4jTzJq02FeneG0UQt0MiagGK059+6upykuoX64/NY51fiZpdp0mZNKD0vDFkiMe0VBmFiYzT
4xrouIYuo0BG87yCcXo8lHl2FAsF4ugEIVmF+V3z/lXqOxyQhe/Pw59upV0ugHJITJSUaGzsK5Uc
u2IU9FyS5jX+om6ywGMKqaj+GILt0pjgpfqA1nim+9WGlWdQlRUyGP8l5pNfSKX12xrU9ei8b9XP
UJbVFxZbwJXXayibvcPtNoF3A5uue0yOkl7B3jDDyXi08aAhXdfhiF/rAp5pXU16wOqGKOnRziYK
d+pfRruOPhBTQTAhqvp5z6q6LMkOEXTHGPdiaHXGkaUp7ynib6J7SyRjLJEUVJmrlAjv8jpIFdwW
AimGqYww+oa68T0vQe2FfX/ZaFjVMwW/bCB4CZbajRIpCcGVzw+OQdzeTBK0O+bINA+pCnoFNlGS
MvQNOWjJQXTh38tRYnul8eY/6qMqCrA6fqFOhrJBhoMVqKxehXHh7HXCW4A9yzuxywsvTI1KPPwI
N3kvAC4BbJ9SHbF+J58AYpKUY3/b/OTUmQonYwMgJgdvgD7gljJjUEzxrGANEXXh4MCaaWA/U7T4
IPbYzfah9zhEYW2yLhxqZ9t2XpKlDy69A0+Rr3DbpMOP9que8A/suyjFW5AZw6cPnIHnyswOSJVC
NZJToaW0T10L4K3muue7kq2iVSDvFrquz5G1QgExdfaCAT4eboVkr+Rl48kPdUP8WM2zpTUSDkJB
QHPn3G2Btm4R/44m/t2JVdi8RpzuuHtYLY0CCT7uJCrDtSIkch4YGOaCzIwikr11Df7aZgt4xWV5
NcNkeFv3MdkBE41whsEGjh9pPKJws1s+YlNPWAVnSSGc1nRHqQwHzS21b+MtShkZIIwuOaFonKxo
hohCysRh+WGw995aoVFhufjydNng2PCsAPWYdMtovbNgvmXjQ/83dRx1C0+esZ9hiNTas566/Z1W
54cQGlbAgEgIujGSXgQKVcDVIDEscpdpA0e0qQVBfJ+t/yb5NM8cms+FBj4xTzpGqCX1BQ0xHE2G
niqENUmvm5va5mcG9BBvORsNfXJYsPfI56DFqRUWgheSUX+Q/48BgDODPxyCGboJVI7p6NZH3FDm
fQq4UTXsSupeL/TwQT/Un8+IF43Ow/7bz2tI2daJujKJX3muyprqJ9KYwjix6YPSjoKes3lWZv3f
8ATxo5tsLAbl0YdqLmlz4w2HFXbUsMkZndcNADa30KsoWyUHqNmMlRmDd9HDkBXa6YQcOYQU0YdJ
PoaPdJFISPQvCZSjNtRS+0Hu1hFCACVkAcVbp7nsq51vH2WjExJFIvfshaSOPE5yH5Eq0cMe41vC
EaSMFTbkcfmmYPY42wOY1zURichk0ybLSuKr8yjuJUpwIAR8BNhWhJLgyp/LPOFXS0UannuQGpoM
i2S3D2cfWPp8F2R7B7+gz410jryta4W+CYFg7A8cdjTTUA5KFbJW+Lz2IsJpximSbFZfZ8rKBQyX
gXuRJ8JUEpljXwmT4oo1VXe+z2f9LvVtBe7ZN/CJ96SRUfshvKHTFFfc+dd8m8UMMzf8dAZF9A2Y
YSeJaRRnK15LJUQZ7cig1uQPYN7/6+OGt559ZD1OvF1BNukzFozAvmzI1gyr2H3q5O2diJwlFcGc
Pa4mm9Ti3wiIAI3CwuBdhNaxWrsWt8EEl5hIkCqRnKMdgDSeUFgF6nNgGR+nCurvDrjO4E4zODCN
wThI4nWr9iTViZxlIH7hc3L6W8JljVsjysZhSNCjvxzb9fAtcKwR4SQGKTtdf2oh2h/Uis+YYi67
Hu3Hj/VtESORF+6ayrz+5AFCV/0AnJiCfZh/vJW6Z52VdsxlRRmJt2HJHNGuGWZ0613iXNWk8aTt
QeSOi4is1SMOf/Rh4tvJg7iAV18uKlbNDqZhKP3Ht4ek8rFEXlW0paLhLqxPI2T2fOTHgiwiW4M7
46jumSkpQPwSOF4yyrWhKMvIT3aIsdb6NP9WulHr6leCysAfX+JLCzxPm5GxqZtgTBS4E49i93P/
S5a2d/uUI+iXD+Fps6y9KJesS5gc76QEvGL/IZ6H6gPK1elAKsYOY6u9tUYL4bez6Hk8WMUzUyAw
vjJBEwFeoF5nhhZ1sgLY84TJN+8xzDTrbppvFud3zx9IELNtW4lInrmt0ndb3o0BFKAmFFD3/UcA
MCUUH08jp17bWglIIJcGmYrySugvoIeX9coiip9c2lrjgIPaJSEQ+YIJC1JS9Jta0dcRqZrT7Ww5
WSsjadFYD1WIxBsWO1cxcpB9xTRlAHbmq2HpXXaWjRArJDUx/hqAoF9Ef8HdvoQr1iSvNhrBNNsW
fTw38Qm62BgC0Vr8tmGYOo49fbya7WMHYepv44bICWVspJVZObUxgwWiKdpedKY/Yr4FF+KbVRP0
d4PpAuFUM2ixgyH+sRFfnnK5dqvjAKaZRV17LgVmt07I9SxCPN7/Fb9+krTSlr4ZnySZLd3083Kr
o//RAI3NpaoHSzWs32y2emMQzgR4V5S6foNRV1kjeuS6tkfU7cjnZI3y4KsZAqFjz2K9uE9R4/K5
4f6OjXldFt14Uq+hE9q4xnP62qw+m2Iko2cTcCo3Twg8CGsJZ5GumJht49Qh92yaZfgop8qbinpf
SWphU36oTzKl8Nzbsb//gIHzHXoMmZv0kFP8XpOP087N41+bkpZi5nlU642jER5etUpSvX3avaWa
Y8mj+D1ZtpG+Dkl5/giNeyQkzNtS+93kNyzyTrCBTqhw6f9z4Jw09C07cKh/y55JyVIKs2Bmj8rE
2lTzacRJ+dA01RNcyTis8LqlzqLxG6gszKOpG7w2wMD5kqVmLPRbsgWN21xIaF1A+Lkh5BBjbT9i
PmoGx9b70Ikx9eQmz/9Nwvd1eaRjBs3l7DZ+3LF/pXiIpiQClO9RZrJJosEusTqwJvXnFSfsU/X2
2mTeSw/HzZxo6L8ofFR8FBNnriwhnt/0eaCnF+HaiqYXRs4J4L4hn1YvJ0ljKF7dCd7O4OiV379d
hNxdU128zopEpwvOjUfdU3SShtPREVSsafu2pnLS+ZpPwIQoh1m5fAJa9+3NnSgQP/t/4lP2Ldaz
6Z9+SbW9cnWVkM6OJFsVAMfXHEhqbGHfO4ba/9lZ43SZYOVwDkgBSFBGM2xd8qGaobdfB9olJnMY
lR9ALFuC6r6TMFzqBMti0MKh4UPX+wAAB6HMznUhRAHghMoYDSNGu5re2VfFGJTdj7SZu1rzmT0I
Vdj83fGYO11FMLU2sYZmhG65R6zHaEi9lSEhp9HjLD4hOF7st1o8NlqUEpthOn7wISmy4v2qprSo
yFRHOkJj2IZm8xq4SmY2jrpqTq9Dgi0PvIi1gcgmUCWSVRhuNr2GLjMxGvAoVrIgyVFSFrv/E8RJ
21lAJiHTl5y9ai2LWUhVs/O/gDyRVHqE+av+8FFJ9QGmNUbjiVuXnYO/NFkXMhU4SVQxe2i5wCYD
L2DLddtzigLGODol/XJTFFzELsLSO30YxPPrFgwZtTrjD0WMapKJgyCbT4PGqI6Wm0OmnOXcPUoq
BIVmkOpBmbygIWA9UBmf303Ell8EOEqXiBwLebPUEqGz1862//lsBwzuU22aZyNqcMBFAEP9gEqJ
iLYvThPovNQW5wier9PeTzk4n/vV0Dt3pkmI5Mqm4oiWNMGTvCfs/US2XHldGQD66FKS7seor+i6
mYggcD99+EHh7QX9CZkDnX2uV8Xoj2Od9dYWTqXpteBdEN1Wrw7rp6A/Nz6Mcf397KvZxUiVDJMh
/qjrgTaFTCw9tqqRZ95jw1GEja0tK10IY7V/dlcZwyViQqmfB/tSkMgnF0P6phjJKeSdFJykWZR4
GJn+//nXDYBotC7ylhDNEIAla4Wdid73hWYnzJQZidKPOVfQFxT/XmXjFwFywqJ2Hi34ptPFmBIw
e07Rb5RiyEfHf9lPJVt/YP/zA3EyASZ6Vg9428uWSzZeQyEHVeHmp9m7S1QPZ2hfSpjG/QXYEhnd
+KUTTD3d0AEhT68EMZi5H6aj6Rn1xpWmWKPRqHHbjZEuDeKsRi8GW4XdmhlnFdQK89Zvf9dWgMKL
XjEcYvbgGCV1ohOEhxzZnb8n6AfGgkqgVS5bJvuGvKda/sEsEtDY57aPpR75dhaxm45wPObBZPPt
L5muCpeXpBUseuEB3Qm2vxwCf0CvKV37/GUUwvXsyyFPug2BWfL+fM8uC15CBw3Bi9d+nmT+bFEd
kGChyv9RO+4dltRCC/juu4V3aPT2XJ1uEDh4Xxheaz6E5SvV5OTxHrebJ3v/20VMQ9hz36fZ8qVs
08hzFUUiozCb163N1jXfkoXUkUgM7bQvGA+pViHmV/bDFuD4KkOEbJGBlppIA3D25+++nprnVa9n
b13OrA3WckOg2A7tZehipQGqT/9mO61VjhnNy1WpvKQgCUazmX/Ch8ogsE2whZCvprYXDyS7tZUn
sBrJMsJNvM7Ox709O2vHccJVjZyJW4JKccLIwIfjwgDjVINbV9ACSNjDIer+04jI0iffqxM36WHi
+C0fYz9w3E13qzUrp2GAskSf1wNGRZXC10k5SGcl6a7ufqQRzF16bK8KLkaUilZrbt/jviomM24j
sEIuQ5jpArw8+7P9xEiGIMk2Uz5RygFjgEt7MeP1CWAPqzCFWw7ln8hSZuB9Y2TfTiWO/hu1d86h
HBOXcTHfIa7bunBBCjH8ZLtRldJh9Au6d/bnim347is+co+/ATvYK91z3a3y/9Wgkv5gHCwRtj1b
4Bh4n+1fozFzYNlduKdP3v/XMovEcbdrVI2xBhUsTjp9LR39ZgCxDGwF/SYmSZqjYH2TNpC0B+vp
jMJFDHfB1EhrwRKUTWOUU11UZDMWDcp1NLS+LBiG3jRmZ++SzaB2F4wzHiLonv090PXt6VJVmCP7
n6/LG4xOoePxxtBGyIDsWpjJ4ZPzgZmklrzEgQoFjQA6ICY3JHiIlZXPrZKrxyvIRUj63kIZ5BeK
fUSZK0tygq6HKe41PB9kqJ8Be/tdMaPKWm5/iX2peF3kVoz0HFa60QmK3rFLFOxA5BxflWl6Tevj
PaaSo0y6XJilf7GqZQ5E8TipWpmV8r8ggcFngYaT1WOkOyhA03JkApUOu24FckRAK2dGMgBVzoGg
8XD5Dq8pxpUoZH9G+DYDYgn95uek/+uct79+lF9vGO0lTW6JGqAc5i08soLTwcfR/Hzu9f3SGBZm
LD10q28vlCmMTMIbM6N8gWonn6QFkZ4iDPoe+ObpH4RyeAwl5P6GhTv4beCx8XM+hz+6D92wj4oZ
+JaOGZDjNx0pJOBiLCg7oPVriPn6Lseh8qHKdehKdbmVDSw3hUynUkJgp61s1Al1u3sRjFmPxz8D
hrC9qZMsIr2vcT+0oaypoMwpS4ZFs5ESjwgZUMjCNaMBJ9focjrdw5qwOMFL94tCXyQBMbvJVCg+
Oio1OoBIlEt8ju1OZ1MERzsHqBKud8CyUDkGwTqjqd+vUAhshcGSRG+fMIAztuarG0vCF4w/c3TL
q+jaQQ5EgnBVeyF8py8UsC2ryIlPYQD6wxPaPyQmPx+NCWtNAexrqdxMPRLRGdh0M+8bxxC6vbY/
UT7EHSM62LFBcz46MJJV7xcLRfBvwunhq32kcUPDNEV1uIrW0p8pau+3NudEWCaiOfMjvb/oCyIs
7kakFTnuZ0Ch5O7pRZ8x3mb2bGR/G5PxWH7dVk9I0JV6JhslVi4GUYI53fU0CWQ1CcWocBoGTGdu
2HlJLFmr098wEVFZqR0zF6QLvARhlk6CD0kV1maPYoaBiiZI4jrkKDAEMDkfwud7JTDVdw0/mjsb
i6+vrXkTORAGEq3gE4L5Z0JmJ0zYNmxUfi1QS6ZwLy4j9gUpAKOgF/TkI/r/9uU7yvdrcRbQPOKR
tLoRJyj+QH9R5wcZ1xwbgjkBr8TWDdhig33TManGee2VZe2w11wSExKbRdd2VnbPH/bim2w5Ebvw
KSOJfv09g47mvNVllYpPK4Eqo9CYRYOc45p1bYqidXM3a4jAqkvJuXPoHvovlijVr97Gw24BE4kF
LY2YzIfgX7HGf9KTw6GgOCTtbrDOdvwl3CDQyWIFux3AYRabaAmbtdfFBFjLxXOLwisQDRfEe1j0
iCJgSi2tmPM44FPmVpSuQOgKLq5lUr0P7RqdDyB3W3NpX2LaoBGq9T9mGmuSYeTWhNUGmY1ny/Qz
yiHBQ7WcTHI2/jERY+y3xUCiRvaqaxLV9G5CdZxgAOaIK7QqlpAuyoJUQpErinJK/ZNisHqcgRVD
NXZOSOFOInQTIWdRpr62p5r9Y1aaTlBC6F70DdkYdLnvDaW4cZ1raarbPutSW/OdvkbEStf3PbNT
Cdp8OM/oUnyQ5ArvemtK5gpbkJg2Yd2QD2d+T8uGFsSCorXPH/hrcqfzTdgBqeYKqlER9EsToV2R
ZphzmSk7FD7N2/b3Rn+b3OSzX9r5DyQPRA4WYH7pjvzll/2yR8pXP+tryC+oAIHZ6Ir36Q4bUftC
1HrNOXB9QbvqgPOoKgOA+YCwelCJJY8CAxYuPb45ZjuVEYD8yIYT4DMSl5rX0/7qwTquzyf5r0n8
XgZUV+A3bXTctVDgHZnGBaGCCMHukTTx+ffV3f/jIFBlils+zX4ClmHuzL1wcs3ED9o9y7If5UHJ
9wcNB6xrklwcPcrG3ka0R6R44s++sqAkSeSB2Y+D2LjOQCf1UMS6hkqSpNKqgstIgGxd/O24vhiC
IGZchRHqMywdARz+3P9OrHAXUYuRw2OHwhG0KPcJ2NkOFZfqz0pEdZzZHgcSqXVoPYyzf0mVfRun
EDEWawNO+HKtPLVTyo9lQ9UDfikUj+4EPCtsjDYMJ8/Y1BhTdmNYx93FTLI3Mdl5eINgiN95qeJi
BUpmosHuLS8K/6/lCe9hr1cqur2IutALsEkXoeipSTE6x2qlm/dl+AGYlahZFczRdZoxpZnLrFf4
U3hsGc8XOyw07E0mxFJE+Chpe2WON7qe/darvUAilodRpbWOtXWTv5E57BiX6vODGB3/ddImCdlV
deor4Onavf10MZSj9yy6mbwG/PNG8a9Jov+wagyUXLWL2+sF94+8CKTMbDjSQd+XhIzhUEC4Re9O
N2icDCW7/c/3TBe5w43CIKlVF0ktixed/Y8FZzFPsDUk3ZIPNdtLtT0kWGgd/Kn4ILyROm7ULGa8
oY5QbjSYe63VU+YwluY4xSt+lT/pyynhXZhW4dKQnvMWIIfO3OY32Z61zmyja6QSxqUMM2ExODhb
IBFL6c0t43U64KzczOsoTT/OYKxdS0xS1VZJ3MXHjW0O7lsLBK87UWJEX+LQw9tdAOleSc7R8uBk
2NdXvBypUBez8jNie6Wl8+e7vbIXFmbmLTi26ug74vV2sqIfCYpFGuLC2WAl89Rl2DqBK6SpTXEL
RYaKiMfkn/trcgjQWtkeqz8SlTdZ5ZgTls7Nb0f5fyL2Q9xJ7fQQ7tV1nODE27SCuYtg79pPy3Jd
hdQm/SepylmhrmPSOgc433oGDWVGkkahg/jmqQBFCZ4TTw5wTbAw7QYH3E0eu/VYncaKBYZnMo7F
xHerAdYtEMqsmDIdkMPkKXNJCdETwrbSSRDRVIv96IAKoMzs9Z6Y/NROzKyVoPTsEw/SNW2sn9dr
GFG8oRgzzfyMI751G/Z5suCeACM1ByxlBMxsRcXTDV1tLm6NgNDd0SiqPzSuKClgeomEABVRauGB
n6iKj0WroDAV9fw6AvaEOC9Xz7uu6XFBg/qnJ+S+/c+R9VAOvfV7HzL98ajW3wZZlQcEC+FC4GaL
ADCyZnl5BTVncCnxXF9e1Z/Y54g+LHbdSUnZteL50eWU2Kzv39/69xE4UJigsFJqW3YQuk1YaTef
wHJG71Xi5AAbr75DUUZh1modRUAQBJ57cTuO7p26dpbH2MPZQCWch0nfjI8sJy6tRNaHAcBlcJ2a
/zv/kdauUQUH6u4CtrxtBBBY0rJ5Fses5PKHFeApg432CsDgi2ESF8yZoapgNL5y8hETzh3sE3aN
rOdAonrlvl+3U1y1Mrta7CfROWTv/+SetvWDLUMPAeyKcSTCJBcut7M4GC6iJqkRU/769ZaBYbE0
jvWtd+1YRlrbu4j0Avitj+6/26LwF/7DpjX80C2ri1p90nzUWxysES5vHXffKCATzF5nnq7eNXjs
XcWVzWitS/+MZPEUbAhDKeHKs4x4YMCYz4ni7KyPf86m0NOxtc/lEuZAJTSYlNAylwEFVq8RLmr5
DgP14j1N30HNJhpxM+PjuvSKg+kyPrwdar7gwwuzBGLC225/93U7Wiy6qTZDNIwRN+WHML5loaZZ
HInVOsJnLqXuZBg90Hkctu1tSneo4OB8zQolWWbB0NfLvo8XTbBxn0dH38myqyDXRpKrnISF9xDo
rG2bXhQQWKRJXxO60p4E8fjEb5MbAvn3KxcWe5wmflopTkHhU4pahL2eor8Rr+qrOV1bjXv2zv6p
opC4iLgsLyMCoW2s+g3sARF+AQcWMgkLDN+/PzXr1F6i98F+sIi5NCBOz+rNwnWW3P3gnVGwRrqO
AJmUDP91EjwMCrdPLX85Ey7yWUk7mzr293iP8SEU+BTw1jd6YVsRJ9FWwwUI/Y2DLliNLLEXWwyW
ebIG1FrqWN+NH+4WcaTRw9Mn2Bv8XFef6ZNQ2QD5j7NlS9xB/4TgxlS8A6l+jjBuJdRLXR6U0Tur
kzD7uOURB0YzswMEIxhefDYvBp0emLXl3ooBL9RnqgSiw8WPxppHIAgHBfp4MRTzm7V60C/nQWod
sqF7hruYPmSaBwt9HdUzfnQXicsSEAlkNwd6HmkPupGPfG0q3ArDpGSP4gRNaI2vU7/7gwNjWTx2
jAq89NDKeuMaF/69v4aD3+WxiAEDQOHPB2nEc0FosoGSlejJI2T3M+fdtxFhEwd6sLCbpi69hTUR
goSwQQxhJmli9yjqH3anorgqjwg4AUh6sFUNVKiV6gHeP96PJn5ECbW4xyCpawJedj6j3r6pAZ3n
7AR/xHy+JXFaqpVdwpR4Ar12wiWmqMW9qxx2ns0I5PP1xgpdcC/CoxbHBYUhoT+iDQiPMI/UO2Zs
Uuqx8Xy/nPHqYI1C43nZP6DzOULOuP7rzLM9YYsuoMNY7knVslyg/InyV4Y9Ep/Zja2p1H8lTGqJ
h22p6yHQODcOUU/JWU4o6jmjFrzfRgCrzG1CwiCXENsqahvrWS6/F0i66DEWckE2qjU0gHItP1g/
W2x+4rNFUB1gTRszsQ/LPbArashiBUG5cfgozcQGpX7YRow3z73MbvBBzDHWP/T0Mhlh/Nl34KpO
00PFkD1zw+XJbB6iQXFb7daOvcMVEa0KjbsT7Irb1vUgKW/GYbJfL2ry6JE+z4cnQrnUD5b4ulzb
/LuWGDj2AMT2vfbdA+UHkXGP7XGaNU7R5+e6WjxHku1aNQLJySa1PaP0hV49juz37WGFXoh9jqqq
xTCNCOrsHwVCH7IvW433uPMZPnOStf/MrExwNjAc5Zh5gFcJddRvx/gi9ga3fgDZx9KrJ/P517XK
Xy6MKrcC89JYwWNktJlNj9kHtu/5cyfRapGRRabb+wDdQpfE2rK+YV4PWyiGluwqt3eajILaY92j
QCC/ryBmdMmQzlXU7Fp+FQs8D9ATKupzCDwGcDZhTfnNC0oLnN5GSx9zPguRJJeHBaptQuE8zFlq
RfG9enCxHxIokkAb0mEYMRGS1XRGfJHu+1EJ72dGScoZhaLirFi0vf7EGDK3Hrkdz2Uud5h4O0Sx
Lp6cdgtrxq0OwLRGNw2CpWgbC/b12B593qPdM6u5WiytBm5C4LzckHuZZHqd11/qKy2LksVTlOKb
r05QsQC23pKX1AGB+vQ8bWtY8OptvVxsa7UMjwK5VHmgbe5TUyY4Zgq9OD49ppFGA1IR7V88m1co
4zZn3/to793nyOTWhYEPw+NV5mhlYVeBOtuWvkHZda0qUQPG2DwIj54bn82iNC6Sso6Ay/fi9OwD
IlMXcFzutCcvb7d6Sk25vutbxOv5PyD7MnCIRxVTypO5Ny5vFHFCiftaKejlILfc7YaJ37gCg6V8
I2k0FsxteHL14UsPiCF2afjXEfa2tYPuR7madStK1+SNHfkYiMqB95UsMhwNJlXTkKkfW2j+I3VT
H0Jf7AQteaxEfdkq1E/drP9D1c+uns8Cu2xfeu3fmoNYbskuuu31bNdkk4HoBRlMus7tnIChquls
RqVB1RNS2VMdyvmmfvN1j/mHHDXghCfl6QQzWBb+umGGhdRh1iUlYeHjzbCJUSsOOi9Q2csQ6kt3
30AcIxpb9aIUt1SI6bekwTLV7sJyQKjwEaNEu4kWgqd5ufVrzeANenx5rekWiU6UCS3rtnha03Ni
NcVxcIezS4DPSIjMtTIerLTOJZ/00ELpSi7YiIOKI56rArGRj3cy9N3Lh6XZJkwrNubVqOl+KNWv
8Vzn0GFpP3gqyIJXtZFG6OGr+DxSTGt6qkKDalth+5W8VJTXtk6OdBSCKJpn3T29rN8VEG/hUS5h
Lce+qOQy18iDBwXeMan6UHdRo/sU3ilsJC5YK5waOaELqVZ50dww2bANIazqlIdDSUXxxc3IF86r
tsbMa+bNGJsca/r1ZJX3res7EIxt2W3o7rKW273yqhDzDX67cDsIEqd7vF0eKCwd4CzNCh7rKv4C
ScaEiFy7aMtdiE2s2F8+yPtG/bmEcmorjqcWNUlnTVuEc2aijuInP8OKEqVpzqJM7Gt9wvEhonkR
qXte/br//vZXQBVvZvsQEl3ahNzLPBEyhRWstgajnRpjt7BymmSroaxGxP5AE2nZOoK/o26PLLHA
UEFLtwXOKCgFumOFPkQGUdv6jRw+0Cq2ydQ+lqFes9xTNUh5NojmSMTd7uX7Oy5UG/cEr5U7Imnt
9FV78M0MMcT16Dh8a/i48uG7NNktWmfJwNTiGkhLB3a2Tz2du4MT2+TU/3f85hvPO6OPoiCav2c6
in4ygrVEgaY/YI86DAWe64rsNIgdZ4U3XLykkgJmZdSZUckqfXMxbFpe7X1pV53lVsjmbDE/bSeN
VyU/n/y/afHS/wsJw46/py/ZSLUUTwpPT1ehLe/IFWiSfcDGcmw02+BrzgOJzodc9ug+/mPc8hNv
i5PZQJs1dWuqxSRANlHjEJRXZ+Pba2X6Hb2FI4XJ7hND3Dj0gk+bIpIFwSDDxnhSi1IPFbVd9wPO
RyF5B3HXI3QZsTbQ92/qJpZaomKNJg19KOFVsPUCQK04ixu5eOoVl/xmfue0dY1jvHadu70JUW7T
YQc9UE0lMfOWMNrShPj7y84tkqzFOcbP4ptOzNVQw5L9QHC20Jm8NEjLk9tV+GrlJ/OGDs6VJIG5
AemDHh4e6ibkoMc1w1qnq8Ix4+lbK3Ls7LhLwnbiZ6PO7c5f8+HmuHydJ76X2tmuZdPW8ewugmBV
8kS8RPc+EbFDXZe9Y0sYOi8ReWiKUgo9jwnZh1KRIQKf3Ri9T9Bg1afAcysBHmOqCsUJ9ksnmcRb
Y0lleZ2i4OulGwIZ02dl+EWo/xADliLNvMDwSytSUmqN9LFOUui+P2rXOV85xsl43eI5XJ0Smwj7
om7n5S7LAeQS/3GvA0iP51l2TzlxT8Nt0zfZ8+QcMbRHOV7f85Nef26QGVnt5S37C5o8iJi3JEsy
20NRpzL0yT4GMWW8IoPZ4qktwpOVCIozWXQ2oP5s4qIs+OKff00WNmT8O0C1Y0wgg/gCFZPLaqz3
Vj0ryMxcimeDixnScEOMmGLbimbR3Tr4389ALmgWIC166CqNScUtxc0k7VqfNzJZPntjiYFtrSeS
ul5sjSKBVCf+ZXrvuSARlPVgbUAQVAbppJDN/WWDkxXuD/9s0psVk/ognKPR1zBAygW1sZmX/wA7
oaB1FCZO9YN+RngEJNB82GvKRoK/rVQJvTneKZ3VCJ5S2HIdp1DYHkY4OljVb9GC+2rcRHtXu7+M
KIxHhqdZP+pG6pNI1izCJQ9EASDBNXmrvzMIgtB/RW9Lf4PTfgBT8yZ4CVUKrSUIs9fid9N6atQe
p3X77SbXgbn8/wSBawJfktSvqVAXvGcruaeLWD6kLQGmpFc5AfpOnmmE7QUG8jR0DDPh1rOHUENe
96uadsPj1wQko4UOOeR68h2WIwvQEGW8XT1yyoxEm98zTk6YndHHtde6P0F8xQRCbLM0uD0Rp9jE
Ui9gAHxdZjn79m17N4YfBubblM1WtQD1E30xjhqY1G0HmzDQx/uF/Grb2qT6WjmcLNMK10/S18MG
GJS3pGfObc7C2WlRiRO9wo9ws8DjrwDeIB3sannXudh2M1TK3ttFtf/hEyBveJFNb9n2o4pVhAtO
lnu5dAAh1HEortEsTmZK0T2tvcp+uky/mZP742DaOOvIyj19Bi9X2usbSi1TUKrZjr8DBIsT5ivt
l40v0C9VGw7qTtpti2SdtoZHfnrnraacnrrPGvoSPgat/lRah8x3KAAXKxlp1+g6eiR+VOGyuzO9
vwd+VI24XlgviAM6u8Qx5Q+p2RkwZScYHnMcIoQ7RwzdJLpQr26y/MhsEwL1jxdAKHP1heABAcAw
ZPAod5KJ+/Of1HGQ7zJ7d9POJ6q1pe284F01VM997APIQnb/G+9l7mfTXhOopH8QjTmzQZlbehkr
AFksb2iIrPrKFj7X7QPE/putK9ynkRELeszOVcnKap/vp/7IThRcTYYlAfJXLcS3+GeugKCYICyT
pnFSNLm77AdyDerA5KWx4gQM/ea3iNATrm4IWNQeLy//MkZRqmQA3mmb6Bf/guYFRqGML0qKSdfr
UQu6RQgng6VFU9IztFJVYPt98WlCCyzI8tgyrgY0IcKFcbvAs9A5Hz8TQ3NweTCgwNsKxUzMK5Wb
PE+069WSZk8xvmdXgK9nMTtZhfsbq1byQtAVOSdescLgNxpUkoIsv+E0yURBx4Zz6Aw2aUrAiV+X
oJKZ3i8fSLaJyFbrRnbGDxRSPbdjNNe28kvy7yaY6Hdew1988u3GcblhSc8pcleDSrkDeSMEQLE3
7nIE2unTcv521eQmWXdPEcoX6SjBJg87jumRdHUOuyhFPLWia0+gDHYzcVUg/mx8SaRMjap6VGyp
4WfqI1o4pMb/H7BoOkyaogvRZGFsA4cUtLQluchZOvRMqSduPapPlMcbIwmZvvBCUN/gzsgma4wr
+23BbAQSH/D9mXq3WMAmmU4QI+Dp731gQc4E3MOovqxvFrOGIchyFcMf3EJghAu93WGwPYWUYmPS
wnFNKf/Ufi8+XMoP9Pg1K+LpaZmVXBz7q4Njj4xw20A3GM62wKTgGml1NaywmQ8kwaNpBQL867wy
1Ec8s2ae3jrF+cdviUJijoOE5JFt9LSTO8XgDY16aCqP3+a7PLtSxpx35H6Porj+Vu47iqwMvhCD
dAXuh0aeuQVpIjHMOu0bRUFRz8c50rvWIaGDGboOBkOz4I2+DUIUNDqtiouUksKLlbY497sLQgC8
1AK/SRk71YeW7S8+OMj5MYG7exAxKImJfEDSONtAdo2VYLD3dlcB817p4zcJ8ym+YgsfIidw1N9X
ZXZGJpZGG9k16ku6PEji3sVh1bEKk9YLRpsT2a8lry7P/9PxkTXigwHpx72jGdOWoN8/vWX86Y6A
KMAbbSZ++SHPJ2NGkO7z/QW9w+tbMh8of5SkoxgWEsGblsOyjW+MEUAmhLqXNUydH7kObJhBKoe5
6rJDRDaaMw4yQXeG0CKQzoBOc5htZYT8tisBxIhc6D0S48wWLf/Q8DIDvsi9GAkUnq4uvICb80QP
s2VOAkO+TVSYeBKhlTmqMsaw/GyAJHh7q0ASHDJ97mbpdgSM5lM/Cfvhv5VvYhl7njJ0HcaKjaJ9
E6UK628jdwWkzfBBz+YhL2QjDF8wIPKGtON7UYtkEvVwPxQCImUcpMWCoiAiuvGDzXF0rpAaxlDD
NsquidRmqagF2VIoo7AVBXmoz4MMCs4uiCrNxFTwzUyBDU+9Ujir2bLwyntlGWyJzC4tycdfg4fO
LWRiMciFehK/Gth3ngHsKqx0B3pmVBQo8JaTgoEP/6Am5nftPPohpImfWpcR8K5ykakUkaYkyRTO
0sfcOIQT0v6cX64+F2Knjx1uODCs6QiK9RoxcOYKvJEh6wqs0biEFelHYXGT1W/tnC/uQK6lbce0
7jCuBrodguhqds99ZTGbJ9ADyjgnknw3QvkckVHsE/YQm7WgUgSdeSKvkC0frCaHQUsMDR8afUwJ
PeILgPURVAOKH6Bs/u4bqqVyHDw8owRRM8qyVZcWeOy/nh+37gW4Dn2eCO41DGO8q7YPfz9XpQTa
7c2RJFx/qXExP6rfjR5ryffwZC/5DDgAwe7DhR1HbrNXAvV6Y2FAbBE5DR8eR5gaYOCKVcMNfv43
6CswT+4LXlajGUIfhc8pQkCh/HMp6a9ozo5/2/+7lpJjgkOO2Bv5+RyOn3idOQkgKxjVmla+wCv8
UC2fKosAtHfgQQd6FN4ceeNIZqXPC4xaFqLKlzixwAqgkUGj2028oOU6q4gbQmXXopp+lkBO2zvc
XsO/0rUBbS5a0SKt4s7Wt1pl3N3BDRri92CvIGAV/0pAKlPgrt4JCK7O/zmA/iLGfEFX35Ulwfvz
uXn6SC/TTAyHW9c2xhgx/jXohfPAgu/Mzw1YXLohQK99YLmL+pHtYKwp0jGqLwTu4jE9w0QD2TvN
OTECRQgQUBEYGhSa+T6sNK5az3O8eslJ7Hj6aedDZIfZfvZGa/CPVzq0/vKu4ly3xwgBpM7aqvuR
TOZLsgrxObNLUHf/eBILPW7++La7P0RLNk2FMFKXpylpi6OWj/Q9rHaop9rYavg2b4Kv/KRo26mu
Ea3WdBnYkfOQ37IVgV0Q0Zdn/cUlr3cc7b4R68P+EbPb/IXY97r+8v9RWFpsQzyksOdoMwq9SmA0
vY/8syQRQXZdD78U5te/VaHCmJrpDKf64CqpphrKQg/S7W9uMRe6iOSgFOeKEsVKnQ/1mdBFMZOv
KnBAFjcKgakR/viWM/jRnObk+cF1XVGglJRxyjWYNwR2bJM6FZMSMCzKtTiNEhxrV4hMNOm5gRZL
rPG6p8MkTzI4MgrARVQyOyLGK5zXoEmr4bvJkvY/rFglhZ+hZIwhusOBMuKSJXfv+s65mANC6zWM
4Qb5Ela/A5HxhnKC5DDfJOtGRdeiYpsOEyEMpk4HgfAlNH8ZPRSQd+k8pCP11sQ//fh7WJaGqywR
MTcPXVAX1kw9bNBYSvKJruSpDXXaonj4sOR4kzfuxV7OS4IPthc2e7d2hlXCqTRDmeAxYw80NrnK
AY0NuZ/S7Qts3AdketrgFnqfeN9ENY5dXjWEtFIoFOYFZ4NfPKZwuS/00o+cAS4IRhtoZu0NTF5E
ng+RRKlWzVw1ZG5JwlNi7CprujgR0UpHeKs1NKkIy3Eafw2u/p1/0QR8Kj3z7/AyK8bF4qtVzqpU
1ShkwburhIa4yfwFLYqwaq91notEh1YRJEJ+LcN1+Q+XA20gAxdsxj6McJeeB90r8y0Ce/u2E2bl
7WJD+MoDoM/p6W0nL6e9v04Teru69OBJS0lIzy1Wtnmf85kHY8ieR6TVqQNohG25WQZadZUmKYS5
uCZYZwj/u8z3lFpyMixA00YwmjtzOuWCYmaHi5bOUq1U1GeMMHOpG4bRKvx+NXMUERZXDmetKU8S
/6YO1kptT6IN60PlNKrwt8+7ZpI1wm2ZR3sirF2JvfWpxNssBtwa5g6AaIFjb4S+JwTS4Wo8RlF9
NeJmZZvA4es7yWTMzGKPxAx7Bt9xmG8kZ8GzCcFrCWES/b/YtXbc3ndmlTB3e/qmmzaeSoMZBOya
ux/I0EC8DYTJgj/LdAmP9Wi1iaKIfda0Nbg7gOm+upCLhr3Nl0yn8HeU2u1ur2Ww3dC4Js8ijFcV
1THYzDch23tQgRA9hKthphlyhmWvsHPaSt+E9TN3ybnoN3z28tSnoXG9SlDCod486C2nCi+BSccG
ZV++d7km5DTBpTQJY674mK7i4gGimFskCV/dTwXnTZc4+lZb4pg4VpbG2JSdruNDVDiin/9n0w62
JWL75ktE7gmRPRuUZo0GjTEGqv3NWUrOkqaxI6qhv8iI2JBa076QN1nL4IXxgIkr/Vq+SEBp+cRn
jyDbKVnkx0ENcqgDH9ovSp7v4roQrx409uIRHE4JOLX8APlfjna9mmSsR7jIAYN0N1SekJUe0uaB
XAW5JfOc4id3AkNJuU/fSg5iT3KW0nxhsUA2J7bDkmDWY7xQdRGenPnKiampfzsz9qN1/o+bwnMg
YBhsPWalXh4irZOb3d9QlNP7OdFC9Gap9FcL6J1QqPG0ey1/5BfCARt8dpdTUvRJFTJlq62A9StY
kkRJpMbGgTtxCFrdRzdSiUH+lz4YIRxCXISTmuO+WIaNXRAe72Uj+OemFPTg0OZnnfNeJNJCjqqG
BRZTTa9eYw5WI5dbQEkuGxyarsqjQuqMK3wmZL1J86z9BTc3qNB9oSZvywFy2vBbrZ5/O1I0GQaS
sWJ0BVZFJMteGsCbu8sX+2WZFTA1tbTyFtX+BDJMRb2Iif8W1AcqQwcqxEGc/o6SgFV6z4uHREKr
1YaAgpRH8fl8nHscGhs3jlJhvqMfmJ5MhOVDV/AXg+Ylifcy44BAhp8Az/PubRbSpUzAvx1s/Z08
q8Z4Yh51nnGq/u4e/YLJ+A1IvIGaRMVxbAZlueEt1RpULfjwH2W4q+k9+U3F4Qqc+GFOke1ax8yy
RNU4P59f0zLwoFy7Ct4/Sastl97wSiSlL0An5QqEft2W+F5x3GasUy3O1gyG9CM4f2Mb8T0Rv8IO
eDeMBIQYGO48JoRixvxzVrMmYovhgmUtGvJt9i2Dj32nfVeshi7BKF2071SQ9n/V7SX4DWg68tgR
O7OAjRTX3AbFzX+2A/RDsGUvaw6OnZn0FAGLqBO7tw3jv7amx1i4b18iBauVfqDOOskKu1nTcNi5
pdhp/vTZCna+Nulbsttf/zV5e081d/qnDISC+IceGYSRNCjRmrQ6qi5+RoVgO5yqN9PK93tjfB3l
2t6/hqDi9eO30bz7k4MLpghvXIgtMdvK+XqY8l8PQfw/5IpuV2VZoP7HsTx175IBdeIJw2iiXmuC
zJ7IbqlEUP7MoEkqAAJUuR5QOSGVuysaQ0vO6S/bX9CthMGfaHcQ/UFOagiNvaOQnC0HMKbjR+vi
8sXVkts4vjvMfOLPs4rEpRalHEXyNOA+pLJ1nhGbEvXJ4Phbgcqu7dvv3pKxTV+iiG9oDUcO+sl8
zXxG7tY1EB0iHOnjZlV/7EJsVr71LIYBlzp7X0x88AoxR7aw2YpYk/9l7H8dtVzpKO1JbUaxaNho
O1vZ2TjHJLzDO35yaSV5ibX93PE3X3bsPq/J3fNiRYxTk/J+So3p2grASbscrzOQsyQOA9CElNOo
fCXvoepfD0M/UG59DCkF84hM/lE6UbsOA0pyPGtmHrqFNj2MvaWbbCGxRWUVeOz5qaDR6qARlL7F
Pfc3zF0ecOYMsyfgtUfxavkCIQmBgxWZt1zKSwleIMkF6fUKfkVHl5Rw+M/zHWnmeoDBehQucm5c
BaGpS+wcnksWqnwq+mhhFs2FajclNit+VpuS89IG4ElYCReVCRjA9zGgHpJ/b956MxMDe6WMZAPz
6bcrBTcBQPpJJIDyfENuDPsakmKDpc3zYigHcfKYw4ApUuVqx1LLWthfBMINIfHH7z4XdAxx98Rf
1mUGAV5UK3iX6WeE54FlRNiAGDZK6pfrJ9kLZTvhXfT06w/7zR0o3gNeP1c6NVnvWE+50QShv73e
rx/dSESXp+HoHRG7bTRUA71iM1/nDgjDQd+b5MpSqNy/YmKmnJOO2rOV2u/mmmPj3Dk3GwS4sJEQ
iZUfrpr1CAo4tIUh4799G7orUKLbaiwxYuibpaf58KpGlU7toaKaHTJeZVDx79xMBVJylkYRJON7
qi/tyOjOmrZh5Jal6kSTGVM4XF6nJXLDR0JsEwAtR7S2XDw84K7H51RrDUjPO+dtqlLRf+EySSiy
AiZxr8UEybWhK3MYFUddCHlv6vbUrYbOh3t/g28jJHJXUuypPWi/Fe6iNw7v6DmP4cPI9b7GVbAU
oas3UMnpkAx+r3hL7oT4u1jwfZUYT4e2KY5dkbN3D1ZNNnvs9wkQqb0MtVU15jlJ1XJU/GFc4JLC
ZQtRF/gCV4lFo4YAUJ2DIIOzdRaa/GTX30Npu33pI2qq1xlWSdkWD3HUQhJ8Yoy0foEBbh78dNeq
RXCJTVt0j20kC2x5TBu0aG2WboCKKDZLpkG5lB/0jZUWc1EOO316C6Oj5aMOGXFBbod3nwwLeFuO
Y8qOrpzLE/6xshkKJ2wUCuOcYHegWuvHG/JTRt5T5YkWlwPQmMV5ys3e7oFXEHwtUC/FCOww1fSh
3HEVdqBWjUtDxxoiMB05oth5Ns8an6K3cDQUjdZ20frqn0j8BCFWBFZOX51GEcnnABvaBrptvGCF
nsfdPBsj2hzTeGT4ZvUt/zT+CHW2z/pVDo6lY71NGeQzKrM1CvZgDqWrSYyC0za5uoCpK7S8/237
q1epE9W5Mk3AUVaf7D5FucO7QIzbOYA0fO5x7bzV5bxTm8QeZFUmv78KJslglumL1PLQp4+qffE8
k+PSDYs6qtZrZttoXthN7aE2QHace+bSD6Er4UMSP40N3wmRMSnJwbCYLtStXyaSgp6DJNYqUzAa
aZhDHiQaBOpKZw6vurYbOllRWbq70w94b4YnPRxl557m/8ssMjQ7ZhPTAcOVj9DNQoFeDz6g7x9o
vgWF2E/G0Eb7c6Lb3YKYab4F77OAU0HIZ0TIrXUYfuuA0yWb63a72LP/MDdYScxwV72eQN3Wy8if
xbOzklqekFMynbo/5fskCXUQkSESZuExx17UNHUVoKdzAXggT/6St7hwJ56cVsB3rqu2IHyINgCw
bvenFBQmY5AIQntSbs1YMvm0RZT0uWcqwo0oA/y+FgypNVVPxroVklDy7p/O2o/WPh3P3gJBYdBy
Sh05GRrNapKocmqlAfLW2EwfuXLbEl0Qpn3UEBMJKhAKBvAcGxKcRjj9W4ekgaPxY9Vj26H1/jES
0HEyti/Ls3WG/kAL1hMC8JF57GRqrXoD7H7awTnRW0v6oQFgQh/gza5lK+xa6iedGHOIN4XmQL6+
nZjlrEYargtf/Ga4TNCz90h8iDL4ltd8tnQNkKjgarvAUQsIrtfMqRiYgPpX1DmACVSLRaJIAuX7
TTboxBvG8C+7vKC9kXNweECfjOsd5tX/ocw6e4C/M/gk2N6dULwAEixdaxI6sUx+k8mpqanvTcza
a+P78FQeeNYcdLnX1K8KZI8/vMfr+4K7gLt/m1veAv9DgvJAHpc00TvfnluVi5NgDTuaHRLh0YJD
ZH/JzZcSIg5vursYNdA8tQozSWU4f0VlwchKxV3IpzKGukxq3nS9U5HaLe3bQv2qGbLZetjJ6kWD
pHKXxgmnqqSWWponoxXT578keFRPbR49lsmnpYf2b+anVmfN3wKH/oW/I69DTtqVJdiyRwJ3kvvv
K4EWCwv9tY/to3dBLQan5STOBlX35c2c4Kt7V518beMNQFM406Bqdc4fS8ecWqcOrlVqjhZtyQX6
EmOA/ehktYq/Y0GfJfNZ8aYkoRBPq0IGUaF/My0jefpnalTCQBBF/xweZInZDPU4GFxMtPsRpL6C
d9ZT/6uYK1+Xv27mnVEZTJLed6PbRW2jPk7lIAm203RPCLNhf7Q9lYXSHUHYEWoMQxaclNW0colN
TmslpiOZr1pugm8eGykrG+2775y1EYAAvZn3RKBIQ5YfmivJXJ80aw4sw1WIpt8xikmuuWrER807
2/FU1Gh8Er4vOi7DPwU0JRFlPggOc28inRJYHlIw/lUe8xC8YZHJPnnkfXn9F1nDvCbYfuMTpIrn
E1Z0qDp678mkRGRfjNuJNErknrEr2oKsiwdJ4SPRyskD02jsBFuwLf5FLOS7IjhzjRiwNh/jNynO
OUKdre2gWVXNAOzYOR4kecJZcsIL9TcUhXMXTFx9Fk+C5DwO7zRVjtSMizhXC6Zs2YPfil/Z5rpp
M33UhNoEDmUOiSKQBin+qGw81Wqo0QmVPcB+ZVPhEseaY0c2J8wwqsWggrb5iPob7jDfewKmlEGn
FtEP8LZq11MbPCUQ312yk6SA2zlgkBfL/dNJF4P6mLO6o5u6Q/ZeBs4il/StfBZ5BEYTXt2zeIv1
88hodU3A5hdnlzDkZ1aByFPZmb4Hjs60ayqJ0Fa1iWC1DLYBZWVp6Wnx6TFhSLHD5fPJW+LdFzg4
hNBBg2QhjbRy4FCKPfyBn0mDFdZR81y/ZOgp9Vd7SGr7JmciZ20+k5z+eXZGTYT7UnxjoUFzM+n7
YrWr7wdXWV4HJ8j65jGtd/oljxvBo/c7qI+MWK6w65IUyzbF6eIas6DkXsXhOGgSBOvWIWoAP7dq
0a1s7s8O0ovjKVhWLir6fiA7syUwIQNBGvJqRCz9fs3yUF0yiXu4Nasg0hcvHT+080Rf3qM0iNBh
W16ueaMUZKtF6V7KeDLdxHgCiVYbTtcYEbj620Ax857eN5vRwBA9QNspplLz8R5mGERv6ACZFshR
JWbNsmfB0xSQzqJre0hrDihx3QJF4yDCFFhOxPIGxxYGPkfID3d6ls/lfXkeCSMkPVsp6wt3OiEx
fcDG5MmEC3EfUlESOcSnGRz4HHNMRjOoEiWSF3eL77FNmFnyRByzyROrjmpyqtQuB1DST1UUUR21
Ksd4uzwn1mchAPI4f3Sx6SuWsLs1duXNdJvoU5wG34pvK7AzEtQPveUY8JyY7+Thqre8qh7kmmG+
P4KGwNMtJ2f755WiRojNdg7IQ7PJLmq0Ye5icZHVKI6VJDZH2WdzU1LTEm4uHw2mhxVkpxqa6xEN
sUvxjh4XuhriKxI0jYzkIKQcbDfsP9H7rAYxxtC9UxGoFP5lZARB7zGLlPuhbyBeRg8KlwtnawW/
WYsNJG4jHdOEz/l1JF+CQoxHsNmDVD0dmzqgrXDnJAWqGkVWwVKoHG2iXJej62jwX5P9kYiGj9mR
AB7a0y1y9bf4SxSUqOT0o4jLXn+WPqlwLAac8wzgD33J0qxNMHuzBbhl7XoTTKKaFuV7c21qhzes
Kjxyf+UIWm+KTGmETMNx4/QdMYWrvMCYzPr8UIb4r06Z0qxMhkTRlRl3gialnd9sw9JJcaa3YyHy
4gPzJvYXYGWyWlgm7h8zd1Z9ImOGuBiupJT8CCfDlU50pho5jJRhi2XxPbAELzykC74euoVXyn8u
dtxr59SE/I+lwh7v4a3n4HyotDnkeG2qwxqWuoWYDXPP8igFgFYSu47JCUYloLUmDHq8SDl9ggeq
G2eCyVCUQRKh4oBeyo5ncgDPvzavPNAgShGtViJTIrlZR7FfXn8lS5Lwz5OllFJlUqR4NbQxIqO5
SZ3kO1M7znRxgk3WUWb0oKms8K52x8z9G5LI6rQum8DW9i29XY/kgxPCg+CvPVQZAB07H5Zoa5oG
VJgjp3uNkgnpnTsxxH/Aims15RDso22Sn2p6cEl6bbwbVCwUb1JXQFqftHdrSlO7gQ1oVh7jNHgb
2g7P6R6o7n2OIj7V/1BGXI1oAfA4LFg7nZc5VlGgpQgXnK65edT54QpNyMdSXK78KL7OvYzqEZ4R
rIF7xf09lvXEY3g7nnvIf2cMlELRNIpzTDSce+TbyVWYx1e/goNUBcD4t7VXF0/ZGpLYszM8EH3c
3w4Ycap2qlAOce+o3C8UJLurMk4u482IaKsrNtluBj5zMGUZz4eCVbC1WZMSnp73Sa1tm556FtOt
j1FO4aGnMHafCWdBDnwi4j3PYnPRSSgro6llwaG0N5b7kXp30fOCSz/6FkBZaGRmiBuM3fjclZZ+
aKtNZDoETqLmYbPhcKWH3Ew4USm8/WrRkTfqOGQUQ7U1+8yvek3K4cBazVBsJWHJ2b4zJTi71+0+
QJFaxYxK2hAhcxIg4tC4gUm9quPnecQEfcOesHzsWq1Qx1cFM+S1WhRX/StmaV8PXfDmwNpWtiWY
fQhGmivqITV+3Hq29xYm4P/VxuL90EmSOmx76JSfBukhgQ3PITIVHH8L3mcYXPFVhA8S7/mPspPO
iz12i4SbVdUTHEzb2bYcyvCnYOBJyfh5Cyp7PkQcZON3leTsxFJ7DQvJUwFeSNDxEjSrcXC/F8S8
T3maXykZLpB/EeZWHdKOjrZ4idWsfoNM7OxHUiGWcF4LPjGGDdNoS9GpM6TRjEj8UllJW4hTYEC5
cl4Jwyj0tx/1Dsn7oFkildeUQ2ATTHkoJNlGZJj5cqmfnwtYJqrLJQmNAX4sRne0W2s2M1VB3rvn
bCm6x497YdmTI/FNjbSJ0BPYo5i749M/9pN4baCZbPhJUaZfwy4hmJHEu0Vrc+GgoYOzx+m0zQ7/
svsxghn3HC/NRoImVNNqoDy+7s4MWaF44qta6/iX7APbx0TOHi5h4c+pfAjFwP7hZz3YTTnnor6o
dOgurrjolk6KXWZ4SxXbDO7Hp7kE+wU0OwwpEpePpUUFd5l8fiDLj1NKV9ksItkJFUb8G2kxLgdY
Alu45ghhcdG6gpUYlA/RTPoLXFeyF+QJkPnplHec3RSkopIwg42d7vjq8XgDLDRT2xFZglxuDjWC
zciUI8xfA9IygMg3415x1T5ukceJg1AN1z1GgSGXz1wP6Ts1nxSLIKtXaP02udMtmOsjx6cq7Qwv
UwPWUVCvw+AxogYejzq4Ks+bnQ2nxJ9YOqA3jLgv6cHFnudmjl0mUOK/Vjn9/pVRqc7Yeo2rDzKM
P53QnUqAw1N6mBysgzCLVrBA5G+V/zikHfgV7g3xevxZiSpv0p7RgzznQ96ExvFW9GYRnYtsmZW1
RMp2e5nptkqlrskF9VxQm1mK6/ntkQYoC0UrOCidFc3dSyRHGLvEzQal9wN9g2xY2qvc3R3Jhj4N
0cBqKQY1DCvW58cICcp5CozN7t8ctgG61/CORI1+Z2eHHBMYxxMHWutHBqLKErLlWrkwIfj34/Pk
iCRQRKDBXk6gU7g8FVF9017s9C2dJd/AyChACp2XBNVJTfb3dd0KgZR0ADYo1qQ9OHJhFSg+i3cY
TbeGdeQtjy35tyfh0l21BNIAV9IrJjMl2JcDgo+IePV8+URd+Ku4QqmaRDX5XvEHMii7qtb+9lI0
s1Ag+/5cXNpEetFpvR/bwioBXGwcKRPLDJmPo+/yvMv2NP4vbDfZE7TdLXW4QNUY4lwgwZ6MibMS
ZvyamSpbKmwzpfTieEHgh/Agfz4L6FbfqNXx3sLVuX4Ect2LroTVjmT4kqWR6otetKKskKHxvm5i
ltPj3ROL6WeG9qI54TPGRy8TO8FYUvvOzmucKnVMPEvCvwGAeEMplaP2MQTovASsDjQUWGMVUnAY
L0ZfVQGKGQ3UiBZFMXIAjNfWwvQiq88ZVyBj2OJrDBhNBEjmvWw52JtP73Adz7SP8wYejvCXf3xR
uT4gF8yasTKBOLqOwKg7pfe7eOQTrWIAbQ7M4yTGQuIWgt3Nur7FEW1fJ7f2/dOakuKYQuJ3rJ6I
6DqMhFoBmZXbyRZ74nA8NcLdEWaSRqywvWbFckRsstxEqPqDHruSueIwqEc0RAOAqzecfCecn5G5
9bwjq+8sJDz90dw/k86Fm+HRr7tRcxXvaPdG+RYtEblOmAsPKLH2S5q+ZDgDc1DymnGzjgxQ5RGH
Tt03jMip+W6SvwC2hVYQwIvzJDMii84umRbCnOEaaCVgEicGMfehOr6RTzOvAgfmDdAovT1LGTIQ
wP2bXk6YK+RMolpUvoN5M0Bt7eo7Rv8w6qN+GorZZ0Xy1JSpXWruC03+iNE6wO3fciBNyA8WBMAX
ke2/V9/bWtV2QNFL2CyY/CIrL5sfjpinh76WhsxL3Piqmnrx9ZqiiXpIAfRlZ92SYoj4ujnlDO+/
tagN8Sm07bU3CWEYiuz+COeBHqnajGjFpMT4kFMDfyuqlbhffJba8HAMlUdEkUVcbCV3+CV/9hsM
EehaYVOL62ICy8JgC2ROabg0yC8jJHKUn/7T3su6nOJkzLZK3pyjTRCslFcbCbyT/byRU9/4nsNs
xhxOA1Vo5t0QStaXdzHBdR6qFblFp98qpenH2oJ7eoKpmPFjFrKyuluAwFeUNELqHXFNHPc4pWIZ
mvxq8bqJmbZp5pFDOlSmapEQEngvmavomR/bqhoXA39k83GcClewDKNm9c75T3XfhlC/98s8Yipd
ex3sNNgeMF6yWcf3MH8HxExfs2HIdwuXDP3DUloSQ0i2/I0vabAM+HyF0lMPiSbmu41VJAr+7of8
IUJE77u3iRFOLaEDXZp5Gj/TzKBM2RvNxnAbzrcq7JX6YcoXayJXa91Q6bqbPzaFll9CYL5/nKM1
1c1hGmYmC3htc7W6CKj13X7i9hm1JuZaY0RVMeM1XwKJ+P2+47/ueJDRD3sYmC52cQGOUpKzaa/G
MWFnFe6lEkakrxFEYbbkfpbez97e3n7n7SAAvrP068M49EF8oZsbOIfDS904ws6Vi5sMOSAyUjrQ
1ROx2TzebPjFx+inE3Qdz2DXJCM1D9Dld9cSSi7IkXJLBpPDFKjFXg3EDHuStE3lRMng5Ul/11Yt
tIcYTDd+DGi6jhKgn1uHhkYXunLX/nNX9Pdhb0JYGdHCwNo/zC2bveE7tUoub6bbZdxqs6qHo6Ye
yVTYFKroax2OcZyVDomHqv1HOAD2SoL00TRq1vjflSopDpkQDr6oZEotKywubfTW+tTDHq7SxxTs
Xxady+HLLNyiZZj/nUGbOf/gWpaoeAos/dj/ya1q9QPUafgV92PMZbuf7W92VdFBXBxZqYSOtN9P
Un/cffhTASc+o1IqieOld3nDd9buGZObDWhfZfVDm9183LJ74GMj0hS2aqfihqcbskhVmKCthOIU
hiJ1xIJjUWr9fYrs0u25mGt6W/w+MRDkohZravfyczKu9MwYuJG65YKdP5aFlbENTV8bJys2TWH2
Q7YiAAad1uCONx5L+WyWqAQKMDvhpA82QxbuQMiDHP8KyfYIJDvSPaJF1DGQMXlr0U/m3eYqis3n
i/H9Qes8MMILIYpVofPfOeu0Z7fa6dXWwIVMOmYp6qKfWKIQImSvQy0XJLNhLDPBy9qd0wDdY3pC
4ZDA0GtcfJv9faKpVwH/WI7pqh8BG/1gFVeag5WZAV4sfQN1GQ9jvLQ+6YWHZkU8Cst0Z85ZwEKX
BC/9Lem7bXCohgnQpHGEXDfVA/hOLjpHck5//xQoeTGdN6sZu24ZSpM1a0hOEIUG1TVpu/70eAPI
6uvNIxoDyD6fasTK+yKNCYRy777iqunjQXGbRzK3TWohjk/gNKTMDX1PsKTfmsa/GSpJG9+puVEa
EnYR3Kl03dONhgkBTljIh72dT+xKyXXvw76/pwhvTGiijl21nFojwYrHTc9A+TGqALBc7V16AbEs
vCkAJqNvaTKedoYjq6qJanWSDCZ40mElPVimEDpELVolVk0cy4YsiR+p1Hv8mCxHQF92tUZqMv5z
Nn8oZhu6tnIwYIlNe2QKZNjSg3wPll2p7bPkq9Z9SZI3Xde8/sDW60QfWQnir5wLioznr+3h6xDh
EUeSlvXRp3CaWsJJWjKde3a+7ta1P+50/CsQBj7wqZvRf9n/T9VlpbaoxGLDGDCBGS90J6ZXWkuT
HeYZnPgXvFk3eRC5Y1xJWNZFGxahRuzTZqFDdsZ8c9e78z/IClPCSkzxgwij+sf9X1ab89wLB0tC
dGpH/ak7ei1IVIN5cc6AEsmid9+izzmzre5Hk+gLxAie5wZbswj+EZqm866etQruAYAA+dYEzhoq
WuCYLEx5NEvwca93szTrAGLDxqKHdEnN5HlAZ2mg7+oMLHl8s1HBrlbGj4gpbm9OEcoBcFBHoZEf
IHDzq2UU+4mIvQEAkodv9Oj0tx5A4MtThhW+j0OXNM2Xn9FQkBXd7Wm1dijxRy41rZdbbeozZJtp
xXzaxFJkhJ2Ls2rnQJ/NzTYKwl1i+7Sm4E5qsAwCke8pfNiw8n6eWWkcFSduCspQGTMwk7hd0N+3
H3ZmCkeVUWPzkD/eltFzEDOFn/EY6nkCJBBL8Eo1ZMzDF5GjEkzwn0wxjV17guWoxnnuGbyM3jMF
gduan6/mHCL0c1P9tpYlos7M2sbwmMxHYjCo9yJ/wE2+mT8N7u1peEHqXZYsHhjepOwAfZq7z2Jr
u77EROpzmgIMTOaST88Vil+NlNymrJCWItpkuNeARb7GjhTgmT5jWJohRAppAfkRLUEh12w/CMeN
6nH3j+s3JuvtjdYbei7CvBT6jOAqjUNhFGbylnsawqgxK8UgDUTovlsU+JrkYas9LxWEeQ26vIkb
CZrQOMhcSpuvHOiRqfyJhPTja5ARKBDAKPksaWd1Imc3K67hXWh07D9rmcLracN4S+GfI3ljstO2
C7yc9yHIpbiod02KYFvd0cLOoMgIAvXQ5YW0JfHKzZSDfCZjjeEq8lpRsg7XZwnN8FWP/v5lVso4
ZgtYi2wK2p6WkLyHXlOcWPT1z0v7Ylsq34dCE2fjm/oPvhrk2t0WutZipIjbd7NqoTpWdVFrUQMU
bPQz8cNs/IsfGn/9tC4XbiPgySMSoyrnpsHwU3RfyMu6d19qRew4HVXUhynOueiFbETd349q3bVA
RTz1JpKVgOuL+XQS5oAq985kZsIHx5T1Ohg6Cd4bnpFD3xkk8a6XyRoExZ3gBtbL9AV6YoScjeYx
2Sw7Ec5nQMcwpZn4tqS6Co0WSzWggNGu6girAPPdwrVOI7fDNyhhAVNicHNsfNORl1K/Hdq8BrBg
2rS2byCL0kMMNIIUC7Pp1ASq06hviduPmfvVBsHGe1pW7D/Ki/+TP7NDKTTD1jMcn57SPCQGjvPH
u0aFEIoHIVv9H/4j/SPzfC+3jbMcJDLuDGPFxfiL5r3c1LjUD5IdxUQEoEEo6IA5sI15g0rUI7fO
6rw8LYbqae3ZZNWuoLOV1lb48hFGB8HPQAU6IMa279Reqg9N3qh9r9/Fy2aXccFpXbvjCHNkvnj3
mRwKF9TKhkRJekMgec5pXyhXZdeQby8do7CuAZKw3Yev5wQG1yTzy6jYtshBR7lHUriNJ0qlmn7w
laMw75w+vrVH8dNl8NuJW/Cs6cZgMtumr/UkOLkLT4i2npXSmer0FXxcwrKvsJBIo2n2e5R7nlIK
qmzhs6kmxLHKMvp6ADW6dvNFMVLUUosx4uUC04xJA/daMOgnd6lTMVz8SQ7TFTzuSwlN4yc+rDFO
IPq7IbxL72O5LFqOwwx3eGhvhO9Y8e3fOPrrtWcLgKm6MPhhA38NWbWyM0RjPiAtAPiZ1DPfaqg+
FbuJ+2m9PF6W9ZTmq5XixU6LhHyefEL/ijHAzbTKE9iGbxkglSgAanbF7N6qt6bw5YBUZYzDk8VT
LZ2inI4POWbwiRUqye4yfXHIybTXb/4iEdqGOvQ1J5CZZd/fmU/JNHqqE5/cK1i3wGvVqDga4L5J
gthDgeIMexl8cLLwhmZsfc9nKIC2CiGjLiRZN6IpfQi0N25J7BY7YJHD89XBFTFIdHqRHLJnaP4M
H82VnORPumYPJDM3PfPuKAZic4SUqYbuQB3ACyIPI2pN66rQ3rR6R5DsXfuwVPnG2SUiLJ1lUytS
nbUAoLoos7r48vfxi6oi8bkEgQRcx+k47+SK+x1+GIhNP52GZO83Lq0s1QtU+pYSuKrfYb9p/u3G
y1lD1SxU+226BQpdXhsxnciAKaXbxk145ID5w3rzltBrpzisBSnzyhoOLPBSBNtaevSUsjI04Xq/
4Un9O5Xj60IUB3jjfjIi8K6A0aDHdCJy614zR/rwnQkmfDI1INZkhgTjSXy1Ky6/cx8NDc4lZAYm
3+QA509Iz+hym5HkOp/ks0OCkzprQaGuhlCb+hiHkD95XZEQ/RlNWHMy6ojhkFRdoBXzioke3qNt
LQqpiyTu5tDlLBwoc0/kcs5MlOwDBXycx57A6pKd1WsUa9glAPruZrbr5hRiqtwx/REGxkPFR5l4
aBVBtQ+MRTILsndf9YuL/c+HNk8yZzXI9BDOqMA0YMbPqvfIsIi0Awb3nT8SnGI5AGtmuvk4TJLV
zuFMBwYD5FfLFIaNibmjkINH9FMyzp/QAqFuMVar8qPmvOTX2KJXYU9jaTBBDmw0bc/UXRzKefxh
ITWfEU/mtZ/P30cb/snagejtj0RvqFi4dBew9pspx/KPIfixBY+s5K9tTF+tiZevmrKMFZWcmRBK
cijWNpFj5exf08jqrFAueNm9PWaEp90wQvB83fD7rkGV6O2MrjrjZ0jOR7OZR7OUQdxjRYxROzA/
y/BF5W2Tld6NmWZ/t/xpURyWT1CgrXBEJo8YCGuLArvPAP7oP67LWNLvDAKQ4c5n36OBs+bAJHki
EPT/L3L+YRHXev5qWmiYYzp+2a7IEm0pXpr28ZKnbWcVJTmF3ILKc8dlT680pnijbxEpg+/urEet
+BuN3cUac18VuUVuugk4IB/dfNgKhKs3lkq1ApeB36AzNaHgO5tYIiJS1pUTN2OaIdHJMGsmkLND
Knp3UlS15giiioN3FtYqPgp+Zs8jKssCufLE/WdrapFXystzs8dyhvVdGwBXBjclcwVfi3iAPe4A
QWodfxIZPNlmeE5QuIiIJ/yURTTNxS7D1d0A0xpHylgZ8jGkxuIk9G8PcOuiJ/mzONmq/8tf/Hx0
IgPkLf6lGP8cGAJxL6Nkm/Lvc0+8jqPT6T4JbPDTi9eKX6aV6wB4OcRleRXbjjHNz6A/01HdUTv/
W1XHDuDrL8/qsTcBz/adLFGPV+IrTlFDL5CejzEOxepA9i/FOjFK+RoKh8ed1LL1fgSGghZFM+NE
eLZgjKt0guzwW2bn72GWRgOR8aQmxEiKWW8I+aBKDTYWzZMYiYWsh/NTfjumyp79WUsPuEovdzu8
/pgcMEHVrjGPrV0lkL7I0ddM/1PGTOsv6GXmucSAjScHOiT29LoCkqUSxP94DEpgB1jIum04Cj3f
aaxze/yfTe0beIZ5k4mL/y6qS+c+L/sbun/pmuI3LnjI0zVj6RQEwcgLrOg010ps0HerKRS1ZSwq
xOV6j2XYAWlQuqCyk3flM+aRSMN36q9tEublCdy0zqhnCkcN0RzVc4zZWlF6MCj9IcFkIHhoqSdT
UrWvj75pGu+n8yWIiImdDcGa8xOitipxxCErs9X4Gn9B6holqXlasz8k3N3BtlZZV6Wc3S4zz/2V
cF4bVkVoDFWJPk6RtBenRx5ZTOPcGla5/eiJwEExDcJKx4iL2iwnRsV6fKojDD0nqwAUYWI/+/Si
8f2ueSXRWxpeWArkjZiTmr+9JGy92uIpd9Wd3gR1XiUFHpAg7PCIAhVptRyVYE3ZG5O/lMQy8Ci6
idHpFjf06511ryIC+hl3dVUf+pV5cPlb1qFlPkbq0ct40MKDkmy4laB+gas9RhFY3KT6nqBLNvKG
jKvv1cDS7chqNY4PEeZwX7tiwP8nKfkD7yn+UNUJqSy1EBNS15aLFQddNRhDJrVoQASoZCSTRvAS
2OL2QkDn1Hytc7lDov/7Sh7G2S45MknynhpmevA5ZH6a7SQO780tbM3CZ58T8Yy0CHTZKvc7fusu
VysYvLWrZcQeDdQFpVk4Fvh88SnUB+vDlZ5kvmlRwf/3meXodu9yIYDbTEp044txQJUeKvgWqFgm
aTJB8wKT+v5c3m7nltxikomqgYVuCEU3EOSl2gLkuHM6LIghEyBEYri307Zeq83oSG0c7g6Vaek3
W5RVwhUzYYXerJZ/i/wrOgUGXwH+t/bSX3fWvPGG4+N/+Aw0F5lmLKkLhtxuMHlPeDDJlzYPnpkh
fbV7ZS7kYdWAbEdik7kLg1x2ZxTmpyEKjZdS82Ytwjs69yHiUt9zs2aeSv7x4xBgABqBut6C45CR
rxnHD8ks4X5xMuN8ALUVkpFZhxVIpZMJZZgkOh0qX+rR4YKj4ZoAxDmkvPjZYc+7gQxRT3KnZFGQ
fgCp9tmgLBG57WO4EDjj2XyVRVFk5wXCpSl72pLf2FI+httkP3yK4vCsTtU1djGTp4GtMlfdXXy4
8NGI+v9kByCg1NFuEhPSsMXkj67lQ/v64L57JGyY+4HXGLI1bFuYQe46JOvOKDtU66vcrLiZudc9
kI6MptyZ8YqsXkV1TcbsoZeXdvLDWHJDO8cgRHqS2x0UevynEe3ZqoM5fAquSdgYYVchF24q5KGR
WEUsbX1EpTE8REo+xajJgXzs/7/UawxXbTAEiD8QCeLeP3SDgVGWqH5GR3zooLhSUdK2gMHaWH9i
UUMX0OWBH6Hwccr2xIa52gcWdqzkKy+RlxuOqEh7TgZSJbQXQtxek5b5r8QxMajKaKEWs6u4z0oV
7MgLT1SNpDHNQpuhiM4yxsgKYIQ69C9WHxzCMjUK8kW11OQkycZsQeFumms8kTW+ZGBAeMJOKC7s
pExoFdg+gd0uaKugwtPUhZEKVuxwGlUgHgQwT9oQ5jFQgByARBXdspDhpdCXa1NndLo1VhaYs/In
cfyJ8efZgAo9P1yVE9cjqdBwI7Hwf8lVyVWCqrmrYS/C7ldqCdnHQ9IxSnL4npV/yBWsg0P71Jrq
NE62BcYPmjpr1qgosB56VXgXG8YMuVm4hOjApEpdwsM8JZjTUI/+c6lOqmC9c4ulOlL2dOCgM9FY
GVu2n3HFamt6zBQ+dxwY8xCbS6UXzHSlifq5rD2z2RkSQZPxqIjfh1hgHu6YF7igZ44dFeNsv4UN
sGHerkeNpSSV41+MOe77Rf1gtCG5/643EkBtC3IJ+YSfAgu2OKK92QOtwrEFRQalsfdhK0sNs9eq
n5fFQRAZg3nkw08mTdDiXuyrIgHjI7wSFhuDv1O13A3YwTmPbunFFzpCKLONGBYPyAvqG2kvo1Qa
Wds2KK95tz13m4YqYomn1isWNtuCcCSNp8+XKzgSkUjbvGwyLYcRMYUSm04Ipm81wVlcKcGjv9RI
/u6w0lb4YG0TdWCLDLGzNMO1nljK8KlQrTGLw9VeQtVUo7QdCpQAbgjIE+7dR5ZF+CAafqxa2VR1
KBL4FsN9VQYZ/QJ5C+x2BFjn1YY3kqnWUeWevdoZQBYPhnAnXp55UftJcNDrDtqxD5XhOz7tTo2x
bLr65jdkoUhmRustK29cExuhu/6hLNGFIdvUiPHz28yTQ737buXEVB8cFJrREmnnq7P/gERwuc/N
WcR+2s81XPK15IwAozWhdy5KnEo05IHTQ6aD7Lq8C/gXTJD40ziFu/+UFr6x2qFgT6e7dmHVuY6X
EOlQJUnG3+C+3kekFOPeGBZwQhvKQq9A+gcBsvGubEvRYlqcN0wfSaUToAt/UK+3qbCTPk4mCB4v
wTPe30rAnIlMwMdEXrg/AViZ3649qDHrMNiVKexo6IGF1BIKm/sxcU/IZmJsvks0sPlvjXqxActF
vTdZnE1s/QDbfDhfNPKWLYPNUJE1k5zxb1V5Lw0WH8oyXDqxvpC9uP6T/3aQOuoPNyNOU0enNub2
LCpmi/qPt7ZDFrq2vcu4rA882PPo2vOpkfJe/Fu7ZHop7TMAjX+6CFhZckGpLPKKLJg3O1Pn89P0
nD0i5OGmmp3AZyvgZw4u/Rw/Hjc42AgyPUSOsyTsLtWDeCPxFORP7wu2HbHIr2cuBdiqlofDIrnU
F/Pjmg1XLsbubZEqR3QFgkvw2yzitPhVa57hyg4YT9Tcu6/fgOv4fv5KA7unTKBLBtsUZm2KlXPi
PWcV/RVpizvIVdVdxE6RvqDYIFPIhM8Xgdna8g/6M9pzEw2ZWHN+Zs2PT1emmViOp5lsdpm39+mR
gTA0pw9mmgA+KDvRuQHSyFbjsG5fWxBoFB26xqYh7ehQN+ltJZC3n5F0V09ZPxkmh7wTD7TqBaUb
s7K49ScFUAuhVveSPZr4+yO1RgS+F8cMRnfw5PiRrU8EVbqkEPTdjfzoV4Jsrns9bK9m48oBiIvh
PibcAj2QUmzHrfFJ9ypLzipI6QKLmUVOTuRLqcrNpblrTMCnsexVVtf/Mfv+Vcx/vz3hMzB1c9/h
zICSLKI3m+1D+M8OKBZMndrOx2x0zxLr8e2gcylk8lRVZNDjwaLEK/TaPiVN6gWBv9EA2eZfrIcQ
kRtvFpV4TxSf3ksoJAUNnlIaejnV4MRc5T/NsL2awr21MD6+8vdb8BG7Ucxi+qei+1jtrQVeiprW
kot/0yPuTcpOtcvLvdH7Vea8IHUZASsRg1RQuaC7u66Ng1W5HuGEnLTCPPuGNSi5Zlyj2IT4MrTE
kBTuqqhKmG3UCS+m9mmFl2V/cUR2KejsiqXegENg0h6e07gcLAZoRvArDxnaE4VSfkVTa3FNv6PP
s2LO750ZWQAsLtxmoU1OYYbTd4o2gXuflIBx4tyBKZfbuBHDqoRcFF5DbWS5vSp4EDReJ77qECLy
ZV7AvZEAYGr5O2MBESBxb5CiWHjNAe0mWzCDIfHNz6us/XIAUk12spAINqny+vh89GSEHFcmTTeh
MECEc+K2Mfb9j7Upk+zezZM0KnUQ9hn4SMfqLUSWYWlCBM06fSu6xSyPE14wLlvDFEWBqljiRuG0
o9BHmUd7efB1AJF2HrDIiRpyRBrWLH1gsZqPs7kZtm9O0v+EmbnIzL4f4oqgfGNxU/cCsWhji9KO
elTx5x01AiL9Od/9+i/IlBALwldGFOg8xVzvCG5cJl7nZc13kBcG3/U+Jc79NQxSPsEUN+TO12Vh
frxfReCe0x2M9xxbtBii85k4KSGx4uujI6z6sgp/tFHHu/jiPlqb7lr5QUpAKSKlHV+feDsXhX7R
749peCjt46ElGB9D3JsGCJLPkczdooCz6RrL1GliD18WKUO1mwwsjHbujAVjLZprExi5tX6OGpAZ
6A7TMSc+/rC3BHM94J/g9G2zdaAqBg8cXQm8Xi6FfzvsfCujfnd/r7Ni7I8wjwuqvnetFSMoIZpx
L4KM0o0uNdhQIjcj5KF/2Rvn4jFksRoACIU84KISaO+iVqIPcpIh8+y0/FdoAvNQp6ZcH7JlLllN
eFRvNZzciKfAus1xahYuWPBWMqUUaIZyjti7AUDricrUOxyO+1VnS5tJEwMSWSans4bqhhqFOTLu
rSiut+3aIkonhaNylhHUVVd4jhectP19qiHn10Tjg29/Mvwn6IVTXVxYM2iYL/UVrFp5IgqY5Aae
2EysYRv/rsnfAjAjPp6sXp9syOkleurZyzlpthN0r4XxXslKdpoKvq9XizulNbOFZ4bi6bl+PP0f
P2TT5+ebZI9Ah1vettKtk+07NfVq0vkqJ9+amBTl1Qfw8yEHEngvAGoc4RqZx52GsjgRw1g+2rXw
nJlE59Osbpq1yeahFOPXFnbryku4bImnWryEEbOwqYnApuAInnnYwtvJfY63vDaOP/U2iD8em0IA
coGiggK5LFJZLjC5bvJYkaKvh8+bBrKVh0WIVAdl32q/qycKzD3x0V1VsVUcUuthwl04NAhab2jR
/8fJGN0lAk28WdNZ56nA+o1w+9wSTX58IPZhR13w+xgD9EY+cUYE8qyDVEeoy8pKrqTMrYfXBdBd
gBaoV6lPy/7SfMdVFo4suGzeHOaairoC+jsKReCo2tcnwTf+ZyRtZGIrV06aEolJ+nibjW1xA+Jc
fp1tZCWCmvt9u1hruWsLGD0l8iCKOzyEW1dsOMxy6rG99B2wnX9tiH15+Oc0GNUJPsh0AdoG7K8p
auMHm4v0ARbGk0Ql/HCxsAuq32AWo8La3ZIzXW3VzGwN4wjR2a+UGyqAvul7fykA1xdgqZnG/vXB
HqtTllh5v6kQ6cG1/sWFsrOwA4zNohE+SUSIgiqT2co2U4E+prpYAT3NZ18VE5xbtJpGDntx695n
biUm2yXXTgAULTiVJ4PkO6MW+n/yidEx+0+AeOSQU9c5h/V8riXOphEmYz5duRvt4h9/jhMPSpQT
m5KloEUYPAevcO5bSMRGM+yVPUAOJFdkGP+e6T/uUZeg0ZVR7F9wYcbHICP+qbmTg1l9owZPbt2K
0DJ5D9sm80LSJK2cM3PUQsIe/5lhR4foP4S5IALFR7v42jIchrqhoztb2Osdj4InWW9lFLgs9u5R
DTEjVMiZfMzoythOkG1iUfrwnnLaCs/CAAObg8c8DLL8UiAP/ijwHv8kOG/0gxYiMfUA+dbcgmNJ
avcpwcOb72gq+EyYbTg2QG3fTB8oujIeOlHX3FiIt42GEgf7gWcdKS/ez+FxX9g2si/AbdiahrwL
+SfivKMNMZ3fICdUi2kxZ5gOVgp3yMmHDsIftaDP1iD9GMdKLxYN4a1RGUx+gslE+cx37Z4ZpnWu
QovoIZVo4wGQeXtMuL1VLrjzX11nVYIq4au58vt40kTsxml2YeNie+5M6INbWgqwDoArx7MxbERE
rT2urvYZtIi3J9QV7K1Uh8x9YK54nZ7nETVYB/ik+U8f9kWKsFrPVdSf4/SRsSJgRiExn7W1EKiM
J/fWiUGiRXv1r913PYnJdc85uVjKCYXbWlZWT3JA3FpsR6mqJolim6eC6TWqmqxPsmzJV1FH0VIF
EzjfJVS5fzV1G0FLOpmvZrqTUIXiCywiRLvgpjcrwjTuWrsh+qnI1761gAAkaLMbtnDdjcyg1N53
TL4ZGWijZumyV8SVQwvvBKMstitf+7IGHenIxuDEmtFGr8P6R9T/WAXM2jSS9CdTCWfGHKwm/jSX
+9uHQx3eUHX0EFw9mKT+yEK3Fl4SzhTc+l+skWbneCNtItrvvQoro5FtEb5WhVLfzQ/3qgIKkKLj
D537hg4EaeIFyzdM3Vc32XG6I3q1rrzWMJX73AUi1q0NRV7ggIRHPmq6YnmmgICEcT+iDCkg+WuW
hdPKFBHSeL2maL4KAXDpewlO8DwL0RO68nCMRhVDi3fX0ApGu6B3kOigQJb8Li7m29UvsOqu73uf
NDmu27Xtcp9DLPtLKPFZBbsdLB5TVuNbec11NpI75mwzZ9nVUaFythOL5lF7p6HBl1qCPkN/NjXL
3NlW4nEAV1AWClu+Jh7jOHkBiiN9x7k7qkY+ymQY8jaem/oaMEvxeIGLnvI+xMOUCxgkCYcWlmXr
DabetdHAWg1QknPlvtcPpHCpXI6XXe/BHqowom0bGcHJuPg/VBfoU5FAavRhcvzhWUuZhNw+Fsko
LiUat4uZ7JZ7FyEmjlqJN78XNxr8p7EkiHZXZuXMcik+iNvxRVjJT/IwtYNTEFCurnEvAgOAM5KX
tEedCUR7xtCgVVBqKFpGqYEzJ4UfP8dKPeBr3bLkTmljUOoa/J8uCji0fmB5dpcbKZMPLyH5D0fz
nu4NcAekL3l37NBdK19dNNyoRl5WnL2FachFbFJrUD8GPwfpueNSJSNCufXk77rEcftlYQ+rcyBK
wnDRldHV2J8uZzp8mOm9gL1LprbDVToZBHsRvqG7WnKOa13Ir4ohIgLgoQxjGssQ1Kx0EYeS0hpk
DUzWsjSySK4pts8Z/40wuJT61WLqqWQHtk1a20143loFWkAIvI5KZIgjtCnL0kGRf3l+P7qY2z4B
LeRU3jvOgCJ5bblOK9gbTWdW8qGPF3zb1n1t9GGc1lqPCC6i48BFD6TWQqAbgCzBfnFr3xuhrPu4
I6+alcO36Q3J/Ah4lsCzjBP4g+F0YNKqSuGIEAh0HMSTt1A2gYPGMWy5B6oGFwF2qfbu7bOtwIg1
Ig4BthVoV5aEp7DCOuyWG2B3qVkk1vpIC1Ov5ydnVbGcDVtQmYEAfAf37JpRBa9sFINe2CjbYgp8
SpsEXZLlaEE578J8i+V6Szb0D513uYEe7x+tZ5BzxsSGR9zt1PIQVmhiANfG+Q6umKSqb3rDWFUN
TaRtdL/PFntEUgeZudVvesSaOhm1RpgTLIfUin9qDugXoKrY3Fs3VuYYMNnbx/iU5ju5WteuA1Ne
wVGFNLxvR4+QypqsfRiU2L1Q3086VG7cct+PYWeUR32pUVILKDd2uM3wKjTsHZClrvB8RYd4FZG+
AJTZlfyfPxJtPPvkymMUItkvmsQc/lK7KGAfwWHDkHZQiRJiIFtTwxZLsU3iNfb3GFa7atTTENOL
McoC8Wy6Nvy7gV29lvswmJ8sc5vmvG+ONH72pb2eTx45mdiwt3svtKvMJgyBqj8fFjiqsAn0T6qU
sSKypd9ZdkTaBlpV6cDZ0lS13qcBNZQ7G/BjFegzRJsnXKSDxLvFPuZDOWDK+lHm722N0NugnDp8
ajRF6EyD7r8SOEwNw5EcPhe/gkIuiJq6maHz/a6NH9v2b8aIBHRRetlDSshKBEMnOL8evA1L7Vdj
o4n1ExHhbUza5dtQ7NL4lI02sX/r0H0tD7m7o9CDLIhBBaprccg2dPVuV7Im7VDlaqLMHeeoe4nE
cAXTwaNjXewRuP4Gpsznb60lFz/Q6VjE++WYeBZ3hMKNCOmBhHQzs6dD+x3/sf74ujMiWN1NQh9u
LZNo3KJRMOC8oTqk/1BRrgiCuhfNiFil/BNFKhsCymK9oR9ryOCAhr2z3wcrdULJTjkrP4cmUa8b
ZAYVnW0NcgshTbQYQUNHdm8SNlp/bPTOHcFRDyCbQgX8Ovy+CNiBGtv49jXn+Ynduq5gkXGnkyA9
iKroWvsHSIlknvds3okJenUTHg9rm1HLNEh/x6baX3rikqaxHZ/Dnyv35JcIe4CTRGgoVweeM7Yg
hqZiX43QPkp2phDJ3re0TNHEAbjxvr/RjyvXL4nE8HlSdTI0yDZV0+H4ul51MYd7eZ6ZhtaE/MLZ
eRTYrYo5U4xp+Ogjf1xw5oR3/Nf/cp9NpCoi+NjFlarPGV6+3dW5MtOZwegVaQ1qyM/hJmY86ZNf
RJAOySQwRTKz/btbe478WcVABfMEv5p44ZK9k22/nEkAILyiYvYyhLKUgZVDZcYl2Xn18tInJD0T
r3veJ1A3CHcrqZWXvnMrm8EKN2bhktKjdy4rmE9tlYEYGRul8dnCCotcUzJLleWKwYGdfTBwtsC5
vNV7wLt2G5FtAnnnfOqZcCKPmO0vP93vxjTsAReOYTrHmYf4e7HaSXe+1cdrsFbUGJWR07LKj7hx
tnITwbq6nPOpHePA3Okg3fjlq/HKBH3dECkxzqz+15TaLaY1Qm9ws7NP/LS+x8aujrC3oWqIas/3
nwU/sTxgal2YgX84n6++dPsxyPdSHZQ105UnDcRbUmrH7LLKWJAzht6u1jCOm9kvURg/whkCDaiJ
y4UMGMM71vhO+grUvOLxj+p1ESl7T50Cu9wx2dLAV05TSgGKzrkwi6KfExMj7Kr6ledrcDf6aU73
UFdYC5yE8gEBv562ZtmFMlDu13USGh+fI8dwAJ28A7fvw5BolwQwhknO6mvxat0PLrBj6GdljQkg
RNoM5vfWeccnF9/fUTS/BeMunRsV8ChrI0of8YEOS96sN1jdrewMDiNR7qeULBreaAgSfvKq5+ME
h+kXBWYeF74U0SujexbNDYCjpBFyIR9v5TgIh19+cy8SdeJdAYzTfYPVbxiceIO7aQPcqD1IPMgu
v2Z/Y/z/oMFe4fMKeKtXW3ddJkJ8MzZk2HcHeLxVQilK2mZqLprAdBipfc1pACcZczWVLIIDyVdd
sonScgnT0rtAvH19sFWeuRwLrZcpA938mqU8GL63sb2BI5P3k5DRTzGNiztIxh46TM6l0fjX1Hs5
98uD5xzXK76M/8T18PEr5qVZyj6PBiqOKtFRq02bibx1gY5FUj7sTVnGs3vUxZHnwgLTjZ1hySAz
EupXA6TPr/JOX5+/kU0Fda4D9TL3dgJzNOF+FKP53Cb3JfWiHCtc1M7cP1NWOp5sDkpDgnwRLI0U
zC6UQIhar57JRKyVer9mCzrzGBWyxKUCvfFcct2YhWvvoEq03WBYd6bcO8/IGd4IhZZBXQc1Jf6r
fLJ6ohowr81qTaQKGmu0vmbc8iLVSm32cNlkygjHzzO9Imisqrg+YUN51oQ9X9b4dQa46kljAixz
CvzxUyR8zzMfiPud3pwbid2QxrGo5UJPtjFUOXB3DZeOTGSZnN3PuhrDmgCfEON6+wA/Lqfa7BCb
iTNUyaTZn1I3mCx+BN0GzTVkA4cA5qQbGdxNwdN8hSi5ZhLLOlCStwGxt/jUqYrKocLeLAU9gKPt
SnOQzBByiEldvk7eWjOnwUe0xYkMKbG/AZGqM9DjVWkP6uqUDQojNA55FrBsTVAYf1BpXq4Niz5U
ePfgsi7Ao/eN4GRzeJysJ61jy6GajJlBHjJnaw1orj2escnUcZrOPjCkTdRoX7VC1us68e2cmOT8
wGWawM2bMSbwb7zxZTYZz4TRdKGfzDAv4OvbDBQ0APNt9bf30IJ4MPI5TtRh4Fm2uOm9xW8RaYf2
6JIGkDA7igUTIsbhp57sK6PtwCyAliEiqJTTdgot9RjLYugqU3kRovaXMDNtAWK9b1EXp5Mq+2ys
s5ZZLOclPDzsMFyEQ5Kgu9C5xfjxH4m74LUh4VUeU6e9L65m/yvZSTMPSKKn/64zayc7WEOwULrV
+bE8KiqHBXWHvA6Oh1C5VxB12rp+mRCFPiWyjGiv0JwGYaOIufznBclZHhVIbBZP/X8RkfZPMqmk
Y613rOgVLudcWjvZ8JEnlmgNaiWuAwrMwSijetqgsDktliSxI+RseysJjV1y7I7HT363DgB48mIH
Q+26jUJubVqWJVisc4gis+9jzhjX1RLlJsJNMDnj9s2TX8RRqqi0y5dVp8liWvk93+/7RT6fQVbM
i5ZpfFvA6LJwzwqPWSmOhd0qXQwLuwsksmeyXDL1ZQ2SHmWTry4ng38LC6eRSKFpICOOXBZ766Qz
SefJMsIp93OuBmKn8mFpHB0qY0I8aSJE6jz3nterEQvG1T+/QCVJ0Hc84peGYeFXQureUgTBkXT0
u/iuLEvqHn2B2s1mOWBAly4SWKFjb+HrbtklqQc4/ObLpycfaeTB3Y/43hGFZz1mlneagVLHBx2j
RF0ngbHoTJb+u6vFPMbWegfwcR5eRYopO2yMreswfkXJGIxwCCoUJQJIzqgOVKcE9U7olLXnIpTj
27Pet332i/O7uy7OGcvScRvQaiZQpVCVkeyOi5Ki5PfzvSDLxZxWva2ahZzo4CpoboxZXqv3CZmd
HPsF1CWPjtbxG5dMr+DM9Kb6ljibmp9S/7bvdRYxNv0Ma8VTsyM1yHr5/yfGBMjMx4F+ql4yFaWC
EgXAI9HLGnyHx/8wgY7k/nVgeQGFqPrw78lti/UTxp1DYLbgfm1Xvlbk631N7fCgJiG08qayBvrc
9nE6kpPmFJGBg6YFRMkwjidxpowbeyxOsaGhTE3p3W2TF6zNY1xPCLqv+CHdbYRwLn1yxZS0OozF
einDUS6PszpsmQZPl6ll3v9wgMEWCYrwzAq+oH99N9SpwiC9y/NsvgvzZWlrTrERiah9VnRvpQ8l
RlmRcgEgRqJwMbp3GhrGb2GXOCbWYhVdLryqTCdHkNE6ltoWJEXe5W4c1pXiFoPToKckTyi5BUtD
oR7Hc7I75s92Gc38bsOyvbDTIka7lIApe7Dh/x/Peqc0z5CPdDkvvJQ20S8iBp7UPlBkt4aJoIpe
LJA3h9VajrLbFoWToWD0zSL+k2i1uU6/pJAcLoj9j5kutiiqxPoRsUITU/5eYfbtp05RZ4mafwUL
fN/ChcCTocz758MNzXLnTcLONRWe2yUgmFLI9GRR9jnbKtA3F0866J0wWP/LDrnbvD/jrElXBKuU
f7hwP5H7fvdG5dhfOAH9vWxnH7imYbFfZpXQWkp7T2rvu+KKf3b9aZPACbWkTKNapdkSvnudHXQL
msSNxcRTQQgceyDXG/R3cqNy0bcqf9RjzfbOS4Y5TmKTYQCSi9V7Shghlkzin8znlbuuWpcrqfDM
+b3+2S0Jlz1ygqHbAEt9zqP5Cl1TVu/ic1KBl8UAJhXaL1mEhIgJzVXUptLdFtcqL9lvbU1S5wQO
WMNsNVITQpVblka/wiiet2bvk709MQ2bKjq9/lr+MFGfOolUSDjeU7IVdG6X1193/D5udgK3xVCd
oG+xgJgX/lSNpqyJ5O912FRwZAgNDkWIldwoO2QwjQ7/KqBEfSfrcoSBXKABeGj4mwYOhKK6ztQU
nSNUY7QMLqVIOOOkfxLoy73E3j9ArsUdowk4uKsDS/9FY2sudKq0J3WwfDOggIf2JNXz6LoecI8y
dO21oeHmokKq+x4/qStq7wxDEgGcdK2BqgfX4WxuPm59P4D/lUOh7rkdNu5BCcAGXoiJvehwOm4k
aGucsVQXdxosQbdS/K+4NTEIw8Il1lIk0ZaxOqgRn5H3emG18Hu0kP0NsWD7O2iLR2jO58wSsNPu
tqaqyoReDp5Zihtcy/Ol9dlq/Wxp1tw0x/BIdsAOBfA0fcZ/r2CIFQ+UHKk2d69nBmK2f72xUR1/
YGSVBLvEUBd58L25zYvymO4G0lIY38kqsVS1le9M7SuKH2hpHn7gm/0cCE9dqmm/ODwqiR0uNEDO
KKpoEs2qdDh004LwezNPT5txx7TJdCkJY2mLMEVGWMGPaP7jQeS24Nk7OPZY0ZlK0Arhwt6+NRRS
0V1Ztln01LgZ+tyu8Urx48BEOsg6Po3We/qTRfIUYoNnSUN/BMM0AFSAMukkvUqEkq7wXXJAdJ27
8o/iapL6rRpV2rMWCh5wSrntPG8Uxony4tm7INj6HFASB5LmUAHe4/WJOzbxyMlZJv/hV7XMC/Ut
b2EoUA+CAz6b7iJp9wAGERM7/4Oqw3ZlHhJp1QjJynsrsHZAb0eh3ci8hTbOPsflPg2csxQWYzJY
HeflzmxvsMjQmq6VK/UHg4vMDQivp74fZqWhbPmSm+cDob2isN/zX4Y+MNs43QrMjW1Vdc/GHiWG
JXMZ/dj1JKKPE0iD+qpq9VoLrjJExbSeEWyJ5wp+o7sIuoSSrFt/QAvgCHwUxqv9FFHBEDytDZ17
hpShjTd5XjLTjLy4UzPyPzw5b2ftFEEnD4Ag73vw7EHlNnONpHSPXwCrH7oqxQn05vOW2zTuQ4Jg
6o8FV5lgYnborrfbUnbQxOi2CMzID7yDOqcfgg90rnK9H7WUn4VsyIiXQHV+oMfyyeYBttEZesY0
ELhifZytm1I2TjRrp4KFik0jTMKyxM0+NSyW9TuU9bsk27UIy5Eyx4X78H7wngTuU4gtOr0U23ei
aXq7dZ/LeeGJMQBJpMIxdbClGaOvW+42Tnb5tFPugnDYTiGhEzANS3Uta/DqaEY9ueLlZ9wW2jnd
vmtmaHrVzVaQqV2pDc1n5b+pZyvb2JwoH0qtJF01qDvLtqn0hdIEtvNaUAVqktWZ2olG7GrZMgNv
l75n6fz6ZBx3Thn3WPPV/v/fKZlzC+DDAWtseL1YeYu7me8ZPyGY3oC9DoPdC1S2zS+ExdaRXC4l
Odo9dQHvyRdMhFDaFa99AHDRXlPOamAT6NLNFfIPXiBIuQS0SgKfKsIzNWRJYAZLFc11i6ybYWYh
KKF/uxpg/qTCKDmpymcTKPOKijZQxjLV3pia+3xDwnZnVMoHeWf1g2RlGZOVsNkEc0ZmTddV8iAc
D64mZtldTLq3tDgSkWDZw8m2Olz1DIfhG2n98sQ7mhw1uPKqCYuf/m5tRSNe2otLx3lwIXo2n9dk
tJi9hJDzYk2jdLd0c0BXXaozUJhroZprk2nxbHeTJbbKwS083EEnaQI0Uu2hLUjZ5sKQYZlyz/FT
1pTf+md6asuzAiSVwYfZD0Cm1J7KIP1MtOIbItH3LpYcjTWia7S6Mspk8ajEhvbo9ldNnhRNMiuv
6NDahcBni0hMvhF9NGp+dDcJ/Admv1hID0TrHPAyCVwG/uG3ZwHHhRelTI12ijNCrAj/5s4n39f0
jEjxhQlmPLBiAnHeHtICzUx2R/B2wt+hlOKquZuD1VqxhqdRWfE+2rASU3DbZTvEA0LOTCJlp4cm
a0ICLzPYYTffVwotK2nS9kCsav3cnEQfIH5rR6YfyZTFgC6Ri+JsL8b6QexKENUuAnDg7l58N1br
kbIOFvW4igln6UTAFszWzr2C5LJRnurS7ntAqNnbLVhKTxfs+c61CH3zymk/9df0l7yfItwiQ36v
ejt6dM39b6xHlDvEpSc/qBYst/xw6SCEIEkhCgasTg40chTyDBcZ9ib1Ao7p1MAr/o9VH1BEmFMU
jOy6FXjM5V0/s7dbnMwLEF4a5q6U2G39moHTd6vgaQDNohREdbspUxEk+VeZlSCZ+Z1za+DQdtll
lk7zR2zbMk4xx4L8kszrBKkt1cx0DqbYoW7TtXOA6x5MM/RAkRNIeq3a5aBi3drvBUZYVW7PeJIH
qeAGNgobM6XqYsNxc2IXhGymolvJfYYUBFuNlVCqJHVHh9JSHSVOU35PGBmoLVsJKxJ8D0tYpfpz
2gxNvLwxhDeyaFKQS8xQ91tuZmMZEvlAdjAV9g5j39G5pHiw1uxtwYxOfzFdHzTAaUyxCuAsMBwP
8s1q3ERV3QoMVe4f/leQSJboJ0cu9jkZKLIeWXMqowSWfyxXSekselrhw2WozKmHDTuT1tN8tTQ9
tkgHta0EgVr0ce8thvvwclAKzxRgQ8pF+l59IAxAZgtZFwvs2W9abiaLc6g7cg4yVt9wI297zdy9
yJmN2uJtdFGKjW/NS1ixCMgLXA5qZVCAqTi16IbPbnSL4hj75+TetFws4UinIkWl96ZB5X/+2I33
IBZ5iSXQRI3FJehlVTciXENfnjZk+N2hk6JALfxamSXtzrVmED03WQTnkLJSzZTw8T/TxiTAUyX/
hGQV2KzIBAWRGvs0olrSwfiK1I0tZneBj3aoXWTWg2rZjbqvstYssj+/kQaU1NosFWwquQhbmu44
XCHjSlgWK+0TaQWocKnlI6v5lLUBUAh3M8+e8NHpLyy2A+IstVDS+Z4VODb1sgWCvz/Ta+HVPRNR
2zf6kaJg8l6AyRfaJkcoxtunTYSTJULLgwNCR2V/MU52LBzTGT7HuNSUY2petDNmsKU7b26q/FWY
hMt7c8TTYRg+kd2zBQtjCAeUl8wPEcUtPzpkv38K4fwbZND/ZWqmYKgzBnNYaMWslg6F7eL48PuC
hnrRP4qzOY3WL3tclCQTl3Tu69KwwUDOkTaHpC3njJAKvrvSk+TLQ09vgTmEHcIjVMWLQ47trDIl
uY/5PpPLCxEo8fohUT2hGN4p3wL7/ZuQiBHYhWs+PP/AwlbN4TAFl4qwskmjh/p7Jx4wQVtTklqB
HARImhIFHSxtwKxc2od1kdEiEdNFoVpmmk5mdS+EkTm/F9LITLWTqgqaPMzZqc6NmDtInOsr5WmM
+5cfGIFSkXq6mkk690/3FQox6ME7Vax1clPodzN7HKV1ivkV6sx4oSBtql8Q0lMtr3bLRLxu0qAq
wWDs+dxHZt+/E6UXUv0KQUmnqsdYwlqoi8XIK/5ri55QWDHRxpPOel02NsygbreCXkzI8Xr8pSs0
ZW/WlLK1gDEQoFlFj3BncPWVShR0EK/h1ylDUHgqharN6qLIaSLae4Yb9wEGyGiWoFgZt5x86I8s
hf5UmzyhrK3FcJm7udBmrM9GatkzXWgYxJbyglaz0Z2d6CGaiw/YnbINtKgDG99Ys9BtDuf945xu
885Lciw2qYSSCD3uFqbPM9iGfbOpwZDK28FAV+8Otuadkk8zdPkmEYT9gcNgwd0iW4moYlUFFgfE
aWfkjl3yqEDawBtfrWrR8CkmE22nMj/7lrJ6FG1sM3r2Pend2J0fxbKLaTMeTZNQ9VTBd70Hfche
3LSRRFrMRybfl3pr7berH5I5W1JeXSmU3VIxZ2a3HoQkJJb3h7gBYCKvPjJJTEoRzNMZ+39q4Ihf
Rv/HSqeaNuCb1vxB17fYOJs0N2Nt6o5a/CQgjkJA5jUtXlFU/Y/emqc3rA6xubzIB5U79fdz37bP
PgYldZj06I9wDjnek2F06astvIssX/jzz3EjEB7Qk4CNnqHIqJ0TAGYGL74XRgkLyyXWyPD3Jmxo
7b27ZT3X0CXPejsgkHOr67bFFkxLAqwCWYJ6xXrwjBn+XplTenoI43KxR4wRCNabOnj25hL1M4fj
Wku6SLSgviTjMqz3qCnzIj1l9ryMxybz7opzTO8rT0iqt42CTYwseqohWc56EQTWISGwu2pggQma
88AEumY4WIvPZWlr3X1Mf2Nat/acU678u+Op2syn37hDTFVxBbDpCli6jWR3yIY+bl8uPslmEBnU
CplcHiWYg2+IAicry43Qs4yToxc9YSY21IGOHTI+rhdJ+MiBtOBnddATgiiLH28KVtAfMcSZb6BH
243NUZd+/9opIT5aSTAVCW5U7DM6f9d2jTDfMuWHW4UVCc4Z4Hbt3YAje3et04Qozk9wUcloR6p/
t/N76uhvQS28hG7mdIzM+a9B3ELkHoyKBG2RoN1U6nT3ks7yBXs6b601cfeK+UI9h0QUK+RfU2fK
+NmjqMFdf62QFsKOsaPG8XhEGb3UPITWXchO5ZW8503n4aUgyeexIsSiU2rGy8ZUHOFdIGtMa8TL
Hgi4mW3NEZIoK1mrug1pGH4U8nk4vfUfcVE2dgjiR+yYWTY9dg8YgcqAERdP6briKzBGSABE+EcR
qj377WxnO3bnI7xAftLQqSLu2Aenw0VrfkH6GuTlX/3GYihhO4JaT/Tg5BCBys42t6m67i6q2Hgr
QD+bBf+yP12h60AR1uuMc9PWLs1mDfyu+/HBy3PAO7rceAdDmE9tj1xdDZHOJxIuvSMwzyLhv17p
6CNa6OHXC1Xht0e/24xidhfDW5iw1DGQdht3MHjCgXB9sf6+wezHcyK1riC9vyQBqfK+5awlMYQw
b+3fL7ejjjM6ptXey+jBp2Vq+O2t9ic+lMsxgyN5DdFVp9JKOn7PW9Q7DX8KrKXsdBSp8NdEh+JJ
tX1lUI4TbuWO3fzUWrjh7e6H7+nRlZucgrpto/MVQmzWdKjwi/KvTzXKo9vWoqCrhA4meh4t+pHg
so8+DPv+HhlO8csHmxllegkqRmkfA1sv50A6eoLraoIPMQxga8SA3Y7MT2PPxcvZ064fX75dqZ0Y
UK6RazdjgDQuyZTLt6CbXLKMHkk3i+Ad5+CGsnhy7Su2spXIDF4UY1MWtmJv8yB/XXMZxTtb73Ta
ZOexmjw5i4M195jIHAa1N0PUIBWr9AC52ZxOsl0ttRoRU8P6JmSHzb2Xq1y/eIuv2RxdZo8HqyeO
QL2FZuHsH1kYatA60RywaTM5xH9m6jlOTg6wNJYaQJgKrQVHUk3Qsp5KGyfh9XjzYN3AcUsu217V
EpyD6VJjAHg+bnqBkMc9ndqIUDEcE9SzYY+Y6pPMVVYjcFWvXc/FZLyIjnpqrKTptt0VhCuC/qqw
x9uxmydUV+RK7fQGNDb6FXwDto+Rpq2EW+9CeHJ89xgppl3KWOucUsUpamiF0WdQTsQSFF1SsmRP
9IUwUmzpZnKRbRR18gFSTfqc2zNfMnXpof2w0WPjdm7fnCo1ZuvWQTFwy0NgOFEHcblsfo6m8Bdg
Ss5mc8ct18lpse7d4lHZ7kYDn+hIp4cSMkqVLS/VjfTPAqq60bqr3feGYZq67BTThxbuCeTICGeh
CwR/08peVheIctJVlKTf48QLvTkcTJpIwNmfxH1OWVqWIBIiuKVAHlqDvr9zort7RgaCi2YGDsbU
3yJWB0dojN9OkC7HswJl4jureQly6BkYDwB8yhiR+5yVweCjeD3dW95G82GNpDwuClyCv5jsbOl1
FZiemAVM2EboSFSWg7KdtTYlYy8RIbZrl6PioAqNLq3Z42BKcQiRyBTNVPjJqFbEkZ2Bwb2ZnPjj
dqRGCz5Co8mLgidslWF96BSu9bxRjV5fcskc2tO/EnUDs/eFmdfm64lJ6nm4IBDkUtWPomVve6Q1
C8t3GD5div/8xyiygcEtboKXozJkdf2rieuydKMkL03cYXgKqkqG+3J4xq3B1Dd7lDwrhXjSG1aL
qsrarLIn3Ws3iTXQeLv9TWq4eKXagSLAKdGKAEYsPQRU2qleiIvddec5oDxiKNAradctpEp5G9om
filp7a8MYAc6dP0ZX0jVZgz4ln5iGmM2PF2OHuZFsgBLnhv8NDrFUgRHEQrzJJt95POREs4JWmfF
DcqZz6s2OBIj3q3bTae8VUGr+Kw6nuWnLuuGzn8PnBmBfIDz/8ISB9c5U7gDo5TKlIv4QATHA0+3
b01U5y5O5N2WcClQIeYwZlvbCfwXZKTakB27pJS1+qMaL4Lk7h/wu5b8tBet4AbXtcouFNR+QFue
2TT9bsYHZmQ8QCrTjztjgrWyN2UsC1PwOEt2F0eTsSbn7kZ0eluf60IVCvxWg6qpYE12UYZmCo3z
BCxUczssZSOaC5VlPZ5CbCFrZ5zOKWh6xlPFICvBRGLSnlZZMFdj4uK0tioXCEao0Xm1u9j9jVLs
RK/KmNR2eSySbxWhQKWv8Oo/TPvdcm0E+Gc4ZM7BVN58f6okxcpxqSaWPusXEgFdLZ8G2ILgSKz9
KfCl5x2V3n9QpNwC+kV4sqnTJg8I9LMUL4aI2GkSC29GYQHF52GbkXqHdN/H4CpaVsgFN47jzJqA
BnV7vI16JC3YZhzHevO8aVm17/GBjUKJXml4c3aeIe9+pPkjbP+/b/uDqUgZQN0m0qEvzQPHBH+F
irC1LCpHDGGfJn7FxsfE2yNmMD7voWXvsc5WC8jDCdJHEj9atH1MRXH2QQWvRSq3qE/2oBw8+19I
dvDpz07MKylR99oNHHhqX48rwQWzlykSIjdPINJ2oOx+QMQ/gDWyK7u/VCY9s0dCBaTPi6GSETan
vqdGqsLc53bdK5bjVMG8dRtBf9harK/xOAds+zODgyx1DXzNDLCRdd+tQ1m6UpIqd3LY+AB8dTAh
QuH49lSO+BXgLyJVx6Lxrgv/oFE9nDiwY/1F32jmwqYM+kPbvZXX4D6cb+TqaA1++1d0WY4MzTDJ
F7sqxcAHK6+bFWUeZa9x/Q4BhrlsCU9AGW+uv4Mys3YKwb79Y+vj4GzjTWBPpkx16VQhUXOF4K6M
cqjEWCrVqYYT6CbFT3z8Jvf8Of4eFjjTIXQe7wBPlautwxp8XuyNagJZNfm1JVMxOpuCVPcQbRqe
zYUyHzEjEsujKZAjn9EgPqzvRFGRd8sUzw8oZIDQCJOuRpS3gOKI+q3VVjU2D8k8jrB+APP/yoQT
mevzDWDbQo5FeNjyrex2xa2KtKdziHRJb3IJfIPirgQzxdEMxM+aUXnvM7mt3h2k0OnUClm+6GvI
Ggav6nhL7r70VVTglAAh7cgjnvP3RVFuQkJ53ptKrfZrXhebMTal3UlvxEGS3WGbg7840HqvtNMz
4d9/fRB0qIjgztj5YaMUnNjJRU3MGdRn1jD8O7Aeh10P5z0l7YRCgXg9veKnCuCJoY2xM6y4DHf/
ZHMpeiQ9O7pBOiJCiFukUPINJZmqbKiAi9OVL6Uwp+kzTu/BSNaGpuTx+8CF6d52QLqDQxd7V1iL
EfO1MfZ0L1ba+kgYhSV26UOAW2745QsU3Vit2DVJ6cCMgVk0au47YclguCq7I08kCuyWD5Z64zI3
babuWTIOlr3ynDKMGNbac57Uztw/bO3bGx2TtYSumi30Pw2KPlBlgxiSht+cEYmaTGKYReYOi81E
gF0wnykiJ6WSdApEj4hdVrAO8dSgpAi89adoupey0QHibZBclI7+dWFbz0kmkWVXl2DVwomTrnMM
vSs1POG6mX8LC1AWN4dUrQxp2Kf4jm7jEtOInG597Uqs9NioGbgnLrJjKdE1pvoKBsOTfXUczhfj
D+fO+1nYOlj6ujSJQZ4rbNt5eIUw2i4oPFjyXU2ukdqjzr3eHx8EMdHrkC44NZID2a9/GTB9p16u
elBJ8ySkJkCw6ALIJlsZ92vuzGpWBgKQxhoGuxr1/9dWSwPV9oeeMUrnD2jxQ9p5cg3CLlDXdLaw
ZrhSdKOjwltQEX2YWW4oHhqReBzmpXh8Gc6vWbPFLRA3otnPOkuSSfaZU2wUiECUA7tIzwHFH8iZ
rFlrFjoxG/7TDtanuIqbnibDySktSGvMGleMWYczucHcyxBAqUXKTtjf0vjhtMuLVcXZppQjZpyt
x1beQgos7wDMFa204bnFKDwNTO4DabH+NC7PowyOwUtDaYGOAmTUFr4LmMCbg9pco5IQkIVjT5ih
BCh7+GZB88PBAFjfwI17psYY+qP2viCy5VV+IVe1/R6ZmjV5wkau2gaD3G1RN1vsv8NuhEZBJ1wR
MQmS9Osz0Lua6vrIm/KenSio+AtzHpYMvmfA3VhPjGRes3rbgMYoZ+NUGCbyScDdVM9CEcIdRP7i
7MXj0cTCRtSJhg6qk1iW2a4ng5+YFV/3zgahz/cyTtdcWLysoQV04U/ei4e8qGJIIRn+KmIYv/Xy
TxqOYNkxrzXfmlOg59Gnmquhc+SKIVWEwVDfZnZUJ+4OzCKflomsfYHX+ejgghifHuTQdWG8v6KN
HIBVyfVjV947Sgkjq7P+mxVJk0MQAZUT9Heq2Zy6PqwAvAqLZKJnFo6zo2QdTzlD8QMvenihnSrE
OC3REdOq0tzPUT5TcZW9iX7pFcw0ea6X0PgMcxlSDCaSBbTVKsNQPt4UcG2DWR4zL1YlxZCaD5RO
nkVc3g5LlYhXPKS5Al8L1uOH0/x28XPZyYMsrcgMxT+OisZYoI3TCcqAqGgYX+xkZJ5Dv4P4t/Mc
Dq5a+wG5y5lYBrP7WX/29lBFNbbKArsiY0t8WWV1ZfS5Ez2YuC35gKOlmORRfxUV7Yf0eCqW1YMf
/iSlqERu+ko0FcIGoRQTRquKWoebbBPbcfj/oaOMoTdvLsstU/dBFCamcVctqH/hXD67M6flXQiR
ubRF8HcQ3G0TKJOvI0WRnqSD+TCFGhkW06vVxTfaGt1cszcPAfMG+9ghxgL+n20XPqEbnurjZZq+
Y9ki+GeAtCyVisf858LdbWhxs1ELdVFJU5hJw75c0nqftLlHGR9miyqAdphIgyzja342VoSVyRHw
MyXEIJpUMyYJ/WDt0o7jWwPw7Qa/Rz1icYA06JoF/JRYIrXWQb9Zl+iT2fW/ze3HeVFplo1+OlHM
KBtotgbmD7D1fQnqqCNgvFTsyLv5nqeS1UL9Hq6AUHGRFc5w7yDWvS7OOTd64E09HgUU21jK9lcU
t7+chpQ+7qS8Ebxfk2OvXtTlz3KKG/C2Szl1Ted/Jmr9vlYMz+iFIxW4vYfhr95dJyGBrvScOTSx
F8IrqgE/upOJG3zw7Ewx8KS6X6yhB0saYzN+SYsWwTZj0wt6lP2MAN+m7BBN9HQshgotP2l9SI4H
1Or0b6E8aMcL4EvFtfe+B4Y3VAz78Xnbne60nJ8QGiIkR1N6/inGV5KrFxbzmfeDRRnhKHNETwv8
JbGxMt8/ZjGiKfCgL+XY/KTsMMRn+ABrwy2UGoVU8l4m1cmo/56GxJ7Fw+c1xz5bncs7JWBbzAh1
GF7e4RmjkebITuL9vN960fRjZJmsmTVPnnBbFuB1rA1KhiK9UrVqd25bcCwr8eUEkroDaLd2ongl
uAaJCoMjipG9XaUhfsVUtZeTUaRKnc7p2gmsBUmCBN6NxlMAqRDPSmh8nAGIo8CfoMXVA1OjErgV
E2ukW4YgSAXudxItHABqasVsYydLDTddwaIIhe028xvnIOZOppgRGVzojJDyy/nke7UeCVFEpr9i
W+Iz63zcrOhcFmXpZOPZo9NT7sK3U4TN1clbxU3k6Iv8l6NnvcsLeA+k6rQZWX2Gj7r0+YVKGr7z
syi2w7hr3UOrp40quh7L/qeksxFVWEFGuz6Vl3hIBEs2S6bCs9dXl+0ijVXnbBAyjozhhGepDdxf
vWTcFG6wmJ6VqFRFjqcqa0GQMBbfqDe+8apE9pz6nm3wxJNUd8AsFsqwEgS9lIKICxfaMa1+K8bj
IoaU+8bNcbgA3VQvwj0r+ZdLlkEB9DvNCK6xw59+KXOdF+vSm8HDKVlTrl0nWRBa03apG7tgS3B+
8Iz7LijtecUehmmL0fRhcyu9Iq7JRpvBgslCoJSbcNhJFQXhwFmTEYyFl8TqDBGDsm3TDpS2+oCi
giPntWQc5GLYOlbeyOepoSa8CsnNAGwIQw8N5XHbURxeuQI9PnIyIuQT+seg30veACXFxIf0u1Oi
LBiW1I9plxFF2HI5GqL+sag0l6HZUI0byetrl2vwHCjNr0CrB1dWO1MToWrCAwpAa5giPGZxJycN
o4cfHE1zp/D7N/8bPYzG5imhP444o8ceaQHD1fCv3GeduT7e5o5EqtSIBixWKOfiA26SThRxGMWJ
VYr9HwUeGt/44WwQue1brqr74Y0InbXUyEKim6/8UTKIjI0Ia1J7HfAH0htvSrfaK7fTdaz1W7bx
yMNptu+TMpIzjBq0rKng/niQpqBFkYG4xjptjfa7iCn0AAyXVt2ldHf0GTCnPXcChOmYbfwNAtb8
gaRJEsoG84xQzw9IoC0eW0h9LYLKYq1q6xgS7lWwaMoFy4TaAyqJp/KCdbqysBJXfFe/guy44xwn
3fx8Ic3U514DY7l1jAGLabM9r6YfGbSmRRQqgtIE0yL9MhkUrVu3fxSx7w6bqybjB1I1xs0ikMh2
lbIu31s9kTDoRohL0n1LAixB0Q0D3PJYmmM29o1iis6btGd8ijjuR8tY7uC7wmxV5bmnURmjKo41
40jti0OuXpSroPgKhRIPXGVXsSTmAoMUZtiJ5M+uSSBsa6XzyZSCOrEIA9mFytJcoXzOLTRHubri
USptdBxTzfjKYYJoFobzvYL+CnhvouiRDTvMr/H3BNmq2Z20CXYkX1/Ni8uhJnkATR6Js7T63ayj
C08HGg7mqaRDy97mqZhPAFWmZjHehsIyF7huSADPoKasn9I/5b1roED8JoCa9IDcsUdnmCKa9/Og
KvMoV/b3b8kOKRDIlS6ptz8OppHypYfWQu13ze5/Pr4475+1qboRdF7n7D2IXDXC5NOLVY3eFsgE
/cxe9JqfxI9XuB171I4OMP8j3Bu8nYjMfM0eYTqX3gQE4DWDLsgSXPI+HrAWulBbfJDkojHUTB/v
SD79GI/Tzkp9Cznc/W2RdNwqycm/6PF8goprtWxZISfkSh07gTwmym/gvtMBn34XXnga4CYKGh0q
iIk9PilfM9XCSXi+EmOeZ6eEK/O9FqqwMNKcg+iAU1fTW6T80M0G1tU33moMza0oEd8WfmMfTkhq
zk8STkufS9oadgdSW5zTMlMZEQs0kNDFp4JLtZdORib0HS3Upc+Iev7gjhub51LBg36aCAWxLQhQ
DS3q9RDymM0OyrSTey4pds3XxP5qIYfBCh6ASKLGzMcmUEspRW49L0Gt3M9W52pHX+4AVYzE6207
hBdKJVDfNeYHu+IThQ8QPoubkqgKLa9k1yBFAMSmU/Q1Sm4bAT4ihIRlKkhZoHjRZ9AMYcdZHfM8
mESROB1F4fykpiVU5igUYLK+1SXyz3/EzjzvFy7O4RztZe87R31d1z3TRQ4K3lCrXy4WB95nPl0C
hOwaMmlRUJGB8izq2NgYfvpP53uY2bTQNsQ1yh6EtyoDWayPDrf4Q+MDCKnB6kkLLpxycb5d7xkb
k0qryvhsW/vLEJf14m9OA/DpaMXYukwm6sjtmp88q2TB3M/iFiIi6Utxp0q2Wn+vHlICBaorpN/f
U79LEzOAf4Z0aXD87clHSH10DKlkW68kXcAz8btGMz/VXlUzgZpAiCHxkbCzwhhIHRTJ4qHAEedA
UY3dOzoHBJ+9IDt0Sxh/1oVAx6CmeDIVTglPDIoU5G4kgxY1XAfwhiXX5gZJXUjDkiYZnV1Gs8F+
F/y7X18v/xj44EL8wpdvgZz0+q4R8+lDIcE4IMPDYYjYUION1m8FU0gO4VfxKanSN8sgU//SO3u3
e2nZUHNMES2TU8YdTiP+KVvTBtuQbZU9ygPwtdXLJvGSMTbHrVrgMOfK/rlxqmY66W2RiCaQRtlW
pBea+90qBNr7yyW5rhvJ2bG/ZRLEVFfVKanxl81A2jIotf0+QJnQF399rHL7fp6jS2b3pFp582Zj
ObSqYt9nAsRU+p8v93HZBndiuzWNokF4YUKywjXRQxFGL35k1c8VBYF+FtS5yNwTohwVzd2B+fwN
SYSZmar8l0Qyo4xSY7anfNajhiLe/WqyWDU5V0Oz5vqasy1NXL4RbrOexyMu6qi1l9QbQmvC8JqH
Meqw52KPMB+MM0yQ7u/hJ9CRer1V2qHnpbAAsEHmENCMpQnrSWhqR/bzkD1q5V5e5kgQW/YyWQu0
zABs25S/RK72X705gTUsAiNVZlsTryyXQ7tWmbOVP4AEu5mVbXYhQdd3v0yNjhPWlD7KevcPDTsv
gFSnphCPLZhQ9BzgZ7t/7qcxAXJsMM/mrvEALj7k+M2oPIFK4JtrqH3sCl/jlHhPlhuFvqP+C9iY
D7D+EhW0azmp3bqGW47mtnt4Acew5rJ9oyL/yU+Gvg5mSpZ1XWNQCFAtYFM+rkSAMZBQW5irGwi1
ZxbSsF4wWpjsuf4FDPu4RzqcJKZsViTQEiDs0LTmISMNxPi6253YS+ReaSrXn6smhfQ4bbS+t6uc
JmAnnpQ5SlklRmsgRcFiwPOsYRDzWVXYZgiDLYaIfJUapqsjtu3jg994FiauhbuzQPh0T0L6O+7P
G3eC03UzVWwcpjtxu21yp4ucN65fY1TYK4qyxj2PitaSLr5J+c7owespbwbndqyYrMvJoHU+8PXi
goBk4MBJB2cR2vLTBr68lnh2jqiB8k19v3t+Ge6mM+oY3s8PBk7F6imYelvOsbbb28T6yktS5bzB
76p24Tt1GZyc7Nk4RAxixe48NZtlgMyoYd5OIMWITmX6klQeb2n48L37aygZtKHd856KwvcYm6pR
S+puyozQpM/HU2bfWQzSxL4La1UyTvvdhkEEYUEWOYVQe1vyfzFe9KSOdv12z2QluxgZsorifFRu
Y0/CB89sHs5LGzVnHQJVeM9RVn6MkAfVjvbhAm0fxZTRmi/+KPmyj2704+6MhDxYlGYkMvMQdubC
VR1LEqsDttzHMQaDxxtvGDQbbTHuSPT+eTB7iqCVGQiiAITY/Qc89+vXp5L2bSOaBN2avAGCk5lt
xVZ3euGh5BDUu1cIKgM8Iv2Lhhk8XUzW03HyzbEGmQyQbun/SttVVQiDkd63dY5ghXzswAfk55SE
HZMezqSDK5imd3wufXqnqAbS7HkU6ft5DKX5fryB1Y4JBmdnjA+0+bozzLbc+wQwNmyhqHGLfflp
ETLIQKHsfHxAHMe2c+BfWFj1oXjbBUtf+gwfsb5GaGHmI8JPgOpiKTF1N/MASMT494rPQ3d/rc05
kA7Wr2CGw+PfO7xvx48nlQebPkMob7ua0FGzCU5+pTGjhyzUsKq/fB2ds2qrHeA+3UPl+LFpSMDk
ZyKbL+Wz0/A+57Mktr9iISljnh+ZXuLuRk55iatcwxec1NIHmmCZJcC1cSSmSokgV3TTygKfoKzq
9ggajhaGZDDYnZ9Adc4A1L+8GWOyJAQTyAcikkDmRBVUsIMQyDkolhN/u7PoWWrf5hn+E++wN6a8
0eKct35r2+hFY4HlYGjD6jsg2eET2NlbKuxlNZo68gHjToDFS8AAh9QmVEHCRgPsiW7F8F0RnQ8C
4xawBx+v0b/4n8lUKk+CQq1wJjOMXTAbJadtS/6CH0gQvsAnKh2+H4O9NbKJqW7eBAQwutwHh3M9
ihFnElLQ3F0pE6g6oRhoDuleUHpUocR5vzA2PVgzZNK1UV3SXAFes6KlTW9DUkT8rbkgrwpma2uV
kSaJgDq2a6RVxsDXs8zpcsNKbIlQ/4zf9pUz6Q82d+pRVoHRFYOnZesaOhmP+KvCL3HHg9f+z/hT
NxESWjjrComs72cHeZ3OeIanLgXJG7Z1Iz79Xv3SLVoo0v1+0WwegVJyK/pNg1p/Inaxfd6uMHI2
4SgHBMBQgpY+kYuuiZ/WsKr1iImzlwpt/TZX/arhufUntwzW7nojsQ+C94n08fx0rd+Ym4EQfbms
USuvhW4OSNkBvbA0OAA91fCjaTwR3A3s5h3i9W+9zOFnHz3pJ4boCPgvLHu85DXNKhGybh6fg9KS
jYAcPhuDs5an2uox2LzDKCta+iWO2Bb8NC6YxJ00vVVLHegTDIxS83GZJj62fygIHGeC81vgoYyN
kj20/toXu5Abf+JOTtXQT3sRDX+6bNsq3+Nyq8n/FMckRHz5xGvB++DQEnWX9viTjXtvaJ6BtVZ4
HgCSosd1FlYhST6Ye007BwJwrHneGvi61KmPM6bq5B9aQ4e6kXDu0Rletf6KKHIZy0meLYGKPIRY
q3lCnIPJbOkEGCOMVbRs0FxqBlRv2CN1HzbHtmXw0wdtudMzvU+qaK+j2W53hFHMtVZvzEWtJoWK
WKy1nM/sLaZDnwZI6i+4vHnNMIQ8+PE4x1BiKw+6WBczgHMY3+wc8LWONkzVByOjQ8nOcfEPC4d+
OEupM3knS5Q0MCWnPwEHicWaw6B1kDg0SdvSKd1OqOSVF818OzajwHZVbGQadDKPaFnMsfTPFUuy
gdcJWef7CYz0vmxKKnC0qQcSqz2jxqwScBZfH6a+WHMz/yekoObDMDPfnNow52dkQWsPwGGsty/o
9iNUK1aWIrpZt+f1GDHu1kFTreKFT1rmamO68YIOvttVuP+DMKtxV5UE8kb5LVqUWnMoGNGKULhA
lkt8AoOg8pgBPPD4TybGsZDWjS1FeZIG5T3UN+F4yW/t5h39+/OjP031xImlwYqZwMJwZ7f3B9jQ
YfIRbYelKxN3UHMtUxSLXiHJXDiyr+7yUhby2+DO1LJRMQRMqFjSzknxodN3UT7trPN4N2FNpGPD
2fIM3K1jBRzN6rW1oJ7GV+eC7DfzMZUa8qDQFnSfhNgJAr/t2DEPK44Gu0gG4NwDl2wygfvgGUPM
KQhibXgKScN12Wu+Q0we4dKYAQOb2FhgNDpO+Uncbx4VVkKoRLgFo3VYohKBbsomf7CY+JX3BIvS
g3eNYjo+RtUjJyI2As2X/C9J7AA/m7OJvclQb7r4Xbv9bblxGcyxNeDjh2hGBH+2EqVED6Oqv4ED
PQjxUvNqtkg+hJtDPImOfySwup93euT7aove4UvFBkM0dhoT9I9tiLeN9+NfHYotOv2nf4ZwaMN0
eno7Ac2WJM1bHslAmGiKYZ/UAWKd+dAaguT3fQTaSXUTH9ylP1xuFgvMObi0VkxePHGF/eD9sPO4
TMMwX3Dpt3kjK+P+ZbHnjkr5wsT1hP4Xa8z9WQ7gcFIDtb7bK+qLM7zrGlxr0B7sUck2M/lzytLE
cbcrA9PEisdUi4oEyNeQB7HgkQBxkElegsF0vuRvyWEUmY5DZD2bTk+m1uH/zZVWW+NfrS1nGMnT
N/rTb4sn5vayhzM9XBTREFHNfsA3OELnKsPFBj+HVNIgGgIST5wZQnlvxymQRde5N23VMP4EXhSk
ZlulPRIZPHXtj6cADzJE1ZsVVUKv9kD0FBU6CBGjxEejMBWv/w7FR1CEdUY5xhix9ZiezZfe2gAD
j2MHc1I7JTglhGtoex7L+YyQl4QtFW5hCX1jSfU8F1nFi7gRLLXV3ai5yD4u7eoj6rbteBASuRc+
I2Y/k+CFNWjPtzGjj0Fqneq5xr8Vk9gx8n3fT3FejBE0oMn2Tvoasl1V4u7qRZ2LErWHeuVpSnMi
bL5WufFt1zxHs3OIELvdrIEWCTg8dKswkNZ5oe8KTIXhobMqn8gQTRUORTo4zs3iHE9aXLVhHnXg
QMMxea92bwrvn1YbFX5ImTJNy3bpqSzMOhD+x80xtkcVCmU46nSIZTafGQB0HFxWjA0GsZrln1r/
CE8msaxVG01T4VeT7M67/zjV730TKng/xV3nr2chfxHSznwsQXvI5moTIC+W8l5RLHOKYxsgQDpS
ItBoaeeD/uFtMijHpzWeNsK0ntTe9SU01LUauP8lb9I8Y9nKmJBOP2I5wiWRng6hUeaojiEoTPHn
FBDKEaUiX/oYpBKc13NNCkVr5OC5FHCzBqaHyatqarpu5cjDq4wX+XcB8fZ6RfZePz3JA8cVNIoW
K6FIphTzLm+takCnzd8F7Lr56ws63WthXqxiNFenxgGaBSir21EYCa/y5iWdKoUJgmh9jOq89353
bxBg7CghqNyO8luOrW7iMUswWAOd2BFD4Y/I6yCGOpJu7ynn+RmA7wJSQFacYH9aDI8ss36P916s
ncZjPgS886GO0uElyOShidBRpEnMO5zNdrHPSNgyfVIX39wWWMe3eOrrJaiCaqI6EOS5XgrALCbo
0Q0vsDu/ECOgRbU+iEXDih7sws8RPi+CwOvog/6dQH9opSyDYRorKOHp12LUeZKB9gJP23+pFg2q
eRcWtzQcNNTE3JqZiODfGk/tmlSRK8idGWd6E+N+ZivP2y+Wap+tFl2jYxsuta+VrvO0IdnsmIqv
Nbdqg8Vnt80Ab/nfPkz7Uc6nCf9k7mxl7JxSH08rwdtxa4N9hV7qZ1CQYx+Tyri6bskohIq6Dm1H
Cs9yDbVxBaBeTr+eZBdcdLdRR9IvpaT0E0jmkLBz9SRyJRoaxZeeVgl6IuN3/whFLp8ozdDKc+6J
CHQcJ3yw/iJg6bOgyvQsrC/L0IEDhMA47MW9uXKWyb8Vv6+sBXdxmYhRgxsHkb9zEixTz4nstN95
0TzFosnCUa68f2OJRIrKUY1ZmsPb+NXc8m3QrR2G7iz9AWgGpndJD5iwbfhuDEQ3nUsqUs9Lji2h
6MwXBE2L+UAO21B8KtrHqqskTwm9Eg1lzKMXP/g6dNLlgppAz7z5KIE0WIUS+ewo6pcxZyhefrdk
f6CCxnmns0h7hWJmUE1Ap7/iidjIwpPpfSBRQDuI4PYwChEBhbXeypdyQBzCJ1d1GSL3YFliojCj
OxFE+I0UOel4RBC7elp4S5O0R7ecXC/N8Pr6cdNCSklz9lPb9T38gSLgkmjt26OruMfqdnCtTAPq
JUKS+HGtouMaT8Pi7uW7WscmFBzXVHKsFey64tl5guEpItLMPWT0o7fwKtDb+zo5bzR8vasjPzvV
4jRoXO8sWThAjNt6pPZV2Ed4Ql55LiG1cYosJUNGHJ2ayKAD8b6m3rPnSvxjZwwzDIO2T9zh0vV0
uTMGBRNBNCZR61LPis7d+ukqaNySbH36mDwkvQKVVesZqIhw5+ZDW8AJqEaF1i+vAySOUY1rGjTP
oDupJuj+YG2FwLbymdwCM8HvWoayez9IIuht7WaZIESv2fevksQ6yP5COFmnXJaD8qOavWGW1BNM
wvp//PgXEvZuczKR8/VmcHs1ryTXupztLy1Dhz2AeaXhbRG16D3cqfj65+h27Xi7VvDhUrlHfuk7
nayFTroBIrsGA3AS7ADnzTvuMwhVTwPo4z6O14KB20VD9jGFqphIm1BbrF4oIfnQqSOYsEnas+1P
sWf4IjfGyPF9+3usr5J/OOS4kT8N92Yuq6c1g72y5CcdKjMiOOLxGG3sM682y74cWNbgdoNuPQdU
MysbTsftCzag2HE8yRH8rnVfd2Jeadh3j/Z+Q2W2Tb5wtnOeeQUvfGD7P8JLJY6ZP0JD6fAjKmK3
z2WNXTymwhPeY7K8XMTS8Wdbc72OcnNe+q87rx3VYgDoHZxO9WmCTj7pqAad3ncMQzsVUt2+37aX
+w545xJP6PObiOrLm6HybaxrWnthH9tqWkRPWCtlz2scVHRKP2tqgG2JUmTzNPX1nNFqZSPbqsZr
+ZGy3CmDSpXqO7l0+lJXZYI3yLy1cstCR4UE6NQNHvLyUISVB7Cj7533k/crFSe8vL5Ed1GPY6aB
Z+dFJ+nWCe64XxjaPsae3dreJia2RNMkbKAbBiQnO7VPiO/MqoT+LUtkeDtMGQICWhWAjn2K9HuV
pysZmku5KT6mQ2B96pmiEXgHdGQzG4T8+mEh5m9e7XHZ9EIqLoJ5PABCJpOlvNuVtNhPCTeZm66B
8nFrSI3qE04poXToEjSD+uWOKsG8SMm0w+pZEF+aUtAhst+WQuXLSis9Nha0CP25EPTNXdl96nno
KpQb1ox491zfzN2vu7iity/BU9uy77B2MLypYqFtUUgN1KiXYa8GP2oAzHUNoZQxIfBkpv6V3OiR
t9slqh0PtyVVxnjIhlNYSyx/IDBYqJ+xiJEx5dgWBnX/DobmMOFezTauGHnrt8QCI3nN7jcS1RK9
oZIhsDeYil1XXlz5vDKbk2w6BZpeMgrbPw067XRSxMT3HrLVU6mCaz3rnN/OHeSeILRnw/QVFqgy
NAhN8DZ0x3l45IRqgx+GhZnOU6v+q7KpSEgFzxGxBH5uR3C5uLfqtgKKjgOdb4VsGjhwL9uoJ4pL
VWTgkRFtqJUU84kqT0ySC8WU98oTtWWNMxl6QFl5CCLFzaYJtENSh7ETXH7voX+MAcCKFCfIPL9a
6im1x7O7dhOEYLV0QoJtCnMPFtS6U5aVMxS7Vsm560y9gE6DTy7XFJ7EpgToNmeqO5QnfJWb5iOV
hjL5RtZOVuqE/uaWHFfTxjPES910RY5er4S3u6qFCpktatc+2UHskcJjvvPpFluUw7LnZwW3nYVg
o2h3DnLg+Bmr2KVxjCEIlT2GQqNhcnaYc4ypEvjEXt3EeOYRtuLosBV8posQdz0snF0XOyXvbkAc
iJpyF1rEmBJ8EGLKbB45IU4oDr9aXVCcT07z3PSs2rRuq/wSjlitZObmNu0Pmz26mAOA3Hl3BaAR
tHoc4hnSSMgtai0I60XvzZvxZ070ZByB8wkoh57dQ/5chIJMH9cBQRebrdOFVKAHtV+BezKIWqdV
6N7UI53RiU+HChmggdwehT/4Th+5J/wnpOb+O7sUZJKd0s4c5wO/pLWzJPRnAhoZv0Sk203wMHP6
YT4UJXFwJKYGpP3c8WvpzIsaBHCeok66Be/BrAGsAX/CameshoyZqt8JLDN/TlGtE1X7vJ7vTwbP
wivYGY+0km64CuidQy5LRkPBoxGENbQZwZjukX2ZqH9fnFggCBhQgzkszc11ggpUBnpf4s/TcxRU
1/ab3JqE5F9EMUt4dcEfgRakA265Grpn0OFsWw3RC73V7EgBKitu1Y6ENDGrjgrP2QtHGQp2b9rt
I/S9nd20A/pkgd+I5UzGMJgV8XwoMOMUdTq7yybr4ily5zpocQUv1n8uydD7KII21vh7Et5EUb0M
S5/j5xYY/fqp+XwfYi/LuTFrGstaBzTjvKLJvFxKjieq7foBQ3wkDjelwiYt8niz7ctCqitIB4hk
AvPjiCm/mfQ77kWxokYkKvz49nslELKuzqqGSGNl4sHVqqFBGX34zwP4f8F8WujwmhZw3mN0/bzR
nJ1sh3Ke9bOnKF1feXH2pXxmv+lGQAu6Ltl1E2JbkEHwLVapnKU5BT8CL12WiBLmlYx1gDau/3Ll
KyW+4spLhrMXLfKoobD48K4liEFvHY3iqluuJFcvml2sXOaqtAmsVxGnoVe1kPH6LSTeTls8qhxE
y5pN7IsZG1sNKysYcOkGjnbPgN8VIRhm7YniLWZ3QNJD+Z4763IefVBJKmHzLteiNpkEZabaYHXI
6aV5BaiqS2wuN3BrbvVNqjwo2ULTK9zNFOOGD/2YmRUV95Dn2RY5lb30+EKx93DwxBPuJCB5Du0X
bSiAoiQG0cSZdsbMLOOWidRpzktDa/yyKgnebH/JVnA2aGHUFRME1VTrOLq5EKl+YgXjvdbyLR0x
w0tgDst5T2ujJQGoaZvSD77YAgbVzshYaIS6sLxH0aEur81YiqK+/WzgxjL0dmwndZ1uuizG/EhA
0ErbawEUDAVggHPMq79Fa/DjWvYvGfnZQcAzGqWOjVp6nTUZRGCVixhtZXuK5+50zXf25BBen5NF
tQ3hCX6meKOXaYmliuvRKEFmC9PvXWUW9/1Vpv9RKiK+yzN/Mwfq1ZxDDf4n7KtKbYMFaKbLyFAh
pI9WUWFfbZkZpf83c4ykmCGI1wv24Lc5RIpizXlXmNisiLYoGsOF5n2j6zIDazP/vfp6XE4H2knx
j0VDjfQdmtzjQlaUZo4FMA7xetM+8PiQgAIRQpByVNkZfEpB3TIF/VAhG73Pgl8AdsrUvTC7EXir
KEU9yw70LoB8jdEY66ErhzWPPrZK2BH//Q7AdlTfusVBN1vPFBHc0PkuwcyNKg96h9+CFhJxQUyG
uMY6nMc/jvFbSzms4iE8T7v3rHN4k+MywdHP9RJJWYWXk+X8CHytfk984QxcHT6UMWxKu0nckvM4
Dzn4NJNEVY7DVItl/KZxh8Qny5lA4iReqgKUjNzfPyuG8QYY/BwR/BF+3cDX2b+jzH4Iy/CHM8kD
C1fSKr1I93+eSg4DIV6ao5C1bNFBrz8s3JXrPNvyDuCzGBHCMXvA3xar1voomwWNqzIsmuVtDMVb
FY7DAjZuWTRHXLtZGepsgzGi+VGkIEs4KJEEStKo6H1qrHvODd0UBuHTqJwLLq5t5pKyJMU56PZH
9TyG+RtiCqbfpk/r5ERj/kZEDnCtr5kMQgHKeUdDx7R6YiXGRML+iXPDw5daaKndeVa+dId36czN
P1qSmZrtKF5ectWwpotC3WW3/XF/Q1idZgqWK2lkc+7gh32A2g2e5s/9ErEhUP8ezADWkeJHDABx
R/mEjfgdKvK58l/CW2RZtYENsE9RLmRmxWVQfouddWG+IlnI2c7knvI1ZQG0OKwvbsL8BvL9TyGO
KshYB6TDZJKslMvShnE2+w0mPAus72IC1WFEA/Hwd3wcI6bzIXY13XTX6HdgaUD9Swm1aKJQchQx
9LqWPW5QWGhMbX+dDKQVeG6vR7JTHQ+3mHJcFj2saukbB6vwnYMeY6AfYZIpHK2bQnTrombFEusk
ClHtykG2xG2Za7cd6tEIdoy6WM05mmgByXQpDnOgmFshAmZ9s7eVKsKySYMV6pkv4BJjMHhHCouz
jXZ6/4u4KUargwL+/5luyUPruroDRq92hq7PM5u6tC3uqMCRSO20Meg6SXmndhRGy6i/kD4J/7Sh
W23mzzKWv5OC0PiuaKSJ8BSp/UUtjiAWw3zmnFedEb/KBrzfXPua3dRH+wgab0VNwxiQ18+5fkTh
sP9PC9sd0qKxx11pCUcQFbBbvgl3gbbV3Jn8ph281M+s5SuqaWPn1PUCsSu5hGAGRRVIWlHUWCFH
rNxwZR7lAPfK58IpapdNSvL6eZ4nbLMcVYWJaRpc55Q2Gs1S7tpsmPFShVt6SfyEpafRubLzbV+H
a4sXlJepTKk40D0HK62jvcvS8PyyIF56+i0AKKC+9OXNROFINWgzQggeqYHtKmn+QTbJmIzGD8h1
wkDI9tigqRemsDbxDJZmlLEBN7Q9k1HZF4QutE2VnfeVPgajjq9PXToap7TSlWqyweUYZDA5wDY6
WAKTGVm0zLq0NLUwQSO+Xj2dmMHK/bvbnFJkUYX+uFpHZknh8X3f1n7rMYFYOBGu6u9U/dbJUrPc
2ogL0BalBZN775rORBnnj2j1+gof46dkh45Kdi3czto8TtweLMgK/GfY5GYGPuNuujY0LmzAlHSs
dQpjjTPIg3MPz2G32krvIGoSHZRfPYbLs3Hi0UqBSIvv3PVr/Dn+ECWWqWZPXHrrUq+PB5iUrQPP
pkI4bTbztx+sIkEYNHcorHCVubbF0J3C5XWS32/rbSz3YmJFJ23qgWnhtOuf5KihPd9qPzFOOdz2
htfFvWClsVGHk+kzkOpDQE1alq2dmSrdDd/bng/EnUJmrS3UfYAmleXo6V43aksNzWaLTSYDP7Bt
oj234PV5YiFwnHvrflrv2bjbk7SvwRBb4kuhxAVYDS3MY194+M7AtHkLTsjLVYaIU2vd6O0uJcvG
9Bt73MyF9wRz++cYkfjnRC3/q5qjDudw25aH773KwKTvqYHPm0m+AGPd4AEQ7DbVYq69TFREv3jv
pneqZQOFvka4lfokrtSp/A6lkFkp6TZY0ZMGmFnxBa5KfxvugtNMh6zx4geII1zd4ZG4wHiA6d71
1p3NbMRzjQPECOjO8TSNeeRJxFFotzTlC01yfFiPQc3NCWKsAhoyftXIhtKqd1iSB/j/ri+Y6Exm
coyj/Fd6ovoo5blglPAWrnt0EbFHc/Emr0XVECUp8EpvX05wMjzENM1dO8C1ciPoPOUXqwG9IliW
LA5M6gF5ksK8MoqSwkZb9XPTb7Sur3Tb5U4EmPHnUwmQhHKVn/iqqtZl/6JZqyqSJYC9TNVxQGKW
lex/3ORZv5ugiLwg80uiyyOB8epCuMbH0gSHeNFC+pYxz5cga2OpqTxRSNjibsMDU7d9yBEgA63Z
fzNIuN8PJhwakCtZtl2LCIW3iSxAO7e9hTDjn7CyN/STB/DZZfBSl2dXVTrKK0ZM/9VOoRNjwy5x
PipZ7MuqIX+dvCW5hAEomU2YRU1ZagLYCD8RYRnOrHyuxkO4uXyFmTiuAFe8ZmlDv2GWxGI+aLQ/
TbhiPDrcPfM6T8D6oL1pmg+wNAvdLCpjAyCj0V3hDJ+N9Nyxi+lEnBbv2olUiYVS5l1EFbGISj8v
VHbAOtiwO0hIEWjt7teWEHjXTvmUnQRY4105XWa12owjjz73sblxiLxaLgc6sJRQjKjjW6Mje+4v
Ua0mI5MsoOOkSdstxvTwkImL/N0clb2KxFppCjK3Bo5sKbikgD3nxy9S0SHR0QmhH8NY7ffa3wNw
RG8GYCm/csWpbvTqCYkNe8XDHb+tgCVNNXPPRZ8nVJzFtmV/TaQNhJ3IsP8aPrifYHdAuBtgLQjp
9RgDdubGOcluMnYzNYDVF5uwaLosmWwjo6rw+GOcR6+AYIbcdjPLuefIaCqFsgxt7rzPAf9v9XND
8+/fQw4LOH4mbcAr4havOxkL1a87pDxM7yrrLHMV/x3Vm4V4JGPqYDkpqwJEzxIp/0QEWHtBKYIP
JyMAZSqnHHWG/yEayeuXl8fvyhxfOVR/3wYSmOJwQe/WJ/C4pnYBEhX1de0+h8BjB3cq5SIcoeMu
w+xSaAAfWYZUDuMNDF6DoXGlD7P32CcfD0KbL4oS3PhENfogj/z9RrEDVJeu2c75PH2IyHrZ9nzW
Of0YWNcEMowgRAc/DX/U4RbiqE99d5Uls19CL1vF/drzKVDWklmG46YQ7+QgabCKMP/spUc1XeIS
2LKvXyY8XZE62LbPFOsOpm2v9czVeOq+nBotCRUXgB4E07QDo3fxAfIHBY7xOm3UAxyzCIbZZ7oD
DxOELpCwCQ1jCJEhWD1yqMn1vGUi45grvcSQBGMEDpwfFItxzWW8jaitigCMq7cTAMP37feaETUH
uhC5atntdc9b1RFivinC2onKDgprUGrgHBOVnkh6RwiAlzYxVEiC/J3cV/pmPujtOpgW1s1/YMtH
QCZogV46tbkEQpiYOBqn+u7kihrXjsRAiaZgPQuPX6snJpnUxX28WI6db0XF0Hd7T5DdvuNUKqqY
4UxhTJBqpCP+k9YOT65oHImjHnmztT+6tJtSvQOAOYeRctTHdxAv/AkQh0kEfjF4Z/JK3OidzlCz
toAqLh1oOtrzWNGBVFWBrgexSZ6YsrZ1r1aIq5fOuDwlU5SRrVva2kbFGZwMUwkdpYWRgsl620aw
ObEV8rHREx3yImsL1OCE0+VjU6B5odztIjuWDGr2uml9rSt3/fFH6OGqLxwzTNhbdmKuwh3EobTY
aFZAKaiHp0YkOZLZxsPS6+6ipwBtAOan0H7kyoSURWa6wC+Hb749fzL8P/ardqSRSTHr6ckqMxG2
CMIOaa1+j5RMWbX0uDAPCFKmFx6HCHeARnzw4TMv8SJpOJa65KJ8pGWAH72TGzyC47i1+U42pFd1
oOBuUKZFe0fsK/3H3/cfr/xUql210k6psQ8cJo4NkEzuZPXkCLjaYe+BJih90EbOdOaeifIVLgbr
aeyPss5ncFdq2wUAT1C7iWLaTH4uUUHtC1YBcJybblo8UsdQfitvHjLdGFq1NUxiHbA1t73obvKZ
FOReq6FyNhChbtqNlwLd6H0MAukCymlGJSaPD/45M9OBRWsXdU5m+Rw4+gIt5LoEXjJgfNXUVRGo
AOsSX/tDUBEYcQFD+g2Y4QT3OzOwWmyN02pkQLGr6cBIJAG2HU9GO/y9H3TIt3l82ZY22rFI0DIF
He47sX1EFcBX/mPa/sxthQRvKPm2jFuFs5v5i1n3mXnukPx2y6iVsr/JGjLGcxc4TTIn0Yl5Wf41
f99y2xQBX1QjFcz9mEVYaaXRgEJiNMNry85m1BSU54gGkfFR3YHH07GDqEMLZUGsjVbkk/O6s/U8
kqk/+q8W8ImM41aR4JCXIYZnxmpfCTtjC4unXiuw5TsqWLeC/18Q22/vCkXUEPstFuvIGzdqO9W2
RZS/Gz69QJABI6nIdGtY1OEIDryPwrVZMcH2boe2/QkHqCAzLSI7QsCwpPM4OKEZ6qp6XyjfrGn3
j755pYaIgUlgN46/kpoP4lQXhPk5pzE/o2kXeR3mjLwPOov1UeORNNiR/geDH3OXarxSuROyO8f2
mvZcbzTKLtFmLOSgU6CjrXk+z5e0+N3X+4C0EH0f3x5syDfmnoOO9orcGVuXPVJG8E1qQVi4ea5s
9y32zKe9l4ie+8XJ8tKawMkg4K7l+06fc/oNVz+Kre2lpT7lePTglFDSQQdNkg/hYvk+LX2bcI/j
w4aMIymCaVKi/T0ViuWNHPAEUh1eflLjzkna6ijlzlD9vHF+feUVaDc9tBfqFvFJqFLH6PdEqcWX
M0Nr7gDkBAcBNHAauHzW75hoquKoNCyNeta+YqLP2PlvCZ4rMHhIX/bqfJ9jRmsjWlLnUKxETqG5
ExFQwWrWLk+Zg8I++QrQ/05XWpheZIxywH/i5NiC4P/KLjsetiy1eNwL1wmRn2MD7VNalSovjs6V
rVWAXweqqMXqXJX/yYTSYNTw2cxbTp2H5XpQg3n0KKP9OjmfU4QD+JLCvzFwSMyE9KXz+m05KMAI
IpkxixLSry88LOtyBynsjHMqWzkwN+RZ+W2hxrv8RjIaVAEO3hEQCdKMYmdXZXF9UN1HjEbNZalC
mXyDrZ7Ja6Pt1yFpSVMWv5rYNHuYD98eIF9rG/PU3+B5I3I8CBzpGbranRKvYXytZKYRM4GYQzod
/OLlmNCYBS69KogpkTzknWPAGxXCsVcpXykFxbP8njkC+mGuKgrgisL8Z0fbIOuVw3EfrhTy0exq
HzQOoG1Xr/EXWqVO8cE9c1nUtrpFPXrIe5JxeFBRiyDJYsjSdxu5yVJHjcVPgJPhnHCIaUzvtBkj
d77Kf/tVdo8mGcvKIv9ObxiJHrL0BGRDX1NOtScwKG2uzwl/MI4gIfkKBKdPqjuTxbbPTFlQuy55
vWhbBMmIPzF7fl/CZEsWnntVAlyhTchlI+YNQm2XloXUuB1khfWVCBykI92qng/u8b5F0MQMNtGH
aNcyPo8rOwqXEc9X/RXvGtypDA9PBy9tK81x83xkksuYdGUCZTZtefqGC50p8SKRZJ/Pbz3CAYkQ
n6+DhZG4nFdqoGx1klAlxkv13IfOIAEUog4SnT1gYRVxMNRvjchXPDWZIvj55F6UBnfmkM0G1CIz
4AEhQbsxVfxxO+1WCKQTd1RfouNE3QcSkguTCo0mssbugs0A4+Ihk4pF6cXER/7fkiK8FPp4Mmsm
PsqAq20u/tEEMZ27LbB/n8UAOc5AwtZGPcQSgR2LhNCGd8Vvnmy1RXE+/WzdnxpN4p505bbVLCFr
HWwdDRPiJs+H0PxH8xrcOPlnaU8y9Sx5Ny+wyXu7+UZMwDAEmKt7r6/nB4KlAP1PwV0SMVBphKQV
vqDUhR4L44xGi5GtnX7ielJWVGAQ5oi5VboqO0Ounpxe7XeGAUNPSeH332/yLyJAUIFNwv3M6N9L
UQdAn2Z78DInO41DZYMXx04UrYx1Ox0/QXG7bGs7BPDPOwYmRW6agn6by6iOc3LSq/447as/EzXW
2fwwQ4GRvtiuylU09Oi66sdi75pcqA1HGfjp53D0VYojXAMkiDuSNPvLubtPNw3kiYY/wL80QhzF
TJiaxOiZDOa1fI/c+2sTfy8f0tbLDfxTkPlthtLaMTMNgDVRMCR5PaiJmv/tNiPZs5Z4FLVHvbFq
vgyBoaz8XO5kcUZas+SEXHajynde3EWy0ZupvibFEFlUsXuRReYw1GQsZlXx0iOcxqchqqs1plgF
TAQa4P0itXsHM9uFRCnc0B0MV9tjCZ1zzxegjgu0cknXoksDdg3LX0VhVWGaYjN/6F39tamEI0WF
J7MhUCIQ2lnjCCJglUK02DTHTt9xU9vM3hoc2sWkWnca9XdL98wWRXIcPUNMfylrDH1M/4tSdNBc
UKSOvhystPcES98jOHCNB5+1h1qXZdZllKBdjazturGeqT2J/75eYK858zwpm30A0BzejuquRsjD
1+Y83JKpvj/AD8ALTSz6ToqJ9Ji1q1PXQVnVqCT0celEVXqiHITUogHAWhTVrAP5V5RWFJHlLHxT
U8FDlBaw7YZ5hM0DoGyFgiEx5fLNeMYLows79PPqYHVMaab3bn/BXMtaZ7jWndZOzOI+54E7S2p1
fdxaWsRO2xNbWPXKfIyK16f9ZSzcZnO2OYZWzdFDTPKQM0yYL1IHBmHkhCUzNWWCSWLQklaRJsdU
SGjGHRdLjnJqZ8kMEFzbcjpWiAw+1J/+xvJm4+NSbQ8NjJbgDXxIAtQe3LWWNGTx2NOSi3CZDvY4
66794rSaAMhrwvtkafINZ3rSdQW11XfM5uUy2efHQAaKBuZeGGPpH5AVGRURevl7zAfeVJd4xyMl
YIK8O7M7npMc85gxdh3Yd7YINA9gunz6xRYMlmtGAS+rmWn/cRDthAJxfUc/UOfFvLfrVYR64PtG
utgZitGdCZhLWfCkHTxd3WvF9udGHH/i2Fbv5mvkKjJdBO3hWRLHOchq38DoLIPmT6GPgwgFvl6r
G8nGdP8s5Y91IvMWhW8UnQdtA5jgEbIfimFwHP6dMLgCm3pYfC//MOBG4eFXX4IyYXYRIuTaSgxJ
9QE7eh/L0onFWdi6wx0qH/rKHBelzk6tIowUWARsGBm5hVQQpAHnTDRLy2i8vKyp+i2slTefypkw
UdXIdFGKjIEauftYWy3VsvVmnLdVbSHJN3Ms4BdlZCZaxhWbHV6H18zgMJGotlhDPClv3Gkn0dfh
KKO3tivmgGRfyuo0GgjuypEoCjEO11zM0HfLaQ/ud7iv+8H12tvAPOUvtthPLAwHjGHz68kQLAvX
Co6ATagcuOCQApuFegM7NeAX80sMvjR+oVMENctyTbCzsMxvLuJQJPQ44IZBaweAEFy7Fmgi5Tns
CDh5Aqa9F4MZTSXPF/u+YHu8yI4KNaShiyMN6vHHgTVPTEhxZG3OcCfEcpLj7cQEAfL4iYVeicAA
07H/nCUj1VXsTH/+12oJY4Uj1Yf34/jgRCaNs8vxi0OpiPxDw0h5Ip0eSePbobVvCEclG7H40NXk
tm0N7YkCuXyy6iYCEvPwDCM8vj6O4GTd+DDvR3imztcsxfzU2DZ7T7VbjK6y3Kz6rQP2nMJNpUiS
t1DY34p1+OKJnDD7y6G35bDT8oPiBkuZslhkaAIbqXioDWY0fr8FomvYqNp3nyQD43/2KoFwTPXL
joZrgaDXksQwHu60kA/DbzJIcryBWiNMClLc9B+0zD9RmGh+Y7GOVreRCEbdI6PhePdcbwhA12Go
l5yQpLgOjRmFVp/uY+NvfReJtDtE/5xrSaspMyQERm7JfKmDep+0zw8AARFByS69K4GvM3rxyP37
/GVN//JefYhIXICoZt/Fdct6bXjOpu4tksoL/BZD/q6sus1UhmdTcGsO76oZ0+oxnDBMqPgni8DZ
4rjaEdrZUF2yDbwOT6JhdJoZLYboOXL3LbK8LX3919ZuB6/CRk11GKMkvu1Pp1utSgLXE7YNGKdt
8szzCrijMvCfAnD95ZsEcSZW688NV4gJlc7SJsF+UpE+K7f+DJ3EuyOOGtPE5TDOQHQY8e0AD5hR
fakMBG0wehOBLu6qgEPk7wcdHM0FoTuVTGf2R3IhxjS2CVm9/JvKo1FW4+8jjjjpOxiWzDBvGTr3
DbpN01SsvAf9/gHwlM4yL1qisrp+d9KagARbxyOTD1m3EB9fQB8sZ1+I1MXoSmJo4pC+pIjk2Yl4
lzH/672qimTxuwbYiyjA2HAMLO0QlcwyZ6iiGWpxBvpWJbIYDaxJ2Z49nhaQNEsRBax6TnGtCdzn
fJCoQ/5gcdG2WfKofxwYDGzcxB/bkZp/jPlvNr3uuTXDFUEnq4OHO+7DU6KtWo3wLfzzhq+K7reN
wKx9rjO+CWJQBtVhBQ0fbJmxK9FfCrX/onOoazF+05nDMQyBszVs0PIy2au6cR8mG2CQiFt9AnlE
eSqQSK8lMStv12xk8nST5aI+D7+8NXMchdhN8KTgydbtBg8wToJYHo/8PJ2tRvmkoiepaTapZJib
Gd0mbGfGMmvxZEX/GxlK3430tQAjlxiQfNpAbSwsqiE6+Iax39WP2JaD7lq9d/fBgobp1VanczSK
S7KKf9pFZuT0QyOam15jiCnToY2/k0lf3Gh2dZYF0cNhenw+GvMwfGlK7o6S5EaH11OYN+MC0+rb
5ToBIJaNXzUykOPrhH4p2xIncY6BiqdblP2HylJWLqwxDpoYR42pfEgyJDZa6SQaABGu/ecUihxx
lB9bu7eYqOuZwM1hisTVxALLKAETKkjoD/YW3PsopJZPCoh9bRJt1UB4qJ9lZ8zdik0yL1HfmF7w
qo1v73ZUjwliK72dR7ktgzPo3xMcs4BbXvYV/2CyV7Jn0LkAP7/JBzkNgvylFh9/kcyTPTa8mpLF
qrK/FGRjafOLLi9MBHgHADNzatEhfUPCITqjgNZ7YJ0TN4Awk7omzNMJZI9woevwUJMV6kgI3/en
vxCo4Dn/qXGg7kL7QUD6Tjy+m/J1Me2eeYe7mUX6HsYlZA2a1W465i88ml29DrtpEAOYxRTxgvEt
TBDFHPNFB9Fh6PMEYhGZON3BmeUvankrupXLHQKxHOFVRSXULZYfz4lgnxZqv1LssMg6g8kONo3O
2oAqzbx1yWFDmRzVZFnsur44XaoIwtw++XGjXpqfaC/rx2MFwX9yPu4BDZoinDOaDu+tXlBKbWjY
w7AnP+dl8Q0svdlCV0S/s29OB0aCOikLcI3J61npt2fDkAVlDlMp4xVSzeZLzMHc68LOaKN7fyyV
1+373IxIYgFcDbzDKHds2KBfHxmUtL9afunBOZUoXxy/YklKdUI/IeVIxjiu+wJKdpfhzcEEd1DA
LtnlKfOdrIhYiFNqPavFS0zFle8jRPRx7IGNugu5Jxgx81f6DFHqDfdP8ocjbWzw+BshcExPwcdf
F0TG/b/6U8EK2bUmwVnFxYdWAZnYOG/NGXblSPOf2NdOFLJmFX/+tYH5+OBq4yjtf4qSwDK52phL
r04ETtuvavE5ROA/CPnkWncPn3Z8T1dOZ7bpcBRVbrkRPhBz+SYjoC6VoWJNhz1Yc3lsqKzsd9za
YP23xbqcguPIyAdGdiOz7K6iGM/ADfsYGqVMswb+tkXS1KpYcBTvjLAvmOMpIlpAS+xyyLMjTD+4
2skJClHvpGsRCyZOexiMQooD0v+uoapUmipRfWEqsQexM//heBdSR/5VK+sCw9cxEE4/JM7j0MSU
Ry0wmkouoW+jDGgkftiJunsNFaYa8E4QPP6pRF4pkskryJGV+ZxslTxBupj1FkH4KKzc71Jni5+F
H/jj7dpuSEW08fkVNw0nPTLfdqsaWEcz884A/kM9UDlDmlxpk+zajbALh6sNXlgI+yVBjOvQTAQJ
yN7p510iXPW9qeeqNdX7ERV6F5bD/2YFxzD45nOpWPkLmEGlF1WdavDto9mgrTzQj2eyTHR46Sh+
igJpu9VkCSiel1SCg30eTGzcO8TmYIbluSbBQYqOX6TRmgsb5pyLBx3GMfiB8a5p8vlaFKaB0lNZ
iuvWQYc6FzehlRAfawf2J5vH16O4RH/mf8QKe7wa4IVXCCyXeetH3vwGKy/OgvVnGxR0pqoaV5kZ
qRv36U5jso7Xxk0zz45KHfxFzg5sfrWhqVotNUo75w75NQ+qa9R6RoDucpLmYCsNeBpXAaRAgHVK
pnzlgU063Ndyy1SDoF1e9sohiHHwpajTpwJNbwfLHgG54PAwZiiciMApm2Fx59Y3HaYQxXCN+6Ir
4ZH/ZRVxJ3P7jAqhtf7e1ncAVcE1OsowAjjlfZTMiqprwIdH7JzAyurEJ0MwUYPVFuMeyR7Da1AK
FjiKFW9Kn+XDD7+oq1DCspye89ArzHesveK1dnWQ7A0hCR/P8cfxynvTtlZ3sdlUesPA+D8fz7UX
dI6wW/g4mwNXHww7Z6BShnIGr4SvhtICprebqWRMhsi/7BpoROb81tvi+/GeArw8jgVe6fIMkMqE
XBByZcZZUM5LbAYBXefyLYI0P4k4+HS5l2q0anH2/TkF1/Fx2AwCC486eIiRLHHe7o0hY2NE/Pjo
v/SXyFETy0maphvCGBmMij2G/k2Ih1Ojyo2oKIeYUg9WDyMCCBXIvKNySvps2eQo0DCIqmdpvAxU
9cgn7C5+pt3T0v098YpLCprystveZ7/Gav2cwgrd62G7R+0V5d4UH4T/MbdR8WN4DObHdTKjhpKg
a6UpyR0H7ZnucuiDjEJTbTnB6x3p0vVGSW9n8GvNojEoF6FjT9S3O8+V09mPVwAZskTE2ow9x43U
A1nszmNz9TljG57yN8l+39RyDqJgZLSXtRqBEEBRDNaOy/Embkfz+fl8BQocGZEd3z1dQsp4eB9J
dgDbfgZqcF59drDljxl4PZvBSdvHEGCd6L3DCtBuIyCCUg5auNGn/pRzJ5hd03DG/5YP1WNxgicI
o3ap9gNTJGDCzd+N9OWFlX75nwy2NU7fyshSqCx9+Ylwf8JHOXlol767ysKOPhwLqQK9KdG4ulhO
vKkUXtrTc9aEZmBjCxMMTeGkZNt1OhXJIHcsVjijpKplpUhSOdKVejIdRjGE+GSTlrA7a9TAgYTx
evjw1C9Lj1Tyi+gvZSD+3lqIN6IEH9kXnOdtoGGFEEGRIAii0v/qoa35Qw1NeJhoHkh+G7f/Du76
L2f3zTLae+sAhZ239McbRQzfbVZbavtA3fW0bQynLKSAL3jJ33wwqtWPObGglLq5ITbeNLkLhJVC
2igi2U2BHLYxyz/kAmC0goXDHj5SzTtMWSzpS+i6/WN4+wnYTONnyf3bbb+MF9f7VQkn3gOkMiAp
/0PJLTCygjxSVdifp2HU+r7gs2v9XBX3UvqEkyZuAmOswJiO+HJMRfKtLBw3u56fsVcbSxs2/cAf
gPqU13Q0aD/NpPGdppTSzT+c/iwvSxr+V31/TVAeoiVuvDZnzWZogoACsvgO+NH4bJMxhgClKMUB
MwXXdEbo3vGZxj9khDNuRJ5Xg7L3i0yEil05yACUBq8qyREZyScJqBpj82gm8Uj5844C4Tss7rQQ
ba6lv5EKVvX6FWRC6w/qYZZQLgGYxVQSrA/o1QwywzxYQ36KJRNNpNWm9uoZGQrPXX3Sg+Y4nG+K
D6yzI9/NcwIW2p1x22Xu4iqf39e/lVDGdm2lWH8jPiW1DJZg4s3N7DqXaCo5uWUJhKwEQADWxDkH
f60tCQxG47p2BjxIzSmrQBzjl2UUH5329shOfHSaMTkO+6JfpymMyf4lfNw8cXYaqPebgFQS9JGf
bboMqU69S1j8n2fZ5iXKepZuPkPLyOyNaZkynq5dq30o7GXwVxywhY8VF1duqIh6+iNpCriC7EPp
n8phx5m6vxmN3Zt1LiJzN72SSFUrYHrseN1HjgOlIT7B8ctDjAlQVO/eP/FPtn5g0E2z03Yq4BnR
G+bqGiaC9YHO5+2zUnw27g/S2u/jIf/M/sQ4Bxbr70kRPbUqpW0BVzSa5uzALBlUvzvfJIlqKNuB
NF8UdwDWUZXq6PyXJ2Lx+fY1cDXVAwH1fbavq/FdS6Nc8ViGn2y9ldeOLVCHDegVa2CVQEgG6kle
A6dkavtFvNj62yVR4/eDhK6V/i8cyAL0F7EF7FtBcofL8RUCFs1ARGQ9Xlk2KuInLd6teXc8QsRP
wou8jYYozwY8aqdgI/pJeWS6lwJAUAtGx4NvyBZaxOymMpYQxG6r2GiJaEnaHH3QmH0VExwfj1BN
aX/NUmDlwIm5+0F2NGMgMCVwMGnGNqIMFziLVB1ZKSaPr5YEd2yutF04ZyYJahCGssiQto3FvPf2
hfRiZTXl3Z+FGq7xSBaMbJ3GA7t2TwjJ6UKKEw13EXKfGpU1Y8ymlCRrsqr+X3bE34nMxnGSfPaV
UhtvgmqMeCY5AhpWusQPHozyDZdvRZCME3LTw0GgCLCq5+GzSLTf9NDntJiGRIc00hNn/NsqEFKU
WyPIC9KzbAVmqXUMT1WNUs2Vd30ieYnM7kcxjxZ5z7cteTuED5l6efhemv2/4qMHlUvTUj0zAmZO
N2Dsi02lAoK0FWnJdhXksLA5bhGgyOEKDk+vsEallxeBNttOFPcPwVhvaYyqSQki/cO5pd+amGsk
qPDt2RO5us6/8n7MruaLiFBKi67OA54kIUjnhfDltSjbBBQZR7fDOz5lJhB9qXk9n2sZ9VWGiKEO
BUYTwiLDzeNMbGzsbMKHbihdK4TxxeyjSFYalg9jGIOvXSKDT2Ae9SQJis19pKRgMeB52rbjL7ry
zrJ8bbPtxn/xXJN9Kc2xWBcaaB5ouAmSPHVHZ6Y5E3I5Iq5BwtanBCVHvqLyd5e5wcLRtICPxgae
+gdtrzT2k5yuCSU8lYICYo4gcjwfjDS5H8q74gX0SbxpBaOAy+xuYBKTdTbvln21nvajySsnr96Z
hyFWjrx5lD82d2WqMHsyb+Eu1HP3o7QWotPLzvmi5g4YoAEZVdJeJ4226fFzKYQKnjvfs0HdmLAV
zVBlPmCiTOF1C1fGmKVYvsCMDk5dGQJTx21zgKA6yR7ELCPva5Ma3WD29Pphrdc4+4hBFvGfZQKY
LoiE6tSlQrgH4niZOYqDO9W7JJ7DcBrYEg/weTvPTkbGMcCvJOeqfgk+8VrlNbYtBVRuU5q2YCHw
/hQdHSu8sQ+S+rGoug7T6mWaUIs1eFJQh5Wp0uzWPC61TZE3SArc4FV9LIh2J+TlcXZU8r7S6P20
RWQs+sHKogTdFJTsBOQnigywN+khXqx668nzl8o9krANNtILiVIbQMGL5ycPBJSLpwprxd0hcEBS
60c2aWkKr8C5H4duLN1V9YxftOAgOCMpQHgVIYwMfqAg6eIDTQcHX0yZu+GphU2lJevUzRxdpebB
ysUipMF1+4mgt1nI/2LyrvdIE54Es8YNJaTxB3+FY2145O4YOSUi7DtNGfTrttQIM/6yIuRirNrf
pZohJYJ+zF8jcJi8+YtRP4lEJDy0lfxLSRn4yJuY2sdRqxkA3WtacAjFiv2w6byufdP+8hOwkX+f
bMUtl5NoSH1AN9NaVN4dwFaSiZ2Y07mkdfFqH+StIfyx96Kt83w93rNhSFVl29r3QVjUH8dvs4sS
h9vJBeR+509hQZFHRLLrrI1YAPlf8o2cJFvfZnZlsaQbrwFOui16I5qFTxr97TUTbrtVCWn1Cumt
2EX9Geuby5WiG9LS28RRw9Q+NzrIZ/k3kCc1Eob5HEPesXUTj4pA5vBDpkrYQUGXYvL+mZLH7g95
50k5dagGTEy+zh64Oligqnj6GDeOLtISQWP/LpoVd/+Sdtz9R93dlKhX5xRvErMC+IOa6Nmoil+j
vaoEg2YRr1imMTZwoefajU6Hnh2kuRsYFWxwKQmdgVRTQZss3CXDp3OI2a3FcFsz1cww/ghP4evu
k0bM3HsmwF2SETrku6To42406PmfWwgvFRcNUyKMqcY0fdCBYGdoPjGkCvHyTnq4GUxSjHlrxdcK
3ufuEbiejigQ30dddV99pZrKP0sfCFarL/DKO3gkg9FCQpRDXOgVfPjkoX8ccgwXTQwZ6vBaxnIP
qr0Q0CbRDYyWXMZ0jXx5uO2MHy3k5qPuUDlWemuPdSRcI4U9BhthJLYzZ9I28/pU58O/+ZwH75LW
saqI7dBQBr8A0OxrDiQTbEyG9QQVQHL+U7TykoxlaZlTK0M6xmLTmlAtCJTxHlvrtAQyD7GL7gT7
ZUY5g2WVli59UFlDIydfbMR4Bkzb9KGnObbr/AYoR5GWEDw/rdESNu0fzBzyt6yWQM5DwYtV3UT4
zBX8AcWJMq13y2kM6g3sTUn3a8vvipNxEl1V9IcyQ9Yms1669TkNfG9YgjQOa5ynJDzExuSD/wXB
OQssBO0iQWD9eVs9MR0iNWWUqBIsWXD1BGbu+uDvECVMMICoBElHXCe336K6Db/Fx46JKTFniRTz
62fVLvyjglOU/iS1TPo06oQZNDaXkNwMLkmkB0yLHvrqYJihYp7VXJaYqBBe78AlLYZcMSmzFtAb
VWRDcp2WS9qT9QTHeYP1za2ZiN94Uu1ygj+9qBALjBe3TL2te5rCooW07DzByKcy/QRxsXzBsXul
9IF7iycuyw7kB/T62dMn4yA3aLUikhpqX/k8HfcGJV61m5etwjP5GW43rCBl2/xQf+4oDYX67/0b
TAxP8nYbiZGdk20SoMsCKq3I3IWLbd0rcDFaF3s29wkXFyt1HswaxBtW49grXQW7gYyU7B5TbtEB
Hyn7LOgmnDM88JNKtSXlIRd/f9fnY2LCols2y7knFj937aNNro9O1Nm3VldNm8SVZZhdu1cmkozu
MHx9FYx/bSxLBod1X42zVTdyAXeMce482REvzGYyqeeGo9o7rxCiYXOCdtFjMV6UUx5a6NrtvH6N
B3OrQHl5lpMdptFmXl7tJHRC2n3o6ZnJqpJuv2W9j4RyTZKovIwcGDhUN3FKFHu9SqtzjHpKLoK4
F+0+QijUMB0Uro8Iy5KwHtj8ULoqXptNY8L0MYxIqk1NAw4elUXWt+yLUuxXnWmq428Wc3UZ6kho
ZOWYSgwHksHncKfkdS/ynFhaZuk8AdkTLC3FL8j69a3Xd4KHcAGLo7jBa6jLxD/sJokcsMkGYw9Y
yDyECM/FHthV1RJnM1/P93cggg9ESHww/cNmS71DJQIqb4ViNvoaWx0taGU+5gK5BPlRQHS80Zz+
C5VD7uNler/sUey/h1zGkToSfPb44Foy76SSBjL1TtrhSAHl/ZLvzDxth1UZevBSvunLiKQeVEm5
dg6hTXdZBN7+ZANSkEWwgr+w2Tpx6/eyNlp7QTcyFuXoczzqo6bz34+K98rIDfjokm1r4Sd3uPQH
8Dl3H4g7sjquj2IVrROaUJ/+wigxXAAX3HXNmbadT2xUeaZAhEmYdbyZIXRfmcLl3ou0EAiXUhRX
uHn1E3l+SSHC1HuHyjKw5EOWXTOnbwN0AxCCP40DU1FChqs7aL2u3Rkj1XJvxy7DPIydOjIXF8hO
wRrOqgez7YUO0RUCx6JnchPTCwCtiJN/2O5E6QEYKAyzPErTYxV9d5qnxqqVj9N+9rnpv0uZO10G
b+XfvVbS+tpEHHdfnTe1npJkfNbAgDDN6aLk/xF9ACL4Dfvb9eGxwxEQLd3u9JxlZhGsqqfwCxNV
0LsIrNBXtwob3KIN/cfuCqjwUtnscq3qLn1yZtc2U22EqU3KfQUuvGefFVeDFO5epZjmL1TWjWtm
QH3nau6boGMEwQemAg5a5sgVAlnxwoTYpChzUkiQH95HX+CD8o2SBvDJAZoAaALqclXFthDFT/0E
9mx02oCpCHmFQ/8ICocRgfwJh13DmaiEVKlLYc+al7o1e3xJ4yBketW+pQoYrDqZF8f9VvuhpVk0
bl7tHcw5zI6CFlkt9ln6el9W7EG91j8r4lkwhL30f7rDWfhj74BB3WGsX9NK4ZaZz5RP1g2xH3iu
ACIqjcsNN51Zby8GUUMsRxV4hjwT4VTlUk0uuMLJV9BYKqE+Zp4lCctE3iI33zJZ/gCHAKDhE0ta
36cyxSEQjLc4D7SV48tWDtDOg2ZUkHH2N6ljaPKSNohSdjwSaXsknv5hhfLl3jqw53gFKO4SEv+J
B3J7kWh+NPBskVyd+Iso3tPSlSTVYmwIDbgHLziqKU3G30xb0hmJd2oZqtfchEf3/hlXwlumq4M2
uaZYIm6KQIxHGB/m/PcnpFizl37qVi17kdGnpdNGOy9pCQeIopFkCVItkLmTPLX4xmQEd/aETavA
pMsAZUIA0XU/ey2B/+iKvcQTD0/2Se75NZ1OM80oul1CWy0xO0o14SsFeiy/7uoQq2yP7MJb9MRf
H5bfNTIpM6peof1tuQkC8Y+6xOCj7J9vIZYvPvOAGul4Ru2mCSC8KFPRMKXaZSZRpOpd41a98OZ7
FpUCTnPAchgzyCvjzQ4gX0Atg1gkr7sHOdH5dK2dY1MTuGn0pxwqa6WrzzuTxXBaFd2/hYocJKPr
X3JcnlzrdW227pzXLJZcpppAXRPLB3HobhGtpuFb4LwHn0kISPRMZmyCE1yQ3gdV+9eTxHmLoyKw
b/6SeESs/YAH3Tk6N4Tb/sa8YU3xfu/4vM1P5MaMhp8C4gybQIx4AUHmuYRDYU3UrS4h6gSN1UPp
FvbR7PNMsER+fah9pi709cnIGJyG6qE/RB/l5q/tHV7G1v6qg2eqQ2gDbNnuKytERPMfRbQQIT2U
IykPO0zt3DInG3NNR1wiEdzdYNTlu6armtZVSXU7Cf4rzTTIvVWuCJGNyFCI+jP3tPCKWj55f9OQ
liMUn4gSWuuo/SjX5m+VYhBWOqXG0W2IaccVHEFGMayFu/o9/nNS4UToa7s5m/ssRBgzsUfgE+Qq
HWnAQYOrAXrWbaC2ipXK77BELVMaxhfswqS9mgm1OgkC3PBWg4RNtTB1Dv7glsjC5lFK/VmCHrd1
1N+eOJCiCWGl1RSoL/V5Y+y1BpI6wCKFWY7NycZgqEjdFu2CPpePVJlAHjj3IjLwcLOoc9Y3b8xp
XomfS6Hgf2IxwfATlJjcDF3CmN6AfektjSfZqNRmMmQ7rNk2vkk7wvYibW/BdU5FIYmeJGegRtMf
Cf5312KFr5kimuKdoWJGHY64FfxcxcKBhUV5dvEUjrxSVdu/A1Mu6vhHOBxzEbPNejvSkNFq/iBx
Dc5MhOwRDB3/6t27hwR53oFL1szf1gf7jN+vqVrpqexPponkS9Pv+ClfYmIoThLMqayurxrs/haT
pxcqVzPmTXBlD4dg56CTCMHmOp8+FKpaE6lfZjsgl3De73BbJ4TaOpcd/JMgXYzz85R4NIN6cO+n
BYem30JeYmBbtAqYYYplVn7dIWzqJZ57kpDt19ZMmx3FXefBij8FYLgBHtqwR3Zuiz90qsgEiMsj
4FgrWXP9/lMQwNrO+57C49K8gqmbqt5eJeQGSYFjyHuFvsYwF7wXyhfzQXzlab8/I0GHwpnOd0q2
GNUumCde8goYgWjbJ6UDG+Zp2GGcqKN1r5ZkPZllQIr2xym0dPZ4rRPIwNc4R88DbbD4G4sv8AQu
Ymp7ikkci+4FJLfxN8Na8Pl/NAxCTBLktnVAvkt6i/j5mbd+Zd+ZQ9AlxnGt0DIGWW7D/e6DAyFj
J7Vv5yV+nmyT5am9qWCAoivcAra44k3TSAhh7XwNNbytQ6J2JN5zE3xkYMJaLW1JwsRLdlz1Sbiz
sjGuRcw551lSrTpLoFakfT2VKRdIeIc/9UixkoXfr218S05CHvD6PcjT1wKkYkeMXbUSPsh2RUUG
snb9/CIZ07LHDYtWL5QAzyfiFltuHpdsQSwMzsA5VkrZtCqR8Nhg5/BTGJTQXgt2Wyj7ufmdGO+4
2qYrvre/kRmvejMh2pAKAcSLt8H6TlQnQuvsW9GDefbggea703hg7QrsfpHZpkJFv9rhFg0qiDCe
mJT8bVOnXwHtpWq4j/CJc32i+ujag7pA2Btm/1EGz04Y4HOIGHTLLjcTJrI4i5beZCbamTJEcpET
p45z0AXLd887JHyzjJHmoxMikYrXqI9hd8BcDK71XCYgX0juF3qi3j5Wm6jED0teDSEONHoGp50E
l/8FYarI8qyTp8V+eh96tZIKF8l+8yPgmtFYnFER69DAvaQYFMPkHxiiB30ovgRniloj3+47fni/
4wUhiCngzZTFXsqGaijFSv6fmmhp6cEuoIR5E5KkzO8WGTxD0S1CzavT+uIf2PZUVeSKAedhk+jC
B04+QYRQKt41NyzCvfG0sQSbtRz9MyTBlcIIvK9+kTaGTk1PKCSp1qKMk2szI399OtSeHCzdw2tp
SRtB5rWhQHBdHKA6oMUhzEJKje7dBgtA0rjZZ7J45J5rVeosytIEL+ch0HSFXJ12oX8YgZuUTFJI
DuLQwz5XiXhEQbcpz/6sMJhcTkN5YZFEE0q6yW6G4kpXXUfsOFtPCoTsX76jV8nKIVvjWR4vWAue
+0l16Pl+ukZy4XQ41gbr+8uYO3tCga9UCaqItasiyFiApkCW+5/UulBNNakoGOxm4bQc5QBJBHbi
5DnRYUl4b28TlkXVddfCqlDUdwrP5vyatiOyq5vChWZuaUfD6ddwH6sET1azsh3VbHE39WtvZNBF
nMkoyzNDZ7Np9LNaFlU+I5IPtxyesqkz14wcUuz3LEohN1EyszPy0sANhDBzWRIzGHwAekUQVpNi
fGp32dUbkQaETm5WpW7+nKEd/SSjEMljxBCOhmAQkoFVKhg/s8A4tcXcgO3ZWJeWT3dy5rnWYIOo
okCpYPz2oJJgAX+rTQrtWlVex2oZemYlcrAvtV+rF1NWzu5ks8j6klIwG5XEshHQfh0q3g2LLWLc
q3WrbrJA45ahAx0ai+L2JEXnvAsyL9VLXscL46un8SiC5EmooNS4jKqBsP3DwCjGRp1uTyPLTYLF
nL1B53tJ2ZhH6/rLW7PcWhKxyaNbVQwHtKaLPbRUVVnE62BNDZrkOhT3JlD2Ib4ftWEcqCQiL7u+
ozqIhr/f3s4rGBFOLszr6KGzXG+5zDq82rLtopVKlgCFB4iyP+rrRVtuQsaG6yGcGhNbB0n6S7eN
ZZAM8LedLwqq7BH1M4KJI8YHR8O9GAvOkILRFrG2F3AtWOGORZ9B4sKj+l7a09f4s6OuFoGvZi50
NMHxxxaUscUTphOJSGWcS7Hp5me+5C+cYon537lw4OHDxmtOZyZ4QgpohsQkxZNaVhr+AhBhpucM
VvmI6EUtfTtP1hmcnwPqbxa2zxq2qCjFQZWYJg62zX7pFt5ZPFuWxUfWkRjOMlLqDfiAa1l+9DBm
0YXnzwC70u0gYq7ncnW/Qr4+fbqsxjCY99Oxw1bPuTkVzuAisKhA1wZTV4bFRbs765rCjPFJUfYL
QKg8jdFX0gViM+p09vcoL+O8e/VW0wov1pXavW6BZAczJve6m0Qr0YdZyzlOpLMiIDS4NEaeQJKm
YUnJepkLamqDjcxIA+kYGvJU+R19ZHvlchXEvQI9rUDVTogcQCSUFtrRgw34q/E/kbeDRxlUlf8R
dRYNinDYk8v7/Kd/cEi5q0fuivqy4A4TODch5RL9A/rd4LtO0htZMsMi1eK1jiDgUM0ysIBR4hVA
8D1cbjpY2oxOXxb2wEC5y0i36HUmTAIoxwm+ODvf/DuPEiyGW4Aa6K9DjGZXWzeULOWiUxCaZQyk
pofWLTPusoAIs6EGzdxO1iL0NZhYXUhUutJUHSKDrjIdD66C6x8CvFhtzAImsCjWjlCemAV3EysB
5nhgGWHgH37vXfUjVsIzgtcd7CFVlCIjCgePM2fIQj6d5lcM1dehWooeyi0pb2+6FsTDbRLdTmvX
ZB0srpGcC3G+LiyYshML3c5BrQUeczmfeVu84JWlIen3NRD19XXWni3U56XtVPqKajeCumbJcZ98
ELZyeV7qnw9WKaTVJ499M2QuMQmV60DnEVb+dR1xtv6pJ1tXD3J4y8m6W4vR9p6GwNPND/86YSKj
3sY0JqbDrpj53RmQAbMn6TAcboK9r2DI3zfosm9UUCDns5DDhO+TEos/n6YDs3KPSWi8XUHROSD4
RUmoSSZpDsTOQDYWuyEvOY8cAOHcpWxnOHBkmXmXVSwhvbvUF/hH1UR7UvwAoYbgmqSRs7zNc3uy
m3bk/nFc49+SKmZjTFkUADrHvXmfHugMCU8iPD6FxabFQsf+v/WPrO1FGvqTgn0DP//LiVb6HtG2
GVlTK4wqdqIzFmVLIkYYAigZr5fa2GOl6gLDh39xiGxpIh5Oh5GOUUe1PKd8RLSC4Cx8kFwScc3h
ZhsvrYNb9cUgP+DWIT2wWKjZOuFQiyzA9T/9XL8vhCi83+vzkrSbl1JknIUAOp8dND4uWmgH1FnJ
nSPBORlFLbc91C7PlZFh7uJPbyImtvuojGTVBRIe8NpfGlT+0bhQv3Wx5Ek1YFo6hnAli5oq5o6j
kIMZzRuZ5tJPg8tB3uViMvka/TlKQVV3f60le44JrRAW8tfmNSx7XU6FyFhqxlWhyZym0Y7BJFYG
gBp0+pTuQy2Po7nnmH8oiDJGbMof6O4SDNX2uPP2xiS+wLUVQB/5+Pc2wqzk8r5qNFRc95Hi2rn+
JoyN5Ljl90e9fFbKyIwrBw4LbXlmR15mbtDtGOPu8vkW2NsWofR928n4nvPl9l6La402SWMw6bTO
VYr3vOkW7jKDKLuy6+qICMvkxHg8Hude5WU4/SfVNU/p3GSVMAeL3+7kwPiEkylTWAicucg8XH+S
lZmBgpn38I1RNTxNGSaoceJxG/cO2O0hPg2rGYyKsLBUsRoDxCAw3a6IJ5by3lqkdWPW6OKzp74+
Cj+4TmfekVW4Tvf6o7CID65hti1bylvCWrS+5fzB8A5k3YggNQFs1dDt2h2+0iAKx3czzYAaIWQo
ReL7T/cTPDcTs2nJgbamiyPedPAds9e3P8KFDmNo4ED3+ZszOPMXsghlkzbH/mOYG2k/kCTWHMQw
LGRGqa/UnIpbbLeIWNJcWkBy2ksYUOj7/BnVuap5D+4R0jh1RDfnsdA9xxN2beIgR/e4v4tUun1s
zIvN3NnfGge43i7PvxZxwkrqBMUkdRN8KJzmnyKPVlFgJtRSUJi7nnXyX+onwMYEoMnBUod0Y563
qdfDgFT0EN/8A54hIHKPdWnhI7/AwrFqAjhGP592JnEKOrjzLCm9ygzN9Q0Pd14QWhZGCgr0+O0B
2tCnPXS8ZMF46/hUol/+tJyaO7s5zj9EWBKwGFAUnHPo3FMGSM4pR/sDkwn6ht3ia3yejYXa0oH9
cMgmCiawAwRW0PJSlvEozFTO+OtDi6afpECwwOqrTD8Uanr/6PQui0hLSq1A0nU8we7rBZw+HQyo
gL+j9Q8WDEqheagB7WXg2D+CXox9w8vUVtpkVnw4fJPRLbvo8y7w98DcOdXBfhTwP3m713ehdud2
qhkzxla+E1M9MYPPP6fjFCuSNSH9/PoSyfoX5rRC1rtM7tlGYghBoDb3eR6TUZFUzyIlVC8bkA29
fC7MmwGtth/cvGi/QKtV3xPo9Mc5iUMLHpg31g3d9FFHEccjFhxrXsdXJD9FOhUxC5/XW/s6Jc87
aDJ1rlOPfF/M477sQse5OFYMPHZhrKRr9g3VySQaSLux79nUUORrDXSqruo86AGdD6WqSwZNgIqS
F17HROv2/Hzu7AIpb7HIpyPbH/htZTaWPbzw2J4mmDgrD5yJspAu/3mWM2M7WdtUtcT3Nefp9ez5
clSjLLM2NDfgJX5l4CRjT7OxiUyGBrXyCGm3RpQmai58JWV3uv6nTQVl0X9Nc0N9MYJvWKOZHzUN
+8ejYDkHJJOtzh8YLCkeP45Urp8yXvt70Tdxvbr80DKoT2V5z/vBnjrM47RcbK53j02IzgyLOgcG
DnPRbGMyVSISp0u0XyHaPYQ++FrXsV8hZhTvyz1DQ2L/nbBiSol28Qviyndk9lxj7DPU6iWAXE99
mOjrVaqHXRpGsfp6L224yJ78xp6OeDLltTsg/0NGOxuAcAkWpzFSTsTv6j2kS6t7ZUPWuZfjyO6Q
9c1ALXjj0Pj/uPiZQNOH76fHBXfhngJOjKv9LuKwttuMCUhX4B3N+QIEVv4KDeWXgMAThB5tqrxS
eVvwKxvyo16g/juO/KyQHn2kne4tb0Uf0GBlVrYfL+e9eZD1zgcT+tuidIeqs8CgTgC8EgTcAh+O
zEKHRNh6lWngV+3qeo7wUMCfEmXsDwKOIa5yQlrTszIrfcALKAQy+iG2YIJww9XET9aEj5iJLL4/
rmxKOLlLSdv31yZDbp3hzDmPbTfOsAySUWpTDohLkgRK3oyEjl/yfOBrLvx59nGl+qvwpbtg6wfY
lvlkWlJbOJBbye/P9cR1HKCmfk7D1KEi/nIHUelgpmudsJHUlGowWXWEj8LcCTD8K/NfpF3VlVHh
epWdk8D5Cjll63IX87LZG7Fk44/XE6tSpqlKlHLTMm78e1CwkaLVgYIjRFd+JSRrOX9epC2rKj8b
1LuW1YXptxJtuy2B2c73QM0zXlAfmYc65CzKIqlBB5BDAhXKPe09uYDLhkdMuKmWT/B+qaTVbGAG
x5OnmycbsdIE+bKsvUh9nHz+GHbx0Gv4tAGQxXFy5SzO3lDmXyit1GTc7PastgDEjAIlTULBZht9
KcFzd4BUr7ymhEMcbkkr69ciJjvpGzlK1LyWfWGb1OFRZDxgun4tuPYfxSMNs6EtrSVLjJQmKfPA
b8DBO/PBQDUS12E3cOqpUfwSzFnBZsKpUWgFCAQiSb5GScYZOjMXycMeUrmYixP8vEcm4mkJ+bH/
7twaNWTS8JG7dtwJ+NQh8dH0lqBTSpGcCorcGGFf8ilKoxLRQ7HPLDEwlUGR1q5Z8shy4jp12/NO
vNdwVSYTpopuTX8/TPiYkL2VQrIziMT6Rur7vNCA7QGe/7KhyCPiUcyY1uipGUeYX2iTCTcpfb6T
pPMiwPrtM3J8MMokiAxka/PsYcYSJ1eodWsfjeLZpeba57SHUA9kPVuYdQr5lzYfUYDx7bA3supk
oUyR5hp1i9fp3VkdNqFbPLcxeFI9At5QmYa3i9PPjmUOK3zkxNsZZBISStI5dO3dwh3kY97Pzxao
B9YGH8diJJqZyuxAnQanh/hqYGOnPLOevX0ViLhzO4IuabYEuajoGIEvj9EY5rsRVneijhkprf6g
3QkQGtcbymwR5DjgNGQuq5/whWhMz+s3SAbjEarMNTGxLNYt0THz/4cSNKoApD0z3mv57rzZ67pb
efxJP9xg7NAJz8+C8NRRCtGbAnm1YFtwztS61nEK/6C40hz9A2JiM5uoib7s4g4A46dCRXuYDWFD
bHw+Ehd3zkr2Ba5eskyaeDRgd8azj25zX9qNs5MEpQmYcRgk3eWNnqonoHUrl1lKvUA4RdoimOeG
7BxSYYfWbo9eig7ltktpS5ZbQJA9o5mbe3bSecXSryragkapUxH7mhHpNexL+zKpSRjDDikhVgtf
rxnvbe2aJ3bdMFd5Sp+5XDSo4eBihuyOfSA/Ex/ideEercN4Sk3lkpRAAf4/lUb1Nxy/kQT0yqeT
BlIDO8I8IPOfO6yW5KNoFqq8zM45PpXLcUUJE33pLaUADr7kGLwtoRQKYqh+6SOrhuS6kt4IpgcK
rDO4xqLMwiVKMLs4A3t9X6CwKrqHTH/oIs4U/HjBVPVhg2SFyiYfUCpvl0oo/KeEzzE0Nwa1O0kk
5y9VT+JWGDekrFN/5HVTMPgF7lsmED505Cerk2Qvlx8sTUvVu/BzGdwRjP/HKpg/ibKVVhnbjBO1
hS140Z7Tk+v5FXnhCY1zvPi1nwe6/Q+jaeD2T+eJKrXmo2jM9M5LOmifrXqn0FY7wsqt06QhugHc
a/XdZ4LZXPf2+WvydRt9Dl5GAqYjeK+PmNTeLND1KAlWAIUYgCIDSi1a3uFjKkGhMchbtcbFbooE
uZ3PgPq4xwpmRHm6H3H8ASamumvX3OUsXnxU9Z02JxN05zER/zu7gdhP46fNyC1FsgjUY1oLXER4
RfGeTNEIkdW1pzrFQMIpbBS+nUju9WiWxXygwSnUhMtnX6zzeNzJRJRv9Uu0nFphBQBjXdMlatfr
gmge4siDZrwyy61DvaLLkjxWGUN5NFRnX/IM5PMlKqVxuB8AWu+UwUu+R0eLhtnouB2s9Fso01Y+
76xQotrSCOlypMd/gwiwK8Qg5b1LHLo4wjUjN6qKW1sfpMvfL+77/4PoF1xuVMBnyIYQgYxW7tfd
4iCK6mApJkthjOtx7IsXYQzzFDgHTJ2MQRKVAmHLHq5jj0550H+4L3K+GEZTcSDet3r3Yc0QvKGJ
bX8KgfEh+zo5PctPszUXwEaJX/9cBRO/9Jg7xiJ0y/YqrsttvKdEmfnErgSikpd4CeUPTD5wr1/J
YfJHihSyvduTQb749s3M5fudSQKPbpxA07vMQB59barMyLI9k5OtSiu32tNKviNG3Cg/T+EFF0LW
9IjZb8YL0kQAu36kQJ98158+yzsPCDCWm9L/6wjMOuMM3+4llq1pG12ZXOP+Yv+/WiZH3UQcJxKm
32YKoL//W7PIyaHVuv9VNGcVVuV8cl9GCOg3aK/F2A2ikKKZX8D6rtnBsvhHAqDGXC7axC2M9ph7
xtR+BA6wG2RgwF/DY8KeUl1rZjJVgU9o8ory4fp9L37H47byQiqx1iov6Se7JYNC7fJEnmvGANiK
3XcQWmKSc7sTbRxewfIHzk1v4QLGPZ0UMrK6skPETa56XEVLhz8dsCf7KXCYJVyV9w1mdAm4e/eb
hzyg2ZVWpl5Odkdf8m8laXXhLbiGomY9pMzOickUMgf6TaNpOlXK1Ke+kgiBxXP/xs8rkgQwa7nc
0He90PvZzViD/MMoRvW6onvpfg4CZ8yHdoTKVWup77CesmMTttUCcI26DQ+YDvQ15riP6Dz5j/H+
xBoK40N1Oez8fZ+HIIoh+BFtLNz1YYsIuV1Lb5SiZvfJGxVBNIMieodUA/aJG0/UbdXudD9nsm2r
am3fFom1n8zDGPAGN18zduloNuXSHYdl0q3jGHjy9DbgqJjPtSDAzFdyeJC+NEUTgyrtw8VlxWdt
FvEQPlUee612wJ+NwKioVMhBZ8Iax8bTZMUGQeGcDAkErTurdvAAg7kArUdPEUiZpvo7aZR6Fb3J
FfIDpsKm2m8FjLCYea+FKSZRNS7PnP+vPBxnYr0Tr/J1xrVxSGfFXlIy8RUg26v16AYB/Dlp6bsi
DqlTwL+GMPbcelj6hUdK4gr4lkKIbusdbiDYR/7XUJAJmGIiRdx/qU6YMv3iidS3V3H7RPYmifbL
SltH+xZicOAflbMz+unuExrZkOotoKGlHI2322YJ0YM/NmF4hR8y3Mjby/RLu13yyuue3wEh2v9J
ljiLPbfsXpSRZ5RVIv4pK7BKeUYNKmlcg/fvJ87zpddZgcruycTxp5eY05gZFf1KUiZHSePRTUyc
JgbbcJuAwLw/gkeZxfANkgERc2q3TW4/oF8tl4ZigCnm4yrXYXhNsQkwQhlb4nLGc3gkgq8YNbv1
iP6PoStWi53FLhPe1jUMM4Q3oznkBtsyY5u9Nr+c6HBergP/5nJmXAb06xgQ8wBhg+w6JaEs8bhI
z4kEXrEkXvwiN+drpQGePR1Ec2GBuT0XofA7SFZsYqvqfvcfT0RJ+dU8/i6TTmvPw310S3k7phWd
dKrlC/fLjl4vUiuXHOk5v3FT+3Z6b/MJHQUYOxVx+6CQ6F6Mn77/Ga4XwU19fct2nxDj6WBJHBrk
R3G4ByXbVPDXHVXnFFPeOua1OWj21wh1ZasfNcPPk2GMXtdQl5BtVdgCwFduIDthRftd6NyvmObU
ls7TExgT5w+kOvOdyfv4zUvScw359BnRTfUjiAhCal60xGRVF82yMRu+S1gsMWLjkBM2VPQ9+Uqz
la2jNonbqj7IIFdhjiEX3nYDSghWSa/RJFBCfoPA/533GJIbufeoOi0kEPOPTkFtZY6wVCuz+79P
ThnuMXo5CveWZRDrv84WHxHlclDy76kDtgKLGAx+LUhAVhHozPPi9G7Kc4JOINJPf3VkNtB2Zehs
bdY+jOYVu6mWZ8dHsb+lOwLFrn/N9k9yewnwwsMyqMbha++iD+7Pm84vp/ZbyqUUyLw+GebHYpW5
dG2fwFT57utcUMTzTz7lhiKFypk3QIgmIGFT13TvJkgdzTaFevTJsxa+1mEt3sGvtI0E2jD1cGaR
/vixjw5wNs+OBTkquz8LpfhHKWyHKn5Mli39IAeaBvr+jyY87QSQ2We7+UwWfBwZgrYD1oZXVuB0
VVxtF+kmbPo4JIBQvgjM6NuTtDRxJvnSah1Y/TUgzmzcQoKfFbmcPmbJVlDbYu1Rb0nBB8+jNzW3
t5TtGNuwt4amUdO5xHBa2lzOncUAejHT5T/OdT2DS5ufcn0VrU0VaZm8B0nUIuokQ+WbnRBhtCip
tZ5JGo5g+kx9pFyuknAFcZrnvmU57HTYGp5bMRWCXqgDyBwN29hS8YVK+AJ5kDndJ9/s62k2GIic
XrVnjgE336xFZQj/071MWTCDDNK78swqnG0s7SxIbdNdJ6h65ao6LiLJ/Crf1/e3Eyf0If8fQWY+
Yj2nCt5A6aKOipZybN1aVqlfO8gxHCZBKQGOq411WUzgWhFTLiPeGa0MzIpyZS8YlDQmLDRo9Zw1
nanpWwBh6merKxduj65LM4rcVu2KYhp1Kpt5+dw82YZR5btEyG30mpWAcWpVMzI0p7VJ5PI9dPkn
w+bTtESOWdG6hM1XWf9BPOV8tFPlaA/QCt6wEiuYF+X36oJPJ413guFX6MOvk4JLJOuDAZ+HbKyu
r1xCibJ1ZBC8y+reyG127zWc+AiFz7DUgQViLdKjqQQrxW5DkDabHRaemZoXTMtTTs3Sy+bh1VE8
DTqGxIDx1yZJ++5/YHXzK/9q15IUwkEPw25mIXlrBlsdkdZ20qxSugUe94S3zC+JsU7pAVnKNQ0k
XLcbbP/UyXK7M1kwHyvj3MVuY/pS11gxgjVCZdAU9IkXPd2OEcm0j52kO8472sDofz/GKceXKiJG
zOyixEbSLCNuyGNs72OO3KyYbvAzd5FsCG2cqSGpMFxpG1L2bhhqY/asTCe6jtvVvUUvHRublIuM
qxd3D7lIE4RV+nD18+CHOdRScdXKFrOIY1sijGK3v0GDDGQ4zOmYJBZL9TIFFCStVvi8ghKZm6rQ
kcTXR5kKB8PV+HfrrtvbepjXHHegH7sjdTUBcs7/EyiGa525xdmoCbEscTQd2C8KLNYAb8tZn9tT
+WfuQwxraur5UqORlCNlFfL3PG3wb5k3HgOpwS51W4ni53zV7Fo5wx8t9be5tNPnxQq/UkVvm/RP
zoefYcUkFV8MbROw2yoYU06PLPNjwcwWkafi5cED37NFm3swieGThcFqExzBa8eE4Nr9Ym0bj/4T
vSjv0RlA5MXAZwh5GvoWhWMZp92TqmQXjv+klktxoYWHKchc+T63fzlx7boM8i7tYHjdKEvrYed5
3Eqp+hNHgo03/iYSyrxtDRtykAJ9CJh3FP/nb2orWM1sbjK1Fh3phlCPwAK05wDFJJFR0VUi/6Bc
Vd64vG3ImxrMjbFQN0SOI9TxitpUa/xKGmF9JdCfbKnZ5UqxhyYeyHswe05t+bxlJHOXRoYjMXKj
HOWVHyJaNteFWWwiJ2WToM7MvgyOLpj9orpSLNPI/ByN1OC5mIgD4G23m0d4Z2AAe4nF002KkWxE
nXmdUvnrWvPXP7XWQROCYFDUb/dMaMeQT9BiCIFY8I4Sv2WC1QDy66tdEPubEGcXZWQAAfMs5473
AC+MaKXpNRz4FcYoqk1mvDtxBM0TwapAoCgST0IbsUndj7VlZsHXAsMzUx74cTkSoKZtslnIlH8g
yHznYxJBnrL4cu7BAFPk0lvExKK5CswV1+/Kpkf7UaVZsp2Wl4269WnoWQ3OtSyAQdQUvis2uC+x
UQjPTonaZ12xQh6y5ijtN6cSfTUZRbvBjKG4zOJ2j9QN9Z2y7LE5w1LSFSevjr3z7MeCkAlqmY2L
Q/T4KKFlsE2iU1hLkhhtwkls3gGEqLRyZSPAB8XvJRgVTMKsaYyMnglZdb6p+ImvvVp5MyipJca1
m8s7cuJxFVEz2aaiLYLmF9phpx2NhGyGssLrDRr25bOJBJixHcaeAyzUKWfnLLMaFDOLLh4TMsjx
7cpFL8xaRon4KP8FYpRj3LF6pkTXlm0T0dCTJtJbIZfCTQPbju8F97ThvtmCsnSHoA4qKB76M969
aoc+ME3aNWEb7zbAR7s14VugbXHFdGx7vcFIkGCxZ2DzN7CDb5c47e0oUWIyzrpZ0J7p1/053ml7
owE+u16cnNQkhfl5XUVVxIeOTkdAIJH2J0nBzk8MtR/XKgetHZJd3hsUexjNBK6QgXkO4Q6jakD4
Nhi8up527kdNCB4D2g2Xak19XkvOoU8q0PfKyy3cMX3WTb9pEwYlSwc1OaxmwLW0Ir5LZLor++XG
aooSGlkXzu+lCEeVlpepF5P5RjoPCvU/MfUoLQRDXDhXYJp+T9gm8ZH6LdDP9S9nC1m28iUoHcOa
qd7A1GZ7QBqS0mcT1n85Nfj5YqTtVGSksprLru4vmKzWhvDrPX8XJ3rHS/mJ6SnVKF5zVBApQXP8
+LavjiGzpjMy3VMAY0BladjrP0IlqlrJtVgT4LMMYEx8Fu8+Q+UDZTKgpVwvpWKWsP6Dboc5ZFqH
i2c2vCKQkWQa2rYSXipc0PDjB+3TuUC37gqX4YjqysklEan91NvTjdN+T1Puujhy6odl5Ck8MLR1
rENX1hP7w1TtZsl6bPROmZFbaSQ6tfAWAvGQt1usbgGStowdIweSZD+qWQy1OmSIVVeMYpFVqDyL
sFG2sAYRTx0sj7mw/asGOooCLqw+73ZrDjPyyFPAFHbPd8vlxehRmjsTGB740hFyI0Ra7VqDC1kv
tCisyyanKLlq0EpVHTUAa+JVruZz1WemAKd52oVdDIymJ6lZYKgmNasd8MfDSQUIBDeVhtJB/6r9
nMMewLnlt3crGub3d0QwMQyiZ6UzZizJPR6TchLtmcXkXyP+aD8jTdoQc2ZBUV7iakVoBm/+Krr1
ByKwgeSObAS9khZ0Hh6nMKdXfb/+skTdA5qEqtBrjnvg9X45uS+pDnHOji9n4wWTJp8952RcIkz3
AvGqOR89DOeZcffJrKaGOlf1D9fS6HJqw0fa8vz1PZup8xTXTnIQO4Ils0932LIL0WciIAl84v2V
fYWmCLpUXy1K/w/7kAsSzRbs9mlPyYL2LLQFRsToSVSKFW6xQe1NYGO4ZuDnEgr8Ms/p700U0q4X
kihFlzbnsuIg62izUw4eVBNKOjMxsZCTBjNdg8leYOz7YQ0uO2XHgvPKa7FPvmqT+6PHIDjLLDPz
u5ml+8319rGlWvPDquK7ZHkST9nP5aFblVdrRuFfxsHHqbd9lJkwRFcXr/a4+mHJ1puShumIPofZ
mRxS2WZsNz4lwJ3HH1AVB2QY3AZB7cvYLaDUP9MOdyOp4Qi4AdFi8Y4bPAP8cO3HOEJhDB7sDbJ9
IVu2BSX3GDVr/EQLk/IL/dGAKLduZ2TgcPyGtE6AeXzt4nE6eArS6s4eQQxDwm59BpfuNpdMhrxZ
Inv64siGdgNqdRhCbpngR9GjePKF2HAl8K1F9GGuSnnVPkwjiFynBelpgRcOqqzPc8ajoMhRmuYf
rjijF5NwWcnQ/tAXhdU9YmPyIcl9M71omiQApTx5OstnC594WD4hMjOZiXE1RXwCTEv5rbyimGvS
VBMPwvfNTadJrwPJaOEomHiixyYepGwxoZIye/ja3L6UmVb2u+jAaEGhyK9Mf3QlyN9CzFXF/JCi
+L4IsvLrtjgPGSS6vRf7dDspw+TKJ7WXhZZjnqU5WjMl8DrjMOco2APedmvM1L592SIBAmZxwbek
9tzH9iVka5sBVBD87U1Uy5aYreAVWU3Z3fv9PFmQhpPk1TBhCNMHoYcEZVmBA99mxVI0FJJ4q0uT
FmbC7QX1sQSRnMaz1Bt82WlJzzPHdSIAncK/Aq/jQGU7MpctwKoOcg0dNX5YDM/91+YNKxyxy5u9
fJ52mebhxk5pFIerlh323z8x8GWwFOB4i5fY4U/kMjG1Iot9HBrgiAUq3IFF2FvW1Q2zRtiXOdZM
PkfJ0jfE2CPJdOyPo28mQ3R8/+D3VDay66G3UhpDDWGb9C+nuc1BmkmL6YlzJRz7vaSmHU0aosDi
L2CGPJl/hu90XZLsZWaA7Po4mef/kN+jHWe8ZI8YilYgkhwFx7gzCX8d+RLo/C9Uc7bgNbE+I3Tj
tRmBYAPPlorvm3BKYpqDwF7YoiDBn8/UDgsSj+S9tpGDixhvZi9rIxqZbA1grV9SDrCAj4xEE15S
aEjTiJyw+BTsalddM5mLN6jLQIILJR0WkC6fVF7LG8TgNkRE2cjyZ8F2eZDreKuHr5HyvZNIKOMB
hvgPwULOabpty594fZdPUYKRdRMvDFlrPypc5F2bbMo8C20HJOQC4V00wcKOB5naluNjGpHGnogE
svlRZbV/jkqskVXII9yQ2yLyDMIWeijpIoaDHF1hnE0oRuVEh/dJNehZLlDOIHfgxcMP71XiLDXS
m7y2RXIrYEIhNfbnNDHXciVoNBgS93RBzWGGh9vI5J2kUjHOSDZSRJVwgSvydvGIjP4P+60+CsJc
It6iKr4QYKrw/BWIhu5/HtGTEEkvkupICMaVn7qH0Oz7NSw6QtSfTJyV0Hz+j2Z6U/e2plXJ4XXZ
YUve2+te3cYka5J9yFQ8wt6H095j0ubiHxITTNkrp5lFWYgrzUwyt9ULFcEL2DDiqXorZESrUccG
Mw4KcSk435P7yX2a24mQd++4NLnZUzF4Qmk0dJwf1Eu01CSyUc1oa9xlMk2zuTuMAp+WkXlrx1WP
QeCL5KKjSbuu59wzT053yn5Txh7eZbrS+jtfkumlors7DRvVLyZfmTuqAxknQTgBNg1D7M1UkUDN
qWGmW+K/hC6bDHgWpeylkXKtf1eC7w11TLZe676NUf6raM50EtBvIasCpa5eQBxVJL9EHBWaoL20
i0NusEK44IofW/+m5WeanyBchT/J97KhvYWP0RBAk2a+vjleyqclPDBOCdMQNvNfp2gTKzwyNTmq
h4XGrdD5uwzMEkY90d7sHGHFSMphf/Ktb6T1uVHAXHkojaYE9kSS+8kYWCYmGClM8stnBKlP+7yX
GqSWyr+6snoo2TnRc4a6XLBD+CzIJ70BdBQIsW9PS2J9tROf8NNF9dZ1zkcHq/2YB6EmvEIsRp+e
imQ3BtwkPeyhqZtkBFMTg/Ul0RuLb4Ysu55/fwvq1c5N4WoQVzvzIWTT3KsKZa+gT5djl5snbwCQ
CFG06zKrsZhuqh1KPbIUMt71yGPA3W3TPI0Oh7Rtei/Ps5IoblaNplYgwhqNNVKbVi8BJZeqL9H8
74R8StYe28yFheHxh3QC7bIuq+9ulQM7U5ppjd6n0esqLGjsqtPCtJDn6o7cBvM2LizXA0irB4dm
QyVyRR+CFzldJjTQ8E5NEBbYYSo/NRsVH0ddP6cmlPAL2cz8xRLp7bilqusdaLumJW6FaEN0HaSv
yzrK4SJyjCci3eFzFduXJHID8D8++mpC4W14GEuI9JTmWpjscwhYhA5dO1jNEwFRKzqoJXtrVc7Q
/flo58gsmiyWk4+MaEJ8ubjwUOYIVPnJ6/mlqmL2dkjxLv7JjvxOMLeVtmKa+JUeNUKIJ+K8AbZs
s2eTnrI8DTqXE3Lav1BErz/vkEehQcfTfYKqqgcUl1PGi8m9H///edZqAoJuH6kA8RaavofxfuKC
Ewg6ChSePML6a2keUQJolsudRcVeT8CikMzqgQuqxzQfwtONtbxJMP6w6OL6M37yKXG/+siTuQh6
+YwwgSpZOB7IVhHDeY646lNQndrXb9BK9IXKhZGxeXOLgckSnDUdp9s6X3AGWIaOJHqwX1S8fi8B
yq2opJ2RvAZ/r1VD86WAi5yZmCN3PAIvAXYRDLcVzBkVK4BwFrenx8CNvWJlzxDTqby4z2fnCXrA
AS9YSNKFV/MdQOpPKuJY+knLZR0qF1rau1RMmjb+Lj2OrXI9FMv6S4OpVJxbIscYgscoSiXyheYV
ii6UB3eeAY5EGCojF+34Kb3DbsAFTUt+mUtylW41hCITDwSvgois/tPCP/qh4WkpfZ+wkqfA5gY9
V2VzQs1v6BuZIWXX+XqNXpl8kXp1JpYHpcQASzrlE8HEyHQvtFJI58S/QN0CJ9eLj5d97bpA+KiI
8q6YMQy4eXl3SFw+eDAruzd3HzEDcfoA+Dvzo/AoQ6VDOTpHKdDoxYo7797tY1pTBn3VRcnKBoai
W1g2XJNL4QXxuEMmIOj6pI2QmuHSEYU8gqirWILSmx1oA8Lp2U7JYNj9HlCwDGCmCyyWA4aYwKVq
LQWxJUJCtKQ/B1aZu/Ogsmsmde4yC4zONQjMLVRO66Ex1ClYnvJqKpvWDkIy66X5tBHcNWDY9N0s
FEp4bk2UzzZmxzv5txPKT13FQTz7a+/3gY4hPEvsqXsPH/o07YDUqdTnj9TDvCDfx6r6delv6tQ2
G7ny15D5Zzh3s8IJgOptHv2YA09VdVN3Lsfs6dbMMxpG+UQPQHqWULnBa63jbJcSIN1i0GOC0VFX
pqiHtKVgrP7wnkuvJj3gWwbIoQ3gRGDGRFGAhstsqBP04paogdQNNDd3ACdWFyDOB41Xlkd+S497
17I2vj5pUggEWAUIkEwtWb5BTRvFeBFKRvITHWSOF225VPUAN4f3FjMD6m15o02Ww7vKgi4jF3zP
J5Jk/HdSqGCy4lBOR1z3z2MQMGqz/yRogNTDVp57/RTOT7aXyv1cu4862NUqMXKGP91aKcNJIxra
ttZaiQqaxypriyw35sbYzAWqeoce7bcEnAZtK71LFWNQwi9rHMlytCkDjE9zmjzGCRApOMH0nFm0
Q0Jt5hvOcToLad6U8PzSjUwwGHU22CO8FXzCc6TNxByOAzGFrRgoEGpgFvPd4U5SWEGucERpkraS
tEMhwplKPTvB30+icwo+2UDTD7rif2UoDFr2UySrK41uRdXLcXEql7UF1gHj5AZ1fy+tEsfscWbM
n+JlXSijRn1w7us1fTGYQiwyb8/YA2Kmaj3M8hqwlei0NeoSI5z5IEuDGnGZxj57CCD1PsNeN+2k
yXo22pL4krp6Qe6Nlvo+/D5TnfXurxBnHBxzZPdozeLvsR1GfdtLwFVlVYKUCUqfWlNhhRtQJUV0
xA+8LLSQs+WNAULOwkR4pEyOWkgx3FO2ARLjJCQMPJM0zV3ChJXK0nse4zpXAqG+U0GOobZivgqJ
wOP1rYpUaFegMtUBYX+UXKU/qZEKVzsObUHS5kW7vhje9JQKDt1/VfQcgHGNXkwl53gPkwwD/Z/P
HTIeYYbNIl0NSouBqqRC4hHzzpgTc2bt9ghnnCwX6C3ntictPGc2SoJ0UZkfpA0aO1pIsG6YnMrt
4dDox3wcV7khqwZ1UrMmK9DAir98WssYrnizsVDhI+BkV43eKhbrZs8NT+0op/ANXh6/bPRNz9wm
bZnCj4YOEbtIK8cO6NJvRbE7hShGOZAl9QUpjVyzY8P23Q7WFfckrvOhgpPhv3GncOC5lEyFWv2U
pVVjZ3+rbLeehSa2UEnBJjr5174BYAYvYFJzkORUEOjt+m2sePDe4wKpLmZbhj7AgBaCB44wMrNH
8Szbd0bFGufoTaX2UxzkqkPNStddOlQB/OUbPU1mUL7m97gvAuacQ+veox0lcjx6zuy/Lx67rKOp
Qw5RaIhaiyMTXoFDCqL7+Zo/nMwe19vxq7gBndfkZTDNGB5afQQ9ePG9VEjF6AVaJa64fXkSihct
Ej75Imo63t5bMH6g2Gyf3Ka/rC+x/aE03f6B3iu6xZ3PbUngr8rqUJ7ZsnHjR7zAcyJBG2rnboJS
ku9D0r9izZ1LzLyQJu1uZC/Y63DH5yst2GB1uQzYotm3r+gJ7qwkqafUL2XYmQcmIQzLMaF/2tYZ
IVdD35IrgiLgZZWqcHe5HD3ml0bQ9kzmNYiK2Yse6PElvNFTqVBlLG4bnkjMbOdLDb33+zO8pLVG
7FBNlvIG2DUgPthCGb2yM6Og19YmqS+VeVmrfXey6n72Rh1DxtS/JM/7I9CE65jfPdGAT+RUzhxd
LXmMyEtK6HxoUzg/+q14N+nHhk8OFP9TCqGHL7IDJIPUoUmrxgNA20qxb32vNPkrlfNR6dWcQAdY
2RsOsZyDp7OYRBniUthaX/Lc8ILHuZOCRytGlvU9r5trIWE4WqstsCBsPubhn/yRptV5hSKc4SZd
EWYQDV8BTtjrOKLRTanwvy+KpyPKTVBu5NQJtsrUG25KheH1UrlzYAQ809jhazvSbWlL1MsS1ynt
YVS+2bXv/bEtZJPOmu5p2Sl24gZSFgsOn1uRrL2UZgW/vvEISgYYAskJfG1tzsYyz1PXA/M7eQuT
7rHUYQ1Lq83u6L6PT9ec5XaeljGcqQz+eecJrTTNOcJrpW7Mv2Rw5KbC2vs/+ht3eBuFDjQ/LtPn
AvDS/2EolkB0Ho7tOmSf/pNrIZ8gQ+zWP5SvpkHjpP81ZmWw2tABFDG7JVsYkIbY28divy6kp8Pe
ocoZ8/EAph7HdQVteEU3i1q/HjxrRcZwjEnPJBrgw4y6OGHcPlmxNxvc8kOy+cM9V6De7HMXaIxW
isKlvDpo0TUrKxeEPgUNlBEwPsABfaGuuARq4wUj2UEuiHxL+sMryJkCa0R8dBUj1jiG8tEcY7Np
okRTsOAUsc4y5iXA+pWwWVTC+IBmc4f015cIJmpBz8+b5GgUHwnBOpRJXA3AVX7Rr7PHykwZiSLw
5B57JseHBUyJ1bS/uiKUbk5/e1zsI+RI8njQhYRTV2Ha38f7qHwN9syc+1+IKaFZbxGznsCGzzE2
s9WxeJJP2WGZW/d7ArP42HFRulHdPVRNuCQsEe5B+l4fKdPUwYIub5UTJ31ZEI3atvAzo3OljgU7
XHkdDgzHo033Orj/nQFqULJnN4VcZpnjcMkLh50apMUjoILxyvbuBD6343ROz41+HOUhqv39k1Y8
FJS7QaW8l5gn0H8fFY23WKxevvNZfJO2aa8iNBXI2makmAESpQ0OkRGCpvndLbxXeQGTay1aERie
1u0JqUM16kmWPYLDh+FuEcAKT0VUWT7QrSmmeABxjGd5Ev9Lk7KxC+LPbalVxOtYCNeCPph4G9iO
7TL5zpQwVXQau7dp6XVsMx1EuElYpKU7ASwcMyZSfxl0oqXEPv5q4ghdPAWtkdErRd3zJpGiWvbF
KWxAtL2iNNculyyaM3XItiPvDpWamtnEI0mBL4SzlJuOXFA+Le9B2ygOTqM8Vy8f2TjuuTeQ/wNe
Ko9s7EnRiMhPrMQl0yk/wOdusjgo1g7BTyMCLJMrXmHGcsuh4aZEC0OSQqxDdQAAO+It9u7CNokX
XB+f3oy44JXLFENRQHvYqamSUMl3i8FLK4jfVXyQ3WiPqxTvQDPl5p3zDatJc/Ff45Cw5QlQkoBo
lWv3N3mdUg20YNHgvjGOIwVF6KnSwI8Fjyi/8i1871cPPLiHGlIQhCncA9eMdQpdjFRBk9cq2ttr
DpJStblEOSCKQFOjmfp21nYj9MAESfZjji+dEEEWUpbZQ4xJxtK3LxoHYaQ9W327spk0uWQxM7We
BfGOM1Vo1zGDksmm74x7wE7/fzTP3Lk3uXH7i55y+16aDXNw/EM6CtYRwZ8TS2GmcjAa9ytZclIg
rdf9m04btgNyWSzK7XwcwD97kE8VYSFGVsZ/OPlaT8n7T5eHzrpxDrIzbwu5Ndr81xDcm+rheRc6
WXBEkDwH1PkqBPRtlNUve3REoElmyCXii2+i/e9masF2yX7cFapFl8BrH6SyCHa4Z8JhtWEI3cNB
DmD5PIork8DAaLwDssXpdKGZ7zfsAKjoD+SQWFUuFUhGByOjmWonZtEMpRD4z1A6heSk+/IFGXrK
7cTrLCNe/uFDtTNMBN8Aqtq53D5S89GZrZ6A9mL/NikSgoon7CKzzaEh8O7qU7NSAjBRU85VmiG2
bR6iLaUI5zn7L/iA87kfiv/+fiplMW9x+6MfXU3oQJlsShgG94jt1jqYZSZWRMCieGw3fvEs/1lP
5ANwzdaK1xvS0VCUOIo3S2BY+G83bhMIvgKZ0vLcXN6pcGxTJPk7YOV3wQg8jWZjrwXpSprHLO5B
LHKXfqvwlIdvh2we6U1y6Wo6gArxpWJ5JvJgFjqQpgERrLKFiJLnRx3lVH9Q3Ay6SnIxFiAVCvhi
+wT9yBMSjaF4ku4EnLW9A+9p0JJ/0jhV3t7UBkHOveuvmeUHIu9bq9lPYWsamTePNkQn4VuHH+uG
hfIteTc1XUowNJ6xudsfxOosnYhyePDtg6+Zaxdynm/e8s4VBHXtjavgF70WcrfrY2MlJXZCT7rJ
OGDC+GqFiQ/xPljkGgsxl2Vm36p9v2eNdr0g/bRd3NNp73AwgwvGT50bUvnt9iY0AP7kX8jU5v7M
33USYaKneiF4xyiPPAL9+AUOI25ua+TBgITmZ+6u+uKB0d87YhLhsLh5EAqB1wbPIc41ReX0z7MZ
xcdt+QFT3lWVPnJqKXY3iANYp9yrjOX3VDHVSq9NTRt90ZYzM0/ZMp6VGkEGgrg+yB2aP7FW9TzZ
z5ixoUbAXDzTqZQd1hWT3MidqNT//ZxFnJpdipxCecXzZCtjtLufZ34xvyQG+8to5jDMlFOXkHt+
7jA6W5B4NxtaDjtxzVwwflCaoFGwHs4VYmHtmLGLfMwh0rE+j8a2xhkg928LnrwBcfWZU/fg5fzM
+n05TmlWdaDi5h/j3kBT/loBSDB0H+bTTW7bYxYYdoiJWGVYomUDjVZBmBhS94yTpFa18+M9nhj8
osSfbEVsDiqoUEcuMmvRF3X/kR3ynBvB/B2Uq6KjlvH1WbUsUm8G/6WxY/poxZaE8jPKdC7Ooo1k
IbP8/nZMn6hrQCL98VA08c+OCAy82fzkKE589af0k72iZlxOO2/KuQKHDERCP2ZiEFOVOgkzFmmv
dZs2e9HXqOWkunscVd1gCIvSilP5+dhClmarcD6NJNddkjPx6MTzW3PLY+4g46WVdzWVet87evLh
/BLqQ9RVMXcONxH+nkVLWtVQJcfGRjnuzJFzGHVNPupLvuDv1zAW6cS2tZtM5qQPqREvkN6ZNqa8
ixpTOjo4YnrmN4i4vSnrn5j4+qpItuWVlMbUwjPu8K79TBH5XQi+QL37Numc1z+ChSw7ukT5G9xI
fsgfEdCcFPUS7XLWPz44Qlisk2/Dxcrv2NCHIzAx9LJMbS+MMrtZR+zdE25bn8hM6m8epbh7gSAZ
NexJxCgycai/BPqR0XSq1QP3d9tMXu/zpwha6RG5gyvVjvfVbxUkCKvud97zGmZ64X8g3K1kdMaX
RoWji6zy2RL11TgVuEaGTEK4rB+HhSqW5c7FYlPwGHXECMXA4gpixr80xCgjpoRnQtowFPJ41yms
Gfco7F0v82gvkLqooxPc+W4EsyUZJB46tjlVeTFXz8t5AIHSETf7PSViYjRtqZFIuXe1qkHPkVx1
Cn6n6Rvn3m8POZpnToda1bwet+nc9et0Os2UG8u6lVAxmAivZA57f6Xef5f2Knom+uav3Gx6gE6G
uieSN7cgmi2o9caTXMFd2LROtgO6x1/iBfekImJWExJKh8YwVjr0g2omI5Ldz9NOaBOCGn42qkta
I8nTNFymc8NMsIxsYZuhHr77+01/YReHW0QaCo9NgIltCyz3DPaaJBKc9gtiTdC6YquStYeDmp/B
jADJCrcrnybWsXWJO3Rl9cR2OhXU7NOKHoEKO6fjDKeE2m8Q7Zvfar3yQtAlzLxZvyyd+vXvlJS4
CD+Mgja0bzBDkNk5bV8UpNRCqIeves85zhQhA+g+oL+ZjxPL/QYqju8VLfMnLlwV5sKdcMeeauv9
12ivWVSyKeeuDScjPHbZbX5Fc/CDAr1FpEuqsqhvtQbBbReimwKAukwwGhGaITMz7yLXC8s1PT9/
YX2EAD0ndD838lufNCVvrzjIwS7L56FbZKpBCzyIQLx6JuRhcT00cIQZfXgbUek7b+ixjICk64Sg
eFyJeN4k4hhN9kMjPwVgHyQDWIlGEjSsgV6H3978skISWqaFvTNHt0kiXDEcRYasRG2q/sEi6Pr9
AHW9IQQv3XBfEEuVqG9gnwyP3OHwX9Y3s+e3CQ7SLpVm9Z7L5UxtXseMpdFoFKsdVyomi009z9FT
Xqxhh0hPghe7oF5n9FSluiFEkElc2hkZADdSpBV1N/khAyHLCW/phC6L/Qx2nDQ1ILRvnpnzIZKb
Uw7OWOQrh3doTBxBmpgedpZhM/RRyXC3b+WvI7RFe30z5wUUWrCuEt3WIQ+QC/0lEOQK22nX0vjV
/9o7GI0VTZXjN9kirZHWuKw1zuVSFrRcmILE8GeUAtjUTx3HORCigTlohpTE84K7thJ5W0ngbYKE
SgzmYawZgDdy5+tK7Q6GIlp2ld9ON8uqYKGRmxrijatNh/zp9f3cnfi1VcBC6Y42BAGliqlexIQU
br1f9GmIkD2GNqTLRDT6ULQpxa9rydIp4azGJnuyRzxevNWT3GUIYQXITfGs1qjnInGP1ZVCQMRD
XU0ORxIVXYyemUQ/IiXLZfRxPzAHya+DUswu1/CMZC6OfKXisJ2QYwhLADen2sqs+3hlP97JO3lz
adLkfPSTWoI6+scD/wVmBrKkzVTZscy53P5lTf4zQi9MyPdNbGfuAtBTvc8N89gfQfai1CKpoRqX
lF39egWC5YxLSN8vTqoOVPpsF4TT4+iKQN4QJUFanNSxFGp6nOzjH1m7tnF6rYkGmhkVikJgyrfl
kpZsDFWmy/lLTn+T8rRETpNhu9zPKwxvk0qMrqGwiVYoRVljePW/m6/XYNNAaFaB37DMDc36wmdL
BVRWH0B5AzG31El8BSswBwQZzVWJOrPBRIRGo8hPxkAruyg2P2sE8f+GmrI5YnZwXkEYcUIrzR7l
658TAPDmPOfAg6n0XUrpFFAgS9Vm1KhKI2Nm+fMKUmDI6ZnslbSEANF4rEstVxPyhO8N1ZaYO1AO
YU65nS0RsizBhIEeSRzBVW4GfCuE1BBjknQ9lY9tY4sNvmWFsX0IHfBTe0uJwS8TtW8cdcXduxKA
hHGFlZHTr7BmqyVT3l0NlWFS4MRxD76+uhii+ZvSiqzPvCfLOuQg6RrffgsNGZmSdX30Momwvc/A
IS9IKQitgPRaVJ2JaRDeiCfj2C0bKaIN7O9vKFQUdFt6TzRT5ApC66XnqzhSiHAsjOoCpDcLsmmg
CIC3VHph0ocrCxPtQED2y0lOR4A7AgZoI0QSNlVInhZlQGx9M3xjiIjK54+FnNAPoicxJRMTlvJz
N8ooSuAmvVqnxbnaBcatlNEO9LLoxidDpwBKe3v0JFquJbUIaQ/wY3g3A1dhhvB8pgrCH0FDhQqT
iuMcQs0e7q7X3Vm4cK+ZXFRrAP/8hWADT5/yzUAcinmz+FkRtZvywDoapZXI2KmzPyHFOkVRE6G2
VDd5E/Bx0cW33L6qNO/N9BKaE6a+xXhpOw6zEF3K7vF9TJHPPmaxj9AImlcp/uhAk0S3eFEmdJSR
GaArmMOv1IseAOv4Oc2WyXrxuofNFs/3vXTHGcuo7DN9LjdxpwEoCt1Z+uk9nBBquhWLdErdKMWL
Pc3h7ZsfLRvcozCRLZXs91Vd17BnwcgZvMDLbkbEy4SQx6NZdtj62uPKVt16+DX1n0dGMrOooZfp
HOizToxRjibxWWUcciW3HqCGvB/GriloUE5myyTYzFPtrpLx7rb+6TQOMU95KCR0Xnj9wgPv9phF
kGQFBZGH1Hhz+OKCa4CGdDCFrAmWJ47r5K8eVtdcX3vJomhnAw6tWWiN8r+BPx02INS/QN0y2IVE
122BAzqX7ngxIL+qHc60Kidwg6rMKlmQVjbSe3r6+PC+zK0sTOLPySzkAXn1ZzTAEevxe6gzNx0B
wLJF86onIYlcVt3zTIzh+YI16kaqc3iWZXQ/aAlRKV0mVSz3XDw/Sjxcn8ggn9xWPU/QOdACnV59
cHafNjH/i+dA0Sa4792eNtxZg2lpJepweJkCNsWGj7MioDNRkkJKlC82aa439KJ5OpAVtGQEuWM6
ZssUeQf7vWefxwOQKqqMq4ganx/0Y7zzy2ULzPXzXqM5AHB9ZbA70JTljG4ZhsjJN49A0/bUJi65
etXhnfwRmF0lQoSentxez6ynOgUi1O27rQ1uu6rWXAm70NsuqjMOGoN+ck6XR4uo7rjL8LRxKSD4
L3qVfcNSKTmGU2pdAg+JnIrX2G8naTed1jSyQWVosPVuPz10dhVh/vH6h6f8SUhJhd6Jk6LVBbv+
VE2FgD13P/qJ+kbCmbXPhF5DquRmf1Wjif3aFnWAfBIGX9APgfPQcsIKUVPMEsS3DK0lRaA/9YNp
pWG1md30BqTGIqz97Igc7HFsOKRXTy7ParanAanPBOYtu9pYhTwyPHi4sEREKhqNJuAaMqZi8Jtb
nxxZjw6NEQmJzAIK8B9yUYQAn5prfqYyXkzE21Bt8DYf5uNysaanTfKwgHuUB5rKBKm6Jq8RaEPj
4kxIwKU2b9KIccVc/lYBRcv9xYW1dE4864sSd+LxLiSG5a3d98hz3CZ33Zhjnbm7GWQnJJSGnBlx
U2JnGPXsbtzrI27h5PSipBEkCOF9YKfQM06ifFUarctBNlt7L6lc3Ukm6fWJTdchKx3yW53KhShZ
eYIp6bYjkotHKuIInxr+Py2CEI4qqu/gbCL6RZNpoTfvMUEVf5FtwFG97svPmnYJjHX4jofUwFth
wJNdp6aWg5nT1l1w4+NVp0mCDeyzmWD+ZDAOz9StETZ9yTWvtksQP5XXOOzhgiO7UJ3gNoqXZ8Ve
a0fWWoz6PWAokePpEM4gdm0mGHAjDllh7mdM7jS/CQHtj8Y79xWr0ygWAaezdcuHWL7y5HSuTFq8
Xiqt3LFtUovspd2pTlz7qeROkTQZJGY3lI0d8GT5rpy+D7maoVZ9qXrfxeUdFsDqxQYhTvM4+eQM
TZBSChgeX58zbrz5JxFe3qHYHpwiHyhO5BfDGgsp7hc6o9r6jha/b05nt0NzVWP8DWE/PIYnPuoq
ViMv3L3UmxPMrLqT16AoB660jQYBg2qiZv6z9D+gvl+g2b0nuYn5zQbT0xkCc/mt8h91lv9Ezf0R
tYOwOpeQGJaO8GD5zpeeLihwv7A1XARI8tsvfi4MLp6NWTWuEjLqsXjFvjhT+LXflA7RsrNNoJbe
os1ggdWMhgWl4Yb5UhOQ+lNkRj7o71K6w//zSrgXTwoUsZKf1LGDHHPQBwEqmExTWldUTTQqFsic
vsNmgWNEKPYF/XoQ4kON/axvF+MgaU3xkU8rj6uSNlVd8Q4CjdfqPxCn0jezJvorBmpe4huZKmKb
LuViEI/wQA6StLAhXZuPbTnvs9nQg8xGXbBx+UN92mNNzUZtSRzlw1t5QfSq7tzOSAynHwwSqOME
ev4BRHUwDBH3NdgIHMyqoVjUrZSJP4IUT/iAuwXr8Ogyv9aG6pkzqEFjeD6o7xIglHccAIGVbUi2
rxWgKUHGOT5FGun9/qbX/EP4dZc4CBDMWBXodg+lhyeLgj8pyNG3oxP5Cfr321KOeLjAZMhnkobH
mzHfJnwLrwbj7Vfabk5MvNljRsOiWP5YA3gTCColgk07jcFgiJaPnbv3E5dNL+pqnt9mOFUn2VGC
KTpt5ylJZvdK1cv06RGZCDUSwHSf0t5E1T5SzNmtYEMI6s5aog4KCTN+Gu28irTDmUKHw6cc3l9m
8/paVQr5rtg9K/9D7ygfyGViHDrGykUyPe5ll0+ms7jKbN8fMPW31s1GJuFdT5UfS4c4W0ltIkC5
HQUrz62fJEQ1rBERo0WchfM5QjUUR5QfqKY0ZuB2iWkkq+jb4E74TumPZHbXhXOAlVuFgUmd+3l6
ko4RzjOzEJECZUBlBJPyp/cX6PpuG9gEWwv4EGtlt6iGnBhFtNMCNO0Di/52sG5U1wtggKE9BfLY
qU06hPkrqq/w/CyI1tIfyxECfNbRloMGVKu0D9/4sNOoUpM3BDeMj9zlcI/zolbiSSAlXwbfzSKi
ZQkYXw53PGLDzl509WeyFivm09EPPHzL4pTRhQ3Scv+FC7RfoXXL6ODJLHsxclml8/pABoCIqt7d
gCsgihYLuW2rjidOwRhmN9OPzcJmu1G99KnAA+u6t4uzVkxehwqhdW+ScqQMg1PcJs/v7znrW+DG
/NixgMJ77hrFvO7Nd7rSUouhUquaOmesCK9yGcoeUgRzD9zZo1aN+35GTJtsmMcjMOMm6nXntAEi
8yFwrg/lqnect4P/UKIxZNKGvPj/tKF2zTdz9Ii0JzmVAxsNYbqlgSZVQHFFu9Dky7oWgxAy6hjN
K2OVjlMc7q6G3ygEkQf49jn+PS4xqz7dkYQDdYy7D18PnUkF/18yld4Vd6NDMrA9quecyj3xUHyl
Y2KGCt9hGjLzebBgwoQC2Oc7kOABeDJDoh0ZQjKPyc8P35B7w/i1Q54CjT894VVCkNwirUGLHiFk
cr8f5X8FWaQH5XMWuIb9ChukhokCpDE0U5izhBu1V63gv9s4Wq0ZdJZY/98djDjCEuzwPtgK2KJg
6bBOKQbta5h52oITI5OhYRSc85j/Zgh0lEqpL57HnFF1JImUN/lnzN2yzjP9SRHRn/ZJctpdQJIN
SIObbZxHHDtz2fS8BWs9/RD0jsaaPz3LELGMyXRebbX0VlBh2aVHiftYSeo5my+LopU/PVBaaE8X
u081sP0wdt0/ySs0S5RmzwiLBB/LT9mNNTCgJXSP9HHpx6ABX+Z7dNHPwXI9TdzUe/3o0bkbjCuu
pkhl0tzyzAapmquYtOX7Wty+iA+e14l+cgMhlz2P4tEEspGDJZE/dLknewyVK7z30kRuQtqzeCQp
GNjbcbGoGjIcDRng4R6uqexvbsw7mI73+QnNC6c61mHuzyPwvWl3Oz+QZsI5Pg27LtSit/EtrzZj
Gvzww1HEMNC+eD00Q8m10dA/zqJ7BtI3qlEHa8rLpEf3IEmN5frFfkSadPmKN10RcpLFKSiicyAW
TElYad6m+7Ck3dEI6sR5Z4PNBynaUSFiTqijiqYXgJWHDXmLvAvV4VORKtz0QN3GyetSew3yVgg4
LUdCMBH4KALpdpCQsplrg63Va91xnjvI+47kTh/TGt9OglIVmvYG+0YtTF9o2jvXcbpW0RXaUtrP
BYsvNo42bC0+QdpWepFMVfhmGBLydrcY37G/cPjOg6IJYaFmsrtmRXIn+UHyqmqwbg732xLgAPjo
YuhaVALuaH/V5r3+Trad1QqUJpn+/8XacsgA7oB74hs1JY4CNoAJx0Pbl2eRmjC3EFJhHDaNB09m
88LSvmV0zK5TtnMgCKU+GivzeRo/Qf0nL3OK5tgdbiM1B6GSb/9WEtoBcW/xCs0ZJmSFYzB5n00+
UaskTu881Fos4exVNy1TLKFAFlw8UaXjWFRI/bSUO69Ei2eRWdBOWXvFDsl5VoYLbMp/TiX2BBUa
zsLLgPml9uzSNUn8vPY8HoigcfCqiCFLPFMRdwdNSbqgdq0JOWrpLtnNwfquZv77RbDQtGrfDELj
0JOcZasRgmZvh/f/intijijBT2BgOvu5p+1NNu6MEElUgZqNVMEYZYbOMrb4NfrrGyI/UiIqfNKY
P6nimIB8/nV03imyzXqJ0r4zdO7xJdLF4Q5ow7uufA3NqSCqqd0x7jLRkkLfpPnLr3wk4ZPhOxxh
yiV63GG9zMsq+TcTbjD5d7sUqGREtfHoCfNZAzZuL9qyEZplhHT+nsije1mnijsi4fNXsm76ayTP
x9AoZx4MoUk/tDaehQUcXsrlrYSJxUTuMT2kd0110deeZYKFyWoLehUK+GVhW4FGFNpbW010u3IP
hc1WBVO4Y2/h1UcXH8EdGTL5yC97CZxDCDyVcokHFEFU/LKuJ7xdb87iNNP5nROsuVhXIsHK76te
DUC1cklvj8p1ZuSGoFzah7KiN+QKuuGvgMNeYJYfOPwrByZv9UeiiYjah23OBt3MjP19z9Kdjqj3
dXHLylJw1U4WrAXCHR8kQfv+2wJnO7BodWh1iiiRzb2nJ1OckU6DCoC5HR3tZXH/QE9OuwIVN4C6
j5J+gfcGdWfduyx5y5zzypdCpZqjon0NPN+Nxx34aK2ViO96dZeeNYzwTQuOqApBnteUZ/2bqQOJ
QIi+xdMiTXfC5fxByvtxlhc3imbUtz6KrzEaFjLdU76nR5xMz2o6RQ/D1NuYoBdM7iPehzs/miIK
XxoKqvrjqYb0RXRf9BWVz3xh8xsbItwKMf69gpRqEv+9V8UmH076LVLa0310tOYoCt5j1sle8ZHd
MgfN4adVB0RKMtFA9VvuSo1mbSpyR3QeZwEqNHVe8Rl2v6EDGuCVtXcTCBxRtdbzIJIK2dUSWq/i
INvlg3Yym3N4i9sxiiBTlkcoiRNr24JFGkGgCHFkPBmYmskoue4OCaX5UVFgGRBIaa5UTXHeVZbb
82aCwLmyVtDmJDPXA47tJ1UZRbsPFo0KwxG9d/Ga+huVaJi21gVDNyxolKDEJqaK05bysmKifbFs
JUcjRz5h7xERB1cvG00HMb7IFo4LOmT9RQ5P4vNVWn8DPyS5XS9GGBv3Bk7+33tSzqQe7p+UtHIx
no4GELx1eFbOcWs1MYy4U/KIWcJytE1AIuMDf6ETxJd/Td73GPgxdnvp975mJVnv/xSChEFs0NXZ
A3G2EwQjITk3g9DAnPDM+iBiBq0dVSXkcYq6tPoLE6JnCH4Tfid7bVH+wBZ2igbtedr0J9Y18kBV
kZ1Zadb5eGMkDIJJdEiGYIn4p7MHnbBRnizX64w+nIvxCKTp9dYr0bn6BFBv/MHoQoTBKjYFQxo6
Kd5y3cQW7rXgIlbvOnuC/ZkHzCkCn/yt7SL0HnRI0gfHJeoTNPzn5Nq37NRIvgHH1nA1Pl1KMzff
QqJjU1+wFSRMN07bsLi/o8pbkOvzrMlEyDY8tMYwd4z+8Zweaix7pTKUWb9g3j9CNMAn/Uv0DVl5
nXEFuNp46rcBqu/FR8Uu4CC5lrvZXD31QlipXLNoLAoUYqnPj4ZhfkyKtKZTM74I+ic65G4VZXTZ
HDk6toC2HL0T+mDbT050VCnHN3QOf3J5gOMmCh2kug1H8QQ3WTrs8+gnKS96b10l2W0xBGMx3XHx
J1XXNj6lT/D4qwGKnRJJVv/D2uhYKwSEimZ7W1A/7Nu1VW3fZXI8JOU+gapZpMmsCrik02HwfjJu
EgG1zKv9/jMFXfYyfau+syYDQPeTibz1aq22aG9b490Iug3M5ZhRWzzVRQCSL1lB449C0X9h/s7i
ICJgw+7T9tsgrtx1Nt/vlApfk2n/le/6V7Oyaga1F20JlhnTg0ZGa6Zdektx6J94DMj+fvlCp8Te
7bqnQLL4hvgf/9R5HS35JjozrNfhBkLR3B+Igr81z8e/VxsBqanbgUxrG3W+TKWEwNff35X6BhiR
IRyYZrYLn6ytjwPhWEcNFPczOsVE8BcRpFVUWl2BqGSUp5g81qKbVHrEAbO+Nn8zLbW2SGXERHAD
cg37aryogEElDkOI5MfaPgpJGfAXIhHYRgyI/jOx1L4FaoKNIPO8OshwLDUDdhLI1JkDKENPT88M
mtk4E6oDpbYF8booPjpj1QMBvGBciFh5jJVTl4wjuIrtVS1O9sXN+VcuaLOGkzvVLZhDMb/zySDs
DVnAYvXukATyv7Dh7aDD6DvoFW3IJVjYoL1ZS3aRtqNvk/nWv0oKzBWi7snzELd8E+k4UodsVDDU
R6AhyXi5dP8QO5LpeyTTrx4XJqfrGG3nOlgbQGGfKhn9I13TPGNeuzQRlX8Lxt6zhtVVHXyaAJMM
TqSxA76CX+ru7oltxCmd7H+XnOxCqJ4NWTHdUm97ctT8BBzqZgMTXezRj3kp7gSH44k/jyeUTp5H
UmcDPio/hUb6TwnBFlg76In1r3Z60qMH2tuEWbJ6+NKBFWGFb79n/gETuDvELayDsysuRWLibk8/
F8jnFnnP14deGXeGyznn4CS12Ps2qPMAhV8Gmc4oSNYS39N7m4zQw297ktemAp9MqVscpy8gv9Fn
+aygS6sdi6Wc5FualKxSzxRDi5Pde1gDXwcQWjutARDUoFLibyQzMUIdCNVQCqUfpWY+u0FkN5ew
vaaLV2+8DX/TsNAFavSnaqsmKeI6qGUo1SRgZHG2bJoppERZU4XRKA2h41DHLAXBbisMo1CgoBd3
Vot41yElU+P2A2AFFebQjj56X1GnuTYaBFgVpoeHFkinEFB8mXzJEI+ZBZXB7QagesxlCQ09/dIS
usU0gNWBWTLlOYA757AF0SOyioBITmhFmB5lmBv7d1Qp3Z5K1YTHQxz/JW7CdeXfmSTuJaxbvG/D
hruwTCGktteEeGTzku+HzQ1Bvyg63HxUm5JUVKHcYwFSzFm8gdcPqvI8Bv4Eo5HOG9OBehQ+rYny
26TDFvBE4dH55ZHKY2FE27H2ql7er1xQ9ln1TEJw5/OArxWyFLjgZ3o1oDj7tfN5W4xluFwSTz8G
R3ygUuun7FiXFZ2NgYPJQXqPYUys3ca1Qcpx+txS44FO3XNx8FCtzpLgKHX8xoHNgd/gt0n1tAU/
fczLaNYv1ShKhREeNFTOH80NocfxABdoflwy3oNHtqGFqmLoT1cB+GZEZPPPNXlNg9dhh9yiz/bh
s5v6LuE9n/k7toa3CGqI+S0QWIy+RbvCT+jGv90B6APgmUCh0InLIQLJv/UUe0EzRNtfPX6OYb3K
FjJ5+TcHS31R4xarJhyav0P4ybQVFpYShhXRoH24bztaJRF0ZE3LoeQ0i3C9PX0NFte+d697GdFw
vykus51KhiNjFBKhzA+GKkVgDzkpLewUjrR9jpns5olNXDz2vf4UFI4IusudmFOaRxTyRd6Mg+wp
EKKH8LGrhZuomvy0QDU05Qdq6UxEW4syP6VK7eiHOu4I1GfPlbuXahBMaYLcAnySimqXggpIOw7w
bnEmtQRTv2HamsYXlL6OBq0koxweJWPoXFff+v+4ls+CXDpwmbEdyB1lcZ1bnOchIwgezB+P089J
lEHtlYyutwMuitWaLpXiuVMvCA6o0vrcm3T2ae8UVZPZMGam2TKnI6Rtp/tlrT5rCqnLBWVi+Uzn
qrVGsOJnXVjqH4Cwo5A0/ff+nPNYVYeJfuL9FmWdygegZvyWT/YsYn7IgQEQG9H5SqwET99rrHIY
XW3YZZb7nFuCNoX6e2oUFW740uv4y1C9PfQbmTuj5guqD9nx5rsjXYneOYNxWLeSm1CH1fxQjAFd
vQlXGqPYQwP8eJt6ZtFkUxqObfy/dIouDjoL0Hyg3vufNyJGHnErr781nqLtXwulFW6GTTbxlpKk
A6u2MdZg+W08WXdMLRDXLr1LcHCO7aVU2iEzbHIGzNAjn/Kt6biXX7BBLJ+pEs3zuhgRfOFFj+UW
UUuQI8BwGuNuzO00cWgZLUuI64rlNEWaiULwQDkz62PLsaMEGHJqV/mMAeSnDzthz1I2xWbF/NdJ
EukPGBZPA9go377RKVbTLjeFnLOl68gx1r/sjvH0rHkPbmX3/l8di4wX/P8PIsPyR1lq96nfVyVX
NWcyWPwXBZSZNSCOREXgQeVWulLIQ2ewazWP+HPvcXBd8jrvtuJvf9bR+FRf3BHnv6hbhxcbQ4bL
GGt4yzfns4TbnUYtQHq0WdXbMlx0AtAxNyaY34iRcojc6M/QVQXQ5hSneL84rDLFYK2SErliVZSI
VBaNmezwGbKDgauf6Yy52OLvP3rVfQkT3D3vyZgBJQp0FJU5fPKj08YNdLmNam1vyUc38gG+lZZc
UL2XjkNASLfZGbmD3Tj5Nz0F+yOlO168QJpuxd6jnNbozWMUuHQ+yEx/99Z/SVrP419IJY78g+U9
lWpMHNpJxz5P9rriuUBf66bvlZ3ATPGvEGDMbhfAl7ccb2dNCrHwFJBxvzkgoQICQLqk5wZQV0AI
hkIbpvUi1H1XXHQoPuXHt6x3UXIhn0+mGGmRe94OcXqqRCmHp0EBs8UI+Lk1e9tJm3r47nOsPRH9
fVc1YfdNYQ5JMqygaiAmYtibkDAeZqtDoJhaHxLl1BPM4sDhFX6a9A4hibeMR/p8PYKRQXPGdP96
NoM3hgNHGVvqIuaoOjLS5HqjWN+o73r1KFKApHRVqlvd+hNUqYZj1/3Pf3VWgXVWBq0TaVHWGcLl
OMKjsM18kT3JLvEMOdtb7xW9ZrjGz6zK54VaXm8pA5tozxOX96b09ApYMaUdbw1KqSVwJ9ikDtVY
YF5s8q9G1ImjJDW8+CqH3wZQNrXBNKsXDbO6AqqmxjcrNpMtmLq+mPBGH1v6mD09CdhrzFRR0MQH
kXvTo3C7hPI4lDfNdafhea487yW7YMEKNW0BydfarBbn7YVsRxI5W2des0U+Mc9jPIXbVzA/l7x3
hFcU+5A909B0Yb+7uXEedVL06sIlmIGeMly5hUnLUBL9C8/cIwuerlyNI6XO5zSbpfG/vzjBlJb/
muVb2pejrmaA2gb4JFQ+TGenoARYv1gs72x0Y4rWRMbXzIzJoHFFYqpXbmBFhfxfnXNIfdXazLjS
ZPZrJqhXMdxG1blyzZTciE5W1lyxmXvUbdRWvaEUo/jOK0bbcl2gezVnnfboWyIwmyeeV2XWH8iv
6mKtIgKo0ZFAWIa94Yc6l5wLHCEDzjOAr/OFFryI/cEnllImnpsO+fokJHXEOs0h71IRVL8q/Vkd
PCgaoqcbywS9Jrft5spRu8s3Rd8cx/1qwJzSxlG1QZVU8ofbfzZXzt4Z2Ilzx/ck0czqaBxp1bMN
YyxtgbnP/hN+h8nUUIooV3uq/oruhcePDpwQxsoEFO0zkH5yH1yQ+kVwyNvxsC1YL/GK2PB25xd6
3/HwggflGsdniEe7gkhUvfER0s5moV04eo+lYTmvNSj5dUf5MdTn7GT7N/Wvz6FZENnYgKunfeX/
NuSI7PxoLKIZzx8y7iZlITTZRZ0VW3KzeW2XcH7IiOgr1X3lGJOx356amfXfZ/8JsJ9CasJWRBWc
UlGJFTYDqJqVwHB6kPNFjSaoEj/4LtAVRiY1FtPb3UNzkOJaUzEB23lxlOnCBp+/h1kTyn02ijmR
v1zWpmxzLROythDiOLrFK9UYi2qRRy8MhVMEmmAeAi+APg/W/InJXoWGTjY5KvMl6fmVcQTZNERi
tNc3ZVcshIo9/nlBTCpxNPrR5BafxuJYBEEkQmBMWD/QXsm0TsxDFPkS89PAXnOKXP3uBHi2T+K+
EPv/RJ6ppBrD8QbEs/3TXZQvCz789oR8eAaFiFcfyD+F0K3zphBFSuYzxGmnBaVR0pd0XKi5C+2m
dEeg+N9riUVLWozYYYNYvftO7ATSPEZDG/bvecYlgi1XU51qdI5e+PT8mNwAfJlJ5znO360pqFJO
mONmD++g0hoUsybQiy54wFl5guFhSY42Dz0G4ttNcDvA+glBWzgyLdmbHH1nK4xCekpEU9u/5lvv
FClvp7Q7LphIlt0HeotCeblCWD6kWX3Vd9vIgbu9lLFaUhahIOXdaDp0bCG7RQZxijZE9u9ocY6A
Wr3i596NqBKY1tGD2/B3L9bEXSKXV51s828i1PBOn8wLQuzMfZuP//DGYTkQhISvZfX1tSqqQsfs
lIuUNcMpwF5Ko6zHc1cBQ3wzzreK+R8oNkRk+KAwtIhy9oXDymfZtw497BsqwSgG7C0H/N6hF+vv
geUSgiqM8NQK3OmkqtZv7r4b7A2+KisQ2rvcfZo9T1suzvHQ55kbKsP+caXwOccTG+kv1mJ75n0s
HYEGzTdJMZtEAgyvj5r9d/cnOzWFWoSrfUQ4hmXjKShnbBcsdkc/X63PjPY50Zkf2IjeUg/dt7QQ
2bjgm4q47mWJN+7tnJdMSRyeGGMekudTR9WQSppyOVvJJuaXghIrK10X+9MPVKgUjggoS4Ifktxk
4MrPDyPa5kqdkYR4KkXDfGFke+tWsAvl+kVKLuocL69eEpax1VwP4kpRZR/gMIHMpiVaDwv+vgno
+dsI0f17B5wJiv1NSsqu4kwyG1jWfGlcZUPY8BkaWmRJmITKKKyUxbHpOWVE6W74si6z+6k4Vgpi
VXzXR5mafM8vDvgqvQch5bV7BDAaaqdCY99T2w6gkgqGmbLCfPcn+Wfd0FfQXEIvU8eArr5VkV7u
ufhVWe0oX6jzfp9UZK7PVDEbrUMh0Qq9uOTTLxZqxYfU136mtwwoUz22V5GtDX3QTJHlPJ4GVNCq
jUkVk7NjXpA6H0DtOTUNX1PaRYkC10p9kvKkdP+7sZA0aifDGYIfMi8ZGwUc62E0klQ/Hjl1ogla
5PvoD3sXcas9Aif/1WeJu44BT5VNF6Ryb1e8SW1Od2enbOL2U2EpewtAbPtnL485iCOBpGrQT/xg
IAf81qvZcDsqWyeouqqN/7MLQTl5ImYpEhIHOT1uS/9hHDV2cDtrcZ874UDBWsE5PA/2WZOwNp1s
E4nxdgzqHrMKbs01WXvFmqEdcSsv523aIFjoly6PuiDXM4sqx41zsmj+yYf/Yagds8JyelcPjVyh
o1bXJVENZOSIkRtA1APrMirAzyU0HIr/yEZHOaZA14q6ftP6m3u5u1563kEKtd7McWpF13dJr+pk
SQTb6GiMVAdggb6Zikl+WuwdohChOLuxj69UBWMz7LuiMMU1qYNKX3vDoT8Yfmji6Fk9Dp7DfCuI
jG1ICrWqyWmT7hPBJvASnAk2/83Ie667Ja6k2jlNnG+WmpejnQMISJ85C+m+R2Vs+78O1RGZGkn4
OpwwkMHvyZYKcnACo5KmAyja8irKCkE7YP/eDq1jWrSwQh5WYWfn2vnsv4bV1rEAkDr8uCjICRtG
Zz8cWUbv51bz+a8Ets5R9ZN6Pnc2kSg3Hs3vw3EjppBnUOFpHonmbA2bF6R+ikDCWX9q680UTrm7
GkvCaeFY03aIXCEwm1fZC4UPz9XsAoZ4w2Sy+AwDeZztkm9oEnoOFYSa0A5y7769GYD1Xw5kZen4
94UUnmry87qZStYs81dTXlUZPrwx53F6KjOfVP1k7Jy7z0nxMKHc0EnexNDiyhgiyA+riN/8BE+V
b/52wHYsXaTYMV0lwfnlUHY59cz1yE0KvxqRQAUodsUbcVCh6JY27IitMmiww8jwKktMaWc82ufp
AZGWwiEPhNhIrHWsnSSm3x1KLBtViT2Vm34sGxKS59SKWP2WCSyKa1hVRR08hV6FSQerYZPGveqA
qiw7JCFtlQKrscJJffGSbLKqlBqIe2gj0HYwqSyjFBfa70y1xOkM9tgZUW2buyn+KfW2i1/eLMME
speDRkVQtcVqxa5Jf2+mgKJekZqx9MI2qAvkOw6vfLQ9YHrhXPb7MbghAcJkG49yonbwFn9P6XnX
NdP+irh1QiV9HGSrTn5gt2k2Njj3//yWEt/jioQQhioHUF8CuXMFK1KazoT41m1DVQi3Wjh29vZF
7xY7WdjywHdUTGOo3u2tiK3tb8yr93YcGcQRK6KQqCTtQ561TebgKdeht3RNd9kiraHw7s/ZmpZi
HCI/nnQ2bEFR5ETK4osegiue91eqFRjJ0hfcb5jH/jb+HYAIAomddq7j/caocGzc+SdmcR3klJQx
5hX4uXrgv7ccIr2vDsqywjP1DDuTp5S67MM2Fl3jFmzmwC9kaOMI8EtEfh8anyA0hB2E7tSK/nJW
iHf9fPSS5XwDWYtOcz4tvo75SwnRCrXLhVx1kIgWnibZRS72EMQMVoXcFCAsw8vo6XZLpvnPADO+
myc49hwPZCfc6AkpZmq1TFQggOPFok+sTMMQx1W0C8aEiz5Cy6SwzwU2pP+4Ih69Kkk/CoGj0vpP
QtrocLCCuNFL9B36lU3JoPVCsQsInByNEfwF10OzfZHr+XxNwzMzWihroufCMj/JNEk2D65zus9K
xSxz/hSjaZR+Rlanb8S7JiPonpdemXGY7rUHlf1dHdE82FU4eV8wcfJ3xI5MIuF/oqSVHcT+S7r0
QiPw50oF0nNXLD+lmmX4revqRHdqCUas4MbaAO1KhX+z/4vHtMMRAMzyiiu6G5QLRf/nZkrIp65I
Av0DdAF+xm7tjdw8AvOMAknywpWLLKWiwIa+wXQv+sFU3w8d5fQIO5JiliU4CWdrzX9H+p6S+7he
l3OJFguM4z+WYRF5qemvREHrpieB/2ukU7TV7yJFnkq0WeHJj6p7t+IXTRhsJe7rl+yrM4jF+J4s
tsL/5FmhkLvP/QNBcG2LjIw2ZN/z+ZLgtw9p9cQKk7Q/syX7XoCcoxjyRnVj4P+n/FXvJ5Xwfla7
6QpiP2qPdl1zW3XIgkMgk4Fpz3eYU6oXGU2iyOSBIIG6+eESnOqpLbaEnstCePSGcBN7B00k/WwN
+OQas8WPu4IK06VoMBNeGl5NUzhbADTPv9cmzSBmsmQ3coRtOBouZbkV6FrGyh8xwznMk0XJ9fsJ
aU9DqF4nooWcz/3E3fj5fRSPOqXueARKGOBjPPkGJ4SUWPmlPaJG5n7azO4hpOqfgRUd9eJs76iI
L48SpO8sYBMEkImZnW+DhAkiFjzEfF7APPQUFnTUYiefywF6QtC7DDoSmQwUV+l/DcnyITNFR/zE
LKeSV1J98r4+MwC/upx3wjs9lxjANAwYxRQO94PQPYNFt2CNU9hP7IF6g2LxiCvIoUlLlDfkp7Iz
1bUgAVnglLtpa9h1B8+Lr1Q0A/qiy7YM67zjoY8NDH1KdB+0ihOfq4A03pEQHQfny1ifoHnFjrVX
u+qgqxkpWhVW5cz4BJbKP2C8Kc1QnVn8K0F5FaYgWkXXVfVtafZjs6OaqA7DV4cq8CqbzE8s3mQp
QaiKK4Cu2sGpelhrtPkPXqGvMAKT7wj6764AHfFQP3Zl2XfUPSInn5HurRT1ow9K9AqmXvRwmgzg
wlQ4WdVg43kgW//n0hiOxTYlHK2GSuN2PZ+KEM4VMIUPtYtAIHLkkJtT2gMoipitQTKHWQt33FiS
uprsaMllVzSJoP+KoPnVfYyo8KPulinIpo8qULGvSpo17FGXwxrXi5Vc04Q9o2ak8tGmssMrxXu0
qUXs1HfQrekXsWDyJ8N8r4xrbksdLDdml1iK6Bdw2+zzGiwE75DrZ8XEzOh0gZ8VZQDHaodWHgR0
uL+aBAtN0uWE6djxEn2JPucsJzJdemGp8s4J1DmlKMD3+4U+Mqj7pUoa3jpYhjL8e4f4/9WbOoU1
9R6d97ZA0WvTtl7ib/mgdt892kGOreaQNlm1GiRtrnptebyJFTNDFq4Wu59MzsW9zpmGOHn7ujX0
ge3/nX5addGfCA4zyVArpnZjwYkIcnNxvCS+Cc0OK/4bp7yTLvRIbPY5LHFuEqeZD87j7TKLx8NH
U8oreaeP/x7BwPB5RjbNaVQNzv4Ui0h/h6OIVdzDB16YmAnyg0/F9LOdjcDl+BxGQcVI3iBhrw8w
a7PPUcGyAu9ISFT2jHFxDYZ7hutIRuVkNNrKxJGWRkIL/OflKHK9YAL+v2QtzQaKdYibusds6C93
vGc/ioBRmdn5HvgzKyVuZYzv5znsKBfYcQaT1ogQgKB4UGteXO6w1RDsRvT2+jTsQPGmwLUa0cCq
tlMyDLYkeP9XZ3DTCYOB0cFwsS8fTIDKfWcme8vH9igLXMZjyKi0RmAbyQLdr8oL3/MUhD9nzGm5
eUGkAuMdaO5VwzhSt4Sb1cYwExikOcD8ahCduWWGEEr955QQIZmN/ELKBRgxx1S+ozVtuL32g+m4
57PVKXfXG+Hz0dIGXB+2ieEru6mIQALUabFuDgsCL5y22LfH0dNKAQYrY1DOJkYjrOl/AFYHMSjf
FCIE8HG0x0xr6PLk1VXBxzS81/2olMguNquJxnPVkayvx+B+5tcmEI7ZI6j1DzCeexRE2z9Nzi7p
L5SUXfbWxw72SPbz0zP4xkt65nRVHxSwfEVkzw14OfqvO/MGpy92u+zCNlpoMo5h5JPXfLwMddMZ
2P5X0uHKl/7t/NxEO+868BLOxnq3Dx14vdfYm1MhVfbvc26uNUvllY2tF4xbVD6FvZHy/UCV+Yvs
4+T+5XWuttlk16Lkq02zrz9nYsFbtGT1VTwgu3SMjJYIM3bvJhxJfdIZUFnyASllGC8KMK8pqp4S
7UoOgeuqHcGKxR066nRmcKj0O7uvzkmYduwXWCEdfL9qbWhR10PC5001OBy27rwNvU0Sgc7iLd4j
Vd3seigRnprsiApgP39be8hSJi8l44ghQY2lU1rDH5wnYm7V0jLbIbXg1KqXyBoX23HCCtlymKtT
IQn/g/JiOyT8jBd+YKsVp8vOwhnr0/gBFUmWLeXMxwD5Cgu+JbPlQV+KBX/HAlfRWl6VnA2Rshv7
pnnmVkOmYeDPcD9a6UvDN++zAQmqt3upuLxHF6EB1uiCKRnmSZnX7OJ/YaOHJiwo7CEPMdePq5/A
jyrSN704VRc3SUsvmj+aGVqembG1Xs8moOWUbad4v0RtQVFNMAcv0j1T9VQF6qo6NpHc/WR413pn
RewcJvCrgIEm3C0sKLM7IWRPH+tip7Tp24wx4lHCrfIqyqYs9Rnb7+bJSwPFOXTwsARM94A56odZ
O/uBhIuOLKVThgc6sZYneGGwSV6TVaD5Rj1/GDS5DuANNS0GP9g/G/MactvSUGHauMV+6BypqTsZ
5iJnikH/QQWgElq6flc9OylQMKi3JF2s4hZqsAygrQWW7+5R7m5bWBH6SMnhXWW+gyNQafZKgc8e
POyBjg+Ls/IOvFQgxFjA7aqWFWwRB2f3Qt2f3NaKy4rKeSxIEfXL6/RGbk5sDbgeDvcZoNRHGkEh
SPOYS2nHM+WXAsIo6ap221teKpvg/Wp3sLB0tB5jCocliPzivJyfd+hxwCiik0lErvtW42meV0CD
79O5oq9vePskYZsacjSq9b4w0eM2sgnR/qlp18D15XeShsnLy2Gvdxo61dRsHVHY1A5J63zkro+k
JWxZcSjG4EHaPAkuKuBgy2DhdxCbcu5LsXgguuuAODlTCzfXd+jNwEQ1GnY0KwJ/+yFvtfsNH+pK
D6/TcfSNvkYN37/Y5bFyr+q5gDl2WidOlbrWCf01+ngQKkL+1VrezkiKL0DH/l0VoVghmjlD3HWh
AiLFS1jQLBG2aryeYcW50ylNq/lNkfbpVHNp4N8MEJ86ukK4i2h2m4XnSYrp5n3dquYThhr0Sv0r
zI7FES0xmYgooEVZPEXKFbVBkEuI/4v+96Y68iaCVuwsiRFMrtFii5iYLx2t7uUChScU5P8DKrtY
EIFfE3m3l1TZoeS7VHwhcgtschXVyM7GvV7y++YbhkDDizYhQ/0RcocnAnci5bnB4m27kiB72KXU
ZFTR28wPU98jDtmYt06BWXdn2O3PTh98/E4AkxMJCou7lIqYGfdkMGxedbkLsG9VnvC4eo9VwY2Y
RFlzYo2aMecuAvz0ElzjZ/BoCh05IpM/HlcuPEjajJBl7I1qmea4NoJ/j42S6j1vwv8/J97+cDfu
wqm46trLaV47FreQDRGIkScfpW+vuAag7Fv+8sIEBlJu5nLR2s1ExrI+VCPqWcDxtDxTVglFOxTm
6LjS/ntlfrFIGOjUE/4pVgQ4BQj3hfQQ1Abz+T4qxK3hDWGHrMx2DkYFpDxc6wvZUS4fV8m1zG1k
RoBamGNSavPtlLXikrFnh4KdARsTaWlXoxxL9XboVfakNk7ALz8JtjVqR5mtZFtGFAVQeGrWayBg
wPasAGV+Ny0oOEg2MW827Pc2U4cT3872FK9Dn4AS4ezSD1EJvF7IekJDnqIfmByUcw62pVhxpw65
NGpWgOn0rCPpel5aSvoi6l0BgL9qLwTuZbgmfiPp2QdJXF3KHN17Y7NAig8gqhzhHJso4b9UJ/Id
ZFAKKQGIKxI95S5+HoCoCsnJE78VtlxyhWYVZJ1fUgFnDq913G3MxNkefb845Z/1KhHjXWZFbg9c
xOPmQn+L8ERgqShziy6b4+UnG5QKcG7GvRD6BCgSfWlu2dI7DANj5z9yUXwRDGUnnHaEsUoAZUzg
Uoh2LQQVrol4u/FAisRhLMF0xuWkS65lzKndO/tLS0YR5BKLXAe0F+a1U8wOL0h9g8N06kuuNdcC
JBUVQgvTxWIv6QVLyZKXh21KYDtrj5kf8ng+gIDzmsCEQQqp2U0g+R5j7bAMHBBxwX1q6yL7PtHr
Xjow7RktHaqOqBjs7JaFCZ8JbSPhgzkS007EMogq86LpqXhMXYfUk69wyRs3AZwWunZrigJzTjjY
5yTRWh+DjjXuPKvQ3QLUvSXuNAp62bfRNa845aysBAzzq8nt0XiW+n42T259/v+uPD3FYCY0H8J2
MIQFehI53VzBCLiZZCZCDMs+WJ0LtaI7kWg3632KBhilxiu8L1FdaHnFL4mGDbNYoDKF3PlKua9V
8TuQf8c/FNEJtIHHdXzUf7+kmK9ujcrPGCl506KNaovxLEr79VbHS0MGtJgrS4zqaxIKnRqdXLeS
Txez8jAvYwZWWn1boP7k/xfIkZMSGAEbe0S/IosvgBJmb2fjjGM6CDSxRI3VmqINmGAW7SMsJbxa
wpx9YYP8neT7uhv/A5Yc2heu7T0i0G3GOFXHrwXephg71V/ybNXeaMH01TR2/ikov8xXsuPGuj8f
sxdqKI31rum6Hwio0n928f8jW9kI+UwaI4P/kWRn6SWezSoMxcLk1+tsJGckyIIiwLuYCteKZUi/
Fk0sHCSNo4T7GvACafXgqxGjTX6jtCsvdC6V+yxBm4LRqZml/O8mZyrAcUCGR9iBHfdKtN7RnHy8
uzV7ofA0TDzqMaGkf5uf2jSOIT1PLcvgoN21f3Nt7DAPwJKit03tjCzxDc+cL27vw9coxC9XCKSw
e+s0A5vOn9fhiX90iuuvzI1BVd2YxsmLdjPshmPcWMlrFTE4MrX/JOfKtz11g3sNPL3UZ7oeVyjz
FR+5vCPKG7bulor4uiZbAd1dNVf196ks1F5INlD+O4ef3MZiZb1BwdDC8frd1ZRaiVxq/2djaqAH
phptXW1Lmw2IUnt8uWnWnzbhH56T6QgvisCpbXHpDo6No85TEkL+s4GgDnA+5R5um2CgQbyWQGWk
ljC9Pf5uS+VE/NbjdgpR0l4hrAesvwQ5WBQVaqFVhA+im/w5bp1bRPAO0ITfcck/B1UegRXokDnM
Jdnc4V1//fDnbG36yg/8q+ITU89VVda1nhlfqI/mz8FSCjlMIo5ckP/T3AKqOjMt1obon2HibSt+
r8S4xGIrBC6A0j3rqdrG/lbsIHrUsDWmCeGdpoCkrTyGktAk6a7hMlQGbLymek8hNNxc4AYS0HKm
mH+t6O+tiISWWajl8s7K67dapp9772jHKSzVMz2mkJac+usxdy2yKMG7d7PU+trRrbOfgvRaR3U2
D516UtBhS0QCkCh/pDRRMWLy/YlvTkD8CBZl4wbqfrvCCyYLiwEVzCaHF8NSFF2uG1ibel7aa/uE
BViqxicX10Nn36Gt9Lv6YDXQFI/3+Uc5mmHlQe2ym+Fopw3eYlVFNd7kf0D9/vDVxsAjm0WQGc93
DbDVG1y8Ww7QMMZi0BouLi5n8mI+d5bCwXmx+T4vzpKtcyQQ9Nxbepml7OblBA3Mg9IulSl8JfDr
dG4qhA4URRybb48/SXf4NRV3Ckthg3EnUM6H3ZVB2mPHKW032+B4uUw35dQ2kJw1wee/Hp5yEzhn
eCio9jKISEAE23ZZhfe88yf1NDCfvtxJaP/AiCWsKKFnN4oqBdwOi68Dbx4wM2mO2Vs8v7GkXl83
wYjsNAbWQhJrAw92H6psqN+N+1as2YNlWmL5pi+CR8VjoktftA5rtlLohvCWmECqk0vgAsEaS58H
uLtMYi6KafCWVF2Gh/uwP+k45w6pWvGbY1RrjLyvfPGKvlATcVsP4fjJEs128xEDEAWDIAlkD3rK
+r40bplYH9ETGraN0FLb4oSGs0UuAsGD2rFJK+nQYWx5s/89Z8R7ivHwNKAcLU028Bd01iBNb7na
VIBagp9rT4wMHuac+h0xgM7TOskP1fydS0sFRj//f2Z+MH0Ev+wcZgH3rNbmlwNJMPwCoaqRewCj
tNDC4bvwHzYn9J/IqFZfo4ohUuf0OC92SGPWKXvVEswCZ4uy51EXt6suMZFcqZ5UWlHewUrL5K3S
vErW4QDrQAy2EZ6d3EVPCOZKubohbjN7i8kOwXGEpUzm8jMXtcHz9/16VkQB09JoZw5KPNY11lua
ThLYFgw0lg0aE4e1D7LdqRtI2xSapcHvEkiDhB4HFyXuvKtMBwv9yu0xkJRjH8tR/MiHeXCF4LeS
LgIVjumntNeBDpVjYqAvOiy8ac9z9EGcFTlLwnesvyf190msOEKzaiofqO/4/HUGqGwYwgG+oU1h
jP5RiUJPNQ7lu8AL2hRjQYZjDbBj/umyNxaSXXWDE9C7X1lC2ZX65AYcZmdAVKfxI9QcyFdbckMi
Mzs++xju8ckcYEZjLTmpg3OuMutVrwIuUs4qsStI5eWjbFpzLtQeSXGXVCacHLnMAbqROn43wm8M
tnraDBORtpDKdbc9zfk/UZ0WypXRoU/UOL5chVFB/Lihrp/kN+ccXjYsm5ESzvk18LpnfpBPJE3R
AVgZ7k3NtxcBoEAtRhWcpH7TH5jvoEg65rHphDUxLEZE1tf/wXMOOe379aLqMs1fWqgfSuXQgxk/
4u8scOc3JhawFTxz4bQKL7Rj9RZ89ZoeaqK6q4BYv80AGbs+sH+3sWztJKhpMPlsHje/yAACC//u
rqzsa/h9SE36azQlSusxd6QKvPmK11Q/IqheXppxl7t0ZfxKxa2ApeLh7fWHJkAErA1AmN81MsEY
6LZSEBp9NnCa0wU9f+QJ8NX6RzZvtgeKEV2JdXEqXMHPZnaMV0nFQvX9NZHrv5rq8tZLoaLbTfX9
DRJ2MopvEoNEuWIHgOKaeXNvTsBkglyRA+88IADKZdIciasAMjLIn1zcjDpwG/dNhNFbiVR47GmB
y/O2fMIXcThPKna39lXapZbop5+438arVoORm6/UmAwm6K4QWx6ps4yiPS3/9wvHmsnjNgDnYuj5
en2AM6p5v62VnY1/Q4kNNJEF9wCj7Ry/q5Jj0l/ZlokSlqTuFfzEDwolnfI1Q53SduBd29lRzNqP
Lkx3hu1a4z3Qo7FvG1DskvtiitwStKohHExzPtWqSb9z80jxKt/Y/1Xke/dI0kcZfnMpUvRtx4ul
gAMFHfWjja8665LSc1p4StZzrubccZbmn9qMh1Isum5+8aP94SBNAOo19f4nGfwlsJ63BAbATnfW
Ufwg0NpY+Svz+SXG37Pw4mWHk1YyOnpeukX1hynPgPFwlcFindf2WXkjZrIo7muy81LgNf4EsxBJ
ZLRni2iomf8RXN3eVa3JeXrf10Da+D/VJyHl08fOaU8Srx8/qkTZVWJYmeLifxDKBj+3EEhdOCWa
rsUJ3wf5Co9jcgdHrh0hI+8lfwqxZhtkmQ6xjo8fAwqJci5DYsALzCAmf86IuqrLozz+rGTN3LmK
Ax0AQlZWPj13LS/7jf8ojOhhS+kx1hhm+wwFDPJsqlaKrv0u19KXO327TV2/JA7DKONWMCKsQAYa
e9AY8PDMSwlsUog8fhJGWMbBJw8cRQ0HQv2SgL+C2eeJEvpkZOgnyWCLf8i/Nr3XoIvBg8b8XrjV
GuD28QovNpXP576ix8hFmeWi4SyyYx+QeG8pA3Mpd8IAysC9QEIWV33kLVpyneWhJ7TeAM4pfTtL
1uBlvhAx1zaNw4T4W2F3dycgT9x+MQj8c7hIy9lGU4Vi0fJFzu4NUA8wmsYHdJzdaMkGRJbLCfER
A0ePiWpVO69P/4c0I5OxM72aeVRocaKZMj/vMQ+I3KbmA9aq90w7CmHhdLRVtOSZOe5EYqdTQJJZ
qMfIOeZfMwrR9TxcsPRRNV2HfFdABCGcSVIA4FANDLgsnRwEhu6vWWVEfLDniBnfkZMbrJY3cYI0
sOCY91TZj90SP1gn105J1v+aH/AOut0tr+Xve0X1RTFIJZilNcWvuk3uF0kKC627OVsu8ZPqC7/L
DPhy+kvpKuir5LjZLo8NKneG7Qn+2ndCoSPAc2oG8wIgjOkyQ3ihHofzY8dAHRDnt8cS7+/IrUJ/
uPaXWWUNjnhM+WixUPQiHuTAiOpxRwt7dv8SPZ00xgToyTuh8YnSwv4UEEptVDpowcFk7iwxDm7g
bkB8uB3d9/qv8RlytSQRYl4+xdFqXja8KxAu2Cm+Wgzi/BzfM061TU/F74CFC8kf3LL4WD/fQp8o
fZa03E/JeegSuFW3tVz9YIIK6RVyTPN9mhY82sdnVtD2SYFEczLjb7M95DXPMMx6hHPjPXDXqUMR
HrbQfbO7KX3MCH7LDkprLL0qonceWwJiq+l2jGM+gRuQCTGNJXaYKFukoajyLaCjo2xf6NUwc+DA
6LTVQDR7aV2aRCEdsNJJtAKat6uRA2WlrkxeaWEiX4OBJgCkFxajHvq5Jro2BSzhqjStgsE8OyRN
LvxtRCAZxcCcn45F7e9RQDu3SOoH5dMMJQt8TLi5q2gw8elAQKVBOIYD7IXWgJmgyYrCOTreKKG5
Le1RPiyHUF9Z05ZukBLC9YuIyaR7SztUuQl4n7OnhtAIYNipkgccq5ifRHoiv0x5N+JE0HSqVGXc
ykVDojNDrFjt3eU+/ui93kABBuMF+gX5u4c2e7dF3u/4EGi/ri+oHa50QQMiCJVoCt+uPB7Jd4S1
C2eVWZGP/6vP3P1idrkAy+7oB0H560yt61AjxA3lzbKHbR6AlZtAsCVkfF7/LskZqydlRlc9IOH8
Mx85J3lU+pdcdMxq6vzeyJoBriC2r8Q6e+ifOnkMCOU8KfDEVV1Ju+5rfdE0ORQ/1oZZv35XZtrP
yheFaCE3szV/FRBCoP6wAOCTHtjMscLm/HZDWpCqy3Xj+xbVXymLVcA87Bf7dzn/52kgNPt4Gr+w
HMqLJt6KHnTks1pv959IjcIpVnfiyGHmrhPGD9J8okn4N3H/Q53HFBu/JkFgqhOyOvijp4piF9QJ
36WqOqgovoxtI9jhcPr7Hq/nEdFnTtM/ssgsOrKJYXNP+mPCEJBiGRltz+fRFl2ItNiPHp8UuPiU
TiVjTbKSkUJ+FwoTrK8hdUJzryvhSFho7/4Uv7mUwcZpr8zHl28/hLFbR7x09Hl63fR+cytcnuRU
6PM41hCf6biHcY496/MxGZ9uHdB49ttOACLaFGLML8Pdil8cIa9kEjcz/6VDX2tH9POuxq9aV0o2
i3imiGYvGwLGCv6c+3XHRetTkvC2j00oHbUnn806dzoNZOjz733vkt/JatF6Zs2X3chaZw8xi+fN
rXSk9674r8W7cgu6vXWs5/bt12RV3PBLYUnthhzYZl+IA+wWCMBZ/MX3OzsXEO4Ph08qWpvw+Iuz
lqNa4KCXDL1gzGQ0DFO5Fza3/u/uvakccRZykj+set+aVbAY7uQPmIAPGOdVj/+SN+Fb6yk5n/qP
rpXFdLyyTQ+J24Uth1CgSJcIbqfuD2rWZuGI81afgKuK8+Cfx5ARB2emoAjUrOBF/iEP7jsSTCG6
zQHIr4ggaxo3kLEJlxsJKoRQKMjm208Su4gGq94zqemReidxmAOxOBX4NAQMX16pl0hOt1AubKNJ
0G/QDikt+hqS0MHGCo+isJ+ut9c+qM7INhbKmknN/Mmw5aHhUfv5Rm7zoRih0fkunQH1Wl4g5Nof
r1x+vvsdAYN0gmkQ76LEC4REAu3z5b9kYX8G1ekPCp9sdiiKhA8STy7RZrO0r0EmhDGD3U7gBRJk
7TE+7rD2/GMDZWAnhZMSd5MWuB34wPuho61A9iQPNkepGnIQZJPlthDg+vQtfIj0TuCpMWb0BMSs
jiAMG4hVNtTwU4oyj/9j4QLDI44Qu93snNn0otzJSX3JXaiadzCdR67LetSWNydobJ+YFoAM7+gC
Nu0R5kcaqZLFqILrTnBLtlB32BHBo3lttLrS5ZcIG4kf98Yl5zo2hwfBuYrgwIOY9FYOc/bNGs8h
Ju4R3aOjpP52sPvWGayt7BwRIOoRJ8V8svAJBua05Z6IeXrq4KBBBsOul8RfNyQp8Wq2ecjNhAnM
A5fTyWnELQRdg2EYT5m5zkTgU81dsYrcvQByHTXWoC3LvcxppgH+0bNBtXpXSXZDtf/MKUS6cWJu
eYJSYGwmQMcu1JJnyNFLsfeupdeaUf4SxEBopXolUGTJCiMeZbd+gx6UklVxhf7GR18u+6lG76TS
icVZ3yM63RkqyrVF+Anv4dmNJuEExflgL+/0phYVAGm3oCPci9IiOhX72E+TaRnFGGGd2o/amdL8
nXpzV+2IdzIQLgUxigJnxL1qyECxdIZDVuqxainYzv1m5wWjXkf9W1yHv7egdBegetFEo7UmVCJn
JryEQFHwhQeSUkgIXII7jiii+bh6yMQ+eZijXNbwLr+E3zAvL9WR4pSRylOfGCN/vRyV8qYD9x75
+S8kte0JQf6qL0W4RXt/dI96wUxLkocr37EKjhtr6PVtPkJvEJX52hs0lO4nIplCpepBK2Fgx3ss
7ZOuT3mkRmOcUhlHJBASFT+un8T69ZuLaAHQr+pr/7LS1/7eoZxZVbbUmwF6s/kuN5eZQ7SvaWkQ
V/yJ/3p0HB+fz8wjYaI/hGmdrkVJPcj4ZBGMklNdQjfltDI/mGt13R5lSjJTmeXM8B3xnb+RbiQ8
60JIM9DcR6mXrJx3h/3BpUxMhy2tQrijj97xsFVQWVjF5OcKnzWQ5iMx9H5RvV097pksAzzmJe5c
o8qE4Avjp1BBkG6nez5Sso8PQe10f0KEQGYeMMNLqgSkwIsvnlMhD9hCfJvGDTSTK5I9e4PgeQgz
v9F0iFUqZ1s5C6IWWBPa7Lbqs6D2HnL7+o7k6PS//FxZm8BumoqJP54VgEj103uK0JJr5tfV/7Qk
QnvHgPGE92amvPeL6ywBtw9rJsY6hrdnb2Ixzu6U5QRM5MA3qpc2RkFzA473YUwkDmQe5PTXT4rI
3Q35/554Vtq4qCKhKdOkk2oOIVTcJDqDYRBl+s+z+YXp7vvHo0ajXD2w0fKRJIOF9vDS4XxnC/n/
oopgbJmx8faSIcZ2acT0psKT6ZAPNql2Ugx7hJdQQAu1Pgdiux3WWaPICEa/lnNA4ONEeuTjMFd1
//1WGqVC36zFt52motKPA4FDInqUUkknlxmOn7HX66jyU2JzkVIJ/cUscAAVwmBKVwYSjkM6IVF0
2Pac93EFCzRJP1zuo4HSG+m7wvNNTbLl+DtPc8lRS4I3fjKQa3VtbVsqlNHBi9uC/zRpNSB/+GPQ
lLPNQPlJTgTZhgRK6NqeKtdBJdIsf3tU5gXFdh/OwljiCqM/oEXdSeOudXGmafQstONVYpzREQW/
s1v75+jHhC2E6bgUMsMYo4b2P3CjEStXJ6ODOZzDimdnmAjmVaBMpwIySHLrPjMNQbO4zCRz6uRy
Zpmbi8FOY1BmJxCc7U5iQqdVuoYldA0dzGVlcNB1LyIoAM/Qmlc9J9VY0VGeMBGvp2j53pSQSk8D
2NMPFy+Ce4NBK0l3HOkakrEJHlajFDB1Iv+YxrLWoWHDWwpjUvd/XFMD9iKpsCe3UA7WotIMJHoX
UwaCa6jS0LmIj610M1hCv8WCL2O3hDjWIh8tAGT9mm9tlMJORq85bOeh2FgOorXJNAV5qRteOA8U
t1ZDHZsAu+SLHVvbgCL8FEAVqoZHjGKEp1n8PWN0iS1+4zPc2ryfqjFKFoX517V/3o6Fxed7WJTg
mG6pZJoxct3N1LGJSjCz7B5Db12kenO1pFxhya7aNe63qYyIA/PBF+LG5GG6XvNVxA9yHle3mkDA
ZB8i3qcm0KasVOL0WcHkE+/tzT8gxqbWuLRQFOUztYMq+OTIuP+6zmczPGSKcwybCvWDc3DBy6MR
9hmCJWCrlqp7YxXcsluzmu6yHsdVDGQPM003Q1H9MP30/cLCfx+BRqaIu4WDIRpOmIWgUM7ENNKu
FKHEsGWV7g1umboYEIY1TZ4UV3myaH11BtTEp7IhVwRQ7JXEDI6KdrqCJzrDAsC0iVlMmFoX3iPT
QD72+1uucVR6rGMoKQF+KDnGUDIz2kLpZLJSDWtN8Bc0tSaPIltSjgFMJvwn413o3CNswk2TCvP3
/ZOLSz8MDaQZ8SiFto1eh7YaUNP2YN2+CrcQco8dd29Nf8CbU/4sQOT0lm1uBX6+/gu4HFyYSbgi
R5StqkSDUy7jFHbwoL1FyMX8WkhX3E2p7hPaPyjT15MyKZNuAPyHwcSiUs0sWs6q+uRpR4q8JlQe
mTeOfnXD8u+0xpvUTCnYyvkLxV1u3Morcd8X3j3o5C0cqNMIQab2wImIt+JZNqKRazmN1GwONMfY
6Lp0w7KFeXdZXh18rBbLRWILbx+YPSVqmUQA5FguHgjtp8bQyYscj32D73f8mEfxvjNDdxymotHc
fPJFTTu/IcE3vNPRNV9wFyCPzy7OPIpXwXnPmZyBMINfUYx5s0Esh6Z3Wz2Y4SnAZlHl2llHI3lQ
YpvfQNy4BHWLy+54ZcFZ/qy1e4Wk0xhC9ARG/KkN2IlhYjjcoDdxZGUBdDpSlrYTTe5POGbNWxjh
P9bCsusWiHg58xlmasEifMRO888xMpEoKgNsXlfbq5jJmG/KiSQwOS7Ki6QQSCglTiQIRG3Rdprv
hjImdjZc23tO9O3vQLLszJ/yG6d2rAtEiaRwZc6/9deSpqRV0bVYYd2TSN5bxf3VGl7xgZKkS4TZ
MYQ818RAll5MnqvxZw4/QVrsN2Yzk6AlDLP14mM/gw5cUfJIc+Pt5gG8zhw+Y9Rp0Wtz/WBHRVyO
uYVkEBn+oXcsjbq9NVxlRwijyB5xR+1Ak+C1Xs2pGIsfgY16m91hr3cyRH4Cv17rYIZpcdi25Skl
tq//e1GrtdLst3aMhyiS+LhP+Yh9cIMkzR0JbsuC2TBO6qVh4ZYoDRGzfiNZx++oMZKRRRQXIabL
abgbUyGrvLQNDUFcmuJR1oMPVw7qLVRTkMlibDJGHon8GTEnuxfAuwdnGIlKcb4XxzX+ZWr1YEuZ
yPPnYtbM0C1aNr22g+bs5OvTrfaRSSd9DrBPlz66l8KyDtDjHWYtz27ZnrB8d5bGZ4jZfX6p5mp7
Oz7ncLx/vUiGWfjPiOZorKiRSmq8rn+8Dz1hhNaFhhujOyHg/bGwcuOnv1L23uL2KYRwUtZ/z2aP
hCpvJR9UobebBudE38KXPG9cjQQKxuwRPFMbdv7wGooBfEe7hbovEGQrQadFBNTphZVmp2XFDABa
r8lKxvWxnoSX6O3N/w8ZUVJYuBp5i+Xa97GzDtvGj+vFR+xJpSdq7BnEPQ3VE6bB4mkHfuAYclwv
c6SCwgxGCXkB9ToqJPq0U6GzfRjNbJ5DkDfL2DJBO0f3MarlmD6UFsieMZ0/ca6S0X6mCTq0S2HB
Cc91CZut8Qa/zKo6u6sxNPxWUXdhY6GPz2SVZxfmoDnE4ZP79aSi7FtdSohhfm3HFgzGBSGneA90
P4VHVLhsYO0ft6KrIasxvXOcjMX+FT6hfrlVu4u+j7nEAW09cc70bc25wJNgeeQ5rXrCQYq3uHy6
K0u1e0KgbivUuwGVmGZNpwZ2jZ8OGIkAq1hBM8X/z8opsYP3aN9RLgwCWtq5PIabNwf1YmeGH5ak
/Vr7t1qrzIQ9wCwBG8MduxfCmUtdEpsrZaurqdkav1jEvCq10CkDBRNSo61IfrrUGMQ3c7RhDHWk
W5moIe8ZQNSsSlkdgOA2vZXheXY9j2wJF3MjlunHE+obsufMa8apzJbssmZBbEx0CYDjXua+MCjq
u9ew0uVB2sjfUjqFDdgaYJlm3GEQVKvGoHKlRo8XrHyH3ZFN06EaThwC6ix73HyM8plHWmJdFm6I
PqTN0kQFrnBjDmZk6wT942m34SHI6i52ssuS7rg6XGkMziod/Fy+qVwwPdUg2CHq7Ts/oTmgFIun
HLGaURvmjNaO0sVk3w4gPQEJn8FzMplF8q3UBg1e/zbT5evMTr8G+QvYn2rc9BaB8rzLXlLNPol4
+XY7u9C7BJmFhUlTwbOIfD/kE6RKPSsMBJKOuP3guVmjI4kwvoE6/bYmYzgXntuwvHcBFg+y0iXX
rc+bcvRp2gM/JweE47URJbCOsRmUcbc0cbUVpDdVvwbs/RGdW2i4PTFMLfteuqQCURfQ7WbFgeJg
PIKHPDNo7G1b+XK1sIyhUFfrH5yPGG+tCXmHFwzVwzsYbsEZmGCFsCxFQOWUy2bAHYk2YcnEmYEc
/sFCpak/vhGeqH0K3D3eSet4GDgrXd+SeaVZKBBNl91LHHC+iW8GG48BSVI8IvDOVBHh7yPPsagE
m+yjV0YtqQ6qeM4lhxFz+6rSg1nFHVTEnpizo3HwDygqvgR4nV38vnedD+LTaS9BHb0Sbv/sIsa/
JaISybgPN4Jp42nW6i/XUSVPr6wYPlxzM2iyljD31281dmBh77XQAbaPiTndHutAqOqgl9+hUaUn
tpB0Qu4VfG/vLGIv5wqR4ciFJR28Ekp2Vd5fd1VGSDOL7790T+SGyq+b6Wztcsg2m7+F4IUCsBx9
gThJWKycoHljEJ5qNmRS4qNvY3I4fCBp4OZScj3R5JPeiyCKByr8MeNTYAG9eldsdsfhm1rU2l5t
U366JRjo82rFyrqQqIdXRGN3LnYYxj8jGmTDJSKJ6PmK6yvb16sWzeHda5yid+HzVu9wdIugzbQl
V5GSjqF6gai/xQwP1Ai4HDvuFp+sjDmshUGiAJ0INx7aMlPmNqEJY3zh5fEpnE/tpzlQDPp6O0Bu
ihAQ6hH3WnM8ZM+QQ8C8Wr9bgVHO6ok6cJfuFEvHXCygs+hIrfE4pFDZxA/jvvdjGf/ajEa14tFC
Ga5f7a1hwlTfTRsDCN79TadLUbM9kpda2td9AqhV0oRSzIT0F6RN8TbZAczERGcoqcmZfFFiGQb3
eIHEDo+T45HxoPgHrkQOu+xWgOFjPsjlZ8DlxaBLhdT/9iwHtqsGoyxmRblZRtjakoQRCE0y3AAB
+cFA/IdTVhF4BP74sq4DgO5M303dSJCHttAKYNJ5tSl6YGnc9//w6zmWkcR13DWG4R9HyVl8KM8b
e2TEO7L8wim82t2rUs4CNdTJ3iq1SmnRHQgRU7wutiuTuKVk7DiyNdz0MQrT/5OY1epQ+nu5LJmq
MNvGg7VH/KkqXhRAz+SHizcwzIAF6YZpe8N/6Kn5n00zXN+VCTaqWZ2xT6cZRRi1d7X/kximemAe
UDeiiPARwqbHacP3ShAJH+EdF5TUbNyJBckXo28bt8xOVtZO0pDlG+AjjqtoSqofOae+lVFef8Nm
HszRsAX3i47QibMgi/QJJE7/EhdxkwgqrBSnzVvBuiC5/x0OdZlx+wAMbeIiFNuH08WI6F6n2ZQr
UX194oROAmlCCXIHBiEWjPuaKuslok/Ib32cbU73IYhOqaJz3Bj9kHhS2CW5W/ZG13iJvb3B9B2w
khsVyAbW8Kga5RuT2PB4d7CfsatPX3lxblewoVaTvuIGDfa6BbEfi4qiDLtiHppXz4EnbE71QuR7
xAa4a6eJj0XcNlnxl4Y+XMgCoezj95MOFTG0o6q1HkOF0G74m3DcUwOQEVMS5qwR4ZNEmgSbk7si
Ev5VEWe7M7Z7UrDnIvVNteXoWki0TKxzdXUheFDq3nq9zT2HvwvLHF/KmQcHxFniJjPqADPo4hzx
lPYrNDJtp+4/8mXm7WKz6mR2VdT51X9e9Is1+DRJv/lp4gGRnSta6V0UDJ2KO+5pKBhb2sGwFDE7
g/FbfAyAF5h7h0oyRecYALwXFTHACCacoXtBWtguReP6DBbRLvdR5AJ9w7TonJE73lh83M6LxYUJ
OrJYPTNDL3RTUtOGyjIBMAoQ91gt686PCBrBLnSBCavGab0jL0xKBulJaSA9VWWQJXr4WlKl5UzZ
KR6pEm9RtFSiL5IE0f1t4P5TRgWALeqiRcQYG8rMU5wGkG2wAdfWbUG+sP4vIObAGAyatfHp/B2V
PhQHlw9uwQsmdA3/pTuREXHRDtDHQN8+8+OgvPdEiq4UQ+lIt16AZauqLevF5hvJtSSDX4Jw9k+b
kUHLBmmksoq6P950yY1yQJOyz8pNTMrpD4PHOiFSFXUqzCduaxyFl/4YfEBMQpslfXW5fvsIjVm2
+8Q2s2eA0sSJX7rlJVcPaNk5pc+/75lGYV0urSk5mzcC7ho4RVlblfTw20dDCm5j4xW1xXfaV56X
Bm0DeB+cTDYAZvZeH7E1nJP4fxqCU81SfOOpZ56+4lL3eXnboWTwe5TGh1vvw9+b/7c9bTGGUXyk
t1DES8eIEw/+K3AcLswdDQ+HqmtrsRRtkgrz5QQH/X+spN2YLRF9OUfmCiVLsUD7cVvmVPE0xi/C
HhQAw4bcTPOvlaU4mvU6eQO0Cx7FVHTzSrvkJHBSS4Vo9z0Y5oQDCd6IwW0QnUIO/F+g2anC00lV
3KttYqFk9a77RiYa/GUUAVcx2qdm9trspACKxTwKd/O57yCYcazvL89pEHBu1sAb+++LF7QsFe08
dOdAuC+RF+2WhYdmRdRUmZkNEmll5g4IWoeGnjOt+8EaWeA98+r+jkYnz9Fjgzy4k490UxbHuZy+
AwkPnqNRIJkwYN5BzDuaVFIYpIe0iyQoEruERkwL2RtIlrdyENIXaPvFyQA02OG2wcs4VGcGJamb
Hhcc7CBGiGUu1hhCAf55UHrVjL9/CxDscH+KAS8vSa+lJjIoDh1MTQv1Za0THb7HaeBr+K++9vSP
la63HdsJMxlcSKZYnjoBkWQTmgIwqv2hCTJTyIhw1c89uTNh8B0NYWTmdvuZQmqzzBrznRJ6w8GC
wp4/CnDhXc39me9cEkeUqCWHX+Yuf5hGCr2bXtaewXPyqiH9Z29QzUewcOOeSUltt6jox+9CA6Lf
G9bSKGQ/rd17Eta6MitmiwN0goUxpOqs7bVx8nQqKFz2ym/pJU7RWsMa+QpWs2UMu+klY/OsBWgC
mWQ8BzIOSy5M5wmFx5ydxwesx3pYxxVSbTlq3v369qztMVJdc0jZtvGgJMpG9Ptu+2hFJUvGzpQQ
DSgBBu6FE8j7CX+7K/7UsXnuUcjj15DTD25/AoySOxrJJgn4XzU+Abg0muST49XvKVSrW16IBvi9
shWvCmOJ/+C/ql7/9llcx4JzVqU90mipTfFkccyGJbrXR3NoI6WzHB9n9Gd5mITpgK8lzp5zLYPc
HMXzanOcZsKGbnhlNYz/h6yK/IcNf6lj09yChHXzMgC+zdvex4uBu9IEa52VLNwY/y0on/Rnvgam
//fd2R/TQEQKW2/kdnjyo08zpey/8I2w8bMLfu9an02bBWkFb3ANbuAQsWXsTSuN+EwUKJTjcREk
jc3lpFSOaQe0mQC0ZruxgEqhGIPETb2RjC+E6dxKWRxjLBjYJtUd8PNf0C7MqTHNlx+dIx8y5nur
LiUNnMq5R55lfbynI3O6/9pTKZN8BJGjk4cVt1cwsbSH0lvsBvI3O6vL/2dneAhazurGN4BersSt
b81frVCdgqMPNtd+SfNHZkVIh8Ym0VlGXrjTtmLMqAdo9MkiUcNRgtrn5AR0R+QsS7IWLJTDuwuf
iMXS1rr7UIJH7W7qGAiuqICTWDmnVF16F0Zu5A6G0Nw9loyp8eKw/De7Fc/shgK/7b7e16JJVdkF
6RBbnQ/L5LRMo/Bn7Nm6b+jY0j/6Cqej0cl6yI4ODf6l/zZ3/nOMFRFYbrjIEQksWSskKXY+6a/O
9Cmv/i8wryELVldGRqRNQUK5ZeHJmaeaXOBSgP+z9qqe4+HXn/BVJCwJnxa86N8r0IX0iCc4ur9A
KIqQTNN2VnbHLsEnZxZ9pUFvc5uovoXYmPyZxuVnPoTyA4o89mhqx8G9qH1KJU4IQSKJeYx8co1+
SoCU6rMbuZX0J+votwBG/937dTR3BRS4ZgLiKLPPTSfGgMp+ICKE9m+adhZDPknG/td/IV426S+I
bXD9lCu8RteiixYiEUM37WtRtrz3Y3tBUbyDE6w2Oo7h+MkCgCB2KKLVHSR3FkroKi7s8Jc/xK75
2dFn1mbJbW9X65nyog19t+zqdBWrNPUWNg13r5SODlgCCbr+GPZflFyG7urt3iAyxKS7kstpmlAT
obBw6JRoH+kPutEoMIJvct4aevkgYj1ltWostogLEZb2UrX1l4MR0mzYtbVmaqzx6JEppfG0h6+U
3WX1IsASW2CyLwq8GW89HmKw8u5mMWUNUrLr1ZAG662EnJ6wuRri0RpnKvrb6+Xdhn7jrvBs80Uo
olWqU2jZv8O2NXu7Td9yiOsddRriWV62DzI6/QGqIwkzbqFHFQXJzYJ6PO9WetVwpSQLBL9/YNS6
+Zq89sikrL5LZHeBtq/Hxmc7yMJUEp7sqAciy76zefy9Yv02dNFAQmMl4yLR6IEYbUoLCoGPWRqO
KwLCkjlqcGx5qXFWz+E2KFL5thqHqpZ7NtXoSnFEtNNReXw+jfL5fxh2aJ4p4rNqGrrvPX+dwaZT
N5Wb8WsI2++UB4iWwnxJVLtQFVOwFdG6bSp+Ja1w1Ts7MBuXed9Rx4LF+K3qS01Kas3mNQNYeYPl
dqxiNwoQY5lB7+IxUYNG3ss7e7MF1l9BUg0BRzaLQY0Hxb+Wh2WcXIJysuyunYNvLi1tZvwuzt/l
ajVr7HUL2q1r5UX9a1xdL+TRxRfDfaYix1jsmOpDeJmcN6y//Oo91t6VRmCzloMeAUMz+CjWMR6d
pZj2Gp9XeGjCRZ+aQoFmplKDqGflYHv8ySXIILBy/UUEBCohyR8LGgV9YOROEic+WltuhbGA5kQp
SVV3/mL3ldi+T0xfOD/Vd8l32j/jyix6DQ79tviqs0tG2hMUOCWpVHkspKQvfDdFFZjJOAVxCayP
Mt1DAilqq/UeMAJ6QVt3HFbb9I/SqPC4aViGfc+GE78E6qYBfYPjsouUD3P0sjJnfTAdZMi6ZrZ4
/neYjlqEl/7hHmxb34PVG19PSt9bcmsq5PeEKvmYBGrA7lEAHuZQN+FtxGDJLxV6ZqSazGgNtvfE
/z6iiM9lpMqb0UpN9X+YH2SsfaMtXdbpUP56m4eivuG2Fdm8uNK5VaOXynwExQrwNoZX8l2ew++P
mtkvkmepXpCI9Z4iHJm05Pd/536DMiNd9fOJEBQ4o4rMSL3TWx5d2OgeGLd2OT80W3vZ6hcT3TNj
u36j+Z+/Ud2lvVo9PTSuSK1gdf1SpzUff64keOEOSo837S9lc/62idIL4PfezHi983sgQPmn5+yM
Ne1GM4T5SKo9kr4mQlfj1d6NdiGt46a1HdPvcu7TH9Yj4cr3uMNl2EExjzMq9lqNp4UqFwwk4E2J
42hLJUSL8g99rus/pw/IpPODFzTgFeu3O8NOgjaQsPQqmL8zvW5SeFRJxhPJf5EwZeqL/dwNXi+R
TXnyPTkUFIVJOhN8LgrfMRsJ7SmztrmK9hubWoHxyGomTw0c5U4qhErgIogBqpzAVPiz8o0KEVWF
34XM2yCpPuElOAbAQtTpmnU0g70DDZP9JG3r6ETgBoaV8WwwcsvgrUQHRLcWJncSubZDR6uASCbO
KE+zefEOQ7KqbqJ3PQO1XH3kUocvF6+MaPgZTCHbynDLu5iwkG7SWBEHRQwevRfPmO5BKqSyspWP
/9MW9fuwTTEc74REaOFZSfxTgqttoDPjrh9Mb7PMi2LJaI8xeVwJRO8bMMm4OHsKd9myN8VVPvHO
bXXD5Mh7CJI4eYHTExGICXQ6Vr4SjSEmkORHh5x2eT6r4U6uEnWyKojfJs8GIfOpFw1HocEgC+TR
r0DD38fwpB4+5qVDe9oVbbMu3GCFS8URuQmQIquNXrMF80dR0X+UZ5YvxRTbTH0PWV2BmBmej8T7
3NALIkVJH1KaY+BcvpUMijcaOKc+uENQ0c+KN3EfN2CFrquLhqSRDkTcl9/RzEZml8jWRl8/hO8x
bvJ3z0eiULbzM7aRfpYhFncgXRdvXJUelEWCuV0QlY8HsC6Xi7GpSjoifdQKsvx3d5pOFiYIdu2Y
XbFnbsM6Mw0MfCHrlO4CPEF14iwx54olDs6yxFtKnKuwUIrmuW6IAA+tLj7xrMGFv9motdnbMF4y
WJqIwSSrwbqqXAoD4dBNZvDIBs/vDdBqgYE5RST2CbgXptYmEkhatD6n9XNfZ0fxjVU5k3D6Lpcf
H4TD+nWAP76cODUYPOz/yM0j/+5PwnCQvbSLNjTUklseg3QaHnRbU2Zu1hM9wkmAFNgQCpZKIceC
10gnJCl1ym30popJeFvyoDQJUVdgoE8VFUMQKBbWyq2k297TCyfWgraS6cqudBHIYvcwSzzxNhDd
Xw37O4EEtia5T2TCrT5n7NrGO24OiWRHvfRUGo6WFGsEIegNqGXToZqMP0aU5UXv8yDSjDG+Jnv6
EwA5flmT8E6GYZP1+XO5MgPAlIhNwer/BH4VQC2eJBwIXjWJMT0Vnz8S2vSnZR5DArjqmo57D44d
9wfNUvQwb3qs+SyjiLkEhBu3LJMG1BrhSgSI5z0qWSTGML/ww2GksXP7Bjq0pUh8nTUVQTFz5SLR
Sv/JCpBBzD71OJWa1SDN7kR6GQQrf9qI1D9ru3Z7ZyCB2PUquPj8gkjjiLMmR5j+o9MVHYML7Rmh
bFeRheyDadUniB8fjb/k/mzeiW5Rw+y5K1Ym/e6SP7aloT9CgrTVwb86W7NsrY+zdd9K95IO6XnM
sgh/4ctpct4DWibHQtVlqSANcqAj3ILRX65gePDnKf7INlrQTBTu4cxKXUybbf6K7UCASlr5JPnN
amwBM/hBRmxR3wPl2hmgn6aaT0lxuXR1jO1SoTVy3QkXdiUQxlM6UmeyZf9Q2T8DRGdv8fiDTnO9
s6vEzIzIp1GGEPezDu5gw0H5OdicyfSNVLeWNL1107UrRjyTIIaohBqbCE6VR7UlHyvb4VfLrMhQ
8jJl3N4GL28biDsRhEESJmff/XlgJUk5yBlwwIAHn23weBTqic/9OFB03dw5/4jiZryd16CNFd0I
eT3/3huyP7twTX7RfpVTmrr1gqx+X28PChSH7sUCg0T1JDf7eXNToBGY8Qu8KXWtRg/IhZx+efQH
WVf9Eijltm0CMHxn/PfiUlmqvBdRnZvTY2QvtWzBoQW3qY3mLCxK1GUudW3Tpn7iifkP7Ajnqji7
xQWIaco2EBAked8m5bPSe+WANdrnEJcQfsMue0pYu3vlnPHxdVML4u62NpgudEEmfNMMeIy30Os5
uRMjQPEWt1aesfAiNWqOk1g3VAPW41tlkSfj7jlXNx6qcKYPwwFEggl8EUH4Hcz4iNYe2YzntTvO
nF6nk6ySB6osqVUzFhSxOb1is4i5GFw9RHUpH6h5DragYP44n7B398PZ27Si7oC0kjHAHd1NTYuO
wfQRInj06uL/V1DVf3LRug51WHMAjuA3Hg9vzT5FKsrUfMsTPTzbmmSxD7/EqzY0apGuUQ4FMLL8
WlhpBj/dnE/ZAt+Pzaesj2n4HLTeeDNzgh0ExCyIa85wOq0oUT8OT4IxUKh1tHxE0blHOcw1NaDg
zfT/43LeuehhWYsAsvfyCcz9pcC+AseiTPsGThmZua1WSx73GloFQTmeraajGZ6eEqDrzz7u2UmD
385ce08thR3LUclAssVWovpi3MGawaA27kdgYWctdbydHWGJw4KXMcfztGYCnHC909hJO0l4YtbB
7y3ASJZ/8NGwLirucAhTgIYOudcIYDG6qwn5iswMdIo5bWDmRP/1LNYLzuwM0Uu91lLr0sog/Pbo
2e5tJeYW1IdGpAybtddSBkJ+uhMwYDg7o9CKfpDC9vCIoux9WkhECiYqXP80I52S4XK8+pUXZCkY
V1mUMHgB94Qlab0BsgNIoev3rv5BnRjlHDY1PR+PVaJ4T/aUKutpy8kOmu+8CWVVXWYNlsk87rxF
xMo2ZYoYdrS7nqP75pHb3wjSi/gkKrZsU3JAy8J6UGA8rybLT1GQ/ypcXZR+kYD3tRg5k7x5F9aI
LoBUOpwbAkzPc9RCUjhAXEcP5Ud9vixNlGk/8IZWb2XqlrpTBiXNZwDpjM5/bBDQCAdz3PRD95SC
mhbnLEcYGBd8HCatQgtGd3tvWIZZRyqy5jI+X+yjyi0gA2PMf7c1HjFVdbFHOcaXgQE2hT/pp2sC
96SYrlJwERlOgFv6dk6++jFPS3/rloPMrY6Zyx969ehA7CVv97n2ri4EFChVzZ1Y30yIA19+69mi
EkBCP63lUQYfGp+yY6R68KL5TVyXWUsod3IxTshmgvwKFTi2vU+HkbTBdIGRh5Sslx6m5vBfjIwA
46X7ud+h8UQFZczND4YUb8vCjGajAYyQkiudt/swdA8bD7+Qm4NOitFoIJQ5O6AFb7/8fAd5jj/R
y4FshpBvPcrd33MyVxYtI3gmruK/5AFaj6Y6q+Wa/ro4UHxMZE9ybvfGihYxs2p3EdtH6KqlX3eB
SbDiQznyG0xT/AFCHjTNIIH2xCzYTrKo+56YzOP0BiY6eYNtLFMH3NQL6swuCY8uMkHVn2cehVvq
6jiWyOIY3D+M/c9A+QA5+sw11BTGCIWy29ddpWfAnDBfONJB9z6Pl7McYbh18hJdPxiw1T14lxXw
uhFh43PScbAAI6IE1qetmvO2gPrN8erAYVveaJ33LNxM7t/X1YpJsthCMQ9/DU6le7GRT5bpGj+Y
TRRyLy6Ymd/H4O4piVo/DtA91YrkJUa2lbRcae5I3hadEoRc9CL5tDO2a6cnVkraRqcdrUIAl7d4
oZzRv//VB6p9yNmwTbChQkZ+EoDjkBrq0pwXqYfDWCHkD7j8VgRdeTpy2NS1Z2CAFPc75A9nyjJT
5hb5ZESdraN01k44zpKR9oivG4ycAgatukyWowV2aYSUbism21KFuL2Wl1jN8KbzcJSkn0w7Izjh
nREMpK+Z1itwNqFcgbtCu16b82crRgBLPIXMv9oD/I4zD/sqD2zsAWtFRVtiVzInVrTJoNcJ7RQ3
ToDdHwafecoUIQzIfyShpj0aJ6XZG3tQlrRLsz3jrrt8BDQE6j0Xo4r0+jtbKWx6lR3oo06YYC7J
Q92Jl+JHrBT/cv+JH7D4kVXD0+Iqa20vXAVxb2vLrgpvK9haNpiSd4kMNE0gPnWoD35lh+ariAJR
JmrMSyyTMJDVnca96qMSpdZL8wzlzn0lGX1VkLZAAQ9FW5mTScQn+56J9USiZ8DwHh5uCtLqDhxc
ZyurR+usAv/k/FDnS0/TiHs5BPQ0eWEQ3dLb4B9Xq/gAlUd6K5zEA68xZ8XTLsB91y2lP3p0bQFZ
PajLnmFBgKvBdbPPdwjDwIPjl8Tq0qqYcrGKRnk/Qo+ogWEmZFiw/g4TFY5F8Im8qplp0DwDqZmD
sS+W45PuUQluJgQALBAD7sJWYb8awPOvBWeyCPgvbtj0djQ6dNXtLHgfZR6xDlohSs69LR9uSzMq
7qTL1QUA5vSAmeoJo9ayEF36ySrqFNjWbPeZT/hGB/4iQWrrQgtztephQIo2/Zl/S0w2ZxZDFTiW
xnzKRiLE5nA6CZs1S+JmFC3QuQIwZOfY1wbFt8Cp0M0wpQeI1v4E2OrJz5jDjqqzyqx21mzc6Y0y
T/KiIEVfTFNfgWWGg2ONVPqV2+29ZILPZueA6tzVSiAe51/1NN7sizmC0alehtTzWTpL7H5drtoy
o1a8bINafXFB6NsB+69xc5Dj3p7mriS6PyxGvY+M6mkQSZn6sJNP4yh0O5YJ4mzfambg0IywlsRJ
hx6RDONloW17ARJnqr+BHFhRE6pe4AXOW8OyM/Xr1T+RlmZSCMn+JcwHJ3bQHpsreTormD2Ktncf
Sjt5dN1FzEAqJmZTxw4sEuU/p2xS92lureEpzC5OzEDTMs2sEdYdTXHaKSp9pd1ub7rdMgBayGuE
k8MwlVMyy6oIWj/9xmoj8cgtnI8RsKNl3avmjgT3FgyQcppV1EnJhy0dqH79qzXZk1AjYv6An16q
PBn0y9ksHyqwkfrXauKDJrXu9HGQwdrgxKwblRV3Pdyd+ecrR/gbdNKXq0aoRx19a24ctNXySJX6
w3yVwHx2bkclHhY4/2xbHfzejdtgA+mpzQULbF24tlrWKGx0T6azROKZZ0T1nksP8XiA+9Iun5B7
mVw2tGhtRldOnsZrR1zAGdbMp2w8PfeheEMf5uEwP5zqxuu9CW+k1VYspxvwPw1Xv20HgNPCRrTr
DFnybvIbhO7ND3Z7E7YBk3FRNKx6FHhneRxUvSQDmNGpynPaHAdD7gwxWCsWQTz/NqX5bmLsrKrB
mgGVuQY39K/1ao35JofjH9hMsZnIo3+yAizy0NvfeLUKq38s4GPMyvfRhHRU8Sbr7wkChUH6UJGa
plIKcBLkZZqxfvHXTeLmfub+Mtin1ilfCuKrtEOQIqSYf2Gd1WvYG9nJiNSd3LHy3FLrCd19mrll
RqiqxOypg0MArBP8X9Os6cwN+ieB4hMdGTXhVbizS0B1HZXUgZ/P56GZcMdKrs55R0R72i38w8a1
CXbnZBDN8KpQ7J0y0qvIf0QLaSlWvtRHxZY6RUQmIEr4ebXcEJDUbtqq8yB11ZF2ENLKbtF5k4we
pVOaLMRt8+/L2JGEtSFbXcml3Bbo2rnykeUslsDDFWic3tPXx5bpa+2vQJ9haSyCGwAZBSjkEQJ4
hKN2qFkLsU3BVF5FwKrJlP1dDRPyMBKMh7fKQycellLnJ8YbCoEN0ax7r07zKbrMP5jAvDe88BhP
3CjTgQiF1wH/XxrL/S82VeIEgRST/tTbCYzHFJf5If8WVKouC4N7jtjxVM27zg1kzy6deN0yt5Hx
5pMwXdp4XMH7tALixLnYxQhAjoSmdMeCxHl6+kYqZJ15kal0QiZqLiAFy7txH9IldaHNNHl8BkAC
GwRtev23JcVBPirKJ5nFGbPC5j1dRbkJJBLjg/eZ3JaxKR5hJFNIH7FNZ/OXB1fZ9WxYIEjRUmff
AQcmVEHUwzY4JwsKMJpe31f2jFg1pheOsNb+vt4edMPPJmwJI5AqY1kktc/h1udgF0WOaeNZfMBM
9YQ5jXuMvPqwMr9hJD1oS/ZteWw80A6d0Ct5yjqkn7qO+jsfD0gvMCYWehk2zVIokVeEeQqBAV7f
refqZEbK9DCReERsVSDNGZdV8WN6QKYUHaFwnuTnv1jOqprLD1CcDxDYqnLcSEsgewB748MCeA90
QcuuLHiVruM5dQUyPVMXF1Lhl1t5XtM/LFuGXA5/fEHfs6BCYvgehpPD8a6aBHAjUSMVwkF+nUud
BFElaL73kX3yzyH1O0Kk2gxEJR0w8iZ6txjY4BAeOxhxLW22ErluJbrLy4Ek58gJUlTPPoW8kqXt
AoQiKAQfw5oPl1P6CTY1zHq86tevlLsoWsUgwUzOfdpJL5qNyZ+LNI4GXWtebbiCRKfxZjDQeY9s
1bSK9iSIWOddWP9mYI7eASGd3t5neEakkSrOP0e6jqqk2RQo59zFqOOvU2N7l07Usn+Bz213zm+P
cps5RuSjof0oCJMdCaxUNsgTqj9dIhFDAW3lSECZ2FLXWLvo2hT88PPMRsuqzzXMxoBWzbLdXmjv
AqYgQIDiaMIiAXxAFJGbn9HPBNkzPr7hC4nKfGIqRvfunc66MyAmu4jxK/o3FNNFEkrWV6U+6oSB
gVyiO7Fda3lKWeMTjSJmj/O2iLXcx27dnVLevmex/Wk9a11cqehgxXrAfbkLVzq8rb+U2/Mpdwbp
Gxk+GSnrq8suWqM8jHOo1r7X+JBQgbFoQ6oyuxHaqriqUL3l6XrFWGWKswfqjy/ftKrGao/SBCnd
P6fGFydzcNzrfNpYLfofJkpynC67iamwmyF1ZKrBJW0jAI2NjRmeKj6BMT/BubdFR0W072cF635u
pbWPugYi+CKOW/LV5t7ruMUEQ3EC0JJfdnDolMd/e4z0YVP15GKIr4JumF14Dj7y5qDv90tU8HRn
L1rOQFVtTtsy9Igtnw+tTus81lEwEym3mH6j5DUH5PCv/Fl7HGegybWdwSdbvLH+QHxAWT2ybRnT
qBCommXOinZ7/xG8j6jWA7wthtR/I1AsZvvS1H6qHET+q0BTjvNvspuZpKBZ50k5xuMx6LzcBMY8
hW87QjWNbvXbmGymq4FvqJhzwkWtMgsIQL74cntHBAxY2Bamu/eeHR4MgC9q9u1HqZnAMtzmfrtU
JnBTu9fUzRBAF0XeyNAVqAYOJ8/lE7JJNDHDenUNQ2mNO0w/ReavQw0Db4NjCjuAKaxjeQlilFqg
btCe2SV5yKYb+V43m1q6FOXmDSR5bq5X91pbI/SFAoduiOw5KHaWEN4m11xSS1J8w7JeMwT1Bdtc
01YrSsg+vdNz9MAWOrVs3qN6MRK0IM20erhSqTzPWEcZxxIeCbGIHrWU4a6nyVFqA/N2PWU+uO+Z
vD5sQxiHEO6FZVsPIdRGHIE0S3LKaOYxFq+bzVfh3RjeUCFUHqvjR/2+7V2jegdjuk9HL+yJygoY
78utCclhjyquQ12ugULGCTV+aY5apzB0zwdI5HncVK0QpDsuBwxyFX1rF1v9Zme81G6/2J2ARovA
fkQxJBySQbzUdE/7mM20030XT7meYbNp1AQ9pZqFyxx6GbaZ0NvAIgMaHuIbmPGgsqVio5UaCWQF
gTwSjeI3Eez3j+M/fS56GAsIT8Bx4XslFbb5w8mxZQyUYTx7SBfVsMZhKmjtO3HOLLs0WUtYH8gK
gi9APbyjujvmPXsJr29Qf6vHHlWfzsEiIAD45sHURJ1nqw9eqEKWjuDeLpEFIB4QMQPB+kh2YCG4
UrjNBZuR/JkYCsrMZYYSwqpqnZG+5O6aLeXoEHEd2htlyWwYHlP5kw6cYj9FH70app61e+ONMfy3
5eXEBTg9V04P4YN136Ebm4385F9GfyxRMBHY4uyit956C0tYJ8CDNgGsV1qFdJoKbqyU+UTEc4rE
RbyBduRDPEtw/ni3cVgsNj/FoCFR+tH3P80q5q5fLV+sKbJttR2OBfYazT1J84ocvyMHXbuK54gB
7SkgqUTj5DsP592eeB1gWBIX/zMlmJBys9r11XzjxFTorUfZIJrFbVq+Z52zCOdiXG8J6H1uG6HQ
+hfeaF6oeU5Oc0CSa14KxPEdnAbAtHghJgrjDQXLzl9UZNSH7USpx4sPhnpJo+E4dQ9be2AaHwUl
2x9V7aJ9dW00NxNPBt2urc06/4Ae7QdzJWgOO1sjiPGzulEfrSbNNcOKjYHx+3Mgf61GUMjP1FyN
zUvMZlwTEqscOlKZeVobcA1aKHib90qhf4F/4rFoC91HEXo9UwbUQKLSUtBN5eb4NpnwHZMkHLEh
cNbS21nTSOfB4TLbnpCXH0jjzoZ+AjkbEQOT67T/LJ9ph7m2cGErDdvL8iVZCLwHwhOluL1VF9Bz
LxPRZpaJzOba2EjhTwDt4PCCbfNnEDM/hIwLL3+V6+xrybWlwUHclFFPJg2ugOAGUDxGz3us78HT
1S2TAG6kczNRugcLBwtBdwuDGETmMl0JB/AYI4ZozXlNr+qq/5tBgbahGBkv1szBmd/FUsV7eFyK
Ccl1W3l5aBAWPd0ux4htu1Ch45lbNBgVH5iqgZcFom6m4JD3BAkSDcIenPuioy8vVRA3bXpRoiRM
f6r7U0GkwvYunxk/XRyfpzNsN2aeh6BLn4+KQ5Yidp2fucSh4xI/06V3OxQaDwIgDgZ6rk/bKQhf
eHSmL+ShpPE+xFRv2X74Y84ZFvCKxqLjD/u1vDDOSffWaPMUCLkPrGqi1eV3BaiTSAD2zl11gidO
gMB9RjYMigT0TAfTCb05PgRF8Gjc4kpNIUf4/iIV5qrUFwcs6+UJEkPpHgHmvfFPH5P7iqQgcCf3
wnXB1fe5ktK88TS9py5CiBcFXxKVpVthd6VR0cbVqqM3E2qDXBlwU3C7OPD9h2YDWP3ULUKtlteX
cad2YuS6leM2p7hiKHqiDcav1ZOzG0trBM5e4wNXY+VVFatPVW3nL3PMx1w5FTcomIoFeI6I/nLB
9tXqBD+mC0GcF02NoJA132zmvjG6Uh2fXQsf4A04Zdb/Qv9tWyeZN8Tt7WiJ4pPJZOlYkoPviHje
yiIaR0RPdniAJ7IUoA19cLiVZEAYa1T7/ZFM6LlQd40AjPq/Qq1x0n1hiqHvzWzqQ++55c9L/IKe
0ioiWyfEY1yr9GPdn1f+IPJiI+6gGq/uKE8Aemzm1mj0IEUWJ8MJWkxa0Dt3LnKetHGZCNRUaF9H
qPKb+5G3K2zzCHAvK+oGcACgTGVBmv5c1wtid+m3QKSuvCTfbJCj+xAB60lctFqhs5ZWSPqn4gxp
NMssekohTq9tPKa2Tm3c/ZYaEiLHFmWWV5LthMpdRXESl/gxQ3UqajQCeZyMHYfzOV/mtvXc4oZj
dp/P5B+jzueDkWU/kyCdpFgQxdacCUMWFzI3VKqKCky3Obpp/Ddga3jFgdXAqiLpUCpcE6yAfbTl
kop16Hdu5wkX+84ISF+O/KgZA2cpn/2NDd6+eGaFP/Ilk6ARqxykja9YYC0GixnpAKukM9/7ir4P
fBjHvwXaaGQalli2cgxFMkqTWBuOBzbhG8/XszQ+7PskK2mBp4q3rwJ+zdXzXmTBmFi4zbS3Et2x
iyO5mYwCnTNRh2cexSIzrN9BHVxxaxfmnScg0wLHSLsahRiCkkuFjJ9bQ0eTM1UQUFMYLGF/9k6S
GhAvD6BhmhBg7GtnofV0y29R/KTcDQtC4VZJUheuNDZDFmQIIAgECIq2AjQEgXU+gJZduH6EtiKu
XVtwJSIRZ0H/v/ZbDqNlH3e8eXjH8wDs7cj9Gm5T+SJZYLQt5+L1FG1qpLCsbeaU+2Jwe16q9aZO
VLqiM5N+vqwOiyp6DI8dNs57MP32JlLGvba9cKxnppk68O3Rp88T32GpoKAoIXRr22IuELJLluy1
gIyftLGvaLzVfUPS7UWuoVGq/h2FGMpmNvXWlay1jfAYp0nCQE9mEpgcPbUmnYkunum8MmBz2rbj
NZXtov8zZjmx5KGuvB+w8kuqJ0qmYxjV/6WhiLfpKhvU62BTRaasqh9eRGn2TDnncgyF07TZKmrb
yF7VOIpVDdSZ6loKd5nLx1KD3SWVY+ltjpClOqXWcwwuRq+m9FGCYKkFPjOkYa7GRtTrT1isu+Ow
tYbtuSMcNd1DaznbhCQq0Fnm+v8KxeazG5Di2x9XecmqVCs2TjzkPLSrD7//cigyDzUSgm3y4lqG
5AzG9tDUb8deB1+hc5ILYJKESBYrtS+3G7C0kWnIoLazlYVb2T96hSQ4WK+MPY8hUOTaAsbyFk1S
ivSmG7FVbXHYcix2gYdgpDjJNGX5JpHHgxO6+uDHZI8rhAw4pit8SfWDSftnPVmPTOXKkGll8LVb
AIF8Ts08YvA4uxWTbUZRKUoQQEKa0SRh4hIoNMl8ggAqnKQ4iis2aQtOGO5gREBEzZTO97TyzWPv
j5BCmClluCT8V5xvufc0UAmOveGPWsq0OlT9MLPfaYRuw8npo4Dc5yglQKI4guO4ucI1WV2AzeaV
gsBRHcg+zXxZt6pdBb8d+913GgGvBMV8HXKCUOiGqo99FTm37ZfRs7c8LUzWLojzFwsXoUDG/cWm
g2Lmaero4sorzW+cOdx/33iDOr86nRZgIrQ+mS8JtXW82p1FQP2I9iFmrnIABj0I1+SOZmcpeKDy
MxDRWUjuM2ecS09c959haM3LTUUK6Txl3qkdhXYUSzwbK3BLWDriE3ZOiLciMhjJZLKlT3YJJup8
FNxTeqkYjz23+P8ggGNML4Y7/DAsVCoDhcfyRGXGcwudMM2CUwWqhdZbdqh335Lq4nKXBL9bfr3V
SOrZwqF8KwzVO4pNwBuxzbzxM/q8RqqYXxyeWbU/i7b7gsks2hbqeDw9Ca+7YTqSX9nzlREzaVyz
b60580VcHMknzJi4PH7F5TCkqafSL/NaJiyjovpCmnWSiOnMEE2yS6adZn1fi9bRaMqJFJrsQd3N
4VksXFGVjnHJnAZ3jKzD6mAbYp/KcO5LtJ3AJzJAq6epaUkx6OxsF/SHqDASxJwENaNU/zJvo2BP
8f4xOEv7DX4pUw6hXVNKj9j990p4cFyxLmanvOVbpl8pr59sgzoCCciOnOqryAvuYBoWkN0PJDWZ
yuURcFzaad67AOuEcqU8BEkgvYlt30FQoYmYXn9cTboeiMUw+85UXQrKu96lXs4h21uvRWo6wTQm
F315kRI4sHRkkOA6plFKs+Xjvx/BMJ3CFC5QOnoAUjEBepewYvUToLHpmZP3DeZ/9Ohegf/VMiDR
6Hhhw11hTS0LHn4Curwj6Z46bAnmZqoUivw79adNJaj8w4Tn0BqH62y/kJFa34uSD/zkgDUa9k7p
WcWPcw//TFHu01yOCPhM5dAQFQFd+Zt3bJkwNaxLqfSCvPveA2margeIvfp+nOecouvIhQTQ22Ut
AIuuGZQITAYmBL4yeCKUP9+juIvkTuHsbF0pjdsaJOcy849SZK3wsIUpbEQGmWf4r2XKzIHBGUXT
C29ubpHqOe4wz6qSOvAjBsImMk95WpLX4QD1GoMqR/DOMmY72449GOCh8nULYw/yxJhhiwzSd94c
m2/6gua4j3GElMkk+t5HTQxIW4P0bVvvypBHUEDVXR3ImcynCoS7IKmlllgrwG7Y+EClEuN0FdX6
VK+pf/mIMf1ByRC67QoBdW3TU5NdUB+DX5d8wCf2gLwfhHCIqWYKyTt5v1eQbO9UmOk3F0bHJWpu
x44U04+Srcb5bY22kPrmm9EoxAHjGxma2OUyKb7v63LXQ6ygu4abM0Y90gEXIzsVNWDRHcmLqw0W
apz1zh2XlzqSChfjCKSsspvHvv0y5ZvRjfP0/7PjocAeQXJdO7rM0NinlD0XME2PskJtFnpfTIup
18cJsaZzEC64bsdgvIeVtqkS/d06wHFV0sgi+VSWQOtBAD0FGA7Gzc06WojcPltnfd8e48ssTFGB
vv0LpV2mG1y60fbJhGB/qZkcaPwb8gpWDK5+97GIv2NKWJhp0YiLKdZhno0q7MbHws/T9H2m3Bau
mCeI7CCWYVCGTWpllJ/JpajvF6Ize2L6JQFFkbPtoSGNydmIpih+RDzXsMrMZFHmtpC+XUVM+YWD
TxtI0ZX8ISOwAh8Z9LwLwTD9BfmRt0vwnIfQM9r2Iv2exsgtS5RRxIS5SBKxHfn+2ChAkj6fk5io
H0G7AmPRE48/fRqdE3Su0qsLKUcVfI6UtbhOtjt7wDNSNppHBxYzYJpjc1BTmByECB7J8pEFuLC9
h6cnt8CZ69GhOMa4IlmaEMKHmZ6dtb3V4SKZ02SciatDLCfJ/oHX1uXNd6olKqhYZezvzM16efxi
5ttezXoa95aWzL8xr4Du8PU+NTgpIV9Ll08pgBVf3pJ+T+7kx72JnkGBqqTfNrbne+umEp69v9N7
uYxqTjvloIDItbEtcBbHBtgcQVeLXXehwTKuO6mnoP7jTUOqY8BEG/B47BiS9dMrO9SCQxegjdap
kbv7num1vHqjWPl1CgjHL8DiV+FgeV4GlOJcX+Y7F+Mt5qHwoqD2Y4NX6MkJPnSp/ym+tz56WkmR
qUJWhtb8oQdc4uS5NNS4xREa5YK+6SfBv6iQIKdv7Tah4yL33CXCxdUIJeg2wYJgBMnJZ+VT6Pm7
9aHoqOb9V8P9pkohCpWx2OvLv6NyWIElMgBxCXSeXblGtKs1t+agfA+UqfIHKdZl82gTTJIZfskc
TIVurdOqOw7y8bnCUbo3TuWT2PwNznzRHtduUxBBMprIk/UfMVEOQVOApp0ZpqHjlQbkrQRhsOn7
JIpRbYmj0fVcv41ZY/Jlw3SJ1aQJO/LfvS/r7Opg89Wilcu5Ha5MmUQ5bQGAQaOH+1PFZScc5kps
3iS5PaC5fw6nChNKw56GLnDjMnUN/k5qot5ZqIciKFRiP7t3I+GTv5WqnyDtkrgRjpsLkr5I1cRV
XVEb3kGHGl9x3W+19hQjAP37xKl1ofeztlEgin/wda6S/NzUfsc2+UVn2FOasdYg8WuE3B7fNrYH
Gh27AKLpYt+tkgoac77o0N07lyxeBqeLJ7ChumRrhLKshu1UlgrgUAXpOmWVNT44hE7AYQ7GN8Rv
EoOm5WzS7YztwMNxCM4SyE8xR71HrUBcFQ/6mrQ13DcI8/aGygkyW2EqbmiZLXtPGWKpvqujifDO
PQeZ/3OjXYPn4xffU8NGvZPl5HtViS47qjIb4+YUYZJLsQOpcBE1bsNvFeoXkomWdoq30lznZV5k
ivxWjV/1YiyM1SxA5P73viF2eWsapoPrqYfzrTUBZcGm19EjI31mAd28EjtVZmjFQnppJM4pJV0L
zlrQHSZxYxExTQ3XPJAIKq5f2ukGJvtUK6VOPWI1W6mCXWJjJVmgWi2F5kAyXHTsv81Iep8Dz3MR
7O/g+MY7Q8OePhGvPPO2mQXVXLniPKxn7TCYwGqOKKZ5IXV95bbzd3H4jkAWj1TNy6MnXIfFDFtw
aNlKXDfaPFneLNARIjExkC+p+1WIGxbO4bWzDsOAlAzri9CU51+JV7+n6gQ6WH2OSqJ8t4Nk95C0
eY2J4xwS+H+lGRz4Z2bZzoD0GVqqN4wsOigaF1IMHzCBl/kVquW3J1vb/4DuiziR+BIaKu69Sr4p
8KR/u9uJVlos8V9IHHJ6+/iA2lM2Yr4WO9E+z0DCvb9NHbM3x0K8Q1TSx07tYJ8UX7rtS81UXtY4
mpHQBbNKpis7ftLLPQxPWw19uwXse9wCfLKo28t5vG3I252w6vfoBfQM4KKivKwPpVaTjOOR5Knb
M6v/ntTxSR5CJZYLAKQ5Sqm3RiZQM0IKy2b4APJE9miIw8IbcgDURIOcQQaeY3nCuLRAtXOmtg8x
1190hlQ8nPes5/9wO9PlId3LoPTdky3M4hWPOMm02qXW3YhMZ5h2V6iqJI7dyWOUKH3KOJbL9ZwC
k4Q9A4YebivSJAqFIUNTEOSwm2lvB6qXQuAn+Z0R7cb8WQOwftkG1lJo92FRh0Z7pPceZ50NkpLX
MYr2NYKecZT6PFsxq6les23qv/8IyIrp5WUvZverAjGT8IBnBHZaQDFGtH5LaFi9MyLrilNhr5wp
6MbGJZxU7NJ0QRbx+nmLUOqBNm2b8XwkNMJtZdRAD+AGSWWvdtzTde8gZZD+7ju8htmnFfRX3BkQ
Ec1LY/MU5I1OgJiwL0kAqVaeEF7C2nwDvUNxJU2aVvK+2IemBxcKIQjKlQtrKOHV1/kIxZqHi8si
mdQo6imNOSbrf4QMXxAxt5Q8KvKesqrVhtZ5AxpisAFyQ1bWgAnD1cCSC76653DPL0INeO5y5SkI
7B3DmZ6cX1o7g/aQZplpnDhkon028ZjLezW8xLpxByUDjrf3PruRDYdNUQIQf9TjiQbLzDmijPnt
aVAWim3grV7HivbqnLQyURz7cL9waJNGQcZeIoc5BjV7wCJ24F08UU31f5DeH1oZnvDoLzwHsEFH
YoetR1xGVWMQCnxmcdrKk6TcO5So4ZWO0BrwXFBusYQxoBTxKO6Y1+Yl7vjwJ3CaBVdfuynnR9nr
z+EjbEldLVUcTdSjmSSGvSqxWfgelA5fK3CuvD7ioXYUgh0IjpziP2uKRLbyG8nhmhPqTUbbyo5H
z1VtWyI14+gA3NQGW8tE4e/4aXibO/9R/ujktnN7ggn4j9mOY4a0/F6/ryza6Q/feedL5T0E5xD0
0SgDzh7di1xNaYbQ80SHG+6L1MrQi9EHUvrqYU6l/ZBDOeCC6kcQfugOpqExqBZh27KtXPwkDNKN
ROknP6fz6U8Mz7Y0liIzrdHBL2qqEoMPzbeLCk3O2mYXDtvi9F1e0VkJAr7ELYOaH/GZh0h97kT/
FWl/sERRIfXytoQf+LIx+1OAJJfpHnUHaYHe29cQdV3T401NfYMzn/2+XPHANdrUoTVJ3MfLL1D2
WU9yxMUspovDuL2X/uDTbr+VbxDeTDmIPQeKLWOhGpq8LxupNpjgnmQhll6QmQuOwW4vGECRmwq9
qA6I5sxRuUxxCQz5EKvThie06Sg/dQl/NRK64No7n87vDed41C19oUjSFI2yIJkHiS5gTfuN6lqT
4icU0f2SWy/LgOMvxy2ddI+dUn8sXaGPNSZ+GqXytmHntwiZ0x/OZ51fCTtLesRw/sjdrfbxSYf5
bk03ol/EJjoJJSP+55z08kwAXgo/LLZV+svzsQSnKjk/FDcYOSzJQ5dyyl57uFxf/T9hpIKnAHrE
FA2CKo5pn8GMgqZ36buYfwh0VlH6+HuD74NWdsjNdKUUJgyvSJi5WkmO85cdfPY6TmHXMMFIALui
yKRTFPe2A1zVQmObb8Qv196w5dZoIrZNPdwcemiR6QDoVwHmty9ufXeT5FEkWtBeyAWy/rvItHhg
v49EpuwMp0czZv7sPPhqkA0vfO1bLu2VhDL4Q57jZGlzS4tTyXuzATU3r62n1DQ05rsYDfHrW6AB
b40VSEB/ul+7JRVMl5Do/VgYM8XCxjUSpXLYvw6cgekPAvicHQ5/ISWkgO0HAcQNxOziBDM6xR3n
jj97pgnA3Y2POlMaPt+rdqAfdu0ZV+9rPX7ToVyiYyOuqJPMnW9ZvqED1fMX8yWnQXeqc1VR5AOT
BmGuwJijp6bhP+b9eVGlzaSOPaA/rTXT3cNUshLXApvJ2HmfJeN3vQQ/hj/FJpZSWPkr4eMwrLBC
JfJpHjx+a53/qwGptPGvsUlnCpDqA66vuzo45wDGD4VH/Kgn1u6TxHFSZjYIqSkhPq5GVDmHnD9x
OyYHb5ho/IHd8MFtV/XGr13OBCmdMxIkSAgeFVg2QJCNCKmF/1CnK1QLo5cVggrympz8/HiYy8Wg
0Ll3cjuJswlpp4rApHHS/tpIiJIelLYkHElsh+7mCqYUV8feQYb0Bzngk3Y9fWf6wm90Of9N/Ksh
SzDZjVxee+8eWcRK6ENGZ3NyeiA69ZmnrNsR25EdECDAzSUzXeEu9T4USf1nFIJtxOtQkp+8o1fM
bYRtOw4LY8IsREYp4o2Uk4z0N29Atakk4kjJ1Obk7ZEPEw2RWJCQZcmcUSVp6QPSEOYP7BAevyCI
9Y669Za/ip+DDpb/Ad5GATby/lusQF9ejShtHuz6B0NRyUktY8vAIGBfhzHKSC+ShAqdAkCqTL7n
kpmhpWecgjHeS5CX+54eTFc3XRbdHsuAewG8HyceTpW4z5zKxkyDae/j2/QZrVjlYt9GOvpYi4hy
0STGcEBCIvlFkrHoXov/o8sgXct63tHvtHEY+D8khEwDDwQoxJquZ+vBTiiQ+Qxz3OTnI5rpDSeT
Cqnf6Ck8qaR/MUeNigkZEEjPT7W+XowLI8cLQZjhHq+7VtkCwK/k66kR3yrlZ1uH4jcYkQGxMdYO
2Y4roGQKUF/xDI+vtu2Cv00w6+ZWNUxQG0b9za91jGWzVFZJUmjEKarCOKc2auzmtCbgN9UFbcpw
Ur8J48oalj3bglHnFI5o7EDM6SN9KWZBcAiF3PDrSUAUungv4hWnWswsDgSR47eGXSoebvmZcAj0
bm9uD5QpKqZNGYo22OL8n4WjPEQOS8+es/ZJUSfq1SRktkPmRwLXU0dvJUbMeFtWX2bPO0By26mq
4FhLjTrfo7qUZSYA6ywvZOoXVGrwA5CwrsgCeRymJ5SwDdSE1/6VXbPYqYidrfMSFS9ty3QzIOV2
6EOLDMKkw2F3xUfQXYV6BawmZm0sdBSrPYJkZ+rPPgAuxQME3h3gnXqy4AshHwHq4Y7ljsp3WlDf
kCYB8aoftsMKhLvfV52Rp1DYb0j4GNfM/XxDNRQCldvO8PyDLrPLn8a4JIfZk2qP2oeT4SfMCXsV
D2RHy6Ffj1DeSjb7bJBmvd50l/TfafiJf8fGc0rOXdiIFmvuJyydyxq5aRZ0KgvdTeMf4XoojIRU
TaZ1ECSlUDAA+4fDsl24PyYHXVBg3CuI3alv4hnWjnRt84wZH9PTG2ckETKdSra3Go+0H/jr/01B
YHF8Dbg7BwSrkmOuvm6KAIJdYIsz0lmNViTeDBxsnxY6TXwaAbwWTF7R38hbpo0IzYojvprFWcJJ
9myoMQ2gBXfKMJke7lzX1rKeJ+IRyhj4M2xvx2eLUvjowQKtZSiADYUCYzKcrbA3OPmjUJdgnc+M
LVLqZ5yfrSdeGNAMTCA2bXsdCS/XJrKF4t1MPjvOurfeEf+kRkdxYpBDkwEiGZ5uotgRJwNSuJJU
bgjyacvpyAtg/OSw9heV2jx8qun7/wF2HJ2JaN59eeqT+Vod46UHfHGIEZkRTUpqvj+xN85Jpsq0
4Ndo9PyEHbBAGUGe4HPAdtWbbBXU9Ww9w/tIU8iCr2xkdBYxrS50yHrvq3fKtVknKzHVyqDxDX6U
ZwWhngssAQK9WYTpO5m93HBa/gu7HWCHR+j5ws+mwpFar11GFBHUBOSUHSGP5XK/Yn7EgilRT9G6
A1URfJc5l3UYEmuFQUqc5OCJPkt+9CAHOqTqSOsPDC2GE6KXe/6teRrpoXCpd3iQ1dlgi00NUoVJ
A91+fDb+HWrjXs3ftaatyhQPv+pqwfQ/Uh0593kbgK6skUayW3BcVOjh6LfFj+NysO07Mxk9rv8q
LZSjvplAYKEB99wva/2AE2iffNz1oBdjItmvCJIKs0W/v3jJrjnAovQISg3XaiCN+i6vpXNwrSbg
ADYylgSvRaIc4W0nLje60kx5equCve90lejMfVkjPtbRAvqiGC0YlpUiTFOP2e2OFdyr9c6akGrq
L9S463D02/WHoi3IyZQicJrZaqm1JTB7o/c7keIW/GhOakw257YjTWImSnG52Nwf2IZxJkWXVzOx
Gvj+5E/ye+usPaAsioiC21o1bP4AGNaM6nIp5Fy11b5v9b0w5vt9hT9aTO6LODouqennm+2AywNd
lH1dqwD3TgN23+xUDho3ImYHBGEdYdmC4MnnMvP7yz3+STcfkDrc216vDtwfM7yyaPA20qidYINV
IMfkODgUaK7J5Rr8wSf5W9GrMDlzm+qSDcHAeN9MpOobtGNV3QBt5UcBh8SY+Nk0aJBQcFaNwVwm
tIAeLyfzZbaT/D+amkI1K6i8nH/UbQPpvFkEzWtui26WdatrSDQ4x+U8hYZiIDelfmXtaQ4ZqaUu
Si4RSoyHkzkPd8QibfLrbcTMXFFrNc1EnY2kx5hNbgKQ9i7PbeJAnpGcE2NTejBHkA/fWhnHRxXW
/I7UhyRlJp/Y9nByK/05Q3nkmbICUMcHCE36sKoNIq29KYRSXuJ0vq6czVLJN8RWc7XRUx8c6P8o
x6BV2GKfdhb/dhrzRuYUucqrYUtO4SzLbCleZuSZlj4F699fnp2EyTefybAM8rf2fV4dBtRQ+FbQ
5OQTbjyID4aeQTOLm7/IdaOoTbBxicuzKb1P3tEOkqioFw7NCgBO7TBgUzmYuHKfmRZH1Yj7NRD9
o5colC9rJWUQN0sy/BDA4ruOkCgsjA7Lv6gYN38ItUDeY/ABe4zzp9tldn5gOZnFnTJA5hQvIIQl
5xoMuiNXG6mnkAKB1WvPvMLIC0y4aWU+DpvE+suyW5myl+PHMs4KMc+IxX9tmDK7cKVI6BUIFlbb
vZL2SgM7YsjP0kf/z9odCyjJLDaJcu7HTdyaQ88K0Mkfn1Qyh0ZOxzIgjfMSOcfZsEjKPiwOR4jc
Vlp8k/mlPXntJaidhilvSp55sWIfzmx34YOhvLvt5/zE945WjhTR2ZKHv7+slRz8CpWO0VDdbEMQ
aAMSDH191PgnOAkVPGJEgZU5xO9zx/6XrUafZ7b/6mCaYVtaypOJqOCrpoCJR3DBF1bDW7NK5gwk
XG2T2+FTPA0kjIN0A/raLyMqzvwjCd/unDnmH7lYX8xZ46X41hjbyBLhxeHqVMPrGg3rUKlxnOi0
CYBhr6ONsFEx/gBS5ldspDwUYlAEX4mQ8K57x1rdFD8FUPPWtqS3cDoL4aHvAh/eboR/FV6+zy7c
oz30+p6JojbeB8kkEDI9BUnUYS/8zFJERqLVSRz7l2SaRZ0dNq0xFOQy/nG3LY2b7/ruMKh6w5mj
CT1pDflhacJ7ggyIbvwF9I2E6aCpFcy6zswUdAPg+f/XgZJBN/WP8LoT1SogHaASIOJuHtEx0uX2
cyLcN4W9bP8jhr/BRAsNjNCM3aIVkRj2gxDothG4kTBQJYsqucp6AYiljP2M8GW1UrgdbLKA5EWU
uAEoqAZdJuNmVqvcU0EHvAzQ1s2n8gJ9XqRHOs+ec4d7DmLm0raNHwQTOTFloFZJUIs911nlwSeK
jhc5zSCE4a6x/wVzj9H6ldrw/zTyO5XFLLroRyXQJnjNlN03y1PyHcE/q6Q0rjaomY38RC1Lot/n
PL6WNYBrvoKOfmXsaY8431ZDXqfPypHV0c79rv4YaN8avmsq7BNar2dP8NjVOBfTJACxungrNqmC
eRSFGsRspDnEp7t806NgPk5ns8tQ+6QpwjFPcUJiw4RH2BHjHT7k24cNBPw6hUeCnx2YJuzUDUsQ
Ly54a6Ed5Fb5UVQJncFtwP/MQvxlNs96VLnS/6XUzFaJEnxQjyW6u9j4uJOnUdiotV7i6lPCd+Vn
kIWHJQB87O88LF/sKYhFh5geXrdPFhoGz14gMvF0TwLLWb+aS5aGHW+J4e8fhEzuRlkqjr5Y4Wbl
tdYK63TSRIIVd4HLGCg8IICb+kxhvZ8gSjWoHT06KrdrmaO9hx9Kc1QAf7AuUgslUh/7Vs+UdmCH
zK4nkbWOgQDDbpYaDmvlUskhw6Agb6baeiGI4CYtMuNz4QDKAPAI2xyyJRGzMJ5zNdlDI+oQSjJl
rGL0gcgWIRoE6Frfw8rfA7zse+jzTbW3lGu5HUkb+owgg4t3o4ZRcrq7nE52vgQd+xzcszjwuq3b
WVpbaJbQkZkmp4z439BnPDazoaens+BTprEsvrvMzfZ07eK+8Qy379r8/Jhmm0Ej85UFrI7ZDQJ6
p5Tfune6NN44gCm89lheRn5liHau0jlvO6ypWRyDzq4qMfV1lN7ml5dx/oZkuDlZ7vHi9pvmSWo7
0eWGPuI470WyvXF5DCcgH87PJtWehsQu/RzaRCZ/LG6gQYooKCdN/RK5ZK6uPeSIIUwUhpAuCugf
o6qGHRYxZZKgzg3aDlAkIFhe+mq2yDidEA2SQRYpX62rU14F2+Tou52E/5YTolu9uy+qdEYCFunQ
z6p/CQl321lxDgO6tIQ51QehoHJH8W3KDqB2drfLHzxNFcyFIvO7e0q0ZvfBRkHYsVOTzJQhV7mg
WL+xegVrN7FrVOOvQ5tVGf+0wI4PS3MKVurmX4mnmOwX5OnHypFgnXhgvOvVBDdrayj8gGfeEnUm
mK2ThfbxgHi9hfWDAJshxSAcNtp0QXx6iSv1BvEtuL486qwYwObU/qdZDd2ARNtYFijxZ0WpVOLG
GPYLDm3GIXAh6Yr/LvPUvNC70G8CPWt15Qe4WsnaJ+i7FB0q+UJFZkoE88c1ByryG1WiEUZLTmgR
dK2fXBpPTsevftduHUB5AlEDJOubcSCiblzuDQVyQ8myusio6RXZsjYcB7wfnhfZH+7gNQWHGDUx
sCeSdGKNWshLrPOJfH0ACpB07vhgG5QURvk1Uqf8A4x56BuYH0lpWTpqdfA9BOpHkKHHGjlcGduk
NDstgusxLYia4IYjadgdS0ABtrOCLLvaihGWJoLptugpveG1oeuP6MZsOjxj9MzMH67FcM+2wbC9
qIouKiuiHahNVi2SJkvRmBbq+liMvHqEk7aYEuYRx1lFfB5OWPWQ0avnNUuy1OJriWUYAPHHgjbh
LqTmmHm/PGPg5N1vFX+7G2FRsYWT0KzaPy3MaibQ+5Qazl0feuID7SgQfgFf+2E9uhF30B7AzMxu
7lunHQSGmrWjkn4bqaERNuZN7uqV+6K1dcO8ZY7qsVGKZhtXeNT36Xyo59r7hrcYSWXSbwbgVqP1
K8VH4UkwuRvxrg8mgc8y7q4SVb5V2lyt/AD+2Zi+4MPY9gf4ymVoEkpPSF5ZSrCWP5z0Lwh2UbrE
moNl5HmsWDdY1syi1JP20zgMnIjIJjQlo3I0boVLEb9R0QQua0AukunHA09dFKnNHlqesFlcvP/A
uAKkwhlbDyEFSMEGjj6qIiSm9RNCvrNuAgZgDlChgFy6hULThqeu9DVkKQmWf+JXpDBrvaxZTG0l
9BckywGRvJVPs0dFlcrxkpt2+n49tZ3cCSc4hKG8gB4ik/9Gy/cywLERMGoXYhQAp+pCFcAg6RPX
weT6vJNGZAaQ0Fr6yPv3I2i0mRDX9Gyh607PpoYj3y0OtlNH6nISf8WPO4Mm+4urmAb06lMXlwGD
QEwMuLVl1J4yzeB7vOfmJHbtDsyi0iHrwipkRGXSvCwE+qMYBFeFfrWYjhh3GWObEEk7vuOal3ly
/Ifm8noNMYPQNHps6rX97do/29bG2SexcEGk2T3vVcNizmCaBCf+PqTdHzO3EOiIOPKlOZGH0HSP
HBovye3hWW463QIOP+ShFetqGtnV01zjzszHFw/0gNr3DOrpkGOu1zWmFxZXYrwgfvpdA7A/Wr14
H16lxy010bQwMrEQFRF38lnIPmpdJ3b75ZM4x3JFhA82ldY+2J7l7LGlYl5xTapCcdrhYXGQBZS2
IW6XSRlrzCxOW7haQ2FxLtT2zTGaKLuwDnKtetHpEuqccoisxWGKuftIciWryTo4UB65nOi+sOyF
yFkdZx21MDv/sm+054lj37x3nOVX7GOqgumzMtCkBkHk/pEkQH6BOMkYY3ryBgb89HyFOBVyjvDL
VGUDfpj/D35zsKdyeq/GzyEYk7MW9jhLNvnZjKEEJTqoyAT11SESD75jZ6mEFTFdBfeVy9kfdLxK
4jzQKWu3LHiyzFnlK08Q3b/Ch2DGIQMoL0xg1VvQiCNcur41B9wJImH8qr+4CZnZ2nFQdbSPiIyH
bATDcTWwv9aP5fCVG1a8ZxqG7GSJeaRWNyRFfLYfOGgiVnlFQ10sFzrr8fPDnQmsgcCqeKfLMcmC
b/dSPtZ0m5VLayPBMvHe4oigTtYm6DstQftgox4L3KpEvO/aawu0tSjtqP8gCIluMASNg48uMgma
H8iR/kbfs5uPukAcER1rT5T0icTRRqNETd/Dang43YIE4qauX1avAFA5OPW67IY2O4YgcmGcXUCR
c9JzQ+yzJQdlQp975tCmQIv6uRGb8dePfugbj5LVKBzM03va4iILuuFQEjMzLgBFJU5pYIceVDqS
9HfJAzykPNE93k/FjrSmXTn9qXt/yYZX/p8Mny2YmAp80pdAALN0fpPdBM8JBvN/a9w/nkeXT3Ln
+jZTX12woTF6cKErJz5nGJqE+VOLvr0hYsLXazKv+5zsCZYgd0GZrhKHQ4bVT+CSa3RliD79JOHg
Vf+7bjdRbEgBYjHAsNncaY8u/56rg04I5CBnt+QtW292PfP6v22OtqxJHf+YypdjzyBufqFCUcEw
QXv3d7/IHUbQDutW6orB8LcCa/lGSoIBq4GMdt62OfQhmm/+4ixUjIKz0JjArpFk7OQ04w8rGlBS
tlsWUflV9D8GB2cbKYGdA5Pto5it/47OlIvz0kehzdyeB2n4CJbYQSon5u4yB7Oni2PZSbuLljsh
dVl8UcnSTV/eLXPtYc5Q87fImMp5sJOXVIpABjdsJdIZLVoM+N5Vdt9PWFOj9sasCWzP6V3QvA30
uQQnkKr7x12caK/JIqJxmXz6hvrS4D8k/P8IWEFwpkFneXpcCrGAt7YaOeJ/6Oa4w+TT3w29T+VX
bHoBenJQrcS17oZ8pIIT+2M27SQR/BTzfq+lOYFhpT6vKVSSrPY2Cb5G8MwtG3uv8ved6IwuQ/DO
SMfmJo2ESZia8wDfMWhsWcWIP1hW+Du976hnNOaR016/8CArGhjaRMc7n06yDUmGZLNSAYQjIm9s
k40fE36cyHFm6/+c5uoPMMH+RfvAowlhINtfB1pr6iOjwwWP5Sz7MjxKqcgdu3ncfz6OBy1/+S8S
5PUAiKrC/1QoOe7BI0AhJJrDK4euGl/Ok4GYUTScrUB0yb1fAFLwdqJ13Qnd+rSNHRsdKjKqNMHP
h6Hk+SBAEQIrA1DZfcD7F+0W0903IWwRqvhlnA/0OEjMEoo/lTNfcgn7G7gyoW4A0G1195wPTEyE
h9mU38nuT3FQh5GAZt6dad1FmRmD2pDUfMiy9hUfkUg3CFX2U4Do51Ks9D1cBHgBUw/Ef40fTFR6
ljG7jVJmf7WUpXj/5LbAZn9Bx70D/IDwdTu+aCp8lpfnySSU/Zulv0gBUxKx8UDgmJtDTVmpJzg1
n+i4iyMM2Wm1RqtX5SJZrHKGThJn++ZwBC0n2jr0vkh7YwQWj2jfgc/GU5HgJyE1BbWVqX4s6PQb
uyaHA4CrzW0Ipktykk1O+vnt3O982Wr1z8FhvmH8p9xQy8DkQv/5fHTSbjscv+MpQgl56Z6CEJox
NJCWZo7FVKUBdJoej9nHzfmFRCoO9Se0eOmNHfKLTr8DVtCn5NNC3Hh9UBvaRxaZzFCPq+Jyzf06
/7z/aYQ9+9tdYzVDovg8VwyHMLJDQ1gbNiSHclxLHwg4ASq4LM2wzi4jgh2gc1JyVCoiTwX9pwpI
yIAzQlBPAoGwfk5Wq1YO7EaLC9TaATYgR8AobQ7GC7UBoOhLt/uBNGv7B0rho6+n/3KgNaYOa1et
uF+VgDjHetIGc+F0c0NZDneK50ScIGRYIvezKyNS+lZNN/pjZi5iMgZRMvlkTY8Z5nRG6MUoi1Ei
FMrw+7SkYP9jNa3YvqWvAINEMsVVU0rtgswkKr2lbw24ICzvhSOBUF+UXmPrCEnS71ufAyalmmWH
hXbaIN6+dPxAWfj68fCQBmuxxLw+SuOgLzSJLLZQ/TTBTGgM9SclZ3LGUtlTCzWqHLwTu9OcNXOw
clkWXFDrjXamqxzw5FyQpVo4MCdYVjQ4K9CoXdTHmNrgCUkepvzoiSON2Pprtebdi2AG21i/C8fI
T8g7aIoiB2KS5jJMbc3zRHWo/Eish3TGbFLRIjr//sAe+vijprbturS4iglnVKW+0te0Sl2+CSgl
wrDovDo3Ek/va3ozgT4iFTvdBdq4H/pWgSoyJVjE0oT7pp0f9hv8ODwvHHYcnLsGCGzSCP4yF3Y7
1F3VZe3WC+lQc3P2iZ4NjNb/6omW7ZwwhIDj7rO0E9sJAZuOabZY5XnzQeRRJ2p5AAGN2b8k5zMq
bMAHOuekQ8WfCkHdWarrzUbVTyTUIhsZoEL1t8wCPRfVAnUy2DrUW6PQtx0xNoEHvvyjo3gyc71e
nu7mK9Kr9yfrwEbr58z5QUrh7y6Erj70+EA0tpqnUGv/VbOHPYJM/MFfBgZV1m2+h6rSygdGLcFp
7TYm/GVIQioAYHU+10tPnGAlLOenNY7AXoVNcnK2uuit/WjYMR2uS+LG4hqDqxznd1fxX73y0caO
NRu9CucqB/4h7H+osN8tEoE4Nfa63rgt8rt6Vr3jTFMhN7VEo/fbB3v8nH37fHZpzot3ZVVYKKXI
9JU17WkQrebGJGqeBCnJGgMewe/0frjtckO+QHqZA1/0GMO0I58flDiSr9LVu8zWqrfEWz26EnS2
1cHO8ozPfvwmic0raOOtHlC8JkR0gOAbSnOXDytqjlAQaEItJm7nDse/w/PA0y5s9e76TC2ASZxv
DsJnMSiLnYPiAO7HgBo/U1/tBBAs0RuFTVeskmGNYMbmsP5zEbg4aZnilr9majqZKLFPQWBLoOxy
xlgjSM1dWFjMkuIBhGGjRyNdwcjrywVYsv7gV4noA/E5HDiFjjWui0kHGEFMSORcS1xfQNXchX48
jb6avTA32wqlSsnLoQ/PoTQFH1pBovxly0Ty9CIv5s11ne7N2aas/tOQpipHGWQpBVaqAmG8Mvhh
JstKejyTPAyjFgngBkqQLXsIbHzHBw07ZZlNvsmAb1x8ocmBlkjfUlzdLiVPevtsG0w7GLGsvyWQ
y+m4TZvdnKr5FnSFAC3P3yoVz2Z/jgYE86c/6abdIh1R5yJ5NODH2i7cmW+QtqP/epZErpQDG+O9
ZlvjcHl3u3jJYlwLgD+AJzH/LOJpYLgSm/FnPkbbSPzE9aV1JRfE6emkkTBT9UawSv2cV45H7fh9
kzrrPstlqiTm6xLt9uJWVzZ8bv6m7AUUrEhspj6qL1jN67oAo/FjTOXHmRwJhTWt2ZK808OAVJlq
Chjxmt4eLRuWjPk9wbLDh3i7bkevHuxh1T837KJw6e8o5vDhIst/LJaiHFEt/jLKzdj8M9+zz5i9
usZBLhr9PKWtp1Xlya4bB8GmiL6JIMfAHrvugLKrRgdZPllMHSGWm5BRra7UOPTAR+SkLVToeMYj
JuE1SjveZkXIf0WR1RVXAypx2iAJTSifBcux8Eau9iBd0iZrvMeaN4TiPPfytF4cIUmc0Cq1oZSl
1v2CNsP6KnAj2z/wN75be3HwnORo5X2lsILl3bMmoF9skElA1SElnrQxs01ZJ8CpWY6kfOtC3VJ5
zdzt9GdHuDSMR2zK9kunwyvE4bhWTtSeO8eid2YiRVsSVKOyS8GmFOowcjRPotkUqnie5cBILfwP
q6FwWg0GpHcI5pEPw1a0WGGe7UMa9X8ZzX0a2ca9CqTeGFkiFEHJ4/P3Y0r2ftLunSSuN+EO9rvH
FlU5sX0KizaWFeKTtYFCKrmSjQQzDvTljKF+HqDJqGDGK+2FKbpyavdy0PdObPkpSELK51tYqHXI
OSr8M0IV2u+iwDjA+YQl+ujd049kNrNN7nHwYjxmVfVqJSnI112c0k1idB3XoFhfR/ebKEjdSiZs
VEh1mwlvoENjiOPB5+L6LFjIPTd5ipRnH9qTP69OFj0YBiCI2Ok22zXXk738afOsT+J/s/kdCkmS
Qh9Qodh/FTQKdLRrLqTQcG00Fk/Isnct0jaq2KCLXH08mKtbTW0zhhrA3VPRBiv9dXZ80Me0V9R7
TS5dLjydeVCG0Mv+TFxjPRorySuaTnvpaByqpjR2rYd06wHCM7ui2QWUTRaB7+ca6bMVOf4F7kQ1
s/4JhJtho+eX2/2mdut9qYJrsShAo+zvwSlX6aKYVr0mKYgPijtTNuzhGpNFXiKQnlC2xok/3gpK
eVAhDIuBrilwicEcjOUlVuuUWwYhpHEimfNQHa76/KSFbAq6Dv+EF01v1bCP8nzbI4ntGt57G1xj
h2LoUwFOvfrC9pUEHkva/JcY99U+bTJ48B3OCZbhYsZ5DdmJKDZ/9os+608gbOZNsF8+D+AW1W4W
SHVrQ67I77fU9j0qnqtWvDDfqROSBrVrQpzG+22zaGl8I2hCkGWTMM7/6B+3lrJewsciV4hFBINv
kYyEkfwKhulK7zpbZMJem2Qudeo5xLvM5AStx8ETTk6XUARDAydogG4nz+2EwkZH4/5UDQNdZcmq
Js0P7bRXTtmZUYbibfB3rIi4fnsRXQ283qkkvJW0ybsSh7UhTyuGSybvl3wEiiHvYd5O+Fw+5Mxf
YQ7FiNbUH2W6jNp6tXb1yWpY14DGOlegPg+cqGHQCiZvTKytlGFc6EiLtPCbzhIxtNw9HCwX0KnB
v/TOFOXDdYJuFB29M5KxCBO0/Xf8wG8WrI0u86fFYqyza34JVmIwTEg8Bsfk8XNhPi09apogfid5
ieGOI5o1HJucagZV8kImkTeePesLOFbsCqSw5i8/PX2rbChAVPL3pLptLvr9ixX76W9hXf73WeQd
4Oc+kPHBBblX7E+uh6+KRiBxBESCfcjnZb0o5SFGGE1YAMbo5wBqr/qfB3+qGHJZUExtaoTVriZh
bKdL2sp42h84IZ9c45ruozFqlPvEiOYqGkLEXip1NBNewnuPo63mGikZkQlVTJOleabOADS3gFA9
7DIuVQ77x6nMoeCooslsOxhpa9tvuzYKE6Bk7pC/YJI2i+It6jo9U0qsO4flTDdkJW7X7tvkAb1P
l26rbNr/u21lx4Lu0MSDdN9Ma181WOxaeO9KfzmzhN2c/+HW7rnR9ot3mG4PaF9MqCzaxHUumFlM
fho/8aotJ3JWA3rda8SfWnH5Bf0xfII0Xf/5LHKwS3ditVJdHPE0XJdEn3qwnFhWrnsJaGb4fjte
VeC5rq4JJovYTzjzJ9MyQY9dnj2HldGszLHHHF02EbuVe7EWrfxjuM/GL0T9+0xjviCByQAmu6ls
aOf5r6kNDomFDPMeARLT5zNZ3GQAf/aSjebgIbyxrRXZIBkZY0GmtDuP+JZ3v5DoVyItyILVHSRq
m/DLcMqnCuLAScbsqOeFi5EknMhfxorqfGYXwOuNSjJxmMOfiiEfGMLV29fweTAnFwodEdo2/ebC
D3XwceVNFGPidkSuUMeo4Q07VvXS62fVgU+yPmg+fk2e116MNjQhk/l5kmBbkfX2FFqcxJhTtk2z
7XVjCvol+T+1AwXnnw05Urhaki+AHjaZaLHjZQrVIuEVrJilPSa+5TBfmcNeMfXsDREO6pZr/PLC
IzE2fZy3M6dXxdD8yDwGz2ttIx/+9SzsYqp8ST+RV4XUmecpnxI0l1Qi5bmY8PEvbIX25A+9q4px
OX3+BaMS5LjL8e9KdxkCkh3NavR8C+RU0uvSSeXPAbqV54lSZ4X43vo5BOnQQmdVmJ0bugLpvQ3e
jgFpgqO1OM7hy9rArNbG+NgLpzi3Pr/3gZjefH6KngeIoXTbOCyvoR/DsjbT8grf0FhFtiVQ4QfM
qHrbmM4uKxxxAJmHAwYg14XCwHBrj5oIcjnDv7yO/quaYlVwZYoP1wYZjiY2x+RouJg9JLNo90Kt
/Qae68XW/ksSWWacsNVcP2mG4ehUsordMck4o5XPGFxPwIhdjZFVLLNvGO9npKtPcYmbv0sYWuKk
ffEFq955phsqV8Da7Mtma2124CE1W9gi8hY53TCg/Z/AkrCDkQmjcaMBPQiWbGI8wIIgdfUtg2Tn
yB/6RfM2FGFIoaAsmuim49UeOOEUnpocIboOZLSCohbgskBukv50A8D5Ht9J07mseqKYa4hvUyOK
lZs6Towk3qSTbBZ+nvtf8yKvjsnM9qJNMuSwwQnNmWiSTKq+hgjEKUjLhPDG5t0pEUPfUaibt6dF
DpPBU9WE7aPk5DCyO5YDaye9UNG/4eFaq09dPQ9pKRGA7vy0BB8S/nZLuO7b+yUJnluhEYu0KhKj
c2Hz+4xItNA1lN2GrT5jFzVQDuIk/wJqa4wBb1fDIU1jgCxY+Mul+PKMEoVWji8v29A0psvEuEC/
fI5SAcnG+doay9LZWtYW1BIUwHzXK0Ta3uqufqmfemUMnLbWYxo9DHXwEepiNZQ6aAL51VzH4CHb
wiMF97mMscoligKr2cKNl9cyAWLezvvleLs7D665oWi/mKWaxUb44pqvIFdOeixOl0F9qRkcEkJH
bQlp3WzZforpnRhvjalD3I8u5y14tw20koTbmIrw5csFLnHKmnHgWFjMGi2X4hDCAi/9zF6nX7Pb
eF6szarQ1dgJpQfRYUgcopMEMKQQ/jX6229PeH2Qflo8csRp/nRZJMSoGweaMLKErBBCIFLIQ88l
tnmUhIoF6ABjZuEe/oXu8u7JS9D8042zkX75AW+RDyRvrYImZIkfFgM0dpEXxp50KKkVcYegO0U0
lTGQfXvfBpsEmGs9dKx2ZfDCnqMITz5bSSjed1KpjfQR80MbajZVXlxevWtHaaAZl7BeF1aTpXut
IM9p28M9eRgQjsK4V6yrajm9oMCTXZP7ClQtoBw/8/Gg7Cb66P9x4DiB0Ab+c7JXTVILQPPnj/kz
dgUZbK3tso8EmVjxM3N3IBvd8G0nQtW+hyXjYc+rgTA5v4jJ+qFBn0PWNMLwyo25WNj9csKj5KqD
Hmqw1YHmgJoMDe31B8DtXBKFv845PaqlTbpa/pUKaGshucSFkWOH0m+IRloW59KDDc8bdX2i1Pvp
p5EAXNYMy/Q3DB+F9Qs5qP73LbE+XQ/7ZUwWFJse9pU1Ab1h/Oa31E0EM1X4O6UXOSxdrNqr8zf+
voM8d/Fn77cDsPn0/4QOrvESg8XT4KIskwH2Lcq3jm/TB2nE0spNEoLbFkm/gf996SoQ8cfyAFQc
H/9EM9MHSeUA+6u3S7KGZmCInwcuMa1nHcnSUxQpRLz3CgIeSHBhdNltcp2S/emHSCM78NcToMoL
kNNtM4SqWrBuizgzn+aaQk/hcdJ+qQIy5+E8XOlxHplvO8SZSQGvcXj/u8Pnm5BeQl4wgwBvhJ0s
sezRUO3sFHzOQYsiAiVaaL1inQU3EcuE/TuWK1BMTqNjWX2uYI8bgHbBFHb3+tRyaG1+5ItnqANi
4a35GQXia9NA/goI0RFx9b7sSXr19PYHnWzUrN15N4x+/+ZjKjTH4T00++cikgVynjj7UhERjJsG
kFBVuN/Yf+mIBqJu62hdtz1BQA7F+XuzLYDk1THmUV2F8s3yKhD1Blp2RCO3EcZXfWEW4Lx3ZsBv
/lLRcsjaTEwT9bpmoXuuMKz/IOkeeqYrU+k+hHVObB10gl//H49X4FfmM17nPPueGwV3Vr8iMiDF
IaQ6w13SlOSznRbA+X35Kd2mN4jlStzZk96IPsBcJKY4MP473uFxnfw7whhU1RzHYBunVONDkYI5
XX+JVsamc5OkYMoXbrJW3a2GztogDC72oZhQgnp1wXc0i6c3HYfXNRFeVbEEJvSOx32xjAu8rouv
TO9DR+i3CMH9MZVG33BHYTWK5pNarAe31RFzehl3E2GRrVz5OhJ35UTDySqcGKzj30xPtPPyxdLL
PvKafqtIDniVSjGiHwKWBrcs+yullC5VxsKpSYrhkD6VDTjT6kjWzo38DE5jzoWb8luME5FeyDjb
a4MDIUdusFyiVBPDLBaAjGK5qneEn3M+dN8pFzFfdl4aCUblMhcuGhAoaWw6HLrISN1lLd2Ut3oB
nAkeL+NUSCfvMFMsIWxV3YThG5b3/k41AHTkMPPNBAnHztKmcOIywfvNrH36wESXbVTPgNCMtsfD
+1VsuB00AwmAvIpfJspoULAZQoxPZOEW51tbVbVKRQ4B+jBrRIeutM2TM/owAzKcDZZeJl+7EVPK
ba8SdzEqjZXMgn9+9gXcRGUenJK506pDoMuqVRz+KFDz+dq20eJ2KlsCHMVZFAlK58XLRt7TkM5m
72X3HZvmdpVp7A6gqkEVhxDOGLEH2aNeS0vulRUaikvWSbjJ9xKyB5jlj8GTkOKFPXF3d6F+rqop
e2C0SCwv8o1h7vLjs+t/MjHYKk1+KAweF2FmbV1pqFFuevzEnh8P2D8ZJmix5KJQSf1DDQS5X0DM
pJECNLP9mLR7t3glpySZJkHxJQQvKUaIhma8Dabk1PQClM/ZvgoOJTR15C3M0cvxtZ6y/umJ2P5U
vw8Y4HA4Ah6p9B1oRJk5K6/rRpDPALUI0Am2UjYZGH4zxYRrqPsA3U2cdtdKyQlZWO2+HoXdodhr
xqet7NvBbPN5fuYssB2/5xvefu0ogefGds/avQQSwKL0/qSTk4EbdafqMTMWrKZ4MG+d6Va555bf
ojdcgqDBMHaLtzX+DxV2ZUdpXWqG5aQLlzB1c0G7OoEGMdIJLE93G4w2hd0ocMzhvszukjd4XhLF
IvG7NA0gK+NmIeStI1W7YNTIU8Qs9rNgeftegAI69D31UYH5v8ZoMJTHHJjr0IAe4IxTFEBKnGKO
y1UI7VqyBsoShXikZPTm47MPUoYZzAQTwLWNmnPgbz3j9XKs/ZLbnybRgVnY5sLzIbfOFsPlwIA9
Uqsat+fiMAvdZJ1wZ/bWZvcUUMkQqISrVo5UJv7QFqtZBEOhfdKIqCQ9w6W8lR5qHS/Ngoqozu2s
HvD9BxjJZ4n+IxiaCEWaG77/uy7NS/didMWVAj5dueQC/FG6UrR37X03b0KbUkkbPLgRKkLWgNds
lqgSrzRPJ2gBmYhK8MaFsQvJlwh8WCHn0B3Umk5mxLiwoxj71IcKTgiAY6/HTCB4KkiRCUr8gIf1
ED/cMDe7QSGYDu4QI2PFerTX/bzx1oAZIJadojNVt5ywaEhJMAVBH9waijecFhfriS4d0T4BwVyH
4mRroFkFhRM1vEE84JCaOSBIUA1QaJcRJ6GEe56y5v9rXxfH8fd+b11A9jwv+Xo+erYio1c2mdBm
5hn1LeQARAoTGNps/hqUjMvoG4tMHR7bC7MRNpmROIETB7pcgDRd/9sGJ0dr8ztCCMhDFkQ2g3RD
8v3PhbJgd28TRwDl9lQzWLleLB30rGroGjedDMrnjkNL6HtQfXAQOqExwTWA/UWbPdL5dpoTMMpp
LJUjxBKV8/hhsQvQcobydushVPJEN5Qrnf0TyJ4sk3T6XI/OuvS3j52AaQdVLMCMQZdQX7IyaoMb
7vdshTwK26w++XTP3BK7EW5YHiOk15S+gQv6sluUKmITosNJ//sCoX4ckpW1RcMXllBv8sr7pO6k
mE+j2WyIXwEId5pGY264vepU0lC1ffjO+K4flT7OADTXnSuKWAxAbN63tsk9mnpwUsy0EyN0+AMm
siNuPvE9CgkAcR8PZZr8TYks7uRatUGKj1/A8GvuYWz0o8CKAEF0Pq2/p86W4By3MBHhBzUVxc13
DvNjE0aIT6nNZ6UiemDo86pAFAzWakR3wJUQ6W6hB4jNlvIWxccYwdmA9vV87ABcFHP4pqRlqD51
gyyE4BM2VIl/gn4VzzalWbFGItI/2rbsJEFPrPgRfLEr109CYe0nGZ90ckweeEM/9RPY/HbnKJFI
40z8eQV/OqkcIwx45Gki5zhpXODeGMFslJjasOPl2JJXcVFmLA/YW+hBeSDEjbC22gYh/IZyIx1R
+fDCUfx5MrlwvA5Jhtd2T7pupoGcBpp+Nd+IcInvdiXXBbeWtB4/mdZW09/Ic0YH0jbZfcJo2dyF
1M0YSczKUon0ZEw71AK3y/XHJvQZBoxdWtA5Zrj3FIEthBiOitZf5wWDpIvsaeI2bI52eZGbzruw
ROBeTd5/OD+yylBKTJz8Xt25c85d81wnX5S2eG8Q7KvhpyyGz6KM0vo2l8qitz+mP+Ml/n80ClVD
eyFy9UFlUw6L8Q6KDkY+i4rTXBjQs9uQM+uwwlJbxV60SlUShgYdEfL8armQJVL/V5JvTFHQpQrZ
Oa53H/LibnmNadJqj+IXE04lK0AwUejL5x/WQO3PovHi+qkvkKJ6ITzfXKLDa5zJoDZJqY8pAa2C
YA77U9pE5xs75CUqVlCDQkGRjYFqZgBYd3pySgYnOj3sP9rqyxQ9BecFPKLJ19+zH4g+GrAxvJtq
eLSz/ijDbI5x992gkqXJ+sX3sSRbxySqkiIxUqH5AqggzHFcSNVLrXVER94Kch3YL0h24pX3ueAx
SiMKjIaA2dWvEbmew+HfemgZYe2v+YPbk1rrInFRZ8EOFoK81cRwiTykwmJIWIP6QrnCb92GtDyM
AA9NHAN1jXXf/81mc0q7lYTX85QYcTuUalPjoS+E8LFol74hyB7OO5ZunVqm3NS5DcNa4dCp4ObM
/PLL1tiVwhNg6vPDUM2bmlyC5EVd2ym+stskHINYx4GuCyE994f02AF2DqPv+b2tt55BEH6wrvJG
X4zaphBMSYypsl/zvQdyNnamefGfg9nh9+bQ1FN5eKbAC8TPY56MU6pnYeLpckEeH/Jn7Zbh9RSW
DaLjOw5OIsFA7kuKd22r1XAThQDzKMytaUNCmn4DX5n4xC1tVPD6VK5rvKctq2ipUhsj1nJFJ+8h
r1vyKHusUUkg8ixc5LNHsq0hXJIWoDITh6vSdNGzeej7leVmLNoF/Y+DNqaRPpoPSGPg1UsSfn3l
LpUXwriMJmiD7l3i3D0RcHbsJfcGEVJrrL0xG9WPIdU+iLQ/EsWUgfV9p3G3IWZn/pty3+3/xkcO
APoVHyfgv8BHNGszIuunDblkiW5aVwReCOE+yL99Bz/i+c6OPX/m3B2xNxdtArmveeonXRLbArCD
K5rTSPcqa+UtuOKS/t/zqBMRqIYn/AW/9q9X9I+PsZArwlPxvd00X2u/ycav4GmOsVrkpOb4+UAA
RmdftZ72EEsRAj1vPrT1jbzBVjTt2TgvA9GfHeB2YgLqELUwm7DettJSOkUvlR/vmDTYO5D7ItPX
eF1p4jzLmoGhrY0GvfZtvUeq5Phc4y/Z8E1Jxn54a9RLpjd3Ssmu7KGt9KTxpkvBTa07J7hfWjx4
e4tulMvXv8GlCuekGuThMmGQ5bb4gTFLvGxYBOgRHmsfYvbRewfcFHX7DesLgXrNlGXTlVV3cdSW
nr9LY4Jv0fTHNF4ZGA4/bbEc6BCXYOQT960hGAmeCn1DJfGBgQmexP8cxr0esvMOImeJXHWKt2Ld
l4251ODbOHe2bIXMkyPdgv7iMh0P6S8+Xqez+UVPKqfy1f57wqqPmrDYtdv2xky/WR83cBfC9EMh
P2s3TUbUXnl8YnTSoH7B6kbJqGkl9idDxutnPLU0gTnTflDQKmBzMuJ/R/F+tp49iBnE0WcLQrvU
UBEedsAK1US+rpTu7qFOWIhkcYftD0MC6qzBN8gja+6cJSy0KBOcFZiaT3LyobgJU6T8J6Hp9BGw
gGBSN6pkjFCS7/oyBCujBqhuHN9nUglQOmjFVDRfy+whD+O306Q7cmhkTbPNkLPhYydE/0T7RECK
HakZHIMw+1RJlFpf2LpMoWzKq5WDM/OFgMR4NVTnsWaGaE27iQkSfGFFF8F01KKCpuJs9kiHNtv3
b8LUeO5ruW9dmsPE0vb9iMZaYpgZVGvfua0tVHMqMD1/lo3zreuMB1zNgulqRUhpQYWQijOhoV/0
I/U35kDm81lxFvxMIPSf/P65LHrD8gn8KJKk+uotatoQBxpcBD0uiZ3td/M0P0TL+CVpFn8cijmy
sP2sArB9K8xu4pkeIpxl4LEFeTxY2mhH7BFOhFITBn8EODn5WEDhFaHWfaeRqtQjnJkMnKMjQDMT
oNE6ude80Ci4c40y2Czb2gIWSfCabONlfGt9HMXEo4P5eYPjvREnUxkb97jH2n/TJZIBgALguer2
UMWYjt6itKxguotnH0XC6NzQzhuGI5Ri5un4IocEJxAPHPox0pQeHICCWcIfPBMVmCHp85cnxEZX
BYpV9DyYtYb1AZSXQtNUgesxSAhUG69EeSkb1L2qTOogWAEd9eStcZACHRvy9Pt185EOQm4IzJxA
K66fmfPvIJ728mmIoPIHulM04W2Lls2HBRqh5iAeygSFHQGxvsHnoTubkbsse6pbFRYOoU9hrzP4
TVMK8we359r/NtmKZ33bluCE1CFLAckEcr7IupyZJMxEc/AHOPEl4GkYhin9BOA6JwZHCiQBtZMz
Dv/P34/0Ads8rMYvw6/l3IXdT+iaMB0GAHKgqZcYx6Jq9r0ovoM3Ui/ais1sthCzWg2bim7HG+ia
A4ebxZGOp5U7ym0bjVYXY0RJUqgnCeE7m7SgluYaCm/hbkzMJUQuAiDmZS2FJy9sOBPgslg4dDXp
nUVSmaN8Jf0z8OSVJcpywtUrCovZRRfHTWRA+qPNt3ZoMcSnIKzPds02HlnTeJ04ckUR8m/VDWke
pK2cPpfIGYkhSPccF1I+zatScxBBowZ2Fzg0Mw20zwKYcml6q37xaPH10ovo9sTA+qif5yh10ESk
Ny2xlf+dpb7jgG2FpXS+UJ+ggEOy36Yt7y6oUUgwL2yqQtS4ASTrYyuTOqYQ/Rq7skTcq9kXK9OK
CH45T8lTNkpcE1KQQszsCZXJS7DSE6olRMdcjgntrIwg3XpkBUPZ9pQkGWSvLBdOID3MS7usgDCR
GGjYu1uJ/0AJtNHUV4ArFXQy9JD5ilmKYQf/WceOO5fHvmNN7st5XlVL5IjJ+frgv23wloWomngW
Fskh/sTH53n0sBOItk/1ekINVg3SfQcnVC33Aszur/eYrRKYXjZ7YFrueWN9HX1TjzurMIJVxlod
V6Rp3kQCuyVe2DM95X8qG2icwpgCom2oD6SNR91LTCJ07wqtZQK31xNFifh7sRccZCswHe1C0Gtd
c+8j+Miy+QyDeIpgBbwH7x7Drhr8aMlmJViwfQhVkMa3zpClv2szCX6ne4+d3+XJtetMPw0fdoxo
P7Tk3rj8WQm3NQn/s0HFq1xRxf1PJC4sSxDo7Pz3DR6OaYhy5d4iR2knJiHO/w83H6Sk0kZRRaWN
NMrUaIeptT5X9NUvs2AfiW4ZUxqx0tKMPNzsdtjUl/lO2dz0c3YSKC0UB+5A1D5AvMRAdtJOpyfJ
gpGU6ImGC7DK+eOSQBX1oHwSrJX5eVOFtAWTfFRg9sEM/y3cacGfn8s91ZZIVnk/i8EUrEV/8Po/
LTVLhqkQXvAbsSMpLRfUPAyv16AGKDWF6gjatMNbzbIPJ5AlaaU0nZnfEXp3UuCpn62hUbKcEVrn
oqO9CEfK1mVcGDe1AmrcvVRySuqYtt5TO1YHU/TViz3cEpmZT9JpwWYu3BRM9jydjLI6xKHnk3y0
hLnsRGWhiXtJ42iAmtwtnXrc6yLQcVFSFyGNpR82fVGTP0djlJ2aOv6IlmyDWRyTiSu9hyRvrYOD
dFEhtdXKm4Ple8XBdr2g/30atw2q+ujIDGhtBHPV7nG7rHtVECI8/YX43E89cATKoV+NXSEsGp3U
Ks16ezYZ22fqGucTpk0wAeoxXzO/8WuXyYjkQS7Ql6fImlyroYi0oNaOlSRfMs/lldQxJpzRUsw+
BW7A5DFjNo1Ztkk3rRmddlyas5EyvM8JAAcogdAaTy3rlwEnoCij/tlIlzarZK/TSz+zLAiNJI3r
ejFh+uf30cTb2X2PN7QfpfLnC3H2ORkXUMmNwN7+D/Fmp5d8+8LOBOV9ea3n1ww+uezyWA0Zn7q+
wuGMgFYvDMIs+ECzJIgmEx9ccCia18Mxfle2sawEbubgI+8XZ8dDW5tYpbU1Ne3fCpXqGNxed/4g
gt2+d7ewK4/6IUBvjdgCyUUl1Scb/BYmuYzTabjO64GTThYo0lQALoIR49CNwCYLj59r097HqG3y
xXRLXdzFxbYxxu5G2sLizAHWVE8Db/A6PPhxqXk4Gt32wsS3qkbhRItP5hx6ObX//zHh1Ty+pBWg
JX5vLp970zk3R09BVVUW73ZNt11z610FCXRMFho/AA4gMat9D85px/uZX/BEfANBoMjRvIR35+io
OX6YupO7gBiE+CidFQUJEW30cnV6eP3hZbRg60UBhlSG2+XVGRpl5w+58/LGiky3Nw9WfAjUAGYx
FmbE83u4b8hnCrxHrprNiQHI8BHmHbc0gFCpoY+P6s8vLqPt43IAFQ3s1PBGy+weGIfPOp+cjWTf
zKJZz+iy5HpK/RS30PPvJB+VcZyqXKbp5su1WHMKWH1ytw09HrrkGkfhusM8XusfyDFJmYnuIyHk
C6Zz1JyRai/kjkOUkQpgX+IgaBaeiBxJm8CdMWrNFMWROlABVrK5jKsxIyYEQjen6RZ3vHSAF3r3
NJ9rD2HnxGUTjS7Q1jp1HqyAkyYj+LLUtzOd7yjYnd6mY0mNkulVZS6vMzGdy+xoxzEu05m9QBRf
BU6EtVxqvXALFssOgF0DAgmt0YGS0QuoyySx58x+71KxFoYuy+OH4a3RNkWEQJPsFSxbV4+tXxf0
i3E7+Gly2TvEP3wyf5NSEg5yEw+wSV6gAXwlchjaQmxFZU3BoEzssggxhz7dBvdetGKM9UCuCAqc
Mtk67xpBHknewcyZNktI4gNJy6uARBVvPdJpRjGHCL7aVGAOINqMFcRNvgkCnfYdhGStCb2cbpIU
xPfjsrHuLK3b2cZDgGRralh/cMkNqB+n6bX1WjjtnLVXN7v6rQE1Gazb40h/X/V9qR15RdZXzHz7
XoJ6BiPkZjl4VtSksgLJFaklXKXF00XmTdz68omo63rnT810gQkYivoCp8K/BcTGSrFZ8xqdxmkS
uV94sOb76g981DCeBqj+mxYRQ4oX6fsISYHjzDyj58xIXDf3FZJ4+MLtW27aNayscpaDKCickFeJ
jBBDh5F324rfLg3s1I78UdRCjdi/lTW8+tD9761PkL1UjdJjJCfJfy8/j1FLQUwqqRMk/eBUrvg6
Nx3wibI/7+qUQ8NF1bGgJyVDVVuI1pIOv3gR+R0C9sP/1KYwxS2BxMSg3vxUG3OqGS93hmYF7PYa
7oWriL0Wmvv8yIMz5lkryB42+lLiizQ9+/1qVHipOt4X3qCz3qx2CjZEXuYx8mRMOVx1cV+L6NI7
AnB0O++18ZuMAl0hy4yzTyiaXDbRttYbw5k+LeksfiZg2u7XYF4Bpi1cA4U6zu1dgpr0Uxu0kKcH
mhkqmZmRbmN36FdnF3NFN5xfotdPd0zJF4MsT4VXw+SAfHizDAnUCFxh++HyttFAytNYlrqqyxKK
p1NMu1kZAx4xXocyBjG3m+wWG2b55koZ7MqQytLopl+0QbapZqk8HSau1tof882SIpWWpFZAAETV
dsHjqtMOM220YLpVfODoS0AJP1TY4dy5wQTG9ySKyY+f+H5mjjxTaI9vVtbPlL7cg+0QWMEvCape
sJ0/ODbQBjZnRDH4LiN7Fv0YWdj5mdOEZnLphXm6fz3+HZgupKM9iBQX9fDjUYzvvZ2aita7ARUO
48zdC9aSo7W+zljVZPJk/dMmiN+YaCXUdxCRcV3BGC/aa23KP2jawEOMSjgFPt+6g68xS5GRiXey
MWwxhx1jSoySgoQVJbecjsb6ceNKOzZqXj/Y5R6hHKUFuj6s+x7/c+f5IGBK8kV2lYPH9ZLctAqa
FNY8kWT0j4xiIXYIQZNGe338rzi4au3iDOFihK1o1k9XgXHpofopS4bZKOKMsiUQvlOIbyVqq3N1
Ubn5UvHgWHTTZ6xmZxFRZ2PJddIQ9jk19qex7l2w8DqLSCl/Qg67ERdWiqyPXzhRH5MUfDK4trk7
cAPny+Jf7YgenT/MimUCj8suRZyXHTYwPBBvt4z5jOH7pA9zjuFpyinT8IZKRD3QlH+NQ6gcrEwT
M+pjbjU62EjPXyQOL1pmaM5WbYtMeDurqOeDNRU0i00enPYNpRYSUlPVzPVg1OFrL9HTEcuU2LjO
zHuU3SzOeJsHR6rJ54WUskD2BUw81aC+0EVeH66Ca5zQSAGtWS4zx3Rwu9j+oGXhfEkp7piGtxRJ
EhBWqcxfnU7YVitn3aJBUVP5fiQeHWKHZ+mQgvoPpTLhuSiJ/fCbS9jwg4HNwkX3NeqzrS0TUhvE
0N/YGZu4ozw6rn/ArsOSbclDyhYWrWErZMQyLCmmWGkyHyL5qIupNI032MQcqfRa33b8Ckk1ZFHZ
J8bbx4d8xii8ExRzWGI0cWMKBnvR1mAvIdJLLzlNmHhPrAqCFjs/zU7/A6Tz9G+EqNZDgJI424Ll
5093R2xndO9m50cyxcA61gN9kpDbXHnMiZv3mJM38/Z4Y9vZxQMpbn/kT1zQAfEYecRvMnyxBsvy
1Fmn3x+Qv+ouEsGjb4/eoTtzaRH5DP7QgajBFy1nlvAJRXFwQngRNmG1LGPi6ZGDRkIofnAE9ELD
CzHhC78JGnJHLDU00KhXyyy7pOyySIFgH/shEp7K9ipaXNIInkPa+67LGe7DWT33+wXwO+/ASjEV
5EgQXmgNxFsN1e7dZpIyL1Iiip3fUGwCz9W75/ZddZ9fnhU3Np+qs3XRjzhem6mg1xZT+fACxhW8
EXW1by2Qpgct4wsm/iermS/akRcC+NOmjeG6H82mVUGc2R90m3fEhT7yzskHa+A5jrZmUAOB5hSD
3DfCg/mIy1m6K5rcKKqt7dVBweSP8qrXxT/Dwv+mC12vSUFVcektyS0EpWrSH0hGiCS/yptd405e
1Uo2VtC+lGDL/vCBhTBfKL2fhemD06EkVKipo0Uo2YRClaMSD0QK686s3uKN4tk1cUGN2RIPoNnp
GhSL5pEAdksl8o7aFQrpgJxbr4FK3eznbFsUiRK3eSzSDkcxUBm+RRb9z869LtlgbRPjz4IJA2q5
zYuYrUgqXsLx6Odw/0rCizlabfregIzHwfiBfLOZTBHq4/Ggyj4ia00uRg0Rf6DNORbBHEWJXk8/
bW3l/DLMfhcuvi5z3x4jYst86VWCHJqJqWDTtlGP9cuZC2gh4lrBmDD9cB8oIg5ezBrOSPC59VyY
TwC3BDiPNmrg2MRxSOODGaqIzyP7KCms1w6d8Cp5qNrRE3y2DpgB6X541RYHsrgX3SitJxmxaTec
93JqTeqMz0CcxDsw9Ke44C/UqrV9TcS9v42j1VFs9WFKQKQ82DYneyqG0s6bztn6XIrLG23DlXK9
H/ROiuHmrSvlB0OkEkhHxlT2JeuINzh2qLgF+XlS2l+1k/R3Kcny6jKHUMop63HkCC5sfqtwviGd
6axfRHXtG64unUEcBodQgizzGDuf0qV3mPt3brQvLCue3kLsNUueqYCc9Xfeo8JyGFSfVuJBLrY2
toVcYVVkXpDEujlx8WvinbQ0yU5uGtci7RxtHgnLVRKEgcZ0yViX0dTHMchFggE1IrENMdhrhkvS
vpwcHbYMbNKJ3O+IxRBphoQjd88lhj9ivcoqeDyP5sALzAaAblNaMaT90hmYyCDGzToGfmANqRZR
c82mmv/JDfODaWzPHnPkDUnFGSuqlXcqpIcBm4kIfaWQsPcM4eA8LVspQtcOuorblgei4EGDd0GG
Zlzx2ANaIE2poiVIJUmQa/wboNTP5CFCUcjNMeZHPAheftvjEfji4BNbOzlEdInaNs+tn8UGRdiF
fQkE3dED6FVkWpUGXEfw4f7bzUy5WVcjSkT3xFpz5fREiJ1s7CvxqscSlHwBNWf+MhFZngm5dNK7
IjzmdWRbRwGoW7CXyWsQeQt+2FVAwoA556nJQlkMwRd1LCLAdgaRNJIyqx4DrQsaJz9K8yPjabGx
jX5FwO466R/6zZ1xTPNha3ZiiAajghI2pePSC/SsgBZQzqyHecN9VL76g6wZSEj63Z+qKjymcfI3
sa/UgpTWr4jCNJgdZMMUCKFN6jU+422HdvoRcEViDXMq8PJH/9Jb1bgzYbMLyqIN1LPxNB03/a7l
PEr9g9A9QYkkmgQ4zi3d9JAdpzZuz8yUIhQLR0hO2J0R7EKDoEtYYbnFi+sMF9KrB7nmwzg0Kcs4
cB+b0n8zH7iHaGZ5zNMluqTFD8YVDlI7/tilj/JSpcN6lmSITF2AJ+DqvGSP6ufkSZz7rnCNO30I
SsWldS2CORxB3BPDrKYp+naxu21URl2NwnMZnhpkKhI6qoZSGxAuWxfMf/OGhNUa7ZuL/tB6TUyl
n6fMIz5n+GCtkuPgZ15hIgfLtv9Cv9KgTbiNdu5DLoXAR6M15vBnwCrDF4EI3FXLn9Km4qsFhQB8
FUiSFaTH5XkM8eNE9QMHf5g2TkDO/j6NnKsm6vVzHFJz6FgJLrribd8JVlqFEnuSMgF1XYDRkZW0
l9ZvdLMg5HdzDxuba0P7AhhWoqbNZdv4Ydbpjb2jC9p4KpaKloI3y8jNBYBI+WxqYelIpVPq3jvv
FYSirtsQq7I+FM5zm/VI6WUZxWAK6HSFt7++AnyR0ObmxdFxdBOLQwnqkheqQ5mWR7HoMBaPMUAm
67ZnCe8+ehAju++NbT8xRkL/WIeJQyh8QqtPNrSTYLBwCDhMHhZspga1GC2xb4aL8tUewFwyR3g1
VMow8WqZmTlkGPAwhS0ywvse/mwSNdfL3fA8wRvppMk/YXKYO2KIZLH3YJVMEEAN+EDzekPk1TGW
3gff9AprffFJ0LCe3Ff9X0cfy5DeboNIRR//5asKHbEvS6Q5E8fGvnk5t9Y6nbkLmGIt5iIeOunx
EZO+UxI/gzY90Cji9rX0p0rjMqbgTdiQsBLKQkOWAs7i/+D5ZcXrGTY/CtaLvqG2e1X3RnUpcjMr
m2P68l6HTT07ZlMOhUhBq41utTT8hFf6Da6ZKVfCEOlRrvsFbYoKsMKG+TOXhdAS3w+al0qwcDyq
Om/OtfJLcgT5CyxD0zP94R1BRqncxffg1+qKIINRgK4KOHTDZrrNlaNrCEQCdNYKeHos++L1n9sc
TAS7qho2yXOX8WOUsH72Llw8id1qpJAxrpQJC3mzbxrVER1c/xbaMN/MCAE+dws9TcmbDHIvkB8B
PLTgTbaBwe8k9brBhKT9LMvp7hQT452w9vZuQSYxw0GLSWQLF5d9WpYbSqdxeECjt/l6nmR73xit
rXZSO1ndhEpgJgnMrmrqYFB/B2j7G6kq9wz0T+yRB/uRXrf68iKmAbvNcKiCG7gq0nYU0tBSPQ0f
bHxSS576JqHpVCfWhBfAOMzRcyNtm2/+gN+Dk3X9/lytMJkcMR38N3rmsWfb4w6e6kqlmQ1bShda
54aL5GywXDHU7RVOaIDOmOxwHhK18fl5pNRhu7YvTRm39TzHImanpbnLMcmLyeKzmZVo9i0pcCkC
4VzybqauWxplGVwKGPAwxZXTRhTi37xf9YBfVhnAJ9PbOi+Px8sLljnbr1mvRaHvA7Q8H8fjp6be
027ikwbY2DlarC7yaRMJ1TUKt0hOH7daOhMyU3hYkCJNUBFzqYB6X/kFvKA/nUHj3Ul/B2CjeXRR
mV4FO1IrynveifbjKVBiLwcS3AbWGFVF3bfHpVKG3l+YxPHaSGAThDZgTpLP3Ue+LlwG2fJyEUQC
7TX6qD+1xehlQf3H71nnG0tOmympAoUKryvlpRT/SsU8lPSJJuQBDgoBB8OXSP87VfXde35Sf24q
31U0OrAUbYRg8kHbRh/RfGok7kO2F9AnyVm/ySREsTOejO6nWcnNBMOlqJRcDf0LW/JXBhIqjqBc
RYR2L18jn8gkGkiMVpcour05u6hW9NU8jKvXGm/hurpt11XT03/et7UBJFjOf4Rm4GZOI+yooPk6
G4llXrlRlstvUhd0X0Du0YDYsbIcH731z7wdWDLfA0X5By36uMtJY88+qPY73wQfHZTmdR0OoAlh
u/4sUamN/XJtny42+kLmJQ1+X29AMS8FjtNGff84EEn7+7HBzSrHPuFzlwUPEQBO9KdLTcRZezqB
FA3VLjuVmSSNwnd50QsjoLNdOQOTjfAEPrd+NW20nhgg0gHo9CJtAmVgafLBwuGrs7Q9TXeAPWRZ
wd/sqTUDFSTdGmJ0U1vHQ8w7NeJJ+2bmSs7JVpihzG/lU8+QhfoRQm9V26sjnltlG2RDuwnTbyWl
yvTgzLOW/JKzDxGW1tOmcCNFHDSi2hw+BRqIAzHgLhIcxB+Sf3QRL5ri/e9mh23z6a9Jr9B/+10t
DbuKA35ssNZY/YKvorau2KJyBOG1r01zioMk27pg7zCfi0dOBSPyf9aQb+U52z/Ppb/nY1Yl7ekV
hgzQqydPl4lgPBq6P3/X8zG7wyI936bE+DRt/yi7KzDTeVWoJ/XWCRIlrONWqaKV3oIhLcmqfIo2
idZ6BkehaaTuNaCe8oCxNcxvf/lZKJihX69x0+z3xMU+1Iyg7u+3LffA5MpnIbWJEHn9jchydwOF
HhS7OCn5xwBLKZCb1vs+1LDu97DO9G0FHZ81jeokvm2liN9UXb8cN1gvezGneJ5pbVVd2cRh7Dkc
ky2Zvn+8XVIXjJdp9C0knhiCBpyTMoHdZAFmIWM9um8+LQq2nnNZ1FrH67kZoKGbOJ+i2KaaEZ2k
/uU9nff4VZ4Wzrkf/PqYXTe/pGAFRvj5PXOyDrqdvqXsF+i00EKeYFYQjfCnLN7XQIvYXDrTeTAi
TKNMKzGwi/nVa2FM7ndvyvz0IVpvIk/WB1ybmyR+HoTxNAvgvV9RIwTMZmX9hCBzQSJYiB5/NcwS
SNpqnL5NcNhAKuv+vzsLxvusd0E+5IAyNcvvcjOt6h6pa0Qi99xTZ6LuI25FcJnpT/Y1hy2lqfw2
/siF457WGc6hC/yiN71ppdG9GfkXEaG8SLk4kl/iEmkUMrA573TdZcBchOAYSv49YLh3W4rDEIKQ
zVfri+be1icEe3/v6qLg/rTf61dlN+c1gKDCCro+n1KAPuvs8V5KXInFbFVdU7bG3oN+l8IZJTIZ
DnFP1MkKZ2UB/32Nnff1LwNtTi96MfZSEYTgWvmAd6hALyY4hRuwetCFHwxxeU+zGEPge9yTORpU
xdE/JaFBwYgBhsvPoiBN79RLxN90pxuImUHGqSBxxHuEzXPXr/fV/TRkBM0K86uOdesW1GcGgnkp
OorfLmHO0sqoDIE7RIGNLbR1895MbnPzk8CIJJeNBriljPsAC2nJs9F/9a4NdoL4YO/ZbsPgZDKg
ysbleCSrQrMKlmD+3tsbA9ty94a4nowK5Q/E5RVbsRi0FGVNGQE7psOPHN4ZiFujEn6fYZdqWbkH
60Lka/rQHwWxSxyiWMiCtZR6YPE8fkpFEufBOA+BFSQNlwM/udELeIAmxKIkLGhQQnblxzQJYkqa
8PFyZwFrCMoU0OuLwDm13R3Yp9M0C0n9BjWF0qLZDw+PEagP0hLC/x4FqEKxCTT4/+RZ+1cO2cVy
i5nfHeHy7AoOCwmMtc5yyZUvobMk3I5P/rc8H4MT0Ua+lpLFd9PBE4R9/Ns5SPZA9KmHqk30Qu56
n0CwOO97NG0Wq4/ULIg53DeWPDGM+rdy2qac2cEdTxdUEkOEGzC9Z+amKHtBnOx5r1Lr7Ol96HqE
kgWiBeBiTd5mxlidcIHweK+7Y7IkzLTuo18z14foA4lh3YmRBdcupeQv8bFvj82LmuAZi7gCk/o/
3RGY0yTDxiM4oBVL7A2NL2mB7ZgkmRUO+OxWNdY9UMmTZ/tP+lrX+cRzfAfqGLA4Ci0f0FfGrGtw
y54QUSDTidEoxUGqzk+yIFfxIPMMcDjTghHv8bTuCGK2nX4DOlykJTdSL5JfW0Ck43CP/9gwKOHj
gJPx1hc9KUy/SjVBrcA13K/WWebiG1FtGZHX8+OVBkslfxWwYNlpt0/W59OU/RQ/htMgxGhqzHEA
W1t066NwWUA28/lZ/KtFGS4K7HwH+IQdVWL/7otBDf73blOnlHKFiMcHwLdORpRUlPIp5HVj3kFV
La9I85v3UU3DBxVmukZNGSQdUik+70Vb46lfyoWXhjtq+vH8vGi0Ph38L6wvx9BbMoOmnbAOQqUn
s4huSnGY44Hgk9YF4/cRwHbDY1fPASvxX02WfA16V0oM233IeXduHZg0zRcZBc9wNcz91DJp9mnx
JDB1dBuIBX08Kpy5a9BqjrUOBzXXS3/dFcBUhE9Sb1kwZD+S+eGefKbA9i1jC3xTuURXdA7wvcy+
Cg280rqHsAmFTwnGrt+N6qfJNobcLAnrevb3Zg55kVo2zkNwy8U2784/eZr87gLY2Ck3XuHrptZI
hkayMMemdrSp2y2Mt26Ss7X+/0P9M1RVAxVg8drGYD0gtsmZYJpKe5P9mb9ce02FDNQE01ZzTvMS
UYY7c5yqENR34F9iNDnnYUTAZDle214xEWOYM0ByB5q9ujtnwwD1rhwLHaxQmCFQzmPOc5fkgEbR
PEItvvuo4khuiuUZghVmZwEe1x5xcaT1Pty023+DPZvUHt+T9yqa4CD1X7aPz7+t/ibbV6r6XbK9
t4JHHKV4qSiS01qm3KNawSU+2+IRwGd43XMGCaVDkMTHP6FwmHks5wNevfKK7J6QYxDoukBSpZwZ
o6OlfB7UtLD6kXD7r/s6CY7cxRsZIwt5hgRR5ZQprQiSrl2btNVH0RoRd5dJg0kH4QSnt5ptR0bL
P+I+YcX6KsJ/nYZrkGt0MlyUzwJcaxltP5NUNqLOQVzO1ZKpEI8a3GTogvFqOmV4V98l5GdAUsIP
MP1P5g2o7MvvTuhsWuvLvm/vWyvVu+u8VScxjdKp2JDLd2SLWS9yBTxstgNJ/bJJJ7BsXzw0LFGf
ksKKVSs40cJAjKC/jJI6PZg6jJUywTOg6UfYWBD8kZqq4iUCJ30AHH9MhqC2rAkEben9hbtf5Su0
B8O1fUCnTF/0YCtm4SE4wuZtq1i4GKJch5hn0hznCsNrKAjY/kJuDb1acPNT/77If9AtNX6bZZ+8
7V+Uwgu/nuM7eo3tw15S21ubPPhOdN6qoM3FVe/NvfhEX4xYq4lwH1jzCK5oTYzK1L+5P8R5xQz1
abXBiigBJlRLX7nr/m3t2zrkLik0jnhGygAvlhKPxxs11mnXaumvcaJSGlHT2NYvWdMkvQGzb5Uz
ALzGEeE2qzHSexcXVgf3j1bcxbSuKHWLWnPe5rETKhXqahjdHxokxt1T24k7hIdOseNSoDHDBCdp
CLF23U+gBB58WEQQBv5UVHV8humch7xOKZH63MsOdjgzI98YNH/z5lx19BuOOHW7V7u/bRCuwQ0a
Dac7hxblPX1/giTdMFDuDav1g2V++6bjQUT2rl46o8GLmrGsDYGyDKs4OnOBmnkTMO8L2KBN0YF3
Le9FqaNMEVMJIOxLIsp2/H+AkzcMwlUD5khtbUQ6rpHTx59goYU8VINS1tkL+Y4kd9vKDswskC97
EIfxginyxaTWt8gY01fmlFO4d14ucaQgsIYphKHDTOvcjS9wuTpn4sh7W9q30VgNsItuFI94MbpL
dYjM8yQhDHOcoK6ITkoS4UC7h/EGkXoiZ1QwUw/nzRLQ6y5t/UTgYaeh55IhhmGfGoJ7j2wvBXyH
PtY9e6WHY84p036m/gFA15BjgQQxLR+Zl45K+Fy5gP3k2gjvbTVkUwkQhoC3Sl8ss7dI73Q5A2Vi
TOoUwnJAr4XYi4U827Ql2xUozZUx3p6pypz1Vz9YFCTdnI6LmL0vPOTSJo6GuwSeWv3zedDIfbd0
YkfXuvlBfplIPkK+Md7NY1ZPwkworCirH2+Y4GjojXMJSOG8p/sBcxbYGpdrS3uYbiL6nvTV2D+K
hGUZdORvXhykUi0zCyQfmFVOvB6cIdzzBd1KSlT91Nw7A9uQWIdHnmyTXyPa/9MPijSh/MogcHkX
Pt3+VaCnWRMUm293D8esmyP8m8bb2YaE2feSobPjEeloG0WG3yX4CWiJQDi7MKK6OzWUFr0/wdYy
6g/4TAOH8r3W+QzJYhT17z2+dHmeq1zl/66ymhVgHjjcHFClbqRTxgmH8HFbPzd8FZvMlCu9MvyX
6J40Jv2SuXUosY6eB6krA0Hq8RWELL1Uvi8oB/UHt22krCJuuTO5AiwGkEkwetCvEiGo2g+TVeQ6
5ynaWG5vNSofISsB56uyVlO577OcHoid76Omu1N7G1Fz0KkOdJxyzsldQuoiYcCtOF/rh2wY0IVe
sP7s7V9+9nHFwRbJ9jmibEN2IS2+7pLAB737Ca4iFXe4GqoajfD6YHyQscsIMI10Ze0KR420A1Mg
Xn3tXRHxWxpbvj+F3DD6dTGMK0ZltJUaZ/Wj3Jc82PlWvR18c136DEg15rDmZTcG4ZENxxaFCEBG
jlnz78KN1VpnLeVY/d/Yj1e2cDlcdEWyJTx4l3T7JTsPF6rwGtqAxvl273LtReWAwXcFTytWG8BX
czSc2uZ5qjCyUzDJx6ICDDbvqLvvzF3k7hakq4u3UE6+6tkC2YKU6g5AEDsp6ax/o9ybTuHlEA8T
JogwjZ8xyclgiCB9TnQoWws3nlb7EfXiQldJ/2caWWY2jYJ7vCfS5t4W5M0E3Uzy9ndJJtR/FB0w
K5k6yhqxSDtUMIeFr/5KjdBZVAa/HLgejhuzaKqT8QsZ892vrlqwfe5aeM05TFhK9UZIfDJSPMdz
NEWoF54MEnJ9Wz39wfqH8UtInKMVOSPofSL9Va+YWb0Kdnfpf6DLmufc4Br24kat6aCBG1yC4PtV
jW2bVahE4Qe6rgMOMqGrqF4ag1Dc3dU9iEsbXTXpxoM+oNuSCyQnc7LGl7e0mdP3+i7qUu/ptAzv
73NL6b1Z8YmiL2Wua2nwz2QUBA0N4boz7sMtKB3H2/zbMEt+h917lRr9YHo2Fj+TGW+4cflwWvVC
YQGgGH0kpG2uMClf4Vz8wLC//Y4Om6XvzxE3IXLFFNIHKU5+E0Ov6J4nNOxOW4b2IVQGoh2M9usx
FcBZ98KCjkdSUnoLsZbIximffGuBxL6GrUzzaNbJfjYo4aTZOIr3BsLDDoJwtIepmKLlbHJQhvqs
4uuTM8GlbGStg9x5Dam26H7z7Akc1hLaBzOeJWuqQDpcXJ9lOdE9mUwfQWOR+C+SmGuhiyYXCKZD
Yvdt0uwwjSrvxzX7KAkd4tJbQq7EIb2DzCql0Ic/LDrQgy2VlJMV8uxkKmGOUw/z9vQPm6aHO/Y1
+5KoCoICwOeVC3z3V38HYN3NzY7NxirCxT0lrp5DCSdalJVjSJOwXuodgqmHm9j4cHYyqMyjFuHK
uq/ARbRKn/oq4/bIw5VZCy8JKu9h3kcSKEAjgK4j6J03PK/ZjbRN3EJBitifpVdOIEqo433aFnd8
k3VsHPLfwhFE2Afmje88YWP2SGyuAlQ7ianljQ9zjOLvo3r5pMI4cXpIbARb5aA2dEAcWNoRuF9Y
hXp3wXYiA84ezZRGR52JR/OUFiXAWCpFFC8rLqUfwu28HIKZTnmliezrghGZFmPS8hNjahFGKK/Q
Ut1EaBgrTEDj1EkzKIiyvqW7HRGZs3RjK5qPg+f4AnuoFicgX9anVYWwRQuQ61zf+JPkFoPlEM9c
+mtFyr4FILZHeqxS9otfNwXNhT3+Yu98lXQmhCebtCw+xgwmi3CcmqgWosmQXkGQY+nM5lSWoCMm
P6xScJHKvxFJTIASQKZLmJSIYfNZa7lSqASi6gKKx9ts68OuHJ0EIFRfv84zZwP3qhh3y2b+JFYr
uucy9jLNZpAsT1DQUubftnLjDVJz4sJKk6MA9TEk4m9PyXB3N8Y5i3A/Dx0B5I9t5azFSNKwjfMk
t3Pm+7C1/egHz/eWmGnewSM4KmOp6gYZM2x7lSKm4zFy2OZe6+YpxGP7umkaA9xBEu0h7hTgjLLh
E0LJVoSw3v1KBqcJ/bk+XA/8tiFViwg0QmVcDga5OuoiWN+T2BC4yJxVF/6NUjsz9IVuvJwkb2nk
aOw7/5x7zugY4+xOevuqhdKrdtMLoZCXjFz0nfqkPZFdcKn/TmJ13/YJ9Yo1jf+90oMZYuaa+uDC
7y96dqmMn9IgO5cJbr9eMNvp3cw/S/8jA/BzsCD1bJ/E1Pxk8+5ozVYyRMlKilpe6KF5LhXH/deo
VQEadvnahu/+D0AtfEQr8219YJAQ3Yu+mj7aBPG4cujSoZA0chu4cCVEWEG+0qi3w+VnFi9fIepE
OxA9M9bOde+N6GDJBKj/35hAjZuhQGxU4DGjZFZd6cDJCP6hsH1RybBfEfxAnxeUZuGEcD8zIpRB
WiTDV3zbMT/YOO+s3fkFyLZSuUE5dz593cVPbkp2ATN+6pPVisIT9quG9y5/hc+7WI9cgx/yY0dT
IHlPZEFkfg19JZnl/dbJEDOiUUEO8ohMayLfzNiVBvLBF5VTLrmzlj2tg9KkeOAAp1+abqPkEjK+
jicr2EZuLnAWM1J+nIsPrj3Qb6SqlWNoTTXJCHjVllCcA3DR9Vn8BT1WOs1+k+EIgE299QE0NAem
7iMBfXxXuQKA6msqrKS70cPtxDbXGcMg5dDc0jlqn+yTU4GZCY0hhG8Q1/PL4vtUSsYsnWYE0yEr
iwNpRKVsUO9LKJSmxOr0pVQj7CLC48I1zfKSPlRoiyDgn7mlcdwSVBKuJGKJ1Hj5uOHLMn3Nvz72
Jf7xq9Dz7x8NuxTgVsjtKTZHkoqY+q4cAacKqsqlXUxMc/uTvLvjpKxdSzqTwI/qEv19Z7yXTrPz
1SZtBBgiPIU51MhGFJOzsvFB1dx4lgV2BF7aFqH8dPkdSgcYPrqPHZAeAtHpHRXFYF01EtZ9307f
2YMiSOpZPTX5lxBCSUBCYXmgq/S5kKP49IL9uz8HLlqS0Q7hDwOnflt2/TR2iyyG1lIWIZZC7iKh
6GJY/DF4MUn6QvJaUIJ6849xoUEORH6mthnQTeJABv+pT2QgzVGRRIJBJSO3eeR9BS9ak2zAR2K7
FS7wdZYflzHkDrhlmE8kuf60pDF7J4Lqzwgw7pDcI4Lde/Qze/epJUDJwSxwESh+C7SFK54WQkwk
5ZPg13QqczYASnexJ2cV6lJdPrunML3Wa+tBevPnFWzPqX+nM6m1LgElMVzS0PkGzVzNoyhFQf1c
RqB/kiEaurJXsCoBPnA0s9z5HLPzoie5LNtcP2lRUEHldsNomwupTHZq3xHAN7GYKNQ614mbPlfg
FHHmOwbo3RagIMG8cJUywr7Mtuk89oThB0RWF0J11BEFO9LoKn8p1kh6/A0zhKxBKjJWf2AKW9ed
Yh7YSpfQsRoOE3O/befkH/XwhN/leIeJMG6+sWPQY6kOKNUQz2rpo3UmrEGOA1FEpBi3CkEHQ+js
QNww5aTttfG9HU6nvYDVxF4RvPalmMZCQNBIRsMWP/4zDQUbjBnXNF9cwD33CSAOPsa61FxUEzmw
m/zTYnzbaXebUmYe5Hw/Lj4QDKBlF15lSH2Qw+/L+2E4WfdZIHqSGbVbGYul5G3i9FOivsy2f0F0
vGn0qyhs1AZAzYbc1kY1drTipg0jzTDh2YMFCitxlar9rScXNIu57TODdRQlzZ7YQHbV7fRGzjq/
a6jq/xRR0SXPzfM3q0FpaTrSX70CEPlxrW7gp5OH6W8ePxjkATkJGxx1tQjsD/YeMFhyczIwKEf7
+nBJIF5iNcjOhpmJTckbxgHcWEAxcqPU8daET3enynooeGySi0Zmt89UhEp9HgaGs+Uj1Kymb0H1
JaWpG+1G+V+kW9IVnv8wToLRVVcPLhVYaB/t+r57VDTqowtf3xUT1HCFGyVOqVUTwCuVgqIJ7G5U
qwPULUPRsJwCunlw82ms3pSva9gkyPr85sCWm3fuewZ4yxdhaHJUCLYu4UUQvTYYEjCjV9IP5k3r
o9NiT3FYKPlIA3IlCGpRRH+nQ490jJ50OZX3GyMoIHcKiFs3bzWHQM3BibyGtNUpsWscKScJhJM8
wgFIWkiR/Cz0ccgo7+hiWkb8Nzdac6z9CgbGvh7Wi9Ib2HjNdFGIx1vpdZh5tHliVcQILc78BIBc
Vcn9193wyYw1io1qDHmQaJPUcU4LbDHOXRVZqrrNuCXBZaO4uxf9ObQMF1iTmeErkRNDcPCN+wL2
XgMq5/QOHCYbh93LbiImB6Gixop1eWxxyW2N/qdKsFPCiFCPF+GNXz1xzICEa9aNur53ydBpYBDi
D2wfYCfLrdcJWMzofX86M4fxWCbNDpOljLj/suZBY9thzPoQ828Vwq9Nm4esGBJ313bimmwQfGes
w2SPGwJBWCyWw1bgdmdZYY8l5CzNTW+FBkGNmrLtALE3ZCrc6stiYQnVpKa2e5V38ZQE0N0HO11m
Xi2OFBI3HYtw/WU5DhPxi7qkcBesYhF4Tt8qLgtcoYGLcCxRqP7vFZIbClc8rGOQ2nEsjVFC6Cv5
nodZu2oSKDq1fUnlG/u7S+WsAgC9XBUpgarIlGYgSNx9OM9fDCFHtMxbRuH+HZ4qQdQhyw3x2y0+
3D/YFpgf8C1Ovt9fT0CuTXPuhB/xn/YqvZCHzdnmiz7NEDBMwyG8v6mtTlMgHJndMDtW1WfAzsns
o69DLxGoMxBEdT7h3vZZVHzd9SQwLIi/Q2yn0yL722iem7qgweyGFcdmzfRsCAGacTCQM7R7gKiz
eeK8e0mjuNJ7OUbFSQkb0qNTctUrUq7xr5Eb7GfZQk5Zsm6RtTo9PUusUB75k2uRV+Fsdkjb9HTu
A5KrpIp6ACkwnnNlOMz/JZZWK8iTWvwm8opvYYAqluPfSFwwjkjGFE7yHqRTJ4TDmJO+KZfxzwAL
4NyeQqtfq7dbCUFl/DFyzXAA3E2SMiYyhUzWFAuIfuwM+Fc01DvPkq3/r6OlqJ5bNH1I+HXv8INt
eJKMpbE/sOQ8K+3VGrab9embkSXomWTZXo9nr27SwwcGF7ep24KdpvMTrt77mkEk1FaXKVeWyD+0
izktTP7BCowv0hbSWpBlK6FCtJmY2oXpEfGL5OOrKrl8abumUBGpDEw2ueHLariwt+nzGMoA+JCm
k1Mi51pxf9rLPhk/1wUmUwvBKB8Hnye5r1Gi6Ar+qdX7h7lg+JWD3XFaSSYUoXZX24zRBbXo4FZH
akRMY3c75kCmwRtvxWgTRBFd725TQFIoGpidN5jFmzkh7d5bWUeTvTrI4lzyYa1yw2egwkNu2j09
isBIPJDBf86jr4R/qs9Kp52jv+ndwWS7LdChp7v1qlv7mTuEgLjzvmUAZ4iYsH441T+s5gAo/7Eu
QlVLgygx08e14C5y8rgaKenznJx3smuiTd1YoqLjwZTVvELqkUM054BYvmSTHdSIARpC+XFzxY3X
TlqI3ylMuC378PW5mYxW5bEoVwhtDFQDIcvjJxNESQd6C0s1XcLJOyVy3oCFXAEneTai6LSLXhTs
11BnUwS6lxe2bbuiiOWXUJ2uR26LECnCHhclNNZ3pGdNZkkYcGFdRXC99uHLNoAd/9ux/YnJkera
KePMRV/RkFJKL/ZWH1s9Bw25VgWk51Q5m8yhj42kWchvC7CeJacTlfXHg+R+C5t4S22YJA7torve
nsuxPILIwHOi63e10vIDjPJPqadJt5HY0LNL2TLFiRuY9U6M5Z5pe82FzX63sSCcEGrOaF5X49Ke
HiOxPY3iWaHwUXZ4nmKTeExzsmosueYLC7bD8UbljgPbsaqxJYlGGvEA0t3/KgDvaZCBObfahe7F
Ug5R6IibDCwBwS+IOkp6L1t9xY19ZJTAn4DxqlZ29NdK6sL1IOBeCp5o5llYc63Idh+xktqGz0ht
Mtd2oI62daP/lRJW6IY2UHsJ6tVpbB9FrgvMwha/fLL8YVhfOTg78P/hruzoPdlKCHjU6uYLAKoL
vRVIsk6f5Xbi7nFsrP3tay0ipFIEK3Q64DD80goj04NOe2sVwXraUaZty0lTl0fRrLVrZZItyp34
MZJ1IHC0W+bYy1rntVRrfTEpxoMv/FUZplq7XH8weMEaKF0N7uXKFMNJCgEKpshbej9E1QHPqUfX
k/UmWYMpV4ckyxguoxwOUFkmWIR7+fz0XNni+6t5DIE3Ve7007RSxgG4RhYKP9/Cl+BmJJJS9jg/
cT6YX2Le+gxFkgtzZ15mU3+/7DOzj0szK+v64016vWWob0Fj0bDzVEIn3OTJvCJSMqWPW0DaPVLQ
uxbFv0ElbOd0JnCj69YePIXmjQ1lh8hezsVFmo8Rjy5TfyMLazcT6RbDnY3YbufdpNmi2wVstsmU
o3PvlHlynE5TkC7CDWx4Wi3G67cPx9CftqD5ZbNhzHKYN3pGPIGvRcHiDjcxp8YYR96D2IfS0GC+
+T7ezGSur4AcH/3UhTPnmUhA6Z5162OAdPUiTYxrlW2P3gGxg4u28xqPTa3cXZKD+X5Y2OESR3f0
WoHEc4W9hWVc3VOh+3FL9AZ7W+Qh1e2mxtS/KMT15iKPap6/1FpGNBTqug1+Ss8mLlXqPTVpDv6R
XMqVuKSScYcLkHFqjr46y7YD34BUfw2eWCqVllssB6t52RC6t6lZxKWpAN/nO7KpqTLJERUxvz2v
qAMlpB2wscQcssm7I+TW/38015PmcARrwEXkYBSVuVe6grVoyhs0c1So7IVXKoQCYbims/ZDMWs8
JFNfAzE6sRkokUxNg8Dd7O0rKC7qufjBvReOKATTlguYAcI9WTOzygRU4DOWD6cKZu3uFBqjY/7q
9Gh83AKRjr3E2Yd70kKs/mUMHfKF7WFES+ElVOH/5MX5d3ulrWnwqXcIij5nGKF4854oU9K1boBY
0kTM1jUitmqghJqaH+Cg6NnXK4sP6no7KXnzK/rYNR/wyvButW+dTS8sCHPt1vSigci8S+luX1yo
S1YGAFoqZaY4JqLQ+BGxAlGGAw6yPd3uByl/dzwx4VeUOblibFYhjvr68eA1MiARKTropOI/hlwR
va5JRVt+BdmPf94QIXGdQwcrB4V8/NNoZAUdVFvq1Nkgy32jRPfkieL4ZJEVZkSHxP4ttxweT6kD
gCDH+EFdZL+pAy5gojdO47j9JDkLKLEjJKS6scLrqKIG2S9exSifq5FL6PL8GPx8JuCWyVRV3Osv
RikWzSYPqqq+aqfKuHF3CS5AodNsLTDLGz7RYUxKXuPgT5LCLCgQqrUEaI1v3dsXG3UtR9Fth7zO
HuONUWBa7pHU2Up8SPwmSqPpzdJ/k9u71sd24HZ1winU8JpS3MoHTVsO8e/JB0/TYOSRt1WojExX
2jZQDHGwn25woz41QURkbDoa8ZnwPMNn2MJp5MF7CwA0MFldN9qh8I0amtGSrA3G4ct+6G03q/R1
A7tHufYqXnnujED2oGJZHxNN39vpLbkCTOQYozIP7UjHxUxnLzMKlhCJaS/Avc8vqms23Hq/dTkQ
Qs1fRodtFv0mWi+hbKGT2reIu8byDc091FNKLbhHc0yS0ODMnAYsY7Pjm+qhS47yD7vpodGzp/GF
+EARalbN+pKOX0KCb3uqwZ/gvVv0yAM1m9QdO1JbC3uHsRjiJIF6Bqsm3wz0q8ZpeGddEY+Ai8xn
A01SL/FE6gqUjI+W2XOp5UWIi8nDnE3KOgCoANR1Wn4ajh/wzbN/P1YYsRMa1afFDmXaFaMPLDMt
8vv5CP6m+W5OFILafzikqEWldISEMnqB7VkZTIpeLTh8kKxehyW/IMOVMmW4A5JtE39TVxwX5hu/
4M1EPaGdUGDmlHlayfBKu38NT0jLmYe1VkWBvmqaGSjEM2tQUze0MIBJCeySuL3uxQ37aFzdOHRQ
O+FNVy7hZl6DWAxOTZv41EzSvcdWCszj3EnUCukb/fTiREkBjZCQ5JCpIMY0uficUuX5V87Uwvhs
ahZ+rYhg4SSnPLqTZGoW8jmGA/ywTk9++9PcUIzPlmmwa4YZGIXtQ0aM1Go/QHfL/0x6aWruYeSk
gsQJvZuCm+5hv393qkYknXdnmvwLCAHnGcM11p72261Pft3ACj55X65Gkf+7iJDIEocVk1n7dpE9
JnfUYvVeJXFUdxITzkqHjNIYz2eAx7GWQtYNEuLK6vcnkhbOVxUPLhZhc2PWJDu1fMeK/gOd30ec
YM81qhnQ2INbmHSgXA56E6w9Xmcsdj7s864I47qB3IFXPNTPruek4B96rGWTDQ8wO0VhAEZialhP
228m3cInZTFdRPfJSuDTAY/91+X3msfA0AiZ7lGovGaAAlKrpfl7KcQk3ToDoSBGoLyidFoKDWmz
InPomYVKsdQGwWT3InJsm5t8ZDYjw8OY8f/jIt5Nonmk5uWJbRzgG/yeN5ebdYLecciiy5NHxlso
hbLmViYiXOcbnsh6lzbWnkWkmMtxc3TaXo5wHuay/Nz85NDlbUNTzIHFuo1y7r49uFnU4UECs4zR
g38c/AeRDyFhIN16U465uRfDYDwR89g8QVsrA7HOk3mNDr3SwL1vVei3swRvZzc7CwxQoE/UkoAN
+FpZgOtgbu6LXxEWGQAWBzjl0bRd1ZEDABBauLZy6pn/1gt9rTEi13VOAk4eDdo2dQocImWsVoxz
WNsP+pZIrOXo7kdgZrPvYo7aKUxWtJQUTq7UXlHLRc7TvXUWVbaxTXMrgD4vccO92pGXiZIvJiQP
zSbI0rbJvl/pVvVC07MCfcuWTGu0UoMoxIek1DxThSFIGxxn4a2lDaslHTAYsUmpDOuFjFfEmCNH
zJYjfI8nYYXtDWoWB5TDXRiQG/Z4cX3T9nY12mITolTAv/PjWhaOwcTlo7+fjm9iiDzKnl5/mlQC
iN+er8K8PKjkvCG/xJYzlAUaYRAU3Z7hSDQPuGH6uin2sOMQZx+SzfpR5DdhVymvucCr/7rhYcgr
8txzvnDZVq93KE7HVTe8UJZSsMzEMiLLUHf0IWZZmF26nHp4u/oc2nkYJzhRLdj2IjMoAl1adOBy
ulr91a4xQy2Kmbrt/ETN7KDA9F0pzXHQQHZvMknHrOdq22JIc2cs6PYaOuz156oXjnJGlUg4kj5L
FwHdQzo392mIGG/12qPDIFxZCUWaeZZdLrbdcCvWdl5xZg/0ksrERyNMjncUGLyYfytfMO75bZfl
HGYTXoUkXGV5ickXiNl+w10RdBvXJ+D4G/ypX33ZbIanCCrGA6X7IP/ttFxhXxxHw20JC9smFwSX
fwQf6PI2MNJSwEYOzVmf+i30dGmkM+H9Py0y2eFRmuxfKnqcjAcCVDIzjSmOOp4BHDxhqK21XaCI
X5Dxq7XB3MOiOiCxMmEwocr4u2PHxW/0sUOCoJDPw+cdJyOjAAM3PQdTOBMFBPwXZnghkwPXN8kQ
95rx+vcDBkhdmr9Hde91pHB3bxaYc6M9h5u6aN9rvDXyMukcOQ0jGR8WW7+CyRv/77IQoUnGIirn
XdiG0v5tQLvJV+EqBkLQllxKagj8rslTxhkH3GkrZsybJtQ5JsasMszMvAvAFivwb2fpc0mYCDwz
BbnzCmL38WNE45WyT2lPruDemTG8foURRJDMxRlSjl/5v1ZhdoNOWohe9Z9KKb6MBnYJdYdYLjgW
X9LxqsdY0WRRhL+ZNKiS6CFFZqgBAspGajTwwYHTtbyS/oO350XJCKvkeAGg9dvDcB794gME0ijb
Rh4cBlB75aFOdvxXpa83/NdmpzipSdl2Ha7aNSMhpq5WK+OnR63cYxIITN0PDu7YkE8lxzkcOf+5
xbeNUsfTWGLn4qaPx3i5S9w2iONHjKgDBzmLUZK7kZMdYIn//CwKet2gR7Go9vC9+B84JowAB2hE
Skz9/6jXUHWv4vW1kD9TzBJhz5C/R0qxbBhye/8ED3NadjOvL4M0N1gUFq9sSA01rWUGJcF6o3HX
2jvPulHy/1p7SUJrCy2m3Zl00tzv7fHnRpLzTeNqfHTuAEX4Igdr6OuckUkcCR57YzIqOQ8iwrAe
c+2NBLV5uG6Wiy0fqdVnkxpLRZW7B/LgmAKTi+N+RqDFs9kPRmwcs0cx+FjAK8bjAck1ptUo/N5m
qZsUOQrzMDJHSECkqg56//ILKa4pOcFreGodfaQqN9Bw/mNco2INCGvjV7ynz/LARrBRL7oJp72j
tBm6jTBWWht0iJ1EnGV7QVKpHEQ75OzDHLOjXtCkZsB1pVmV0WSO9h9L9EEbV4ulwWWS4ynmnDdV
187a0X0j7tvmyPOp2wWVILKIRvvvYbZqyFbX0e4oS1NITEL/ToNaoMRDMsVhQBjYO095oWxacxV3
gCnZrFIG4M2MIWW0dT1NUHB1xCz95TOii2jcQdwSCf7KksSlcU+DWSc2NrUSwm7O5+0lpERqLJ7L
f5w+LeT1yj9picyWxmOrAr1I4XQcZviDxE3fLtjPa3aPw/jcvliFyWOR90+D6B6swiVv19c4Axyi
TbD+nPjfXXtmoBk6TEO+wBbuaBU9hFWym8cnHlzHAFcrWqUI4mlJ5vN2UH1YWSKzmQbv0yhH9fGB
3H9Jk4/SLptTdQtvakjEfv/HhnuEgc2ICggBDrG88sLhZ9OTWBrdWl9nkWXkJ6pzFONhBhuXVPFQ
6J++R4yHDAGEOpwURSak8enBqVxZfFMcm7/eo0Enwqc2zkLQJfUYEH9J43HXN9HNawZEssaqCJkO
qb7YLO5t7WZ+p88QCshFHl0hjXQYpA3KnpPH23y+0fKKVv9ZF6ZgHE87ZZtrRhEYGw4YHJ18NUF+
Awv5lNnGU/e/FqM9DogD1J8LhbBv1LZx03IWRqmHQFD/XqxHy0rY1nJjbyI2hiAtJAXy4mYwJBz6
niD9Y3T/0s98rschWHApREuF9XGuUI1uKdPrKtLY0aHfA4edT9g1+D+F2NhxRGg+G7JJlhixX+nw
nl5eKSp0v7MXuysT0AyIjgfrAcb4ZX0ynd6QnD1Grp10Iy6xQ9OPee1kZnmKlYZIvoD+qYs8JFFf
IPiNFQe7/Sg9Xrswo4QAtSETfCfiQHhqaQXU/paPGCayVoItM52oJibZPKcyGcp0D0W9LLdTUJZ9
nAPaKL/kKd6svnXBcht1gsBjCt9sSQPjYcNxzu5bUmggsOk7yXbL+PeyaclO/Lgjr07i0w63yXlX
Gpzn8dP47/HHyw3mLi9DHTw3DVHwCmhpCnA6W6GVZASa4FpGAbfEHdSZkqzUP8WQ67OsXMVccXj3
qWauIHAah1YILQjhoLo6faTOm0GX3uFeKU4UXM9Xo0/Y82ytmH/i4rhSDcbc41DIv40WrMcx+x6Z
rPYoFnZAwrPDLFluK3QsMAnIMEQ0FqR/yg0hIwvfLtU+lXYUseYfaTfl8PaiyHdewTjptPPG1uQm
udJ4wxOe9Bn1004asWdx8w+DgDeC1X5/Wt40fsrDHCLX+dJQk3tibWLO0v4nqYeYfmFwVCEvBhbY
b5qCGribkNFMsql6xVQP4rGghjT/dW34fpFpAsGfNidfwzz1CC7VPCQLS1DUNJ7SkXab7ZXhAdi9
zgCpUwpz+plLRpQrWNm8el9D/RiUuoY5IqfKhV4ItFlPLa5pUm35smluOa7XZu32EqMPM0xuBs7N
9IEmYOxQQeWgxI4WuVq8nJ4dr28BBpvUuv9AGJ1k1rv4k11G7VvHj/5p1/+Uodbzqr9MLxftx5Qw
k4hsfdEvrwMGcxKpICt53em93yW4hiXMurO2Fr4uSV8Jijkygi1RI+fjGThtjIXOkwl3fQUMjVyd
Q8A27rfXiba+/4pXTJDUfnDsnofPypXHrmUk1WC0DCMwgtVfeuphwpAM5nPNHNaUU0MzO2RpmeJV
PzBEQtN3DE+lV/kbOt9lRoCfXUExeMiIbgE8xhVllbwYWBFhvucepubUU5TkCWb2xE+QptsndL90
+EEEGg3L+bOQyV5J1ztGIB4PpLvj6es3EsnjQ08D/DfVHVeIRSL1n/+xuDFnwdeJj33rjhrclkd5
RbRo2kr0atjy3/1MENGunPfmuOFFkzHo+XJcWUljnle2q8CK94X1kott3bcYDnv44mZqgnc390jd
bmnq4jq1E6XxQZCrrI45v8WYd/C3V/7z9GIXy8QWBgDx5tXMi6xY4z3J0TEKIQn/rh2eu8KLVHXk
KyUY3/L+GKAeTqFBI+38ZKivBO6LS0XFBPH2xtXyYquE2BjsgabBHgZUAn3Sv+G8QJGX0cMDGB8i
eblkoEy13Ol5Ilhu3Mu3Un0HJ+s5BTDT6w0WFj70aOKItVmZKSxonrJ1PKo8d2JL/mSABwk1LLts
Cjg97327UdPJvqDxWIgUSn8gOmofN+FPpLpMyrHUKSSh/qk0mAvaiWGTHvOBXI+dRwCWkbSldDwo
hTiDdBcbn+MQ077KRmdx2gCGb71bL5GhuYccl57hXyWCHSXOGRpUjQV8abF+8MTYGUIl3VLX3SNz
UfDdmVC1EMxPSbZd/WESTPMtQa4dAwaP5uGlJvjCf+HoiM/ZbwDzJK4yk22gn7GumcisfHaRuA28
QyxlWLiCOe6Tg6p48ccGtTdiA4wj+L5XorQfqGQqnRmbXbZFe/PvsQrTAUkfQwl5f4SZxkbOuXif
+5864bevGF44oeB01s8/4IbY0GeluykPGdZuWcTzBmONnoGlDAX17hxaDfXl9FiSq1Z7P+ZWYk0X
ubN2CDoFO4bMz4j9hipP8nqyIcGAF25MbgDWueA5dPQBNS4VutdyzdxodEXhlbqxWCXofMPb1zZ0
uMt3RUZoHO40h1t1y+TNdIc3/CYxbpaY/CDBlBFDTEBSLOo3jUDhqgHPW5bgW0N/Crwev1vuO5Zb
Rp8ceRmergcSZv4akYIk8kZckrCwd2RfY9Mra3irKNZlS7fiz9lFFITMIh09B3I66sN3f6MkBmly
PK6HrCQ6g/y8hoYv/Takk7+fGPChAeCQI61NVpfdkd+t33tnXj02M5MasUTjRwq8hn7GNZ7R0hQZ
b3kDWHY4WRkDWt4mo4QKsj7jtfgzkgCm6RKeaOdWWatP3W8QEt2y4rlpf49gOIOfONlhPsNzc+Pc
A8EZdV6gH+kuwey/ipDNjPB6qEdI/y9Itg+3VGwbqqZTIvL/uNcNyYZP03K6ZWQxpwu+Au/N2sDf
S/VCxEpQUT5ecRJx17wUFvGl9EJ/7X0brCzZBXAUOzYY5hpAnQY9qfrxVqVZGu4fHpE/uBT9a2Pu
2E8W2LOXo1f6T2fb4t2cuVQv0PVTvNwRxR97O8WCXAjOmrdjC8OtYk4+deJsKboEbq5+hhSsTool
9EEy/QdCL2vXgIwGE6INBDkWT5EeEL2cpeX0W41w2VQHbYLXEtVPKSA/V/9d3ZMuflsm4xg4xz9E
RWNp/UCSOWbREVLlDvRVsslmGm0G4+AOs6Q/glPhczevMY4xcRknFl2yZDLuKYtZd3ixZIktyKU+
R0bgpTMdpW52jxYQD/EsUAIs6XfpM8DqhsRW993Tj1cwHlki6CNJBuiF4ndpX+s+MO+TmOV0TGhy
/frfGVqXFa7+7e9Wfb4Iqj2EVTDmy2dgzyVKDMyQpXbIOz6X+D0bu36jheGvMQCYBEvBrmJ0Zhw6
qipsBqOQWUlysv0V66M+yehxdKkD4NyTPx3uhG8cZGQDjFYTCFekV1ea60iP14HwnpK7HnSKRxiR
14hTQYW3PeK5pYhtnP+oYSFKgGW4ITCrz9cS1pewXQq8wBupunJQ5TONBHrnaOJncdbtc3xUyqIr
MbcqV69xDjzDCXpbI3TeQ2/Kf32eoSA1F0AHQzFjxfEn3Zv6XPAA3W2yifjyKV9qXUO5XWHO6Xze
kjJLtbnpJeg1w49K8fW9Bz9EVcjABLovBN84hHXQomSWBzWYdqc9dq28HCgR0jUZaiVIR2bep5Pq
IGMJs9X+SL+ABZoG6BLrl9bo4TQXh8FHsmw48tvZ6tPrLRsVgzajfg4JewdR2rEH8mgDFUbUWNwB
U0EOLQTZTQjJL8uILDYukrsc3RXvTT4rhE4EcAf8BAJqGMonYBMSAkDLOWyw4xMNy0gaTcvjmYCV
rK7+CBe5sjlsDXOW/46Bt87rOCSrpB45IHt75bPTK9iH8SLW6pA/C+udORptKMHsX2ziaxMoAtsS
TE6HAWO6mmcgDee6edAkVZU3HMu3hLBqjcQuQHvXPCVnMVs2rYAiCS11IyT5LPOKS6pbmsYmIouz
LxxrLwhBr5jYzWAlN3/1qM+8P/sdPZWNg9anyKB1iaZLgo2Kqp4a9OgolCL4GrFMZ0rTvE11T3rb
lHBHlADHD2rlDJRtOByqabvJrPXI/gB59YN1IsNq5z/qQngfqrLNl0vaKhmYE4wK84VjjFGf9U4v
6w1OnBjfzdv3BoQAz8kAp9xfdqHiybvzjQbUGBErx1mRc1zuGrwflLFtnH0uPjrkIHDbcrA+xFIj
mH+PGH3VUKzvXurvdC2YCzLiikWJrDr4vSwOT0MCSSAURpRhJxJYOWRWuMlimtPBP5A2wd5oz7qb
jSAn35doaF2eVAFdJkYgxRhFlZUptvJQC9uOpCRxZBu2RoDa3PzJIB5iOmGkMfdEBua5HyLNeXYV
lFeV8toKucNyYoTOptMJ6F6qorE5stuMY87NNm6u3C2yiZywSn7SG1JwzwXePtbxRNy/BBDEmoVv
kTM/zo/hPZOO7OaCCBbNvDj1sNEFOuCeAyOV8IWChzxKSej4UUFD1ZMNsMdOtho6nIXz0sjQ7WGU
vr4TJT98YDBCbR16BuL622OV3FyOMYXR6dkAy/uKdMO1d+HmYacMe9Ztx5C+hoGd2bV2ztrB3Ufk
XmOfZMx44g68DJqF3ULdmF9312E9NW9SxyjXLfgVvS2w4/TryMSRiCRZ+o/CrzQG6v9uonG6p9zI
lWWbhCTocEjy9Dk5GCfYXBc47flCjJI4iao1qB7uYYnBl/kC17rKZc7MoYYzaNoNhuzyJPsEBhQz
ZCpDYXBwIYHJU4/M9sSMYmTO9Swd36DZkbRHF4HtlQfqdiIu4Ju+NA1C4gbotN7nXMfojZhMlZkK
WX9kHxT0pe05232ACTjnJtsywMnTJqXCaR2g6DjmSMteGpb0Ld8buBrPUsZIbNGq/vYODJOTtyf3
2LbJjRVwCK0H7cP1SbiE+334OmqFC7W5HwZBIAQEUb/C6iKmHxYlZMLWU6S2Z3N4hVtD6xelzRG9
3ZMWc8b/pBOUqB+EdzRySTT1hdM15uhv2gwVv9e69vcg+8KxpJySYd8y7YlYd/9nhQ5LJ+ik2VCD
NSSjOtEPpNFTSDYL1JKdSxg4iL9j574WJ8mDemSVlIJDobmvu9tsZYyTiAPqk0X25kEX6erGv+N8
ccdid/xP0vavUadx2wJh1Ir5BCEvT32zPmZsqxitOZcGvct8NJQYrSUjkjXsXT1UWx/GALnaLD/l
REikC0IwemfyNf03KPpVuRejQPc2S7MO5NrAHeGeGrLmZMMEAo8NU/rRUncD8xQR29RyPf6XjwD4
bqamKuFNRefh20+CUAePKj0hGuZaLj9n2Rw5MSiy+OD2VjfNfqdiYZ4OJJltRu82embVt6kcVDOu
WWvc/aWehWsRAuO73he+5vSM6Zb6eHqww0O7zQL3YkbIcABOEq7O98rSyAnu01DC3YdUtMcyCirJ
13OsQkRDe8UifZLdHXqJ8mWtTzmdufdOqY0nKy6FJ9zhpSxDs24Pin58s0tKOCo30o9p+j0MRTi0
J52Hzz0rRIQrWpgNiPe3NR+IBmUv5bRzkppQbKvczBbisldmJ8jSTisKpqy3ajEaldKT18rS5hyo
rKmf2HSyG4pvemC+lWzthyIIs7inzJPDOC4TB7f4IpHJajpQO8CYilJ59UTPu6UOtoLS65XdESTU
P7kDXsU48sASRqbRCDKR4JMfx6/jIkitliLw5+b3e3BEWeI4LqXtfWXVfH08jlf9qhUmNJC9zN4F
KJlDO/ZJowK/v+/XS7BXrb+gGgUCnTwUpJKwsejcw+yZW15hQSWYApdfPMmOPJ3w/SoL5L2PrWw6
mX2CH12IwFKs66NwqwZkBcq4Ecz21y19RQ4OyJF6gdPsct7EoPYm5ZjGLbxtEn1ccCc2BxnxoBiA
K+VKSqqjUEAAWEP0CIBCUxjmlexckwtZMqflOSVVtr/c03ftdW2BZ+CJ/+sundtB+MvOOhEygTfz
dlsEjj2B1vNCBEujn8iB4+VV5uUD01ES2L8YbcNPwOiFOvTfRC5fgQWdQWvUm5yCjTLec2yQxqWw
+JXQ1sN8mUpojnov0MMOk/329jWM0k2wDsfx72ji++AnKy69f843Q9GriloY2+7T7R6TYLcFTUZw
u1P81N/Ni5o45EXtulmwWQBpAKuxqrGZbE0dZCUXwX74pnlNtbuULmoh4kbH8IQ3cEWqWaJnLkpc
mJ6WlJvCuDrXca1KlYkkrGs5frTklfjEd91qkr93qnsok9V3TnReK38lJD0prPeDYD1WFBvRbwiH
49wGkEISm3vSCLvymgRU8Qn5u3OdzniFV8FMU5kgHvMdZNtdKqrMMlkkxZMO2+uOujKCfdxZ1hba
iOsMXCG0Dr3afhOn3eJdnsOwS5Al2JeltEM+RQlhwVT4h/9Sdw0iRB6bqDR15RrXjA8TYcUk5P+K
qDkgiKJtSt6wcmfr63dN/1qpp4E+MT470iU2EJPVF5HyGmTm8Z6WSa4ynYFqL2+f5yPYgt1TC3Ny
F0wu029Omqbh8VAaZSU2giKzZTXCBsUPZa3ud4Ec3YLq5fHPK95eM/ergO1fY80WacloWX7YD9k0
N0UOM6XPCmqnrOXVctgkgz9bRM31WKskcdojxUsbFgaUiE8XbFgQEgm1t3gENDsa48CY5USpgTzc
bTVR+VYf0ZGRIHo12FPg1kYWR1jXQd9AVEXQbFRdrJGkXvwz52bninqOsyqCPOfEheCGEP0qaTUJ
RUBTW00zq3by41g4LVA0pjCPrDLZg0PFzrh1rIpRmfpvghqQX++vr8sbh5gqvNwQyQp6G0FMT6h8
l43/bFelIaT54s6ulXChsnMgtptHR0ZGEVTBJNL7a2DzmFcyYQ7mr1rENiq1HzVzvh8NjWcSzqtG
HTpbi7njoXMpwtCTVFwdVQd4GEUNCrwurDRLKfwjfxOYDqMwnY2WToPpqZde2E/bctu4iHc1xfG+
74IndSL/c2HDWN0H8JS5XTJd8n77eYwDj715yh6CWnJv6fKvPP1ODyOCi6soJPxkxDsf0q9zTy2H
jRg8td58Ki1VXNWiTZBeuun+cI9K6oFVNg6RxQOO3LrqicjjCVnaTFrtoCNQaO2qjP6C9pCcdvIw
5iBOArwX8+3CMWNOSAEEaKEk+hLUwD0SX/36GS0janJHKMD15IvJD+IuCULaEBqRQLCY0YNKLxNl
WpCN3PF8SK5TYgKC1A5peRi3rBcC8PhqvgnSzQhu8adym0rUD+cCWhdwQ8uqwzw4sa5I+/ZI8T+m
sH1X7sMJbvSXmSjrWHOZF+cAafn6uI293v5lZ1GcNIP6poFPRDv+HayQ+NBEN0xXlYDkAY3P2JL4
PcB/Qc9kaCnvt13IzboGe/LM866THMp/YSC4f9RmeXM+f9O/7N4R8NCl7/IsO7SbUSgvWhaYP+Hp
2I/AJEB67cVtexWJmsOgdT71dCbaEZXfRcJkOLFDNZb12FvmqAq11Z0wLox00sohRGZaJOXE4xhf
ybPXfoQpf5im8Nr1PnodAjOztHvB3/rOwcrI3NTDtcVbZ/OH1CsdhDj+BNvplx2Z3a+L+uKiYFlt
3hYDVGDJwDErxEfoOj4H/4j6I0sa6gTF0NgV0CTeab4Pg25vnCUpGCYE4hzxhcJwwhfK6YhfMUeM
5sNDTXe5UlHLcyLkYqAcynQ146HSjMA1eaD/oKUNQxQWgzblh7nxynYiM0DTBcuYlitEL5P7Ubzy
h48fv1DMCOcOJ/eyV0MtpwRd69KPMlcD4hBwYfUhNNOFyo1gXXETxdFydATt19ddj0q0YSkwWcln
DYQXz7F0F2OD2Qgu2ZXvPOfgjIzZXl1iFLSjlWs/bmH4BkAF5RweTOuUegeAbLi+NUVHTOsREZXF
GUD/NSKyYXRfBoqMjgXxDWUe3d3vSi0x1TRS9nIEbWATPCqGS7lTZkRCBuvvdEEIVGgqp7gC9Fbu
25sG8Dpu9ECJwf3ra8598gC36Mh3Tde/1mmB4VRVBvuRS5AbA5ljF4yft2hO7Ij8iOCBNNIPvoj0
sZ2hStKYJPvK//AkEO84utmW0Adi2xGxluWqXhVpuYU1IqqE0iqfUFDNbm9sFFG97LHQOVsGg9YU
1QOAMYTdyGsQ6rfttigSokjzHJedx+z5PE1xdXTw6X4yDc9y08QC9M/4qUm01Hm+7Yoraefwj7B5
4kAIDUppsIm87o5H+XryGK5Z/roRDmT2b32tpk7lEEWucRssikhLkDP4/F0/FS3IC5WKI6Un8iOq
c49SFkO12kvQOHkLxhKWmVO4Lc6F7ZkXmPxPxMkLOlfqiK+phncgQY7osjNAmI35eW+vpoIIYdKU
yJJ7/A+9vncLIE7niqTZhLl+3h5dt0Q3L8+3atQnmyNR6wQApGZQavHe1k6qTy4VgqyqM0c/O5JF
OCVfueIE2SKel6BA0bW+bCdtpNSWK8e/BmcAcucNqv5chcnNjopDL1dQqFUS/Daq1N+aTaZCnqYT
AVKWeunBw8s/xJLJrvpehYDYTgqfPa0iiOC2q6CXK+3FUsV3eT3RXxcraKX8X4kxegr+QAcJhEuT
BlrbXiaCIkIS/Q3IzF1EHKX5MqfMluNxEUUGEfFjIGmE2mJn3Os3i5XuZ+Jid7hVw/S/9CijiHNx
G3xTjMrTjRY5QrQ9zMGKYHcDm9YhvjJl1+jefzk4aJb8EWrvkY7qFbU5Nps6XfUUUqST2D6J230Z
PkiNWouhSQ0/Jo1FDsVul+XXilWNZTDOtVIC3m3HkCNIZ+nKczY4QEA2aOb9lPIuK9JuBnwcWf5k
K8QGtsYmhvBUt5/4WlVOoltr/HrTum85oSnNzwbtEXmonbvw28cqDa0m7e+dd0DDBV4g4Bcd6fV7
6/urCiW1Ro+d2t5UCd6AMqSzf0xTka+reUBDykNoIFnYo99CaxG+b+o5k8Z/7NuNjJR1HAiT6ZnB
zYo3U1ZGjcrBI8JmWdTxyH5XWmIXVVz1/WMN7DPgH1I5yyRX3wMdCWeEXMarEtILTCSCQTtzwTr5
PtM6h3k/X/e3kPcvqVb00+4VSDWbLtXOIqckah866NEA2a/3lOb4oMU4OQPZtucymxJvvae4hBnO
m9/qY5kCGz+pOpc3kGbPsJUC3Cnar9I3pq2lToDkPoHQ6YSWhqPZslFpXBpxegerwrHSmGw4zSs9
Biy0Xe0eT9lt4U/SUHkzHYksUGEV4q4ANYecfYILy0B41u5l3HQ00I6szlDVVoZ9jxmAP3ligA8Q
+HkGbCpgOsWVbqqqs8aDueY+RF6GvqDtxQP+ZdwxqDX1HLoMR2hbsRUaHPWNe9y/NR/lNAk3KxxK
9tpb94W5akzFBUAJ/dJlCO7HLoOPisJzkhVCeN0ynvBfMZpt0JaV5dzT+fjLphb6nASJVe054U8w
C+FxEtA1u74P3bJFpKuZtLGKwJAJ1fxPLPBcM4g6KwBB+ytlkuJarCewlp+AZqghuTg1gBbQsILo
Ohy80oWZSCgS4n8AL41/ziOGiG436W+YTs9+bmvYYOVYoRpnqcHJhd6Td+1zMIpbxmt3W5s7Yrei
EOx4pmpevT53fTA8P0mh/yR1yTEcICTyw61vulJwfIRVvzPwS4SWgh0Bxv9Z6on2FwJztiXC0i7S
pi5aJXlZ2hMNr++7V0rQ/h/oYXqyYDVKFRUJOC95R4XA88+BprrUO0bueAT5FlQp+5Xxi+6u+L6z
asDN8etsMq5ISnAUynxhKJ+motjPF5KZb6T6EGxM+SZ0euVP7ofPwi/qA5aWy5u9jSdkIubGjO7f
c65+yolklPvoez/ucWdmKN8fq8HImlN1ODIfmMgkvBNBVuzvHqFag6a/gKt62prfJ5RC//RH+YHR
NPhHm5kaBkdvZL3cDENPQWFQxzcO5/Kx8+lZwCFyPIL4FxE6WtvLsM7pXvdBJ2MVMjhfNzrrDILN
xbSRTnUMXET5OpiuC3FTqGaEXAxGf2j0KXTmx+IDx86/olFY5JVqMnq7mhYpOjQwVxX62u16ROvF
Ty3kjHrA80JGF9DVgUBJ0fhH9i1U1OlxvvxgtIZ84cLaHRfY96IKFlooWDEeBOZ8cYRRRMYSUjQy
uau4gY16YxyI5JwgE0yo15etI3TSjAujuGgNA7edoICdOSlrGuEpAtlS13xySA8ej0lhSwYTOrJG
Eax8QhOnTgxmmrOJ4wbmhbioR7ZbORpi+tc4VLsIYJ+irMcYRBNUScinUvElRLeboCVV9jUyi9Qm
0d+1RCZZjBN99SehB5WA85G4zgyPYRabiG4kBMEW4No0KrT/+E1UoxY50fdLlbmf4LfGoOQ5VOAs
pm+DROFCphTt+TLd05X2AgG3p+cihTeHGF+17eu16XC6e/zLu45/z0kvij/aEz9cjI3EQs7TVxHe
wwcCM1lWBhkXuFsZ+HCUa9mFvLGrbWXEkuJ2dkGyZ5VtI7cRZ8F0vX8ar4B3aCkFgCcswLPBrULm
qdOUlt2mNpr5d06Hxs5fgY/Esdic8NmZ2ep+i1vNL8X5xRt7Di9dOWVXSYVi2veNltXJ/6rZmmnE
tcULdG1aoIbVz8cIIfPHI+COf9vMGqmkH8tW8JFYr/vTwvfWJ32CFnlUTjKiBBOjEaGU8h1dhcvj
00JICXGdnRzzxyXiXQkk6FyrII9IkXYTz+DlQCCs1lbJgI/HXEy3JsectbIxkCz1ZHAlVOBhILea
Z2BtFjWT6Mtd9i3VtSV/v76aq6iDg96IfZ9lOfcKgfjOpp1bDqJ61itjPlzK8BiSjCWxAUqDAyjb
JuXhlVX3zUxqC/MtEEcT3apFJhlWP1KJraA7ORv9YkAPEFLl41TDOaTMBckDSyNddKUCos4lmkh7
+8xyZ4n1N3asF42hR6mg2SRViXG3KKdeQovdMniLfQdUmfWFBAvGSeJIGM2s63Nch3l1rqWVWaM3
gUulhCmJjuiRpqCEsKOsRHFBxjRqQFyUv/UReCYMfzpZIcvberFwWc5BiKJ7RGDh70xt4g18m7mw
WNVUvneOiYalOrC0V+e6Oom4i+Djq8xk49qeFO/ayatjjX/64jDzCGgRJ9AjtPfhmkoSW+H+0bQ4
7DifWnECPhyDSXw4eMQpvtkzU/hvU7E6XNPFLNGkB13mCXZSgeXqm0dbUdWmtJUcn64tGOjSzWoZ
AcV7awuIAMUV6gAL7mSvNR9e9MH8GuCdYPw/ejT4sYigukgnsM1rFRli1ibAFGfEcE0AjO3ifPwv
e4KgJeftSyzaCk1tAIiNsMVO98oQFpeC9FUBceO61825vDL6GLrwK+kN/vOu0KqSvvp/SWIe9ezV
ScsMW4koKxvvecMgRQnYy5dbvcwaewU7dxBNhGekLLjNzfWQdI3/uexHnxugs6su5utrKbKAH0JJ
QtXMV1IwQz9e4rLW82lhHJ9BMxUeZCBxMH+Qsq9RUK9rlutjnf6obKn/zxUGTteAc++l50bOBO44
mTjZLFmSf63wLytVCwhcqmd5XeNH5Ks2dVlVBDWmlFZ4Hu3X9GbIk1KFgAubLjUv9yO7Xj3MnSWD
nHUMZz+uLUI80qh0F62ujlt6dXl9RcxSBBxRQdHHFM2Dp4TCnswQhuX2HjwV7DPRFhr91wlSK+XL
ofDnq7IUudVujNWidhSCiZCBbme0Z97Z9fm8Rby+R7D18R2cTjwszJcOA0Jex5zFlAHawrFNlOeS
gfhyOev34kLzEckFFkRVVGac0Li14yHjlrxTi6auT6hrvmwjgjorgdom3wv0FsmObaBN4yRuuwXS
VXl2iZm1oNxf2bo0b8MeUh0JcknYSDXiNShDR9N2w2fKWyDLvDMkSpMtXTPLNyBItdtXCZJNBEiA
YhkWjLr+v4osakf2vfVh49hi8IKtpNk8TbDxMPkdoU/g6EITjmOilQyONB6mXBioxuy0Z4+bT3iD
85P+oFl+l8IvZzA5hR7RqgcFIeNlLUyxynZcgGEn9HWQOaW16sn6WQx7NxwStsZ+Pji+g96kCH2H
jP2NUaMAvPpvZihJxYx4Ae7QrxF1kmUfhRgCzbNzXm9x2y4l9LSyd2ws1cvSfFohGNjq1NEKD3vj
ZGIB3JSRIx8e+oDPDPabqUBK2D4VCPO1LutBAlenBYeFqDCJimpOkr46tIKjnrtpEUHfaVSHawFx
Onyk91F3jHA1R2ZwyLcM6Lewnj0zgIRk4Muas4v33peh3SNGu9dQkSZPKvlwap07fHmkJ5aAakGK
HJmiPArS5INaMqdXD4SWuK3853ZR7NuI/pQUbHQC8+UHJ1RjUfsqJjwDdeTHiWq6PwTu77g/JDwG
seCgVvsPnGtDV0raURKnc9/MrKmd6MDuR6F+XIGvF4qWc/Dpn26q7IsJoFJRJafHfCcmL1v586H2
ZeubJf45M2XR+JVdfBNLRtcRgsLRwq3L2ddTmX6TSWI1HC1j5X3Pau2tf6s31DaUiU1YDj8sjpHA
BzQp79oJBFSJxjhgr6s3g5sx+FPUy0JLHPhhQmdWLM6bANVotHmFHitQB3cjmcZLFnq222lF/J5c
1Q1CkHZYFRrSP0cpvcfCvI0HnJWbEp/qnIHEVCiMs2YHrs/JIjLZ0VBr6ERCtbOnm1WM1Zik+lDi
JOIWLswJkKsM9dnUkHjfeZt073WCS520nGV70rPI7s93cOKZNCH3EyMwBPkQ7jfM3cLeMIUicm7c
UxR5s0pQuCr42a0m8pJPh7ZTM+oEjvCPKSXTquSkLUtnyYAiwx2fS4KiX+dJFxxHJKnhFcvCDy3X
Q3lt+zA1gSdoLO1G2BkzkjcibFspTOww01f2WKXU8pGxwrCZrChSGBxEDY3YaY7qw/UcBmFeiCP/
sRMkr7w6EZt++L9+0W1EkjwPztGP8MFFExjFHb8ZnqjE98NeKjdNBlrlFOoNmX8f0lgsA+4kQfpI
jOHwLsMYScM6tzmwkCJiDIVKasmZljGwl1E5Oh5hRnrgpiwrWKhOBZGyaU/0BGswc1xF/ig33vSA
WU64x4Zatwej/CL3qYTJpWbt76J11eudmgAthxjYIMCaZO64U5hjEc9p9cXgzxym0vImOP8sFFSi
Jki2wyQD/z54mRicHEkXFeUxFEGT7yLIKomn0PxBY6lIw4vV//RoC1MhJOod40HujJRhh7peEGPk
iiX2mCed7Gi+1h35cw4WPpOCfyG7mFklTAT1Vk/NYt2jmWErRRYu5OgsVIIknIE7HUFitfgLytz4
arBmP/lldIZqVRATJXZ9/mKSjL5SCRo+qT7lyygitUauYkKeJehyPmtidzJVnJJEr8y5aNfdJnCp
MVNKXRvSi7zUOjvdXw86rkT3ZKPcMt6CZzYqlhoj9lLQ3eaiXAREQ2kOUGnCgRk0jjQ5B8Kd7axU
AyRQMJ0e6rzeRM2YY7lSOKnpveBQUwiaCygXL1onri4OtDWT7OGKakKzd3T4lncpRl8zR6j7b4jE
JIAejV0OjWPtW3xV8NcPXtEhjfT6HaJ/6GwhfXqPhaoB8s69pnDcCAN4sLRkXz4LVgn3rU090YnH
ShyQ4o2HgzEj21X1tRrcCGuMZK1XQnUplz1E0ns6UCkA+l5iF1PgvHTwtmWs6SUncTiBMdHX+Y2o
VRND6Npon1/2jmrumlQVplSEQpt6pZx9+a0tI/fArawDTeQVNNoJaiFi6KLZ7//iP1dNFadc7SR6
9122EvJZXLOpKoeE7CvNuIsLwhNOf7Lilh6Y59U9g1/TYopey8CyaSEgsXD99FG+jSDRcqeZjqSe
yx8WLVHGhDjNy854gl+ql7GAQt7GkrBezMkB+E3fpkPTIzeNDvgWPOcKqCW3KnpvHiIEj5iqk13R
GCU6PBOWYGoVayyw0ffPepqkbYptxyu7d1THiQ35glqsJ+r2wdNUwi/A2oZ6o60yMxz/4lWPPb4V
bEiR7Ir2UN2HxUQbnqzLcDYkCAgQEOFi263RPdMXwFt7bsFyXhzTy0IEmFu7wICpGgLr1X3Oj2ka
CakVhCci0Fip5M2f4X/XqKVVdFre1hXAmUu/k9J2GjM69+OsEztZ9enPGFF2AMUvDpFi8Qh85avU
Y0H2SxEQVL52iI8VGHc7KA0ND2BYW+lWWcpueSOrcV6ME+GDyUF7956w9nKCRQPOiEsEeKjn7wDf
Pxmx5kn1YyqSMR7ZlMCotZ2kId1lFH25wOvREpl5lRCoERHCF9AgDHEB8AGavlutmvAxQV4oHSKi
AF0Qvc9ft4jY09ZGKr6nPfpB9YoeLw8lv0rcPPpn1c6nhLP7Wv9fw7x6sgAl2OENsZj+BV3SJE+X
APQ8EZlHIx4T+B9nl12XJxz5DEW1JoKGGkWCJ5w8Pdl9UXr8+AXE/83Oyki35xxOMGJDA2eNjsIP
eRFj65pcBWp9Rru2TqKgbEstL0H01p9Y3WMrMJCoEKuIMhtxxyD/Maf6SCLNkmfrTkm8diCWO/Cc
AFzM/kI7QGAuIhAS4GdnD5CDZzcnYUaOjLpgvAZr48GM3Cm7dg7rAuA3kEbV9Ug4F12UXRM/ZGcV
/rOGMMSonzCw6JtET2ZFutWxoor+G8UF0UXwsGsnrC2TLQM8iAygvcqE0Yc5KMMvBhFcnyLvDFBt
cIGncPPCOpVYFYLCaTvr6QfStr5qBJ3V9kGVfCc2JR0xoNcfCEVvhcT+1l/dClKtZnBgl6t29bz0
3GGw4gm/J+AIpZBCK/6uIKZFcEJujPM4l8/fckxXf1ZYxiHJFwhV9kv5RJ+Y3tuzkyA322vegu3R
+YNFZvsb+zqyTP/66PLEA/NyVbrJWsFbweZN66keZ9h0eJUshTne0n9CD66XhXGGI5hxlfL3i/Ur
nb0w0jzGqjWqipM2zAXJkaLtAyW5HYQ6m1XxH/4knyxNUTLo8yVx6LK/S/MlQXcMnI2XOijzf3Au
0TkRUmY89VY40F0PPg77RwPfOkzPU7gkGy3u3pRkctwTGXYF6o8yNQmbb+dgWhRSjy446LYZ5mRp
iaOmRWljENTzkVXmFN3x9/sS35QrBZ7+UH8LfF4rJIZTpPAUmbA2niaGPRczqDoZ6KKPMmz4xazb
PE/E5IIBPzKK/5gctAfaxCvwuLzeNJURIkeWaj7P+33Iws/GWohZyenspVk+L3MT2Bh5Z9iI9STw
+QVHXwWBinrBC1eT6LxUSecrfDEdWqO5yiAtLa8yRbOVbgUkGbi7f8gZbfyyMCtdgixXXvfAyNO9
OZpboISMALvYM3JG9bwUsIQSh0amKNRERJsmiL3JW3whHGlXng9pIjeEoPLFPQOANKq9IxbfbV7u
EYQ5UHm4+HjvKKYa9eSa52/hTWW2v6agPR2Jkw047zXxzpMy/R8u8zRk5r4h24sKhxfWUzS5FCVb
giIzA5vzaq+ncQsIh/ftscrs4TZEnO4RZH2Xi91z9+nJLOWCQ4XUo6BC8q5Dan8prAyhpD8R7WUL
F3sqzAKLPeWsFXTEu4z2WITKcYusegKfAVB1VrTvA4g4JhPnPMAR00VwqsDfWa96BrvCdLPJuwKB
r51CBSLclLwZfLQGGdmunxskA/gEJSKsNRnBfODN8luZJnkzuoVJAhRh4wBYlvYeQErlLX8KAxWh
mLTk1EyLlZ/bBkLIKIBzTLg59Ir6+ik5SvRDyjG8XOqlAFmDz5oNseE5Hp4PuLg9YeWX/v1S7qo8
sYAHJ34JNNFVUizni9k7orjYZxTiUHP7aG87YNFmo7+wYlW2LRcVBWqH2kcLgtDVnAmsVDCeW4oo
8/bPhXRlQSq8IwuQaOOsNNGJjNM0ioB346iWavvO3fVqvYukUc9qjPzkZ9q4n4KZy6idQCPJH+3k
rN0fgmTsKeMIriV4YFE8BswPk5nF7iI9PiVqRlJBBKPCNaBikyZajs2soYNKWL6/7nrLB07jKOmw
G8mKaM/soUaDH2idsDATVLA8OuMj+nk+Lfck+P4a27vipoufT0wzA3L5Sns1OXO2s8mx13bMSWxg
I7Iv6FnQjpCV4du4F1PnX4vE2VH0tEISYwC8C2pzWLtkV7FupG8fIEk34/FDypKhbZ39LCBcE5as
z2ZtQ0nvW4W5slBco0m/vYa2Mj/BkMg2e6QwABH0y8cn5602vPghPPsxkpNVr/DdWzG97iTY/C64
MwNKKI/EfIHCTPnQ9b1TtemRaaJQzj6zNOIMPjmqpRxyaXet3celn+1MW8Q+QLjzuaNNJxrSFCJP
f0Gzl1CoTfL64NDyIOz+vZh0etSoRRoWhcm6vrtRVFua4STXGTaj+aSB0RVBzy9wVyLxrrXQKhDh
XBSTGJLFBUl373BItTnaqLCo9blPgVBBjzPdVby/NAjHwh2ziQHZOkOWIvOYeQ0+OIgdv5E7TfHA
9PqNb5hIkXENsv1wtZpozcXhejNn8xHsLHRsKq4QWpNSQxwWHIMP/AakhLAi9oT8/jcTrbn5RbZU
yg2WGQqGXZXjLyFbZwp61TOBieqJ/dDkice2smitkdCDI0n8AZnuOEHsK8qSnpwF7q7qUxNxH1Ve
tP7jG3c2sXVE2RdHCYqvbo1gXoVVdrQmyits6YVR8cJnJnxPPN5II7ZRgdeNjwu3+By3dSQXavFG
PPOPau+8QEeog5A0KUtCi9WUyi/toV6HKnKcI13ACsXOrCz8TIBHlXJW/0YwAoqSu45/JriW1nn5
iaNbJemODT1HQvSbXfzRzPc+I60CXAqKWqTcJORQgQAmQfyI4MFOeABZthqTQzoUglFR+iFo0Ib0
zOBLr/u7OkxTDUokNAX3o0VDFnVZSKlSR5Zke8flgqKF0Nq1+VNdQS+2SKi8QcNqTH/bM9pHn55Q
x655d2jMdQ1u+ZyMKrlibQfcetE8fz0YVYsMIWH23BIomCnAEbllZLxJg7HoydNQK+30rl3WawbZ
PGURtd+8p0X5m2BGirUrSz99UemTC2i5Av0wc2VUtQ3axyLdIDWcCWe/v04Qiphuc2SvTIHWRUHO
VtZGOsTp5WbaCKgMt1KXpZdKbxu1qQxg3GvuY2oFNOHeU7DrRd20uI8fEqc2RoubK7zt022/qs6t
lOn+4gYlz++LqB2wFlf/XM5VonkZ4q5OZsIvUjnTdKyMpyOPQ+uP8r3LEcK/qMnbOEMtbu0ogVws
zc/3yQ09gxeNUgdZVNGJ9jneEKXSgbOmaiXfiYTWvwEHHXHWRM09xcizzarjaJGkrzmZfRwltZDx
CZATkbv0JH5teGqBfrWxDwL+k/2UhRDy3Wh9LO5lsVG/dDQtBqgTvPhwYpA7aznEsSNpXRntXZGW
C0H1b4GldYm4vh8FgTyfAjlbSeRQCVktLP6hcE6v/bJtxKOYKouh+Z/XMIxxjsNH7ADDpVrvowxJ
EBhFWpQTrPCtvJEacZT8MxhsKTcb1xnOp9FaVtekMhrcfmr/GoGiiQMcQ2PZzZIzPpZcvZ6ffCiA
NM+PGf13tMKosFHfBsFbzj0aJCnnMZCxKaJ39Tbya3irKJwDB5fs1lAG8N6ICr08KVm0U0kWPGrb
BRSGgZTIY5uNcN2cZbln3W87lUOzUI/GDxLZe0oEaJ15BQJmDVmkXHIdW4TlxQQyhJXQr9uTeu0h
43/HR4FpW3U9gziR4l9uEtyV+KQ5gK2yHegjbbKQhpoZX3ly7e3cu8J1u9C/ahCkXFOYgDjsPt7R
VojoBBwh95eRiaZ2xzrDpiGmlqLR/ZBJg4GStNOxSJEWYWP6p1WUopU4AB/go1n3y70D5AQjZxFy
iki78eCo8EwTGoWjcAU74jJATudmr+6o7NAzNPt3D7tmTsPZGC2zJnGIcbwSb1ybETjBBwrGozvn
dmjM4jWDSsBbXynr7IShl6SEbhR3IKoFDWpnDhuJ0IACUlc3gvPYoxywd4T2yMCLj9+/TFss86N2
dtWiGckmJwO8uiSeUt0ZQ6zqSY7VTJCR2f8T05cMi/PHni2/FJX8aBBPtf5mguq9iWTAN/97rhXo
s0zATmMqjKl8QvaqAQxUT6M7em6lsS4aBtNTmSeu5b/bTZkFSywI7zqLkBKpI6GNfFTmc0z2Ux3j
Hn3kGpwSnfsJWCCOeyIrDt9DRibSObSXsIOTd2g57NHH1Bsl6WJDE7yj3jJ87ekg8uSmWJLg1CiC
E+8ArJ4e13/D2jF9YFEhsQTjOjQSZgkI2US3aNq04PD3dHqF2UUu8Skot6XiOfNtjDPphc8tBL5I
o6WMqNbVeQlXumajoQhARXSlx2J6QYQ9A6IcPFgSQUKgXgkF5agd5cRMD+KKErzFPsNNFdUMYi/p
QJKjsLz/il/umbIlsvicbK8vdDZ70grmugMtMOgedaryezVJFjO3WuFTB9Q78smD5e/DAcC6LJDr
l1BsLrA+2C/2ZlSkHc6k8QYEvSZRV6oUyU2uHMGyV6EqaKYGvd4wVDquixsZ3Rg4g4EktwNaSt+V
3XQ7GmPutBkY/Qv6L1gJwo2biXi49NeeS4Qc3aKE4uH+2wZbDOQmOClT/oNFgdfui/iVRDxQ6/0o
Kkrh1JBLFHst+Q/cQfaGI2KflfNdbzKRuKn2D+vxncUY2h15ugHY9kerCCKQ9GqkvdoR2vv2Lv37
2iMU0vkK0HWS47AY9HpotkInrh9ZH9vmd8UqCeJ3Fy7RomQeac0JsIIJtSKNu2JRtcf96CZOqoEx
lNp/Bmtcupxk1WkrlY5Y7evqVvZvWuKMFM7A/ZtKgFolKWUwk8LHPlwF3MksxJ/dp+XR2/J+Tpv2
VnAJLO5o8oI52EgxzJFYp0FStA4FwQ7O3oXeYu1RaYjmqvnff6j4m8F/qlio026krqJ/zofmDAa2
zEHqvqo5DZFm7r7aL8922KHnBa7zSeOW7l4WmZH4W9o5Tzyp+V1LvacMaP9FVfZKhqqIVC7ybA1m
+F/IkNwJUc2QG8j+b5x7bWU9+Sdg6r7SaE7ijCM2NA08/zMFqoUV4qUnoO9ccWcDANPU9M3qKo30
qeoh0m/yqwzHWgyQRrnArHRxi/XAGq4NFuW9kZ/OpmccFa/jZzYhLSSuwiaEtIFxI0ZNvJc93Yel
QA+fwehckmfYeGXpw36TW/kZghHjy3ynnBva7M3msFaqUjQ/2383/0uYVGdVrHetSAD4GJCxTYNE
f0E/xIahmPap/4FuZv+btkgI/Ce5F52as7EeppIGq6mE7EVmCim7pq2ueeESZ4U6m65JaNpZz79d
cD0f/L553LSvBSdQ4QG/EDO/INOy18rUZFgd2tMhOKCj1hsIGvCqezaaZtPeoc3c9QNFW8R8gErG
xicRfEFIyc/WamG+s72jTalzN12orhL3A2e3jsqh1I7R8HiC9jANLhRif6CO3Jz0mVevZr6CzpLJ
/lrigw6n/YMzj5Z6PD+OmaZ0gKL96CIccKJWdswrE01aPL2qOopKZdziXO8n0w0H9bJzbQq2/IbI
4BsAEjMo54YyL4mOHC0PFDGuSrfIXr+X9vneu162JQP9AV5xY1ddC+SsxYSyyTIGxGoNckl7QEip
JjoTZFRTRx9eNGxlxe4hpzH+x7dMKy+YiV2yjLe+7Cwn7gtPLzksc3fsvxJhGGQSOz+L/ytPPm8l
9+MwrsBE/R1M7mteU5CcVDymUpd2iw/6o0AkjAirk5H+9tGBC9NKP2VqVconavwwtxRskIL/uqwf
GyF2eVZ8IamEX6Uz7RK+a/sDwMBtcAKG/pXI1HA294gjymmF+1OWFFPBEJQ1WOtUt3m9lICm3yXx
8xxfzct6rHDxMt9ND4/4U+4vwSTicpUTSJXB+sRIuWVZ4aUKGWJOiquzBnw1v6czXzL78Gkvxh+p
GHPrh0oOFcBBVQBKBZG4ldg6XELPK4dtcEiiemOX5PfXHIdeQcAODtE9+w3Bnep3V7J1yYg59CCM
KcKvEdTXEmz3hClxEOZ2RO+H7ZCoErCuSIzvaXwSQfTzZx1s+dTR2kYCH9iTve3IZY2aJmkMId2U
7p8ITq59iu3ubw5F84gwn2ESPSHkUBir6e15FrN/o9gkEoQQEBTmb5h7Pe1HAjHG9jXTtvUH6ygb
KwH/XjCDeoBeJgCMPIQlVqEM6xZx6WpUKlVKLpCUX++it/UI6vbTOcIVXZ7cuYh3F4j54nvDYdZK
PCb9C0sOCVmEjyfyMrpBHbM8kzxFLyCZ1YqVDLAMEpV+nJLvDjmV0g0ERcI6mTawsNiGjIvf4yiB
Vs4GHT2+3AL/Nt2beOw1miSh9b4gCmJ7gTYMtl6QqdKhyJHqmBiQQPMgZqvaKP0jWpLsYE+KzUn4
V7FEc6SQlBrVJExJ5gr9LLNrLfU0z93fhY2dZPgQwXLFRifrE8qFofNHDZoj36YZUKpOSQPe51mh
xXaYgU61bUAwlOuHBmJyJqwF/RfDjj3mpUA35MyDh3Y5B3ycKFqr0vGN6SU1orXMsHp7FrMA8cOS
a0AoK2XhpDWZ0ddTwwRRvCgR3ApxEeRUxou1FWFLY9QtMbUan3NYQLUUk03B3cyuu1sI+HZCRQDm
sBWBoU2BOZnuLUvdAj+oGiE2kEQswjHiFqorB+7Fucw+MA1WJnUrFeHjSstbMrqcGhevfj/SF8wz
Fb+SIPpjvj2XmK65/3Ea7A10OyQ/XSTiMj0a0g7WosNH2Snxi4fpaCCfCRQ90GX+zlVfRwPUw+15
ySP2vCUhzhq5DbyJ2fnBT+dZ+FiwLufMqtOM5v+GpAAqKS7cw1o/V8B2sbGYtXHLf28Ujts3ghHr
Cc2kPpZHJU8uGyfZnqcxcM5kT6IOdxuq6orLP1LuBn/OOYJ+RQRcGe+9OJ73+YFDjdkzNMJnUDeC
nSEMX2s4u5B3ZXglBTzrV1HxA16birydV0FHUiodQh7NWtmsQwgR4EGcce1VZ+/nuuRrSEGvgR5R
6GUsjsh7q8WglFamTK8fCIW7lzvYInLnFm16/Kl1FgDfo7q+yAkhzv4zFB7Loss5rNgelQ8uqvpE
KY94A4Ddpq0p/ZwSERV390/E/6AVkWqxtnJVSMkNSE9zCOXzBLaPIT4ZP4/7BtrTciJBGlgJd1hn
rmiOfiiiVwGyiSIyzcEAc22kLT11meQmTjYkLoFdIovP23wum2+vp2ni8Ctx54okATv3PiJFx0rm
BYEUE70QCkPCWnKpSkLof+w6WDpefxJYph2YUnHVTSjejM/l6foS77Fmtu1jNOSednjyctuGvLp5
9jvQMEgezdZIqrGvEuSbONK4z8XhaX9KN5Ek1NKF+3UinZ6esKh3WKsnsO2TRzoz7FYOxx9WMlFn
QpDibxI110ALirF1VIB63U9j0zMQ0jWxgGMDZ3aemRCycJlwOU1J+J1pAptbyXZqmKFUQJYip0lB
4HYOL1UKR4hQwLzhj2kswUE3+U8Nio5QW0pMK1GWPqUdm/Mez24Z5OBnTp3du4J39LTUojNmsqZH
CxTglJmFUGkov6hAbxNTlRfF770OxxwGccPJplsnMvTFFp5G4vMTJBCFD7BcyFVPIVa3zdUH2PDG
GoWFdzZjnb1di6yTE4YhM1en/VnI45nWuvIpQp6nvMdEiqQfRD7TkGFvSfWs3eNCjlrS6Msk54yZ
qgN5DOD4dMsfyaWjHms10w7x+QkUCEAPX0uWVoZc60U/HWKOkmlOxz9Kej0itN8widaZtOnz9hXQ
6ldSZhmb2QPggdDEC+QzHc2NU2KVlqtGSXQGgylYK351BEvvyDWBdFGjHAWxTITxT3GlJ7C3lmVe
QvCgpFV66piNB24w61DzcrjpeDrXVLmecxMuVvqS5JnEj8EtGdvEJ09DiNexFkRkvAkYvsD9faAH
E2ZwPggcAMz9PRbaE2laVMoqztgYFndar/VvoN59mekw1dUUDrvwt9nuKgGEQceHvzDE8H+8x25u
lTslQB02D9Y8VHydO7TRyewJG9iY/HPB0ruCT5xF0WwJGNqBCUSKrWrE1skIBA75D8me4O5wl/vx
4LJemctvquvoDj7LupeWRO1YrJPKJGZfVXrV/De+cf081C9XKPzghIPe2+Udq1//4liTgjz5b6zR
9cUZRrt0aICGpEF6gxhC82/45dbcjlrAO0Yp0JwdPRW6TTzn+qvYeum5xMSkxkoVRerhZJiC46u4
Ay5R5tyac0mXq/jZV9PNrWihL9QNsGnWIOAZVOFS/htbx4RS5bSc4nze7gGRWHL1tJwsPIrGmLP+
uXXLqB2aaLAzPa+R67/1SbtpcLAQkdlggR5XAy1gR03Pn+nIbOK4J8RnsuxVdEhNtVSEat8AGLTL
Qm6Qbf8rYAI77SD0QxAgRHO+vncVCKv66XSixxlIp8jdOcfQbJVCJMclsSinmVWfIAlzGiu7HVtZ
+uaw3w/X+Mfx9jwMcvBMGaFshLSWSk3ErH5Gt8QQpK5/31x8rQHfFVd8DVdsBc+BLWElxwJGLuN2
HyurQjPiscoln1BFV8QEXxYb2yHfE2+AsYYJIf4kRhVNieywAwUk/IEZeIyjwZ/2O56tqVKn5IhW
ZhxXr/QXFTQs3mCaGZIwj7kzEkMUgzsOi+kyfTFWs5upMLvCxU2ufGvXjUjg7sVKytPY0YBj7y7R
joNCJGIQXuCTusFgC4GgHT6p+0R2BuI6XdkEuCQmAtl+I8G3hzr1W2lKjWjHHd3ExkfbixaCj3y4
0GOMmVkGTY4R1a10mo89mKPpH5f+UFo7D3GS91O+oPH3c/YCv10lH1VGTmWeXuK9C4gFMQ8QN7xr
buoeC9axj5/BgQ6P2f4fsH6ESr+LE8BxIPBj71lPU/sqlOifXt5OsPIMvc2fTNCSRBGlsZ4h/pRr
dN/dgQq+FkBE1qS8iV8iT40JRxldxGsiQFpTIC0mLWPnPrQcfyTr2KqDeG33HHEFxxeZDFoQZpN+
s33WXfotTXAFNqI3PLR4oUKILV8o347pTCnBpPGiei7/JeXBzcKoAUA67rJIXYVe0c9Fc/8ENCID
TyOxxQXrEApD4KU8edRqGhz65WqeZEhRTYyyHZSiaBPMd1pi7Io3+QTe3N4BlT/GIpdB4CBlpzDY
jmKeANzanqeZwbgdYMyAlaoFMgl7XM5CFUec/rLxjOhb846FrJ9NEpoZWYJJzBelwz15YAelIatc
Yqnyu0mj6dSBUupd99kCtgqOKtglfLJ/SBkA7+H5ofysHmcS6EZDHjhJpf0KgcRsv+xzpZwf5B7B
hqtTY7B5kFSfUvHtmG3QuUnu9vmOUEpF+7q3Tk8GHg8WhkZoeMzT/c9EeVVvVV/9jiyU2wss6Nxq
tQ36U0q7GlNLvO/u6+ren9lIKvWnJlKoiKFgrlYlpHmRCbrFWGNrz7Wp8hJi9OyVIWbnMl0Ybj/q
6CNT97Hh4grgYWYX5OchBMpt30XxM6QUqaXoajoUIerwz6vY51xCe8zs5ACtgoaACZ/6xjv+xoMW
u5bDOC/O4wXL4lnEE2cK90o5rJtPgTGfix3xGz+7VG69jUlLBINPfMC1NoH7N7Oc590E2aW/DBz1
7B+z8ZhmWHZjKKHLHPW1YNUyaTv4V/eGq1sBC8HNIWgHjyoUL9VA+5P4YdYUXk25s7ZlP0K8WKIu
R593QVqnEaV29T2Var3DsGX6QnyM6Kq9SNF+L4Zh/qUeWbnaqVhMw1wmCBi4bZhcCwMDdRd98TRh
0zwiUuetNb8teeiDe83NYlTQot0VHHfmrURJcaFRcd4zMEeM9kwjyinGCtgdgyEnQhy3o0lHtf1r
lIBBQX9GH/98eMmDZxPR3RbCT7I4Z2xwyxhTmHH99/E8SKzdB3F6+ZW0fbMTUCdb+HvhvSFkur29
K9Nj0AKntuotwqR1ZyZdgFfaAyXWCvJiXRsWV3uFNS8qYoEqPVSWFLoyTcB87J+yJ0uFKrtIT7cc
u05my9w7OH4u37hDmdei/t9lDeEuRSHYymczkyQe1nVVz8gFCgshetQp/r6rr1q4z7RaEdM/U8HI
FBWx5EhB9udG3+wbjfcaVVFqN05F1bs34MEfYt4RLjgpgDXgUtBl8veotzFOsSDJfwXpwYr6fDtt
5UfWyWMmkkJZanmyOTfiUkhAYrxyOcRilHqKtRLQzbHESxWPiOUdc5euyYBh8gJbKTeunuqe8fEx
bONTbHqUdDKQcZ2rYtwYJubNEmrJjHCCdevFWofAUWZrXDW7AGj21mXxGabRJMI6inK/GojmghvH
8FYIvrH6a0D2ezfvrTsIZNye20UURQlrceT/Z/RLRUdGUWRRTayetn1nhpe8pWFASoRel8//gKot
44APgF67c7pqmI253juZNEsCCnp72329NooW6RBVepkmNhY/iEIgpZ+dq4WtwCjuRIqdus0Kp/Y6
yTKm6rt3Iak6UupXGibQ5Miu+huZllr3Sn08PSVOc56g3enXjv6yX7j+x8WjJ7xaFPQYDlbliyyI
ScHwleg7ZrN6JZRnGmhjVXbQGdOcgEugLExrZJCY3jE/PiglluXpU44+UfjUK4stPW1L+NSNcnH1
VQcFL2ibmRMnkETG4yoNrBqPI/vXJYS/JzCJsBvLU4GBsgdwSOiVqzfJHCXGpGIThGM3uxZNjmtY
L90cclY0gMf0HSabIX7ZInNEo7Q6dl8ckz0doKqN1+N+Q4i5SEMd+aCijtb2mEHtwvbg5L9V78K9
Ycm803qsSAHRHbeofCdeFM906ysEszfpA6kbnIAuSDnLjBRfG1iTzPSwxL9mpjn9i+ZwK9bWbM8v
FbzgFqWSrvPOQ3a1z1EbRk4eRSzEhM9GTXRodFWCybyjLqq6PCHXdBJ7dPbJ1JJKqsK8vwy20mhQ
kFZrfhcVvgSocz0v/229Ak/NhzTNXCqhBlFclkRWd7l+u9LehQJ8S2WWBwyOoLyvcaBG/fcadP8f
OTtouK5BAG/9AIuuo5wjEZ4KmQ0slC4tFxRTRDMCAUtrzLCmBoX79x/s/Q/4/Ix8jC7bKw6sKTbB
/HBbnZJ2puJaO+Ssk/8xlQdbzX3TEbnEjF9Z1h18i7mU50cEmDEMbx+pDhRX8zpiDaZRnrnxw59h
YqVmFrMuZCc9Qyh1pY4WG1QGU3O8uq2sSyY+bA2ysfuXXfI8XQ8kkIsusWl65HuzBW3ceZJ8DC9m
S/iR2SYuAgHJT0iSIT+EcwE1FR+8smkDXLoIQYFzc6uitiFdVCWzERL4qqKZkndGcSta2ZbzzrdG
ed3d8DLfsTYH3op1qysCAcuVW12317BLgau+3RHiJfqkGiFck7CN2pSmFhu6kDDhdsw5ctoP+8Z8
ckpC4+oJvKhC5+WVSZv7gbcncwwICjlOun+ETWvNuzgi+DHpmdkF08nmsTfdJIffVbiiAzRkNZEG
kHRP9XnbTOJsZ9/G5RCOCF7imjBWkxPu2ir7AFsC7bTwTLNhjaTbcU+HCdehvKQ4glwTsVfGQEIk
/o3TdDSbppS+WNGM1e5oR+qYuFILRp7QZEEqk3vCJ3bjw8zoPoesEIGlPiABBW5GaYcy8xQ/ljCS
YjOKXV9sNM01exe0vMZ4Vfas6vNo9Rv24ocTfka/FOyaLgWz1rnh3hee4TNEQmILycL4YweGikTx
9YDmSjLKKIWJeS/jmbK4pkc3bIMqEHf0XBVzwpbHXRdSkZY1rY0hLDHzrzDu9hqLb4uJct3aWe7D
BWwJHzkNXrm5RFKlo+xK54QYT8EkNmZv7HcKyz2JKXK1iVfmAH9DkmFrq7vTmgHCAhxeuBPoI/+R
unKCYMV7dsTrcjOW9s84vFMtQf0l+RUN+12xtDS60Xllf23WD3yN8o+cHiwLxSFUb4gVyXQi90DB
b+OCUrrkBQzKtiLfxfBo6uPLt1W6n//tav8IcZUm4M94F4c7+K6dpTJc8kuYTOtnYUgCCrtwP0Ef
28mEm4PkYqxI0IMQ/aH1zUFJz1fpaFEq+r1BzjctY+fmkC/iC/YnYCiUKzd5VicUzc8pmmgemu1h
xmFxJSdaa4oedHP7EO0dySmIijK5KWVQMU+fq8AbPC87FaMO/rRxAc0k8m0Z2KFg6WnXITw1GXK4
fI6cedugSSFry4ogGUjZakY6VfFMSYW3FgOMDl/YolIhEtfcTBTJKAISNhDtFVfVHxuRdyIe1VQ4
ZjclH+dIzv2ub7WUO+67n3heOo9RasnCEYOO1nSq+j3RqQXB2Xq5IT0cJv34ICyBF167YtTdNJl+
wbJW3sfhKssreJjSEnYwZoxCKETDuVThI/p+X2k+iPL/UMDQ0dWFNWqMaiNwlIRh5n+LGHnMhQbs
6s8kjgiNl2UIVDIUnoBULnfrpkOye0Kj4KZnX/TV2XF79diRzJggGodRd1c3yIUsW0WgIxyUPv+B
/32hcpq6ylHgmslzJnt3b7C531gSeYjQbI9g6Fjt+IAnLFK5fCmQtfD+VviGSuc2DSFeNeoRSTg7
eTdHR2hNA6REvVQOhZeUzD+7tvhT9FHlb/e1Au188fZZRVNUdIhGSE7QVqykcgVxfoS6P/vy+uZ9
aWm2Oxm3oLD3HWgZ0xzcn9JxN/ocVFxUE9mARMKREelrj2bTl4eVPQYMhJw8LnsNSdwDsgCf0nFD
5C5tuLNTH8w/EYOXq1d3Uhcz4ElwJvhKTHj+Wg+wFpcKY4En6SSqtcmKKTDDxJR4HMKBVYMcR/tG
4VWyOaqh6e+f8BLVUdfecvzdUdlYEtF9oNL+c/eoTlhXztmrd7KRK0HSDUyRDGdIoEbqcYu1E2R6
dVYOR9ObMpiHhvsmaPK1POXwxvTihNw4b3+JZxN+Iw+x+vBkWhClEof7eBpIh0VThYHVx6YdaWpo
LVbB3GRncEaJC9XGEwJXyqGJMOq3UPcEZPiA4H47dXZJCvcvcndoT/f9RzfvzxkqhnTvJuT/kV9/
EMvvVJx2EVvQVn6eUxGst9K7hEnc6yuSdI4GMGB1tOYghr9/KANwhAlRu1K7PuhOfX5L0RfL/+UF
PtAF5izO7KilrICGk66Tt21psVou/rjArzKhPWMiIHCDYFkm4bHG2c1z9TnSOjw/os9OrZwhd/9u
zeZzczWqYEodff/yRuTWFpPlD4KQYBKjTDD+q8HVirrsbOvxY6tW4xbg4ZrPA6dPD2woIG1nisbw
QL9H3u4AFjqorZiMNjdYURS2I7PPthzVRJ+caQCKw9UWOIRsfs3DxRgiezfT5blH0h4mHj+eOzTf
R4sUJqjOF6Bc42b8LQbL2/zE1xI+5nqET08cRgY3isQCBWRwPXD9hViHK432yGybhOi9B4ItuGmU
wW56Vzuz3GM16SDvFwwIUjigssTtOvCc4jzWy4BLchq7sOV/KCUouabCEC0STy3KAr7ozyPd6+MK
1xeGtmxDQAetSgWWj83t8j+bXdASOmxlOJE0+7MKM/Jw+wFf15VWqDgFQ0iBfuD3eeqDUmwuwoPe
R+V4dE/yKppa15NHMSmg3+BnjzVpf7tTcTF8VCEq7cdEj+IN2T+PWsdD++d4urwukuCYk8MMOpKR
pcgMnID7HWn7z7nu5poFU6WdtzaPAOC5H4469+CUJ/7OlCv8rK3pD3DT9zIWF/1xCIx5Ow1VgwDM
SMhkvhby1VTxSl7mQ0dEh5N+opJy0EhyFSWNL6+8eVtXyu/8z40fdZl+py2Ydi2h0vCGfkX+zK03
Jsx0reUgSQs+d65bGURlyaxVLRiE9vwjseIU6P5YsFkAJ/S4TOhPQZY1SeJGlHer8+vTg8E/y4pC
VkMfifDCRboIPUqo48mkQDYu/bibL01WCNmcDk4mNrQzgLh/YmBI8nraogHItRb0xXIA7Oz7Tf41
34dj3ihwfo/n5m8NSpwy9M5dF5BYpWeMiHglNx/iIsZNXzFGveIHUJH9XWEsqGXa156Tvs9dfrNW
CLjzfAAoowESclnV2Jke0oI4+OO6Es8KHRg/eZwgtYrD1QxoePswor4xcVKwNAorMI2DcI1NMZo8
27eYtGIfoq8/lNM8AV/UYz5rBO7qLeQcTMAbLxn3Lg4Ei+TOUNdAObqDbONfyafY1sO6/SB9Sg9P
QB/zKbwFc8A4vrypVT6QGvyWPWq22kl6RZvJLdn/OdOboL0ohSUcZ4VgQbdA6FM22qwpAb3kwbWP
nZG80LV8o+RnFtPuKExFT4TMf3kGP/eb+cYBX5fFAKd9nkUgo0mVqd6tzIU9RBTqdC72FV21RQDW
udNfXvtcxiT+/ngc7wjfE5JpHXrEWZtTulj5pN2Y1mB4d6hfdGP4SslQO6Yn5vkGZWjD+MEA30EA
I8UnELfT83kkedqEyhovk1uHQoII05nRE5i3kMoTfQhUhBPzbEpVbC1JGsdsqUZWq+W7MvGi8IDt
Q5vmUNTYBUA0M83T19J9lBuKUbS5UePKMI+SbtipW+TBqOsxmzta5UBvlN+VC10z9q4jD5uP1NcI
tCnFUnjesSmoShkWbZF4om/1Tm5vV4XXKJBliJDCq9xsMQdwabGv+MOoRaBzwXVxuXyZWWXCcS4+
uKOiHJafWpIMy+J91N+gKWMiKwjKr8JTrFl+XEWsWq1iNs4cf7LeYanuv0qVTAzjyPrXwiQ5nfgJ
epoNXlvDPcfrnUgwOdtqc+zjzvV2U4V8LEjQqh+CCq6YRzyAFmk53SehR6xPZ4p9pATixR3auwxG
QdPCoM8j90tRaYP2PFbAfDIwKAjLTWrQsHL3UFtQJCdgEn8z3rvGd0snlTIAsOTq5KvJzN0MJjpr
Ir7NNNPXZdryezDCS0MfZFgjo0bBZ3h9KaubU16treYwQ5kaOoslZJb7rfrcRA6e3iowTaU4BYsE
SkOF6JDXLVMlFyrpLMIV+SkMlZdhfuEEdQtDAXmEkoEeLrRvk4h0b0vf/twDl31eMEpbuAEKSGit
JylX1L7CKrKZrfgDgKM/7IJWHQx0saWN9M4OhxISIYikRDeoMv5qqfmOoJiLSlRXVMQ61qfCvhIV
1jFFsRquukD5SkEr1r3VFiTf9/lgQba0dS2Kgc19adjwy4Jb53rYJa0NMPNfwzeoTbH1tQ4qQR+r
O7PPIWKurhbnPRicQA+R47VFeXb0UQ/rasLjg2G6wDrotou/65CRirsO+u3aLy87kbT6TvfSwKQ/
up+Mh/Qpb3C0whS/S8rihLxuSMkY4zz7G/yPuC45wsib1m0VhtGGyrDgG3kE+dVm0lcfDn5AvTep
1v8IDqmfxUkgm4YUSdKxR8FLpbXD6OeRrzkJD/mozw/uRKNCSyD8Lc4iYE9labAhi9ZFQF8M3kGY
Fv/Ela4fFL0CNa1US/IgHnEGu6uk1wgMsJ9urMKy0oUBFuzH8KVVFllLlkNkiqMi7eUhfHzROIfr
bLj8JfPHfOhgc1cihnq1Te9BZ0WxGz4GH3v+/hIheUa7M5pzZefw26ClxbDHosozJhz3/ITmaNeC
ffkznVJlQC6T5eLNc2VAcER/bx5AZqmjTQMFuqTqFw63eqW1fcCUBVlwzzzKrb2vU88TzU8PRrkQ
F6PHTIqTWA3yCTyCBkvUYpbMUoqBXDvXiJtRZgbscP62TiQ8UBl0N9j/Cmq8Py4QvW1MdqdP11AZ
V6mA29F7z05E7Oruw+FmqfMVcdP4A13KwZ4R4YBVNLTnBVokUJI3tLD++GKXPhoo0TUex0iR2P7G
49/G4xuhpo0ExBAvi60C3ftQkFQ+bdYO8AJKE1jWR0ffx8uMIbNByXDjCOr3OzgFhf3r4tB0WeBe
pY5f4JPbeEKRljj20SwKnJoLHu8Yb6nYb8ilkyJC/lKRRjkTdk7ugd46dKtAfCMirKgPhBPU/BCi
MvXvqUozDztrsolAFANSIEhS312MghY9mcFCmzrhFyQTMHRdogOjmsDSn1JV1+TyHwTsSatkrdtt
0+w8KV/zt11zYRigygWAwMpyD9b9bnS7m0ZN6iwhXiVByaRIxzdqBCSeOVv1h7CCoBltKP9Ac/gJ
gqqArrEAgjx13UQkdkrgeKp6haawLgS8IL3kgahOWi2wk7yVBmmNxqUlPx8J4zmiT4aWPiqxj6dE
RiT3Sr488BbxH6t4qPtK5QpF8Wifx98sCorVO9Ig0HeLIsXGGV2uk8NX/kchskDxPSMACvJ07asR
+qPkjXM0sdafi/mxoznkZuGiyyJUL5ECsj4qGjvQLqs6MbPC9aaRSfl5bJnjYa61vkcLBNBKhKGx
jBdaZf7cok4h1erVGNHlMCvGgvShmqjw96SROFOawhDq0qftOpCl/bfN7BvpujfQR8HRw2+1xlh0
MZ3L2uc/c7miWq8orGls0Zbd6pSp9OZ5qV7rX9LkDvVTOikxTP2ykvtcPelrJKT2eXx0d8zBBzUZ
zgQfCkMEViUxZU5I5ZkadpwjHMveTGZQCV2aH7DbBT/N652JhmuL5r1+VyWFyorJOFGX+V1HjbAp
C+GmlJTae4h8wXScRz6YkbdDwTEEjjMfZ1u+63JovGglDqTI+tGzqi+WXTfN4vG8OPHHjdAvWaqO
Nwy5esidjQI4zC0pD52+4qQp+iGuU6rnHj7JC3HMiWQVUYw4YFGgzX6DbvKv6RKho4clNEgKkmVR
w3ERU0/5ydjHS5uPXEPi1IPMdyTNKNXGGk/1eIzuKmy40UQ5lY4oLjDak/on1k4R/FAGlIWbqHne
ttgobg1ZmM7mXTry3axv83lv7ze+pNZe1g8voarf95hXZEOJe0s9jKWyGDI24mbdz5aoelYHdLR/
LfRXcGcX3olQjNKaOTGjnVXOh2DHOSxo/Gf/E+T0vIcR8wCDLqcH3I7QNtfQt276U/ddETgXH07W
q1Ya0CBjO8P5lrsyUk4qTHOBYbVFEUEiLgkYWoRk3KIcDmJj0X9EV8Pu+H/gS3kcUy5C1NfvvZhm
kXJuY74Psll7Qgi+h8DVX38p7X7yEMFRAOmw3k8gNXSeVNGXU0VGw8Aaj//Y3sOJI3aC91HW7u89
zdo+e9E/VlWpsHxXLmqH9tmzl2/7+XOfMvaK0V+9MUekIICcJy7C1cfc4psDEtRgcIe9F0zC6CE0
pRhgunnI4gr6H/8DPOoMdsQVf1X8FDymof4viykLZ0W9118w+3yctwsfGyU3xZGECn3FFzf7BqmN
jXzkRk5xf/lZfwYal9WPLPJ8SaYq6mvnVvm9LlR5/y8WHlru8uFWzmd9k+ETISZORmknorBCuKS+
jTgWks3wUn8o/zo5XKFdlejkONClForw1rg0m2KMRhzms7bRi/F/ahuqwDfcOmjdQ58hnNq/eiR9
n29PPG2gIsLoo6G1FyvQnmJcXfVpIdWBQZprWhiebOMiviD1dMfamer++R09pLQjwnn74EnP3nHQ
ZCGSyWBWe03pNurr85gNc09AZ0t3a2I0q2siWbIYUV+3+qAPioAzr+8bxabmzYBcxHrRXij+7GYk
L/mmsT5IxlC0A/CSDCBwooIafEFILAOHQzfwBWlG90fwEjQ1rAOVZI9+j2RoiMQR331DEghYN7hQ
upjK/yWoLv3rfAPdwrO3Mp4KAukgzliElarwnIQwIjTh+q1zFtNuIcyiljL1XL4/W7vLsMVXKygR
K9aS8Dcxw3S+08R2j41cZDbvssC5Rfu/qTs06AlqOj9Np+1lapxWDoNJgzn4bZdQlS5aOwrR0OpA
O73QYub7sci50nhUwDSrWTlGt5ekH+FgmQpRK+YNvcKIc/uFfVPK4SfhtuD9vMtS2xMocpkXs0vd
DCjXqtmz1+VP7sOjKi3GXgCyDkeTw982FNL+yVaiSLwtSKngoWYv9TJ5XGO+SORFQLIlusaL75gl
TgFD+AzCvo7ISJYwb0WTRtvPusywtoEXWrTtfROYpWGILZ7PEk7LdyHeyYSHO3K3+u7lwotDcbwo
+BLWOhI7q48alUTFvD8+0MXSb6fCEtYTxj3NLE8FGuiVG9Gbr1EmVgpNqPH2EoNEegb+efxQhzM9
+wJHc/JUe7m1OdRSfRvwEQ+l9hk/RX29aMrJVXzChST+jUibOkwbx6bVmZXI1uFemq1vXlEOXF1d
gA8ZmPL/1aR7gpGfmkUfJuheO0vtQJrcuoB/JTDJ8B2sMMjYvxH4mroGiJBy4LgX7ls9Bsy58Vy6
Ch8YCjAuCuwOkTJa8ECCqVhkNl8mDA8N5qZ+hl/OYeTN0F5x/DWTSpCnY/I8/IIRM4o9Kc0xVg5c
sEf2AZix/fo+uG9LitEmLyHzhRonc5du/rsQOPo4w1SmuDCLuk/qimVbrltT9+Bbma8YczWszNtg
1b3RJ1cn39asndqJO+YclGt00mSdwFdw8kzaL5nlq8eGB1Jw8/T1fHuVdcKa4E6moLqZdFDx86Rv
iq9DKHfFTrhJWfpHbId2v5O3qt8TWPtlpCaJDdS04A+WygWVUUJptzwZHNsVSFxsukO6vA40kqHo
e3wXF+ihBw8UkR/BzJORPqSgn/8fOraRA5Y/wdLyZs6UGolPswSwxFMb2NaEyV9dj5Tk6ubZawLo
mqfidp1mqlaeFxNKRoDwoG8kZO/t6rAUdgtAbDia19leWsjqQ0JQ8FKFIFiOXcG89f97Vv6RenEk
GSTQwCIKE7TQFlQc6a+69CUA5o8xF/X1g+8lLF5dLo4rKtqGipcZqgyS8p2sB/eYtWEju+2Lx1n5
IV7M5Qg0cwOsEqK8RKB9prT1Q+ry7Evnh9mdFeXYukfoiWui+r7NlHEqUbsTdHol/10ikugbJO0V
VZ0+TwGkKibQcHjW9NOfwwy0AXBjxFNK+4w6cqWOR0puUw2OZiCDvIY56SK1L6feFhaKKBilEPrs
gV71SYhQivxZtn+oEIAEp56StpWLHe3UrE5mdeYjyBfkGUl7xgo0dW3GoKOtSrCIQSiEhpaLsIha
j0Yf3pe1xGxIn/4QKiGWZcmTr5hn0HaTj/45KelfsFMdK3zzZ1CUONZSYKH7T6O/hbd27Z2mUEne
SFMtT0iwi4oD19FVhO06PD2UA07phr7CKE0P4reWMa1OJVCLQcKdV2Xoy1gE4KjKyVOwu1j0PFbi
ekh8LeeRBe/7bL4lpaaYEFMz5k4Ghav45iMCAQzWvjzqXu046ElPCDyaaMjEuJ7slD9JUd8FC9fE
5yZvjj12hOQzpvwUz61t0nos1pjRw/iVyOczmZRtH54W5iO7RXuW7YdaWN4DKG+cuj1q3ooNVpWh
RytucUbRNu2aGV+BcuafP12vDSzLHjdFad24ZHKov/u7bN9bY6IX5s1nzMH+BgRdNa7xL6mrYcyq
ffQMHP7rENwPC7NiyTic4Ef4d8zgOrSJAXEfMUK3NND8x7OAYaRyuYp1uQr7MXBuusve4CmZExk5
ZRr8ZUfFCg9UJk1xZQVKJMGiNnmN5PJFTkJJKgAfmMO1TNuMoY84+EiJivv5fpWJDtomFKslYafX
WK6KcifRncbM9cmbIej+MXYIN+gkuRjv75tDHu5CIaYwO7r+d0WE2ajsn9DHlBZl2Fxvh81dSkfv
jmSgaf8T+PBt2wCotCPEPPT8Ll/8RGNcoEKwZZ90r61o6j7q199WAD3rsXyIXz5YaYnFz17QQUc6
Ty6L5lTZFSx0EtfBbzDC4zqkT043WJKn4Qqtj1Hd4d0cv52Vd47CRZ1Wk/F/x4khZDCAOQGRn+eD
GEb5/DxRRvl9n5CfUxhUyJIFYaZ0u0l3NEZtMTU+FRPteric7qlQMLwnGx3JzIQUB+BOA+TGFpGy
xHJz2QZTanTHi7SgLiGc0L5O1dDlJnF3KxtIZYwre5ekbAxTpKUkdxkYC2IWFzwoP2xPWlVElTkS
wa36s7fApEE0VX/kHSZZ3nQ4zXF4T5J70Lai/j8hiReuwrL8a3VGFiKNtxphOZCT4PAxXI1+p1dG
dkjm83Cy4CMp1rMn400mDwhEExHQhYTHYaYiACt2Bbwz0azqq+/j8K8hCVHemiGp66BFXQTR1IAG
8PwDETWYWVFUin0tU+4YFygczzE6OVOPp18spkkWQSayf2MsUbmUWwWMHVSeTgcSIiIq5jeA/PeN
0gZTeSYLXT+DHKnVnKKp0jhjQUzgEOxbnrLv/yKUjeW7NTPXvkVdHYX45UR0NMcAcXHAMf10mnNo
QJyCucH9+GiCjvUhZVUuqfw0RNoes3a7ZD8P5nft41iIyV3vwKPztoESIHIqiYndaW4oOgj1qUHz
zwMRZknzFrUYXWt6aYxwoE9akuKlafiDdHRxlLEfTe8Xjai5XSdbKu8/GQ/YVOFKYZALvqLXKoZX
Lt3490hHYOWCwpcHy3qKC/HKNkVc6AH8YQqnhDUucq5Rt7h91UaHs/7e0RHGlMblrJ60IX103VTQ
tY6mQ8kIzjozXUFOdw0KX+K8Ar03FULsT00htWeJJD1jDzQhkzyBCMcUqtwZX16ArV4LSkJMI0/b
sc+xjBgHYgCW1tAXKkUyrKRlRxc90hdRvrx8WoaPeQhfP9z0pHL1JLx4XG0O+KhxxflY46oZlUko
sbzUQHMY/oZTgwOUBN0fZ7v9yO/+18j0JD3Tv6Hp9+BZ8PETZpGgBf6yTHQ/VHSLbfdJqMnQ2oZu
FmYV3vS1MQRRXzSG+ZKONPFI6dDAC93VKe0SUNh0qUFDBX3sQ/qKNyp7IKWz34XVpABGb4aKaq3E
H+X8bwcO394rTy7XuiI7ageeT4gibG6IsiJuDsKp0Ygi9+Oc7P9jewvFw8XUd1/rQsiQ1kYbdGPL
+TUNgf4Ke/fCuGcX2Y5KEBd2h/BwenvJlAbFCekNMfBDb7u/5D1hBsTlQPdQ7vW3+AalalxwB85h
UG3DVmMhEbdjJD1jkE8Vv6quD8sixrssMIhOyYJCwCd5td9s21ZfaaI5A9rz4UcZHM4eoNY434Vi
mAkYcIoX4ym6tBa2f2Nd2M2o6PrXh6HTkCoYltqI6/DvQWAs0+QzCEFjV1zN3wqWW3mEB7TD5N7j
G0gEa9Q6E/yAVkvsL0fC1ZUarvQZiD0M7XwT3gIcEc3QS5wYz02aQJ11Ef5XVpHcSTwpXZm71h7Y
xtMo+f1W7Qvgt1U8+kJeyJfeKzJleYKhyNl+g9IDigvj9r3Tt/82WcKZaJ0M19AE3Bz6Dk6gsYKE
L1T18Cbg7G6djI42OYiwC5qXuVt9ttYh5EvXebcQrgb8SzKOWlW6nZZJmoCC7JuoNsgDSuK3XvRf
Gp7K1MSKwW9dYKsVGQFvB0S4jpUSt/JB0IwrJacfXcN5zQB48eUX5PQMoWWiMHagzCEGBP7VhSma
sdnf4hM+UryxhQE3yMb3UUVLoPZ1gA4ghkHDXqvjejq1Z+A9zM4MDSP2DJYb9iLkJ52WV497rnbS
x974tlhP8GD+ZXwse6BUU6MS5DI5ZPTMyOQPROZRgJ644hbCFtdXpl+8cXKiVM9yQLTbHE45gGNR
i6QGlnwQj8PVd2WjiyHEBB1AuJ+rya/Z8B5NW04nALANciymRywoCfwL06qga5k/vPjtHiiNqo5y
i++lmf9KWOA8gh/gt8yXRIpttp7R4SlsBjSdS8mQE7wDKedEnkS0rMXbGefFY7B0OdTcr+i34dQ2
/SSTdBg7jA26HoaxHWrSbYr3EGpdJS//m4gsymE7WxqgNWubqauRjT3jhfVNBbXHwf+vyxNEjy2O
Mn6hiY7jdW2qxgHLNBPmiv/4EdT0Tg5dNvmP1AkmmCD7foPEwYhfa+Dq8XE7KPv/2fBrloCSkHtN
fikZq+eNiVvqZ7KX/t7TRnV1yGQmyUqQ1tsRh4Os9wcpz3k0gWcUK18h9lbjax76VjnO4l49fTt/
OF9I088N1VGPRKyflBne35QC77NvOf3nBJsQhafKtC3uc3NfWXKPF4X2ITCl4YJqchRZTx24YJ4Z
WVfNYf+oTQm+JoI4r04xLpgjEPxOwnCc8HLFiEYE6N6iok1hthA0VngjmvsJL/HNDWQkpwx3I4nm
mBfgVJgZYsldm0mccDzB442t6ggEvHVDBmRlZKLWvdkKYGGN744Mbksr8NYPwq8vhTRHuUhHDbhK
Hnuc5rGM6UgwTcRquTq2wRH8m2P7qNNvPoU5lWzw7/kGH0Uc5TLjZBLag72YHSn4+KO63Cr7zWjS
VtAXQTmSVB0CeRCow4DeE6vNWZPm8A2C9mN45p6AVccQYJyCpO2Nl3NtsLMw6eYTx9IPRBlew9Fx
9Ga0dW6uKUfN4nJoP/+ASpB9x0NylJqWDqXEK/lXNNnsdG87r7iQBzImEs5TOgaKE+gHyDHLUI9X
NXddkUe82kWdVptC3qacqvz4O4p3G83pmJSyGLLVaxZibD6zUo7XWaDADTfYO1QFDVH3XDid73D3
S9cZebZHDYtMoWD48Ipm8yrDqHYo90ZhX06261l5H/LiWRMpAZCD6sHL050QQ7GARo5WR9hxJwuF
dcKfys1are6rhwPmpO2AiJh/66k+evmQDVOGUVUjHpIeyPzRenNX+KlivudNqrvgbneejgg73Fz/
wymhsMc0RqPQrVD2pIRCO4MticjsjKhhVYYP80YYQpnHc/Z8+pRgO+DJeX7HFmC11NfW2hAgSpqa
aB7ZSWbP+f8uH4jSAS6euAdL8LRymoCmdFDKVONHt8dsX6TZ/veVgUBXEbkajgJj2tsCIcAPDD6k
aB8uxI6vhmg6Vkkd48EraMnw/NwSLaEg1xrsyeYjraSo53nJarhnJlOOhwEQ523haCm7fOqXM5hk
30ZDivq9k372bF4zax9pwj5ogygLWpzTKLt9KUVvj1jL0M+V72cOXETv6IB63FZYD20r4E2BVgoU
GUPfBgSwtImbu0DxLOosTOsNh34kbRCr7gjCnbvAW+ZZwF9uUmLJgbw2swFhjnW/eEcEUmXpwT+z
GMS/obS31V590BymghYkOrkWepD7ilSXl4Zq/6yxEso1YIi4u//RR0yRoscq/COQd+1SrOEFfd8m
1+fcBkN4RSSTzBd3lmI/onyzjQSz3z9Dc7LB/w9zs7NKVki7SBdvONhMBHu5KBRC9lYPnAl6cLJo
1CNzJbTMzjF+NAwtTSAbrwt+2ocVqvxuxP1ioe2TLa9XclBf2+E1DY2vQW84zWzZZgwDsZMxH1Wg
t7ZF5KfB8EYhOTkZZ2/y/zT18k8zDXv9NbS0im8cd2LzIPRp4lDgns3che975H+w5j8HqkDTZvnt
GbY3xnZofjzUXAeO4+VnZCmd1I/j6yLJgamOLA8YjwhRP8Jv6h7hXur0fl2pE3teFDiQ+CzvbeMY
H3jAV7apKIjEZCNiEJd9bCaBjV1J7Lilsr8sVJb3K8AjdSazz7DRE8odAgrqtLslPQCgvGu6CgIm
Dr6nBhQd1FmJb5afoUROlPynx0yttWdxLge5cTeRhePjAIAH7pUVQImm6dtMt4E+95DF3tIgWVt+
PUfj8zF/lv99PHowClLUV705tbDFTGiBzk6x11aJ63IYXBmSn7hBQwyFoIfpaQIIfJDy+x9GwRmh
8aTjKKhJXHm3lsxbLyE0d6qxhTjFowiGeohYjkfHMHio5P0zWmUTBqk130rOf6o+JBjoOdvNPmXM
Af3Maf4hhylHiN86ZVZ7FqKKss1l2rgCxp0Fg+9jpg2frq350PbT+jAwVjdRpJCsy8HV8WeB7CE5
FZXg6sezz0ulSNMAx2ctesFxRYODBosNO0K9fXhsBacwvqwr02uI7I0WReU4affZS+Fwm65Z7jB6
sevWxPHjJgDfqYmrv0TMmHAeeIp1bRttNnwhBc6D/4KKC2eMPSosJ6XhgxA14IniiswCYVYgfTrs
BTNZOb8hm0Vr4IESCXMyHJ+YUQzoXx8RwQOSHQ5PaR6j9XLqgvdFqXdJKUr7Um8+e88TnqaR/YU0
VFVUg+Fhhz4sB3HjChz2DFIg7gZeyWxCHEfEgrKjBpy2swaYdc5yKtxv5Hykl3pySE3jK2NOr/6A
wvojtoBn69n+8ubErIrh2lO5dOOEl9tNniFbrjfUfKc7cnWNevCaX6eFGGM/+0/WqbHRTPbSi/nw
NA+of+y0wXidlXJj2xTittr97S0D+y1gkF6huViFnltCbj0jbZAoAHaAmG8IUH7PoqZq4vLK4XCy
2AHCBETc9wLaK5a8UumRv2tSu2um1dia59wfens6cQ1LhJ6H8TJvkDpcTtUMKyq5bKbclZqHZ0K8
+664ra9Gj4I1OeSOrc4iV/TJpH8Vqx6Qtw4xx4utuTKPr4YXQVX953voj4aCuI42MtDJMIaKlk6+
AD0NkwPp0z+w8zNSInOMiR4f+0YOCXCA5nMRW6csga/oQmiJGBhXmKBrrUsRh4X3BxjM7IWXXC9X
RXAvjrZpTrCKUBhk4KOSF6n+L4P98Sm5LDdKk/vDCD1mrTB04RWxgiW99IazPPEelF8+ENJQWo/K
CImIDpVURokxEOnTCoIO58lemZNJ40zvMgT7mt+XOpfuMjidPZC10CBVd8nPFEx6b/jq6KgXpY3G
L+AWHHyyauP1p8lG9LfeSUznq/Y107vurmecpTWihLRo9L/KDDK9+uwsUq0y7W0ynnUWMwg93ldk
j1eXMmSLL6XGEngecQ+SWO7GEnzIONgIwBuyVcyqXS1PQB1X93WIHZsp/xFBzNU7MjtdNNgbOlD5
vEIZsG0O4Yj8Vy4ZKw6+5DUoZRUu7TYOvbRsIpFQX3oM/VtcDhrs6mLcMS1wxZQXHOE1NKstccPK
VIf6Vyt7bS4ihBQiKvu1tElouPO6smTZJ+TfNUdhA/ONgY0inuUW80WlVA5oeWL0nVilJmTTwKIV
X9/VgyHFI63BAGIOu6xVDB3wZ5IoZ8QzRh7GWv04PYE94kW99FaO1mIEOB1Imu6s8hzG2fsKkOKl
4JBMfabzyIVwFGE4VNJrue0Wp3zUrMk0eY3qKJT2xRaZ/gYPumZky/7fcaE3oauHAq9AN0wl6AHD
Aea2bgxw0Awz8DBDKivawVO3yU7F8eRc/iH+EPniCwBkK2VIvo+2fAAcE/jr31EgJYhAm92iaNQe
7SdKUCDC0T6FC7Hv2e8QuJSbZTIG9s8sSu63RrNC8X2TOFCQIUQisB3GtIP9lHF9tLTAqZRDfmKG
gxcQoJ+zO0oXol6jFxjlpS1Kg516xwkE/A3zYdWB+7o/CenJjQ8e5sM1y0j0CkEO3DHANiuyDJ/j
PnYHpxqmjQfzcUzcL56tMZGrzeaXY/E9d3Q8hYpAhPa9+PIXjSD/6dT+9u2J1jWSdqrSIzwBSBsf
fqE6A+7fDsKUxY4Ocx7lwp1YCzmzlE6XMP48/v5ZJj7ZXHknKu4lYTr6Jlz6srJpvA4q7BUtCFsj
ra76f0/0f/2yZrU2G41Ou8FTZanBGbOBFVo22rDkKTfcH0ls++t81E0e08q09xHA1QMfqUEauO9a
FpmST7HPkEb36+ckqzE+QPWdTQrVVxtscJSkZPYNAEYqriHQZunpzTiDDk7NkJ3OxiT0aPNctcje
aFi9P9WWOCfM0w6oi61njierNsA5nawW+RyZJmKIwd4+2WPjH+iCLLnMQwJZINoS7rM27eJ77Wc7
L0V0r6+tjMd+V4VcGvlKECFDw1q3+WPietfkkDYMYjx9MUjb4xeP6DliMBc979gFEC9SJI9DOBTp
pTC51i2JC05ma2SwW6k6bp4Gu9r5/yXknbjeYPq6rvKjjjGR+pkGTsWIFrV7UgQtvP+eKW70cY9z
itVR/0GqkK5FL+zzDxynGMt1OyVue6S1vs4LWDTuzjC0TElDFGv0Ag+gbWpsfjJFKPoiRF7axJGc
2ayY3NYO8p5ZkKuJ9WmVnL3DJgwqm6kVrDLCGAEvgU5RWxC5oRgGmvNbQfryyxZyZZ+fTBc4oA/Z
uvgpD4+wYOVum0t3Jn/KF4fTjGu8Av4S1mbEf5uDm3SDXKl8fngb/QgYIuq8/fH9cTKs0WixTLLR
H8j+zDY2/igGaMhpiUgr12gE6z7RWKN6vKp1lNUjHLgssfKjRQxmnmT8oytvQQj0xtLpmhehkeqL
mSxoWNn2cjYlTkM4h+QJZU/9mMpTk3FchqGfZhxPDGvl2QsqcgwoGdSq+IIdrWvOKeIwU/au0ZK8
IRy54i6iRu+nkS6KstOcpQKfKVbD27LHfsKqx4p9xATUphrtnOSw8zt6OrYOEMdKyWlz24WTwhOU
HVPVrAA+c61iYVQtQsNTyvAKl58dd6tALWCXmG8yLdE48L5SyRm1a8xJkMJ3eosjdZj0/HtagJL+
MCKfRRWoj1/Ocr/X8HoTOaMi/TOx2DZizzYosfaY76K6FzfMWb5dMzejLdx8sAloWaJM6/F57fue
FYZz5tL2AN4xgm/iVh8ndyvIu8zsS2zb06mjYyFx7bjqFTQ77xXvOgnCXg1S3Y97hnHJtTG/GuXF
yGoNmjl8zuBfzwi1p4yRg8TVh/of1KiPZ3DGyaLEwFnd1DEBXrdBzSfKByMXdvioKAHkUkJDLafQ
p/Pt2fJLZpPIOPS6q5wUNLw5bFF76hgSfs27XX4DvshuZjYh16tbJqJqKb/2Qbn5WlGAwJHzWsL8
6Z4hiWGA3gJdS72Bx+poZLrnsyCA38ZAhv0qtZzlcpZLi179fqj9BdY4UHHtQnI5ahC8FUSC87AS
axwXCkMRi3ro7UXQvKymTOrQ9vQOd1fk+bX+SJU/4dkOlRcybHQ3/eHp3caO9kPFWYOVKwsMGxEZ
rtlESwFlGkGiZaVOD4B/UeOh7MHr7k/GwU22en0llOgKrZoFRyIyOlaoiMt30/Z8uGEcFdRWNeze
zj+0rjnw06rP4slChkFEzMvaPIL9fmx3wuqtNtR2ln9VQMQ9WNUHYu8yD+QRbk2cDDaUgSDPwS5c
uyigL8oOOhtEypTpD92+yNmSYd3wVYdfTmFuQAW0asor8R+BV59DkPufzfrmAVVIabCIBlEkZrDm
c1TSwPIsLptIPrKnviT8ACwHlNUPEhbvT7FtJgWG1cyJv4U9EStispm7aafqkd/ufVZUN7m5cd0f
z+7vfIF78LGuVGL8aMblJrZw8hXH8v6tMHNGoxQXrM3eyHHXAUnH1B62tT5zSGzx9iSIp9AZQYP/
oja48SH9ViIn9X2cizsXu5mGcMg6cLkjYY53y90aZq87sJRpILQZh28XOMJzdxAm4aq4p+5WoQt6
T2z43HmNcjBKTnmpUIDtFJC4XDpEb43sojqG0BiJvrzWFxo9DYGvxFurw2q2ElWKtd9anYVSVmYO
Jn+HsaWYaN/5HRdOQCE+ImxZkK2c5EOegY++BBX1aVj+uILHTgufkoYFFGRRDAO6DJzfFqQeDW3n
++e4wT+lZ/WDmX1FaNZmhA5fvj8uxSSek947oDSQoV0oH/az+jypvNC6BuBTqWBNyoXaUWpawZ5Z
eOCMvCONth1ESD8A0HJsRnCQMEtXDbwL9+WFkhkx51OBJDNt0ElmaMY8TJ7m4dpZqyAxxbHN03q9
PS5y0HRrC5pOJIcV2XNtMsTgiqRoacSpsv4MF+BG0FNuTKGICvJZjXTKGCUcMAnDyW5PBzHcuzJJ
sR9jWxl0vSfPXkKS+u0mlO7JQ2Xs/UjTe8MDqjvZ1fxwdcANI8Nrv80HoOLYYYfBAyBVTIjxI1/6
u4/xzyiFlzwfTmS9ZNRdji6xVaVTf5wojxHEnvKf2/CVxfmhOxs6yGnolt5QbYn8SCoV50RbEP1D
qiVPln9qjh7q8sRQ3SiLiAZrs03xB7u/cgPw3MdCBREGGtMYe8/q9ibJIcRNgVV1yB9sYMHQ2rj3
6ixoECNCj8t6xNpRYpzWxBXhlSog1XuYXLY++G1jNT5oGA97aYqqz/U/hQ4ohMffYpPaVOAYR92v
PvzrEbPbiKqAdWr+NriJh8jc+X2OD4s1WQj2ONEhY4JPV1YUtl1FtRIFMBPqu3XWRm1hi0kotcJV
WTS3rSFSypChK5/lHF0AcY9Ykv0ntGt6oBwVS7YKWFqsKYaSDc9W83yB/ErVaiZ7U7x+ljbhR+ol
v16yRagF/YCGt1/YVXW2m9faVBKU5dt7MXLLBsJjRKJqRjS0dr1AtOMdwUtPz+lbnMl6KrrKF52U
YTO8e8Ak+a65ehARB5NE5c4fZTzn9MsiGZ7d0EIJmTiS4cC+nGhtA84YeVaPmBn3uCuwKxxd+ulX
kh1FjT7jUfV1zFdtUEEpw8hj981yDtVboJBVic/oiRWKqWAGXEcA6k9Va++tA9TLn8xgc5WgRihk
3lRPE790ih1pl7jqVF7n7kEjEW67onXwg6arOdSq6YIVQmlAh4Q/OuzIF+Axxo3tq2+lgBsCzrm/
cL9Gdgzu3pJ3b8YBMU6Ii/7KcV5xPQZz0DDzP84s6aCidsVkmNKE5NFjaeeOICDCvJAfhMbfKnKM
JvoYzOdKGEez+yfWWSM7oS+h8UWCpp6k/SxVohqpVQud4Bj69jE4vqn1Q2CoGW2SV/s426UcDpfn
tie9GrCWAr0XXpTQSOLTVzFnauVjjyW9Vd6yCrIE4dXrJPQoX39PLg6khvZ0JPitsio14GydZ8I6
XKaUyKOnAVkqCvx876PIwFjMXnr+RllbM5YlNDNDTY25VviCifcBOqZAvjBs/MZDgBQfrSoTgblz
NjD/yUi4Qb0hUQRvrCNpwD/8qu+Je5rp7axkYO2/yXMbtyIdsEM5uy2kMLu9nQ3AKVTPud4saL+l
xO67eg32ZiU6gyncFOJ1ZVQ7Seo0KDSZNwR4JUs5JReKXEhiIjvSRUsYoBj98iKXAMUD7qbw4iJK
z1F7qOj6gHth1pzSqVIRCjHx8TG0ok5D6wy5WrGKPeqY5GPT7T1YIVJbGlczoMk42+3WWch8QBl8
b/jrZPl61N/JhXGyC1jmHy4lm5TqJqNV7K2rtylg4fFFGDQPAILQiY0/nVP/vyAitCJNXq+fO6z0
233uQNM9zawJIunZYm/bocJvHUiFe/JsfCb4qHqo2uxZBZ73i4t0ZywddXMCMEBQa6jbGxjqX6ap
j0xTNDO08BjTJ5mEDcmnAYx54ll/+87YhQqSdZMKNrw6JhT52YVB55FtIJWlJTdhLlapGRfk/mDF
pHzbb4RYT4WGVrEkVngcYMU+5LcBqUr748BGq6T7PPDRqkbLGrq6N1rt+awQOuRrRqRhJrGW4V6T
aCuKhw48PJb2uNvcvhTQHiRx5+42o/xpm4mP2H1CLKYapYBpcW1mw4yWny2dQJzznlJlmjj52b7x
ct1b48FdCEVAJZAXQYwAR6GxxKZmIZgo+9w4WY2WxYCrOg1EEwP2j8egezgQsTxqfnfiqIVQTTN0
ApOa+z67KBX6DxvDZluqY++Cmw6nKig7M7gJkuDYNRG+d/mLAggkZBjXn1IN0nw4NfxYLui0hjiV
uhsmf7K2/64wmoUf5RNSm5JTmTdw0sKLN2f3UcZcSXGv5yXJ5K+uv/weUY5eNmGxiM30O+7YOJr4
tuvGTM4CX3SiO0ZR79sDn1m2XJ8rKs763O3uJouP94u2c8HWrLJ7650jpedCVZxtP6jsg7dgzT1J
a5vuRWzdIENEpfQunv9QDMQA3KFCnXvcikO8riLf/5h9Pnx9QuPKVViAlmnGkUvKR+5a6QZiCFvH
A+5myo0incw7yFA8RAL3jBv3Rg/DaFfEC5VHP7VkybJGMTsU4exP5fe6sjjlMMMmx2HrEtcnuYAZ
4xYTm4pbq2f7ErkQ6pPSdDIYFIzjiQhX49gfJwfk1OwpL1ncO6QnWoPFY149V9qCvfJv7RIPB7hz
2Hqjuualb4v+S5CC3nGs9cY1UBU2rkGNb3OwNoGFnYjQ5SSwsvBH9MScYfxqamxdkkP5xi/Hdhg4
jQTwwDj8pXIDUFf/c2A8vGwvCFmLXxhIi9XpdVBWd4N/ZbmYVq9hEx3j7qULHmW177hHlRN/Jkyl
tWBW9Yi0du6K6+XNDFytAO1neRXHpeW91IN1Q73KT05tgXlt2kcKQhJTT5hhUxBIMnSElW9nBCel
preGRJQsc3bHw+DD/RFcbaN2ZqGeCcshH2DfUiIEK8Pfjeat9kZr7pK2k/hHgdf+g/p/NbYhALGC
B9RZY8c0fATgw4NtRpQx/ukR8El1IiRv9vPRo4lWzhXHnVHjO/IBaJIDjHyAHPMGJtKW9J5OLKde
qrlBQPpG3xleoPhpYo8Kq5COqG+kzFVGKlF/SaNiGOp3g7YQCT5Xyp1Bib/ytM+pib2HX9G0sgzQ
ouxMYbbL7eXabDY7Y2qjN+MxXZGbHxevAzk5/gCrSXODXAKn+PeEC+kJz0vY5wNaYrk/h9EyrM6x
14LuvJdaKz8CODLPEV9nAxXHT10FFwx6mjBKT2PSUdiLVj+Fug1ciVmtMJIXLR0etQezWGnvPkw/
INqJSkc0iIkfAUjZqWLYqmViLjVpNl+5eGnQ9VUF9XqLQ4c5PucT7W4GAEpUZ5Eitin4QO7vijDu
VqFTHygoscKn70GuXhpLR5vXKI7gyierODkOAjd+Qpw32cn+cwF3uobErvMthYvkIFLK7CPQGAoJ
t7e2NZduU+vWj55TqcwPBtKohjpXqyxbng9ZDeacsh7l4Lxvhy92DC0A4lpxZOZrzZiJfX5e3EXZ
DbH3yFXxNLOW8sdE1HglYCTZdD5CyCJXBVRt2S4EHMkn646rVhTvCIILcq62QFU6IM6GAJzQAv/1
o826/xSQNM+bSzvmheULEZekNJ61h+EzTBywVndNFfgqfcBPoxZLCbVB1/8xw6lwPTi2LXrx0Z5D
WBTeb7EgGizQwAQdO0TDFvu6kaGGHqhxEcpTl42/BtcEG4O4ktCLz1J/3PmN9Xfeb7y5qMFfsE0/
syKsq+pdwuSsHg4M5x4Xlb/BTh6MA51m26ar3WGDsXJPWAniNwiKtAOjJJ3xujGZmeeGUtlpqLMw
UNJVDYRmLFsg9Ryj8q7uYnei7qdOO2RwdfZvRoA89oH/J5HHHdHQLeNK6Er4za38x6+Ya09jb6U9
WW6x6ENR5LdsU1aBD7odhNppMzlzAXC9qrf8+cQYXisi1uJxHmFPpGTdE0aocdIj0Gzg+xvMFHki
AxBd1hxLBy7lX4YMXCYnIYuFySemy7Vv/3I2W0YtNtOMNreFsoQHoN80SADbFq/PQZFqTiT9e4oA
N1uD4Dpjr9E201ZSfKkiUf5jd9Sfol2Y50lFyZOewkohavuvhX7b1Y5viPdBi9ZXeU1c3yW4slxq
WN01WUqLVmxbPLJAafiOlefHwAi81lQMpO+BYq4RrddCox7qj5+mlHqFkU4L6V6uEv2Ogk/S/uxr
/Q0HkcLC0ke/kqI2pZUwtnt2cItHpmLVRYwieCg9SaIjXCMsYtMtZinwutfXbfhJnebRMYI6ShkF
zV5F1WZUNcWGKQA/w1MkzzmKpSUpyuWlZfaaqJlIhEqN5iH/tZlWN8Q0TfwJlsSqdKCloxEHlMid
S+9nlzCxoyaewy8jvJTEvrg2+xu15XNDnYXfxF4J7eauVfjAHT8y8nosGzvntz1/BALZVc1H6weB
wwFFKa5phpF/Z/n3EjlCCSiQpoStyzpjvrwRxIRZQ3uOPSnDiq1+hH6LXvuEEwjnOit2WchIDIh1
RV33/MnfUdrzvVEbs/slPTwAg7orPrEkvFd8RRDGf0IJXOsizWY9dJSpG6uamGTU+u5H0xocNMBh
Cpsm5CUW4UjRfNysPCkpNBURMX8fVpP94Hoz27jgsggMN3zC2ABAkTGB4dx1JvgbjvO/wmau8jBF
ntg/2pTog42X+InD2P5bOpXsZeOTVroskWCQ2DUNlSLEIjITae/nozLAa52qX/MEclU5Ga1O501P
CijjfN3WpBipY8lkbyKZbTY2Zd+MabvYMcZDksznQQeil+Y75vSJpbYyMKHCIjKp9eRVnHD32X1Z
vvWrF8+vLPaEa1lofa/aJLKUwgn3sC3DXZ8CRX59A+XokJ3Xl8RoZauTTJIzedGlu9Na3hpeTJEk
SX+y0yRE6IA0i79D/pa3yeYvrjBXdOuuOx45LpZh2uYJg/FASHbP2QUzr3S87Ncarn6yWqopatz2
Lz6mmsG8j0zN/Aj9XG9MzuWf/Y9p2ukK1xanucJRNpWLQqE3SeXBBzmQDr+pLTlbPP7EiNgS824B
mcGck5I2LcUQ7Nh2ZdfQOdUVya/5po/WgYFu+xPEg3WLERbqn6XoBzG+9Iyogl5VvkKGDLjbRMGw
6p3/YaW3K6Zm6nle4IR9N4IUpGL9PvbHKFgShy+gt55zZ7WDHjRIJZewmXOe/ntLsoJ+9O1AtBYG
cpyRJvq8zL4aGyhGkqGLLUvQyEPpt0SU/iz+jqXguXofQ+UTaXqpIkzFPaA2nSlRlFnb/uiubh1p
uYAJo0DrPUYzpVae1YH+droaftqLzKi1fhcEf8oREO4uYqzGxa7n/dolSvq6U49LV9nLRvXRefsI
jA9B54s9/IN+Namd983fbuODNqTip6CUb90oIxeqk9yeW7WZqNQL8bexJ3M0g+UUMHlsbh5+GzDL
d/NnPS3ACMXmRd9v940dnMM6dIsuWJfu0j+16yaQIp+dU8ceBAYVHRLmtPLJA6masgHN4EiKOaGb
M7T96fYoXuV7j1xL0aXFSe/IzEs01XrJCErx34bxlsMuUDCLflP7dl2KOncOltxmdZmTurGl+ZDx
LwVDmv5H1ScS3Rnc9Sd+edVsYne0FReaRuS62p4TMRACalsyG7+lcvcaZGTo0MV21iqlxtKpqCBU
oRIF1FX7NjSTPFDYe2TFjpTaU2k9v0D17oCY7DywgGsV3booiPqljJjllHtETKwZ/+KNOYc1JHgA
x6tjoT7lOiK78+z3PTOJAz7dyNytOYH8Fw3CAjjKjvhnI66+3gL7FY0y11/R83tNaWYyqmWrCtLu
1nwXZRzrXnegNPeWqEfY0U0RyX+dXQ4dYeGtOLjdnuSrlshi1M7F45FZwZ24n3F0+3U1RXst4j6m
bfClM7kymW2iE9DEAPjAOOsAPNriUXbx4Dub3oiARx9BJv4vIuCO1DKWYVdQlkxmc0wTNBGdJft7
05YnsYQ28zXQ/7gapR1sVIHyFnxAS9o4ZARJZr/ctuoswF2tcI3kVXGfLBEjwDh+++JmUrOU1LNg
vQPbe88Zx/iAS623U6CkLdRGA54LEt2D6O+DBNdYRCzFS0Y9kdhVlKMk03PRwNPWNl5kGGKxBpYO
/kOvFzhfVKu1fPLpwYUGL+AodY203ZyE61WmF7INiQWHxE/yfNqviYWOTQGU0coN4SfVgysOs3Xx
R7moU6i1sDrjaUP6GiOE/3nX1ZTvXeDL66vPwmI2/Lkgj8m2weSSqjtSN5mn/hazizJaAkvvfTGc
k94lZ1C0uqdFP95HW7HDg0mcx4IUaOweGXgYgxaFPrsPGnxfBunaKQZdmhLguN8jURj32SjSLWFN
tgNnkPrW79UOD1gbKFH5v/eMhY6Vr60HS93F3HViFsU/RVV+3EO3tg+yrOjcBcyMwn9QQ6BdoPfI
676ozJAU6cFAfS8JP5k3b0aPBqU+sVx4vd7z9whi3kvSXCa8BKNEj+81QsuqFU7DRmvrQsphR8kH
U0cXWHklWBsVIKOYP3Xmj1tRAfUE7DeRTsRuEBGQVWeRAMoSsCED3ZBNmRwa81++HYGzPd3tTp3o
j+XNvKyfuxeODiCsTVDAr4bwPWwM34dTZLpvPgUsmNFVjyYSHg5KUyiA0UPwQ9urso3L0qUP9M9F
bK7Gi4V6Xxqm61GLia2Y/5FgQye7kvcBhXZthDI7De/YMojld9GCEVDT/HkXKtfk+IdZekXK40/i
AW0wDc9Hvw9SAzgEpzgEs6IEJhnTZXxGHKtWmVdF+K/Ivqvy9MA3SpmCdPwgzch2fwR+kwCyYLAe
Or9GpcS5qQfYJ+X7Q+56k0PFa0W6KMP0JvIl2xiV7sD+Cf14JHIH8c5DEpV5i5ZwMH2kV6FG83x4
raU561lx8CSv6nbc7iGu01qFThndVY9IgozjjlvU5KGXUtsaROapO5bwnpg7vv6I2omDiCN3AbKm
1/TehmiH69WCkdpz9f0yrM4ET+f7v/ytoXMcVKBhOyULt34Hg7QbIiEtI58/jh0pecw94Bm1wCOJ
NV7nDyPvBLWZ6ttlKtaemY1l+zSrh0iuWWs6C1eZx4q/7W2qkioswBlx/Oi5Scn3oHJy7FV89fdD
YFvFjK0oIhlGtDEcvsJtZzleLui2vEKnc676NpXLqbZ5l063hEgG+x7/1pVbAOiQtr9RzWzMdTCw
WAczs6QGt4Jb4G/l97s01LTu9kV7Ruo+bWifc+VBiQ3f/ZV6CulFBxyLDlTGA8S0owL2PLKVK57p
WjDHNXqWfB15NM5z61TnZVvd85SYIzKp8chD2FcejzRL37wgCdAnKYkoYlUEzqU218UbUTVYotGu
TDmliThJLImLjNmpmDZGH8+ER62S4yj4pznLpy+fzdRmdyD9UW77+jMxUv/igJlHcj4bvMj+Shv8
hymee1DCzHPjFGidjnmCZNhucfAtqJxbk2XfX6cdhhH7bwPGLL7ownCyEZhLHDvjGVofz521om8I
7BcKAdIZssztvTaKcuNk5q6rNZGF/0ahM6uf5ISEIpWrDQsol9KXM7SMgLKVtwnt+Xh3/fTr/Gl1
X1oQCPxXQCxvPSg+aOoNIzLUWj4BhbXNQuP5GsNoHwZ/re28X60bXYPHeU8YyUTr22ilNjHwvxcb
xWtxPL9fdD5sbDoy04pdi/inC8Y3kw9v014ctxdf+agc6ZYjRgVSgkVqLrSaIHudeB9XsTSaF29l
kO3B9SrYD0DpfLpIuUtmEFp1tUc7HVkyP2yIxpvZpfEXDO+vJYM/3dVIChzTQFgJ6x4D7Kh9MZS9
C8BX65+ZAixh+jR2+wHkdHP9z1hpug0v4OluDZk1lzwhqwJbFcL8n2QEzyLwm4hjciI0xOnmCdgr
8/C0/27/AJnD5JjhviC0n4WCADmXXvYm0xVwpu/2V5ELrN8dp2nRYrbRXpr4+KKMmCxaObBjg277
8m1YeYKNiJWJjLQc0ie6ePUCCS/SnPGd592SSVwTGCjXNvwdbiIObhSyjz2o3v83eCyj5k8JHl8B
VFcdygrx4MJ0XRy6yh7hcSQtxP6ni9wVjMgiif5/u/Y6PTnHiCGbIjHqdz4G7OpPe3nbvTBHgk/E
eFRtZ3JjcdHj71hhWMWAdK0haC2b5+yJNRaphRNrFvUfQcsp80pHsqZ9t4rR30iUTuJA5ur+XWyE
QhLGl4M4e5wgnWCgfMgQjRwfEkt3t/NZoJbP1qirG3QGAQ8aXgw9+Zl8oZb1poxLeCy0tHjnkO1X
3I8OP9PAjARwHEcFRbe6IAU7NSW5RWkuaQH1eC9KkcRgG9pHhZHvIu+DNNqF0MNYksrPGJsfQWhW
oFmtcVpDW2cxzEvvXRtybcNW3LjUFzb/lr0ci8SvhnTXFLv05xAnknsOKFDsQvG2PiayDndj9cvw
20N/M7ZRXKCKrEjWebWLn7Kos2Ax4Uv92o75Ke24zy2fSpWCR9SdvvcAUiJHNgrEICzzCV46u0aP
XWuf7pVgPlHlkx4/rX3wta9rgKsl4gS61FrAKRndkFCwNxfvTRS7DsbORqn6oHMkGukb/yESYqPM
K6RwOd7xCIPvZCyBT1M2LRaO3G6dbWJR+XID3yMpUhtG8i+oNXgnTbLHiCXGjOt/hu/cqNpfvT3i
JM+FTSNXC4hSq4/DCyJEVY8JOnakODCX9FjU2a7JmghauMOj6X7yYQd8n7DinfW2urFiYPSs6RB8
xxGIw5pu+NJSoLrKmGdAb6TaUvVuIlZlP2Ueoi/j1P8UvqCYvK34mopUVDwpiqknOmJQyGlfZDQ0
7IvTc0GaZhf/KUpOTT7TCOEeeJQ6TRreM8MpWUBCfkWqoaSBoT58wPEjGxr3AzkqOR4kSnyMumZw
As54KalTTHz/trDAtZCbmnZLnBWMuDUCURjgw6ilfFUnsxkQr4J61h/XO4Wnk8b8dAWWLZV6N69C
t1oimUWr8s6dyJABfazFUZ/xUxDiDncRvoInMa38feplN/Jse4BXICzpMiqk4HJr1dbpfQGX2RyR
HZekG4Paw3YDPwAjeJ+dj6y1xCAXT8eM2CUQfORasyywcB75PUhkbPNQZlC5xmFLP4npDgOvdzbw
BNJL+FeWjHknOfElehtoDWNWxPfa42rHVQL8G9K8ORRG+s4C6AFJPIvgBm+oqsGDvQR/1cE6JWzJ
5AK8xbbdqbZqu8c5CLMIaJ1F7OLuUd9DB60oSAm6WQkMFLOqASI0kUSd0sLhDQ7kAE85cxCJV2nU
46FUNZbHD32FueSj8cjkt0RIubqSMthUXGF1CQ28OgqF3k12SrjtQHO9RLze51QYL7oqG7Zu121J
OmLjK1wWgl5rfch3jsKo/FqAL6fRvgyASibjD6lUTW8A0STkZ/szcDDejUptyB9gLO/UP+6pIE0F
pCD0w+sj7mSf8stklesnk8rasnssOAkRlPRPGxMnh6qhNOqFDW7nEttvVHVLZIvUHpnZ9KDRg431
qudLb7hYJNycLGDvjm8nayjvEcCa2N9BaewPHuYcsLtODfmTOWhu7FdnSibaey846NFE0O/w9xCQ
D5OWKv5SxqumN5etxzY2j2nH48KUuYoqWNHZopR3Dvj/rsgegCTN04JUz5i7h70FatpCL35VsU02
I/wu+X4H++ciLVMUBwa/BiExqFHMbpvdsTpwKfdxenGmMT6W/t+l7NQRUl7hJsYTRJsBp8b18OGp
/zcRna1J/YGNyYRnbMaARo90O9l6zG9o+yUfuSUBlV/zW1yj2s60Gf6Qv6gU/eS84AU/JK+2Pttv
Jk5kJ12YEc5Ag0FpXMRhwg+s6WsRYD4eqnEGak3m5EcXOKgNrXaUhQvliN+6PlBP5gLfeBzVgUdk
fcJolUQdEGbjq5lz+8ATwr1PeaG00NTZgo05YcN8p8ryoVrOcKAGo35/veisqZJ1rx9Bf+LapVEg
bsb8e14ByqPCe8LahNfRdZJW34i6liACY0U8bj0lrYO32QHpYUxvAnCgD+7YXYaK2EE4cKKkaYGI
ghJEMA8nCJ0en39RMKa+XzAEOQf5dJBVGTpWe7bC20TpBsTwHph+kWB0TP/IyxLHet6JAjvI0MTX
3cdq68R+x/8lNux65EKJw+RRlg8J40XSwwLfc0qIHr/QZAG6L040yKPQ55KXexDGVfqgtE8kp++y
G93UAvM9KbfCvnA3YbLrwnxQV2rEQtLinhlInVswLE/217DtLhdUUxsS30fHp84L3AeZIaQ066Am
ahvjNMjEn6uvHTKSGAqsCRg3vEpH9e34A/bYI/VQqu/EgTC/553g/oEhJDep8jYt9rrcsVYCGj2+
sVLCL5+sGC3ULxHM4O7BcpIwaPcJCLNu1LpTTpAK3Wh+vdDmMZX1eO0DNFHq4ldx6btFovg8BUWe
1c4kO8VoFbUpf13L9qktZS1ewLu9IVp7IItSKfG+nJ0GavGQ+ji6sZMJyjrzhq5Tq0V6Ia5l4zEh
uGrBDhkbGtP9FfR0CcXTaGSfokUcloZdhPYG1Wb6ePn2PZRDftgUWmWPCsa7/b34yNEMMjzRP74R
k1Zr2G0vyKO73faHrCTawbMvyy1n/CAgyerkl2d1U5TOvcD6nSOhgdBiWtmBmlbYq4wEQA/EHlM0
iFCbUCMuX/a+2tOBAD3469nl5bsXtvYUk2skq4kheB8HsxVuDZwD12PIDOx4G6PofClXgN4YAkRY
cD+RbgMvVP5lt8A3pCcPMriMNn5zgWC6gBqsRJ4BrJ3x+sGfFclJOR083xb0oWqGLS+/3anoPI0s
2JbI3QTWyReFzRtkfVrTx39emk3UwvXbVvrz4WQYtTxMM1E3dw5dHwMeTV0OPxnDMbeyfr8auvrv
qiafikMmXdyVeuhKpAaiu2buVu4jpSOprgfajNl4Kd8SSKONOz4jFXEN9TiVupfCWyitL7XEksr7
Nbga5fUdDLTrYucyxCvvMnyA8V2vamiE4uoRBpE21PViDMDB0QDNZjThzdh3dfD+XznvokD3i9aE
9cajUzQNhruVK/JawKxdfVveKyt208qUMTlr6F6C3WN0sQ4SCo+XngDsNSBlIHYDFFYrKr4FitzC
Zz/+kueVgVTDs3M2AiPC9ChLO/8LStusaKMQW+99Cj7NO9tKgBDXSGA019MIajN45aTC0V625uQR
hc6XnzcBvHKWdaLLXbjE5I7ODjQQxDF7yDNHgvwCx32zOHPL5MqthUYdO9IMrhA3NzbVEMiw/Lnh
Q5CXaSFkugDFZA0zSt8uM0qwT9Z6qKOwIlqaRbc86Ibpqlqnsb324n3S2hx+t7LnCbH0D/zYfKsX
s+rvwNPIL/LQipz28C/M9WN6BqUl8q7K6zD+ZPhEPtuen65CWnELSIFGAUryP16EF5DIFoFDJpMk
oi1kMzpRqkfVFEiT+0K/MRJdLs+LsoMErHASkcLnVYUgRccuSZ42a7lNDGGgvXb4sWXYSXXXW0io
dALqucRIimIYz9bCHUGgLNv0nUElzRfIW8mvfIva83bFnPdGvVtewpePOwf0lRczo0cm2GoBrI1H
0I2szV2b3vs7//fTukdXPTLk2DTkD9zMr7gyn48W+AVo9fIg5Be8MoblrKhv8RiLhm8W7woP8Puu
BsvzhbSyDihjJnLIERfbjyILLWRirlldU9hk3Jg1sfNoeVsvSo2wVs9iaKV3jTJz9yyvnyCZe841
srv4+GsQ4suqaYcTVpPe9urFjLSyqcnC9hgyZg8mK035y0z8FrVOMoZK+HurpL/l0H3zBLNpHg5Q
pA3Kl9XDYFs636tpAzJPhid7TIWjVMju4q5IILojJ+J4s6EPhOzVsqLlX8xFeTO5GrEQOwLJkdwU
XI6i2MJNAlp1NbQkg6fBXSMapJQ47ubYLLe5vJhNhl3OroyH/N9XBZLsH/MMcchCUF+vpbe2fCZx
XmbE8diio95cGCTHZCcEeCCAoH67+TJCc1jxtNm+PKp75mUgV8GLR9w/JsisSOZ2Ni6D2KaYfcZk
OD50b5LTup5NowSNFwrCAW0IyMwbo7mzedMktsTzNJdNFOQcgO4V6Y6Il6pRHI/YSWxP8fmu+U/I
k7qHw9Kj8kHQN2aDI18fdAfqHvh8ZuWHii4BTy+Yp0a35C/tCnQWtFlgur2ajwiCsVAL6+9uP8G/
6DGawl7vYUHX7fhjFw2Z6ApU2b4MGdpxcRV+AgGJf2AN5LSsLLeAzWwSZN7V+76HSzm9ZoXMToav
dcWVD3z5LUdr/LejuxSoNKKdQerNSwrdzAbpKENXatYXtHtnryh0SsmJyWxTVm3vyvzyYvwY66Uu
AKrDnJa5HQf/0WxoT5A4Ac4BeKaivJ5CGP8rXyY4RQVemc5N3gmGS1iFl6MNp/HjFWMr50NkOC9L
Gama5Gq7S3EVOi+qNfSwE4ifTHuH7rl4/4hrcL45TgIxOv5iPznjgezj30zMeIgWtGT5qwFGPJT6
8N8+lG4IoUkHWa7axog3W5CLIfMUx8B60udxby1VkGdrVwiEVQe6hHxSm9W7MfD1FXcd11DO1K+9
4B0S9gZlA1l+NF9ARuXukfKh9FvLbLsQXtTEmvm3gJLqZy2YVCe5hR0SVb3fM+GXe3mrE1IRgyP8
9X4mPDdd3g+e+5Oq0lv5ky+hJfTjlZfT5nBqGUOWeGV1VGFG72ymPqLf0Ohq0lGi6gyNYyb81n3V
LWa0xSCmRayeyE9beu1M/WnSTLnylgZ3d6EgdiGKZ75HGpYe0Xe8jcbeoUETcAF0uGyzSfZRGBcp
pPsT2tVAGjnOW8EgEIWqFxzUqDDTMrqbtxGSCW22chSzNasB9m6zi+dfnMvymnrlScxiOEg09qM1
CYmoQeJ09Lr4a0lLPzLkuw+9s/nhqKJpA3HWcj3OJCFwtagmznFN2Jbg21F2+Y/YBgbV4sbjYQSq
59OAbXnbqK+0VVPZNtr0EfoY/G+2M4rLDzcNKvQjvdEu9VF8XF9oLz5q+bo+F++JBTk9d/JM/H3i
2lKLycOz2PrdBP1IoiOFBF7e3UcnNGFOI6AJHWA/9Lc4UgG5+CPSf5c7OaYRJbxm+J2W6jM+9uPE
vopS8xAK6KrXFTgiPlpeUaNgoNhPsaTVJvlczrAl+f84nWRIa9s3TDOACba8fHseh4RFoTAhSF8y
ImOXyrLPbX3efNu4EMddOxAosybq8GmKcdLh3IxevNuzSfIw98K4rsebnjxgIa6oakDPT4PHOB8K
6iWGeF9aA1xhkS84g82sEWj2Th4i4IPEph8NKw1aBWJbugZexzD0CE9NHxJYUC9gWp3sskcL1daw
V4G4y031gX1zGjn5yw+1Dg/QIvxuJWY2yV8epfJRAFPQKxu7oFf5aWCssCX5AYpri+WfTc/2dFMV
dzwaCMQ1hFXot6SH6d617Um26IQb/8RfXpZpEeVK1J1efXYQhZBQw7xqs863/2ahXJ4rn/EFO5L4
YRU4LNkmCv0Je5q+rXe+4wWSFYtqcPaikfu2LWc8/siy68tD22gUHEUGQJ0VK8p1qczQVGP0ymQY
uHUaHxqonlLbbt6IIcf85sZJbTUlpjxzOLSjJet7iRsrUry8Xwdq/8U6kOQWkm+q+O97h6Br8n/2
81KE8gD42yXtpQ5JTFPB6sa7uwwHUxniZ6RxfS4WohIDI3ebC84YZQwceWZ3JMNO3Rf5a0ZHAlx0
Eo65ET7/yqAW0AEdqEFqWhTEsPoytQHoWPxsIOsV+0+7VOOndniz/iXv+JiM+vJDitbbCMgNH5LR
wvdQwtPLs1WIoCkSBkjz7lKGu3ybMHNeUBwXEceOGk1qQjuguX15NNLijScIO/swEyaFYzl+ITRl
BhwRZktGDMtChVODytu3PnEGH2Pn2Aqmr17t4XflyLkBtS3fBiNNZ4c9Fa6qJON+pYDsYXM44I6Y
JQo9yqYzAlNpx5OkSlZGwjUYqWTOzlqvBbmxpp8QtaQ9bVZ2pN+oqySn+O4u00hPjjSTshDfO3ep
m0dmGu6UXbp9yxdahkiZUKWOSsazibRr9k0AfYKoIjskzP4pC4FvjWBsoDIF4ToihfuWJcgNUxl9
J+pJuY4j/7tiMwG/mcUUHBn3ejtteBkGWacz97vsmKYfMrBI87P6HqMRyDVsvVmKYbK1yUCerS63
+0cCfY7097IOb2oiYnsCsV0TP3xfc9tH9u5ViqowJd/yMvktrA2md/J3SPLaWOzLYs6zpMHuLmy4
oo7MewzwFSZHEY8QZ0WgVZYDcuY0cQ2GDWnEl4viGpgabIZ7kKejf3X5/Bnn9DBvzYyTJ8Pt4sDu
UU1i8f++bk1pgr/8l8r5bRn5ZAim7oHzhuJiJlv3I3dSStYwX7ktAx8fjYgIYmYxOQkaLvvyUtDy
iGlaL6EaN36IJKhStYyG/K0vSyEb68E172Emi3v+/odM1/v0knBblAu3nQ+yTROtZzy9e0I3VFXU
ARpulpQNin41l5nD+Uz1c5uteqfd6CdVOekfE1nJSEbfYizzTqyi+OXeQgMK31/wKPTMVeuqqMJx
u4eOnslh+ziihsT6RlLxMWkIS0m4P4WNKyU9WA3eE2Bn9aHnOx+KS487I8R/8HRx77H5wX/wxCpy
SKmY+sGdlZijnUUErOfnNKN3NyAzvaPNLjTPwFMi/eUXOicHMDMNZkxT0N2FidD3RZuODXIlZssQ
SAnntx3hNIIqmzN8VsRUyMW6rM4RTXQBwKCQQqgFnmeV5cbfE9P3/qjXzsKEaaUybLHO92ZFsB6W
7KXCMMDZT2rabF3hbFAA7Y6wr8Dl6dXYYYUdOlMF7BthnGbWF5mjj/b1NUn9TVb3oFPGIkoSUVmx
5y6qaeGYOm9YfXhVXO1BgLzjA18XDOzSTypR/VAAfQEd2o7Oz6ZHOSF5Sdpm/dvLjoRg36kQ3cCI
W43YD2BqO8Mz0pzl7XZedUVEo4+4H02wjR5nd6RvXOGz3f4dfYqj2K+6sJoPZ8mky87Wm7y05Ad0
WvOCKuZNh4GTaUQsa1/XT7XiGFANY6gnuRL2nFCmKpwivS1vLl3KFSsG4Stf9qaKa+YNyyYmZYZh
wqYkda+Q/5u3Sdfmmtvrtt3aR9/Gi4ClOszquXzynGVD3BfNf4sqvMnVNojlXxGmymDWnqvUIlJy
CMcyaSwy7VeEOGcip0yA+gdzMfKOGA++sOUoEvHthW4C7zNTjd3O6Hs8/9A3zVT8t8orFSQPCdha
8ELbfQT0EwHB/GL0vVdAvV4/V+mqg6dNhlPt3AtNOu2D9+LknNBxU2R6djggJWvX5yXOl/1Yo8cO
CPV8zjsXhz07A1/AynrgW5kWWzHwCWUrI51qsiAJHwbi6FhcpDW3H2Hy2dZe4ei2MrROq2kH6jFd
0wxvN+aghi+Inn1g1psXu4ZW+cckiGjYlJydM7/no66IS7zQ9BrpgXh0+ke+jcR3Yb/pP5meUWGA
/L/zpSlao1XZgMRlphe4iYSbFn65EQ15jiIIYmKe+7AKn/37YbDq+Z6jnMC6NC268SEi5em3WRI8
Bz1GS8ILeWmvHkHMMt3XzdOJHFnvDra+4UgSQSZFcL3o13dX05tbdcAgVIowfY0s4kdYWj1VID9y
AhPXQY1cmsi18jyzBGNw7ks2bsamP3c7qw3qJ35MZu7gT2E0UJvIJrg0NSMFa0ZgYFoT/+f/juUq
AY7HODU1L37kfDsAEUOntvG31nD23TFcVq+j+KIloXrOvw7FP7XSsvwZDgI4JXAHO96HHgO2YbDC
Z3DPkxqpZMoUZgkDao8DaixSEYMo8IfRqxu6nJmXUr6XkL+8loXfYdIXGnvDyNHONOMNwBvNZbO+
ydoJKguuj644mMh1N2C85g2yguWsFGGH8eHCzN55SzhuDWFgdpOEEVV10ZhaqoeTxN2hotiUAp2z
Nfy8THs84hubB/GFXanCTBupAT6jiIDjouRhN3RUuSTjhRt/cdmeFYpBN4eujZGmSlDNSf/2/LGs
djY5rjW7l7/ZRIjoc70xyoUvuN6aCGdtv5c2qgwp4nJAtCvsM6YjOgk/Hm9U0LJUXDT5LZKoKHBB
oB6qo0otFa4GJorSbj2SjO3zYHRbkAFZMHy2iBo0VReJsMnYBtDEmH36dSbCKKw+UTPKukipFW2K
h4lhqqf10diTTbuoLpAArVwiBCOQyA/4lkZRS5Fr/CGFSDaDh2Q2XKZYAiJ1WQMSAsifr9+pdyR3
oBtmipg9sDGhebpZYOlf8tlFNI0fEqQmxglYWHmXPvi3fNi2Yji+ZEFk+QPBWMpmVX34i+sc8TY7
4N2PWnsNvQsBVNEHNwAQANcIHTfmOJ82gQmseh3BlSzHqo2FKM8jQmQdbrrlgrcUOpcaMokeN2BF
cabHEyHrYzFIWwGQRYzVFPP52p4xqktkxF6UWeubEeVqiMqg75xUZ0XywO403odApbdvrjvzBsjN
pnbrGT2FW87WVnB0xtpHHf6wFrEqej95xuzVj3+az1Dk8DGHTycP9URVFtbyIeV3RLFdlt25szXr
llv+CqKCj57R6LXMxyEDH5uKcNw88xiu2sYPCmnak2LGv6sNF1ctvHu6Qe6dCtiJLppo+DbzMqG1
FW6csSiAroOfpBfeEFihHHElpYmjXmz3TeotEZXiEoDZyzSo0buXDDsTzkS259LizIra6H4mdzSD
GCQH9QCbbuKyc9WXapveNFR7nrU48CNfyTA+G0z9yHyU2eUHZGwmUU4ErttxJ7dKLSdyxb1q7uJP
KrD8z3z0KvhkzMhRqLIaCJmUB/E9gdoEAMkINy2RzKEfsVa5kjbwxMqYSBrHX+T2w0n2mfp2CvxW
pnQkt2l24ePgIrzUBJY2h5Ob2eWXAqC8U3vJEoTOQLCWDhlvna+aWhKTqeHXkULTFWgHKTlON1Yk
4kOl0txBTTjjN630HHjihNbdXVgMNBpetwG8hmJHaYp/TGphq2i6vw2HosSQ29aCuGiS3POWnZYo
c3gJm8IMQwYMAt8uqSlOUKT0U/cAcCBQTm+bkO0mMDVMXiEwCCHlkibiEirO1yhkA8G7LRz5/OA/
83Cghx9l94OWUzTgp55K0q+vxCAjEXI5cLcKgbwCifdu3U1kKi2sUK0g8FAO01jIDE/GuopNltKC
SMFfdPozwUxNt/53nU+85fcXGFObsIQSgbDhNcxG8sJo1ERsb1f7BIljwsXlaAPs/ppBQouzkPZh
kjlofjXhaLsPyft7UcoSvCNne68dZsWmr0SBBuDzCsutnlmVhRgaWSUi0TTfcR1qZ0V+CprukJf+
1tTT5YlC0ldR79+ON0y7KzMYYAEjGfbiSJ7fyPlYuYFXhz5NHhAYHxrX74z+dYtQtlIfaE5Cy9Zg
tp7Bcz6ksnkBC9/X5IXeWjBWXm9zqiI9rGUsccWvhZZTTXAOHTnBbSKfGmuDbdSLxGorprNj3PDI
zef379p+qrQTl2Uy/R0wVUk/xFAzmwE6zM52s+Sal5bBFC/tIOCK3iisMC987/Z0zfg5MAVmWm2r
sJIehARMGmgWdZSKalXi+IcowV5s10E5GedceUlcK6IpYNRzF0uiJwZOlYeaLEYcziIDNLbVrRLy
qH2i9J3EwUSAWVWcNzU4xkTtYYHFEb5Tj0zgBwSjpJg4ByhDlgotYVI9G1Zqat0sJydu+fX0MhCJ
jPdHHJkZTrX/zrVU5bJAUQysTbPiX4dNVDdpex/XE0gTqNP6mGFU6jCuedBTL964E+AxRuQsDbFh
SrKcVERNUhflQBI4uFVkIJII99bq8cmljcovIBBkZmOkBAKj7VM64A/qB84zo5DNWXiPqx6tMOXP
iK71oJDHxFUqDEK2z7FtlebyI1kF8wQ2m1pphjKnGWf6R0gE1uXVPjDWlek84EodkmPz4jRcwHo5
lZ3vvvtu+qH6yOfZfnbcCHmZUymq7CqfE6ke32Tsbg6qBorm2L6e/6R2wkTS0AKWj6fb7TtBmzKG
QCwp3fiFWlusiRJYHMEzcdP+9xvVd0CachV6LMeIqK0MuIH9kzNWMl1VOVDPyY1wPqTGsN4QEZfk
9p/R6Gsw8Vno2s3gd3W4Ubq+n7pr9SdxeRDVzB1GEABLkMilcrFnHiqCe6jZirL123iSKkF2Jx2Y
HjupO/COPussFUJn2j9hS9cx+sDwJJX66rdjQAMvstRW2+Jt6We+22Xi3am1wAWxSM5dTG2kE39F
Fbms4nv670zfvgPZxJNrz9fHbeG/CJGXeOP0zGBq9rWlJuJsOvR58bWVe2mGRpHG/ZnwbmGerOQT
ch24FKu+NZZ7PQUjihMt5xL+Pc/HoY9hm02i/1c46zfWCcnKelwaGm1nh8mNzdsn5C8efFnDSmdF
/YJks4paS3sfiznA9tfcFtOyl/X/Ds7iq3EmJHzxMtL/YMh4iBVjJOJsqLCuPFmKgPKRODDpYT5t
4L6gJVgDlxd2SbWYNMCHzvZJxhesMvr/cbMWL44kyZ8KyWSeUVfl7SQcuIDmdJ4aj4jRTQBHvm1R
61qZ12MUD92661BocUljNMcGRb8WCujjO/Zf6NA0K0BQa7VrPoR9Th+1143NPsLWfpc7Uv7Eiw9t
IQY6yxKZ3akkXg93LUu4hMudRilHAnFav2q4j27TbmqFqlRNhxklya1uXF8kZij2R3oo7apzPsBc
EwpvT/ueoJv+VHFIZMPiMWvaEl0NO4vSVOIYnI470d4LQDwgju2MrimeWvnLArq6ujMfTMJx2RQH
vZSnKp8cRG0PnA1DFPnwrF2ZZ07QuyYTAetTiUuruYp+GBN4S85zAA1Zow3z6jpUtz+P+GCaGMm2
IdoHQeUc0btUG2Ec8W1yx2klqX635yZ8JVDyBBaPO2p1FE1ipivUD03ngb8iBLO4HB0JiyOsNju3
SKQb/Sh6NhO9qsoreibMc5CzGW3UMzU3jlqnJmpyj/P/HPEcfAQP3XO8zNRqnCrDlyVx5fxeNWa1
a/pR+6+Bhhyec03c5bXPTkGJX9W0aKCBcegh0UG+fJ8l7EkrKj8dwM1nbHo9jfoJh1wQFRmuiCP4
QYPLp5uMvaUA8994+x8LC9h2+sD1DElWJxPO1JNMk1G69daIyD5UDjl4nQoOwszwC9hIBPlndjbO
T0XmHXjMmTl+vFoP+RF56dJgqu8221mxOcNfCkzU12/N+Zyl9+KdAcNvSBLCvV5DIbTHffSw4hwo
3SthufPMNh+MYE25iZ8K6qbGJaWjwxRl8qD/yphpSSpwJH7tbvj4gkJcuWLAArousHIeey03J2D4
v74EhPuGMtjM4JBMmmDET/n2QFs+5Kz0aDQ9H6UVwW8cV7KVS3fJIwXt9BKzIEJoEFaUoV90AqZ1
ne+uOLl8/KmsV7UiKAInpGhgIYbNSzouefJSnBu6FdVm8cHHPvlXhmJCGagxuKuxvjbnMl8GDMTd
ACqAp14onlL4gYoFGA5KuLef2MzQsTt/dL8NtrxlOJvglWlNq1q4vvHx1pNWdFmwkS/a6xvsaQVs
Wskx84NKLJwQUzq+MCjZPuyoPbR/bs0tRVs7j8Z0kK4qcuaG2Xxxv10vIhfGdUV69xbmXn+Sji15
LwzMwZczaKBCXyuV7jr7bbTe9Ux+60nepPvv44XcFCsCinOPDmfdQcTKK2DhkQr8UNqztD5bqd0e
oIl4bXJEigODOHk+x2HTrTshBaXDwA3k0S6ztlQwVPXI942qifkcGQY4os1hRxH3mIEp3Nyz7UpF
DQFrD7RBTX+owC8rZlDRePTfLuyicmI+OOFBt2G7R4CFUzV3j8DyxVoSePK3cInONVtrReD5a1mn
tVZGC2INhntbd5jUxvXRLEMKAWia00xAGAlyv2hAeGuRGA+QxA/JgRTyn5U9ZrbKeZH7ry0kLj+Z
AkKV1SuPJ5D0twrYzD/mWhOVY77LWWXjIpQ9CNnLd18+RhS/RFAUyybXWHnQV+1o7d9HlrTCziTG
sGlG1SBIe06evxQEgS7okUTYGYg59xisXadu76luw+ZdFoIIcrNmL4ncC/aviD8n6fuqJx+y7lmQ
dNBKzt32Vb6cfveIFKboZoDbrRw4yh6vkDE1pPc1s9EVBvV+ba9mM/Xbo3RBIQsEg8b/tPRREkqQ
goyre0veegkiRspMZN6C3Okpuwwip19JhR1KnYnOVJwD0Fe0UPzzRSWJ3H/pYewCrLC0u91Xogi/
n1dyGTWIeFuvtw2yDMsvH3MFoR5XyAl++uC+bpixZ+IsdYHU8H7m7l8aT81fryuwN/1/eb5RPvT8
P+fMgd+9dDV1RiFa+5k1lTmUv9Y19iN7PQbeK6htjBG7GbfAJhxgeJoan2SNYVrPX4Kb/4unMePL
Gm2nYkUn/so31CU2XTRFVxE0bx7m691Mim2g3icyTuNeawQO+/ENTqCOwHwouvKerEEJLnsFBE1n
vmmLuXWZU2PjvH3kBPQ5VFMkm6cbwmwmSXXsrrPv0PuEMFYM9+/LvtX+kOYrIAf1rbR7bPMo7BbN
sCt02t32NC5k2YHhttArNU6xpv9tJ9kf1hbI9T4jGlgcsQCKtryxqiM8tCGlholCEHq6uEiIUjJu
ICR6QFUroxUYA2DFORxNNJ1EdZREuy3wHMoLNfSAWLhvRDxbi0fGqQP5CjT9VepBJoyWpbMseAwX
W+25WhwyabKrwPFktzm3jrzB9FomEyeSeX5Qqs4BImZLZ0o4yZriInSzbOle4HicEgrXxpvU80g9
zCtKLsLYK6fdeFe//GO9UJb6I73OdpjBQP830xo3954IbWba0GJMB/GuYDnnSpsMgZzWVm/1/djv
hKQgleEqRuwB+/5D+gQxoxFxCPWOXuOxQ03UIFo4a8wXfF/zVod2+vXsQLrTqctPFUCce2zxCcP6
47lEP40lrVpnVHDzs2Q+koaQI7V+Yc/uciqIOxuZXhjCBEBkmTAOC4BClpHaLCR8kXyjoy3sBTU7
lhGbSYOcaSkk6C5WOiYbts1O38ypCXD0fluL7hxBObOrwqnp83UdvgekTnY8wKCxh4ETTQS56+N7
klN5W6LpWpVgO3IB1OhAnJIKXPEbfTmiXaOqpkNxBVweCYw5BEh8LZoxgKZvl5m946YtJJ+PGERf
H6hOupVR7lQngReefkSJeIRQN2bAPP1MStf0W8zINdcXboEmrW5m9WwL5glx9VvtlbsT2x3ZY7Nf
WBfNz7qPiplrggqQRSN04GMRbVo9Sl2yVs9UxBm+7sXQ5oYzEPYzK7cWwMlA3j3AFEMe7HSW4kQq
JW6d3fubptOXw5vF/34scNjmQ9klqrfILHVuqJP5z8as8J/aZcTEZ1ixwZJZG92iqWWIbEqiT9Kp
RoZsP0iaJLzEQwEMRSXgmwthVzFpPWGbxJ2XDqrOIU7Y4j7XocgEvSt+ulI6dCjw5H2txPlQ8Saa
IjvPnuwdy4uyieDGZEyWud+hWYjb5FSuMGe+t02xwNLBEbv+q2+ZsGNOKAoCBHRwyVak5avtBvL/
qgIFzxBbqg/BpbsaX9XT5Pmr8U2vGjDqZyI4ig3czps/YfoT3+LMde8PBF8NH/bCJAb77uUO3bBF
S50ocJ4xUOEKZS5Ygy6dxye9Pcd3GEwIBuX7gPiXln3PBBZrSguL2SDAuVxyjTL/S0mG4hdk61xI
tmz2JWpN6c7LrcGqpCFbUGYoV1PdSZR7qLOQ+g6eF214tGnSmU31vyyvg8hpHBrOrzz8D+mIMYO9
iTXD32xHFVY0iOvEy/mE1IWgucMsDyWkpc2folB8CLIGay5C58TWS2Dx8w/D6Rjhc8dbmAQM9gMr
DVcATHD89oVtXlHMa/GRs7CZTr19nUTXKuqLxCQGSFYLF2VRXMN8SquW4/fZxGXuRCLHeWft72sp
5ob0OzFjsXcJ0qetmFmbsfbmkG32kit8ebWH3andFKIs/1FMtlL0eEMlL9AEqFr6DK+b9iDL5Cl4
t8fFcqpOKpb5nGbjspaVvO3O7hf37ubNCexfYdLjaqYzYzwnRjW6K6oT90ealtDwiFH+FnRu1Nwm
fviOHVJVEHN2uoo6jFdPgJKeGY6ZNfmQYFwiMXJHoaSbiHYM3ZutU9OiZO7/dmyQaQnkLGbzzp38
u+rymGhfwExvYoUXuBzz/LOa2kCqPCG7QtkN9RjBdY9ubPcvd3XCWgF1rXXLafMr9WusoABRMJ9v
ZNdAywAYPwc/oytt8Ya56jifAaFCSINkdLQMUF6pqziZHj8vK+qGa8C5uGm7MD5oCxNeqbB9r+Vh
mHlNy/MwKBP7GM3dz5WvMuIE4fcyuSd1XKaX77JNAQ95oSvApNHGh0JDkOPzXOUzFYmolzUnBLsq
QWuHFtMPHpA+km92yYlSgKBSSDSfwBTt5hvfV1XUHV06nr6AR8/cCEdedJccBDYAK8rbe/9t01T2
cpEO0igzGpPppOnSLNzfGhZQSauScEFaPHfAiiDLETY9EGuth91nt55P1X8eqx0AO6HSSW6w69wi
c+8lA8gNfUFiN+Mzgf5vqxcGXMa2cOZN68jhBOYC5vWTxTtdzzKzG/sd4RrRYagfVjEZQoITDRS/
bACcAeA5Y9o320PTz84wr8j121hrYgIk8OVwoRSIDWSFlWoiQ8CJ9YeAFCdeymrDjXEJi4bnM5E7
SuhSS+sw2lNVxK5HvjB+bem94DOGjFIoiH1YNd4xHZih4OnWOaOXAZFI0WM0DzOZUQqxQnuhBTnF
zcxQ4MLAIleGLf0kLeA++wMUvAdEFRmIb/t6CsTfMa8N3tYV6hzyAEqsQBZp3boO1siY246XcSp+
XYGvlN1N56qj5cNn2NifHw1KhGKFtSrcj34aTgOF0tEg8iFBjuk1dbEgGrR93WZbYhqUeie4wi0u
89W5ejmcsIU8/gw0HAgdcX9aCO0ml9tOBZF6I4gbC/t3CscJ5o/5Jw+MRbzOjA4pqV6tSKNRExla
2cWBL8RfXxJEZBwQYmWIC+xN8VWsrKNub71Or9d8zBWnYcJW7V/9huKE9vKSNb1kndIi33Gb/LIK
9SZVY5AgWLPrvgIfhObLDE1Yiv9rNkgVMbipIx63/N6AOS6pOmne4Nd3kqsKYbOZI6RAGfvDTHzm
7e9sdVcfyhtuYM9+Zy3pM4YtLQV9jSVpmtJiLtnoNtcNI2Bf338o5kRrRWBVAYbHbADj07QIO+Xo
9SBnAuhy9qdZHxHm4S/kbcx7K9+sFWz2xNcihE7WMg47R+xc+hSdBpEK7HyeSnU4pWrTyppqgBa3
WR4hKbwSwifl3psm5Ghd7zIq+igFXqlVUprc5nE/2I2ByasDTi5N2SkfjLapJyyEaCzee3+t5AK9
w72EUsxZnjO4f1KCyxMEjd/WHgRLQF53Za5xCtL/PCa4AZPXu4SZyzsQwWw+ou5BalnmixJgmO3y
IpYdz/QqcIUxdFkj1Vsi4gnOvg4ajC4b8ZqjfNzgHbuUDkn0Igzkm4nFw+b+6sevjQGbM2eb1FjZ
uyprCyZluw1Cz/adewGMGhxm53wC8XfxyDgD7jiL0lAAKSPCvnHI3yYSKZ0gQWrkPEjzHdZ5qZLS
rss3VFVKR1YSNhE4kBFRH47TzOGMTqLBQxoe/KcNG4HP/YHJAn+F6mxkHJv8kUhqlIB1sbybKnMM
+aTkl2NFq+rrRrmTxPSeS58SWYLac6hccIsNZMCLCeBf7X3eVoT7JGGnyaKuvrsh3s0bPme5/rCH
BWT+Y1JecfNOtu0Iw4l0cxS5zGdR/xzOeKy4VXcUbcmARB2gKuWFLoeIZ01sQy1p4OwGKsoPhhqA
797nO/xzNH6bK/17STwVqjnjZHl8bvPraLhSvWkzVvEISlnYO/cBrvzz4DCuNopVDIYcb6fV8Yoq
JedSvd/bmr2Gt42gIxmQBG2CaTywaGBe/XaAqIvJbcVELeSRqNWO9If5xW/jrWfCku4UlQy3iN9w
CXHDaNSvnIztxM1bxoRkiFm1Qi/5zg/cdmBKr4sQPCEFHhYZtm8N6jh2/qJyKgxFd97HzhLE6wRb
D5wl2rbN9QxuiymzI3kAPtL2StcL0b2HsVQSB7dxpa2eXkqfyk7iTkob8q1eaw/YLI9GhwJhumK7
ZN1fDsBwvl0z4dvbp7Qa++wg9gGvTiq4+dKkGGDTrgxZyTH8GxHzIfZqi1TuO0N9ji5MDnkVUDvR
H5xAgZXBA7kMwm7MSHLzpS8dxXe+Fbq45thapTJ4mBVvY+tNfiTEnZUI0sRyIuNrZhufcdtgsqzv
eR4MYNY4CA5H8ESaLpodP25B5E4MU0KoHUd+8bHiWGtFRUdDY1LJfRAR9Ly6VrEq06jKj8hnSpmy
CMdqlW9gmsDNvd700rbHgBV5/Vwm9T/fdGsXOhhwGCN35O2nIo2AZQVfgKkPsHW8fbvZ2L9OqKMK
ipK/ZY7iQjG/1rHea7O6yLGZcdIb5ZcK20gApbh5vCKkptfDr9WOChorUe1jZBvUespJb7lPLHzX
0kY/dxyJkRVaA4lYt+rtp4qI1g9xW1PMy4wTM2EVANYb1zhTq8BA/6Hv0FHZilfm2b6R7a90MH3t
HOFolG0GeUB07WblgsuyerpTPPyFvYBZDUyouK9B/gy/PSr9TpBjv0KwLx9iKGfScMjvuwqVcXQm
dRhPCWzspyTTQcDfGpyC2WjLOonSGnfp2m8RNJdnQxGAeWea6n7PAlel0onPKCKUtMJlGCql60lN
Dgy2KmH8X/crs6jXi5g5SLkLa6ZBj1d1Kzpe9VX5pQoyoNjhg96H350h1bEHP8W7a+i8RvMHDwIx
v5fmFMjgJkTMEvn8HYmHQAA87nWomyIZ2p0zOh3arl3hs8PGbfvLBWsX+rG+f2tWDcdea0ZY3JVu
9au61DamottbIcn8fYrZAN6Opiqo4k22IfmH/eEN5GLciLDCUdvcC+qIRSn9KQmGX0CHwISmkaDi
ExXnWJPDuMXDxMDk3MGRgcJP19yqAlyiY/MRyIUsNr6ExWRNRFvHSMSavve6wpLdMrjtVAPOxwTt
O0KGN2DBzvsC2UOLPQYqAFs3mfCeT6YMusAVLViVMMPtXPp7oMhnqX0BAiAjZ+m25NB+QHCYUJBH
7C2rO26LhXT3pG8pW+Ou3YS5G1pPAKGQ2igiEcnkzbmC3ha0huVNQ9YdHn3/+u4SZkz4yEhzu3dV
4kHBUm7CDC83veNzvj8/yeOcLOlCf40DrHFAcXbfwBcfGKSQwc7PrneuZ7lmh3Q3P0U1wxsg0ZlE
lxKxFjunP9JsO1QBZEgiP6zZmS7xniGrfuDQWFgJ/OLfiDoG6T9lRNXX9s6pXN7wiiSJy6bMhaMk
+7VMnOhGnO/3oJRIXWCHutx51UAMi7aa/9GXqeo2NOZrihxWbyczjO1nJN/frCSe7A24MHEDgDqm
tl1KP78e0P7UVIt9NO8lBUuaMjY3EFKy/JvrtcTyDhqwD5/lbH0dDjRnhMNW3wQXfHfckzCk09Ua
o2bOdyndiKEekg6JHnTBtArupKt//MyDNyKjyLv9hPRMcsh01X3ghwHAcYEvzoTFX4NPJ5XvOUas
jBnhbhbKvHYbe5oC1BOVCQ5RYLsGMZxAkKtjpZ36R8L9XHS+ppyjo/6GvBRCbHdxXL9oF1UEllZ4
SFyFMRyOnI+cMh8DhAc9Q0wzjH6FE4UclSKR8737B0sqCh8qsFjt0luOdG8eO1JpnMMXmLPNclbX
+RPOb5Ni+GKa0dtv5hZ9D9g6QDjkAyShd8YzSFToVO83VBSA9mF8HgwB/KbgVotoTKDtL9CeTwgY
xTCSD6OA9DX18suDNoDSQyKTsmqXMjyO+mcKUCa51nksGOAfMTZENj74btuzDVW8NJFwSXU8YM1i
Pz2mP6GsHzHRvPS0VIfOBupDTcuuziTdNKKleIfBPxju4CId4RBTffYKMZjRFqBcKz7CP3ntZUbG
Az9L9uRLGM+WZxV0Ai+mktC+j7ksUI4kREqC+RXEtFaTwW00jKg812k/i9sgzHbkFl0QM0iXKOpL
7brbbhp+HgZ9tQg0DhsyY3dz1gWG7QDkDblTkxoNfKnKTIcsnCKZb3GvrcFigvlRwsEoezMXb14s
uVlmfX6mksnMFNNYC8EcxCe/1kW9KHzafhi82V1lewq2P+svNVORj00u+frLHYg/CpD9+++fYOtO
hxskXAqFdzeOovkLA6X6jPTWbYe194EBD8HN7TZ7lyHRwfqAqcxArgfOkSkRzn+PXyql6E55oMG+
+xBmsrQ7EheogEGSWSxlJ0IW7LFdGsm7OiEHjepBMqT/Y+EkNMDS+dedP4lzfEa0vgGeFHWYO96w
8c5Tz3Ra142GYw6CUSSKGH+D+yWWtywJJqg4iZQ5vz9A3LfTakvC5lUXnE3TmLAHfkzA289piE1h
f05jEOzvGYrIKj5vDuNVCqtrR3IUNd9GE71yEhTx1gP+wRdYubHf3RCJEg93b9HQC/C4Aaod0S68
URaY/2BM/n/sQepgnsLD780V4G/S/T/139ROLIb2PFtZQAA8vgO3RsuYzxnpQUmA2AXlG1YqRxWV
Qema/7SO8FA9k0PLoZ/gjfOcKqTwnJ1vXVYQ8z6+KkFs7TvezqTIJFzwEqS8IbJ6ZYVx0vzXLCBz
bXRfhAu9/IgCuxxyMCEU5uyVaJMC8bR6fQo7wSmJC5ZhzexIeaS6tLSNr/RGMbPm71pHo+skeKYy
FVpJX3K0uxrJU5BtckVrAF+HmrAoV7jrLhiLBRrVDc8FvZBUGNqCdzgdNXl5OJoy/JYki0RayYd4
6UhRnEmLLApZfFaNFm0lS4pUnxLGUxbvT7xwT6G4hoFSXJjUjH3jYxEJIILGDz1EHvFxyv4NPjIS
JBPmQYrvnz8JchA2DaE3zVDDXZBR7+6n27WsEWVWf0V1owVdmVyigSY2RVE5ekJY7stYbEGhokhr
/VeSzoBrLEWNEGxsUX8bvYc9hpgh8KeL/RL1+73UAvRKX1KgZed3NlrCmgNoZLpiHeMWQNWPiczG
w+oTTbXWe1QHR920ZYcSMZq3e95G3YHfUPgow6fB2wpvIq49n7KpPacPpeWebypy3G5Y2lQcfDAh
vTga4haiFfU/i+9evdk7nlo5NyDgWDLd9ixr7tKP8nGfMpgmNpocL6gjvvFgdJK9nEz94ZgNadVo
BpOC3v+StDkla11rTuWYumq9dpQtjwyBopDkJpr+tTyy8aG4wEf9yCLhaQhwrfG0hjlF7/wzpsyE
D7YfJr2XsGxnlbjzlbEs/YudkQPXR+zaMU15XyoULv3NXZjxmxYZdbkobjA2s8Yrll396KBfNoUH
CWFCMIrI6Aouk3zer7dWd+y5cIMPKSh9P284RKE0qJUgckxA6cnI+4XeL68EXflL//cu49ZWLqtu
JBcdzm4mV9vFNTn6FyOJEvLyuy7XtUeVicm8wrB5d5AlTRJItOOFM4IkFqQ7UuqkDKBsxvNRb/CE
LZMrHol3oq/PIdJLzGsRlVvsKd+80n3bahgus/9//LcK8BT/lxq6pz2P7QUzYF5AOJJvB16ONDGK
aEREqykGu/Pn9Pqq7cxwcgNOdOfZygXj4NJRuk5MlQtW8BQ2HLH7TAKykTaJbWJJXmhp6jEMPrwv
Ol1vaJ+8iVm3KtNAak1E5LdvjzOhZxHaY+akwJJK98MhBJ+KTyURfiuPYA6woru97+zjtBoWtyp2
HSuGTF37M7qyOI6OBo5hqnY9JxT2IMyVHbZmvdpg3TaE5TKeVa5kA7eed6OcdDRIba5A7jmAn4Jv
Qn14EvCNpjyeacbnQ7hKTA5dGiW4tCZN3s/Vc7pxEsESBXNOKxcoBfstKhgUWK9bfJ99UZEM0DsP
v4APYp3zQ7nncO1gt1UMqxhPoC5cj+Tw9dLgmq+m6wgmx3E8FtJRJwRSq9ZWs6kL9rgXzFVy99FT
+SmOpD7fC7Eg3Ovuqy96n2WZAT7/p1V8R+mXVhcfnJg/xkK59ybpfN4NIbgeXZPjojxwJ5awSqfQ
4JpDRhDm7n7Q6oc7Z97gh3B3RIR7s4DwcSoJkfl5M4lmXz+PpdZ8vWHxsFHnKHSdebROlqGfnX9t
NLkWb9LzXbjRTXvO47cfJFTurpJdR1CJLmWOQkOZFX3kg21qOlNfXMwjppKyjtTAnfcK0pN686ph
56h3vOgpSsLkBdSUjt8R1O4MxIn7e1hvWxjACHcoKhm9qksVOltLhvMsaValBwTYmR41XaNh+WUC
TEv87Xu7rgsllU0e35gC0DSx5K7FF/Gsr7Le01AEd8L97WOgWeVrkSljRe4eF6kwERvas9Qf96Ny
MMplOlwLlrnKNqeQI1//1CfaFAgc676crhrDT+3k+oVcInvQs7s9YYeL490yC+Y0tUUyxdHfFPFd
um1rdh5K0eFyzfBRGAWHqgUV6dLaZAZIEZCle4I8Ysm/lthsNfmc6XByL0iobjC7ZxO7Ikj7U2rc
/kRYuwwgghbQ3RpD0nSnustsEAWO8wNhko74xCubIfvnZXfxtkE60Zk34TK6Xn838f+wWsYWth/V
+1IGBVtrmqqHm/9pw7dr2O5j/KahyViEp0uc6myXTavfIbG2AlwqhOse8bZuUhV6u35L3GskFTjU
cQZjIfPIexdZ/WgEwEK20jyzKVuwSFE/tppyF0PRe3nHispETdG/264KjXeBxDvMOUNPHy+BbyXn
CEcBV0Yg+tcWncCJYGTcaMUepEphb0ipXfHJDUweFioRctS8ZDfBs9+Vu4AViFk/o66jag6sP3Q8
OLqteUzybwPDqHO59WtkOrnUEKS9hZ6iaGLIhNDc2Dh6hkoqtHZjkxJ8MxCBjDT9Gv0WAGU3LoKd
hJJiDgmUcA1/DcSWz8SOlY9stUtymgp7cLXr0ONKrfd5y3A32kihoUBibvCqx8Dy011oQ6DcdKYI
YXQ1GsbC3Zu0LSX4/TFCjgQ2Cx1SGNJY9Snu1K84noQp/R03yg8SmQMtV9LhpcttnSxJrBTdsoEF
0HQmBdtGJTOmPMLpPRd4YrPyx93zz0OqvnM+fA5NB5SZr0tdxmT2nf/CQz91yGTeDUCW3rBWng8k
demFk1yN0VxQ1rt9d5gyqf7qU+M+Obo7DSo5W1GpBknsAD5NbSglwO2oxk4ADEpCzqHrSzkIExTH
Jt/nFLwzo8CFpCq/1vCUXQZxIDhhEHLkM+goqWSK1MEVKN84fFmW6yjDEH933sPJDzevvX6QB5JJ
I2W7KmECJQqZ92JmKgyzywxyhZXIApRSs+awb3+hy3yQjoQFiUrlv8DPf509O3fCWBrCw066+2B/
OTjM3sTfIJQYnZVuI8VZbnaemCa1tu1UVU7+9b0+c/QsxGMhXRTO36Ey9nmd0mxFZB8BIRAubwz1
9kBehWx+IkaX+daR1xKme4T9syHROAL6qSfPrGkQZTpF4tJK3yaFsW4HM/A8lo3a6B69VzqcqZV/
6/ANgogBuhL+wY2tsdnZsoqtim19aMcQBzzspU5A2AaWpX8rg8U+Vhnc/PU2739jkhDlkafRQgrf
mQ6AdlKZ9rj84C9ZjpYCTC+hC87JKnym/HuFLCf1YsBDyv2+P91Mr1/0r4cRCAfzZxA9y627cf7K
YHpgvyadXNH32Bo9SPo9q4ajLckluWX3F2bAyXcMvabTX9vijygLdtZEWkC6jsmHMvrYBHNToNTy
xmCePbVTJKZy0Y+xk5q/JiTQcCyL4MBLH+9MG04WcYfMY+nU113b5OY7WSS6vI36nXJ2goyWlnBh
CKAZc8b4pMwx9vM2oDCrBpgJaoyidFj4UorMGSuTvpFq5eR9TA0GoOsLR+u2wwuj71TJ3ZxO1hLq
mrUxhQVIvIHIDpzaOuQoIhXSSLgwqhjlg37K6q0uSt1clQq/Uw3Dp30C65AJZF3FtfVcRNQLgFll
v2+iHxYJgMvYqy3Ea/DHUC5O+7cAHL0BsilnglicPLGIBfpO74qfJ60x5UkA1HGzYINm3xghMtCG
Ss+3ACKsYl+CCAQIOlILhy/mB1gj2/15KBCgd0XXswJ3bMA4FzadJzIv6BpR8Ee138ayisXUY/MF
AuX7oM/KkyqDPitlzhmGXEvRjglb4AEWyyLkGUX8d82PQrLJDVK372Biy4hGgSKHHoKdYZpMvsOA
GlSYu+GOpUnYzHgQco92OYd9EY3rNVu9IT5QOLuO7XVX6imEQwhAH3qb/8CqVqhRAJR5ymH1XKQP
58wVEjoK62DnnO03moQly+zZ529HpiJvMNwwB8vh579Jhvsx1Q8tHqZPIZoetBcVZkQj8wf5HTrs
VYUtSYzXK/VBeh8cieuHgiau5J4tB6zaNxvDph1GvuRxngOTef6IvA3ItS3p1AN4XrBMigMWafox
YFawdny5UT2hc2OZ3upKirMNpA2YxsfxAXQUcYFgrQMcPlWfL2+MVVA4lLkSTzh05gQcuAsrNb4V
AQK7Oem8WTqbGe9I1lBvat86LgOjzSYNMGY7IVs6WSKf4mrOl4UOS9d+xwetM/cIzUw4hbDMfmRG
SJAkFb1xAZoyDebEgEFG2+czp7pwg5Gfk3Xdxy8Y4Dc3Q7OtMfDDIkF6rzvfWsRa+87k1Dww0Sa/
apUumRpeGpTpWXg0xfi8lFzTSu8pKkprnjhfizmBnH3NYt2SCx1h5En9HYR+tikm+ElmZfsCX4wS
HqJ78YoiedolqQQhHoK4MmjL+XRM2gtI7b81CX75yNQdfyes7Oig3mXoerY3NDPEMe7d6bHJqK7O
/OiDZGSCm66tLW0ccMAJ4Cf+tnF9hcD2nHbe6deJpZhc6CWD3oSkJn8rOGI7uRLmtkUd+2DgMbMX
9qe4DJl/I0x0vSQstdtXQn/C63Ku9bfcIF5OlPOLZQHmD52m8eSddw1GArCz5XcoDRFQxuceq3Tm
iVaxQCpfzmF6UKlSystJuM9DPe1bwKeR9jxchTotr3peQ4wpMNhFkb4LglR7MmZ6bq9onmQVxV1w
8N9ROevAaQGvimO92fA3SqM5STcNeZVHanlLTUUIda2TeydYlyGM+D7ag0WhiF0KkOP09ny9lazd
d7NTrpD9+J/k6Kdp6dE7kL1/Sf64ojzTlnTTWJqAZI8Ys891S0t+iaZO1mYhKIgIbdC0kGnAx6cR
jPnC2tLxUrF1Uhw8d/BggNBDtPH2NGQgAdnez/GT1VPH/LOx1dv1K4zg4x8qgK9rJv3pJxwUa8rn
fVXBZQFQY1UstuyitxrG7N8E05Zu2yzA9Vmbw34uN1rEIFI1GWCTpdZJ2AhiHAi/XXpMYLwUER81
fqZH3/q+AKM4kDBUWUrco02XRUOkD5QFiPXLBIZDCeW+kGAz2QnT451i1d5XS5lz5au35EMfrIEg
Us0UIwKon1vGiizilDUluw1RLGvYlavOBm8+n1irHdE4vvk5JzQJ/jnYcS2nVe1df1Mv75Kv/M69
wqXVMrm0xrpNk9B2mKWMQ6vJADWu2TjZEzBC1ZqRUCiGWvSsOyhniiOBRsQdg4LvVqAWbDQtbwtH
Mm/t6f+oFZEpBhpaVpHVCcpIbsXwLXQqSpVEkN4Ffr/hKYuz8V4zDhRnxnKhmo/OwftIUHo6mHiq
yrXuH2L2MGAi6Lqs5DQvR95/MSM0Suqt8IsdbjystJhSDJmMMBOQUwj4giiBA8+ncoYaCD+XKVQn
vm9tOh1/xAqCXGB0IPelhGhg+NMgbVfNRHa6WVoSmpN4ZHrDXpALlh6ZKkXOQ24bC6e5UXHfqtdt
UTAoUeGmskikfyq8fav+YfN9ucx7c8x3Uvph7/3yX7cjVsaxPI984mAQhpsrTq0m/p28gc8HZT+0
V/Bu1HhuJMjqeKFFFr57ydLt6799g4hrICd0ptoPBqt3lIGf2OhzfeBqWd/kExNlp3pDf78nrpfb
ocNRWEP3s318K5FnPOJNRqw32qyseULB2kVuX/IbZvo6jq19bOEcbbHbVbbRi2hbuP/p25Od9+jB
3lGimsTEjI9jUmmSK+yRvKzIysPqtT2ixAdK4CJ1tn5St9IPpgMPkOms5MPFOYiCqRCbsQv+ZSEa
RLdi22FXls6eRYvs5l1eNVtHNnD3bR7Wab4OSvT4OnFfD7QEEusRHhzfNu8SNb6wZt9ll77Vy52h
4m85/StpXc19cM/dCmHBUcxC9QfpPM1A2OV19X3dCrc9Z0gObCleVtBQi/xd3uoCRQCHFadWuDYK
yTK9YTJy2XnoaaFnRGjdVXZ1twI3FTrHk+1K5Jx/y3EkFPOm5pf5bLbWDkKG+GSdy8bl1Dk6hlWv
aHlyDlAZDA8zgkPTteW8sx9soYyUxXgzLIpHHhUGiPAGdF8z7Trc2jrQwR0/Qac8f1MhBDaHmdGf
7eDjhAmPvOcrK3GC9sxaV37QAiIdI0H3bIfMrBfapyvtZgumbzbxMdMTRH1LMvv34bD2FtIaqWHy
vge5oy2wpK4g1ECNJ82J4KT8CMVNmJsre9wURbXjQKSPIuLbhgV754nW1FIAm7FqpLIzcy/t0/QO
1dqM3u4kkBKZm7kQzTE+9IU9e3jBczG4MdO718IidEA/pAE8j3UwTBmkrhezmxra9eCCo9e1d8CC
JiE2Ar2r/SAdhLFK8VsppvdGHPkTejwZKw94mEL3WVpHYDAEek9Fodvi8sCvG2CCa9Bda3KHQU0W
/KTrIbsojPJBBiPUw5xzWgRjRN312KdTMJVk9Md69/moHGLVgFxRNJAwZG9a0rD5iW2XyunXPjuE
EOdavB/FjWLFqRMgO3WROacriMxqKG7YajRwV39iP8dlY4ksvFPmvrdBb9UsedYuamd0IS9zntnk
KSIAGY5DFwflyzUSlnVn1GevQ3a/AxsvOIvXidEL9Z7m6O47Lv9aywRQ3z7rxCFuSx/nKD/BqVFU
O6Mqdn6EIllmMlsomNwRntnIErGsMBhsH5XExcC5fb8/HghLX7QMw/HYkpynF1BZx1I4DoLPlE72
Pi8+4evp7FX/qkaTtrDA2muziM9ssgVOv4SC0DdOdVxe/ShOa73BmQs9hzaUMrPppoLhBnxV8fVW
tXp9xZEOC5JsueM7R0DQugDibZogUadITYlX7wF1G0k+nZka3Vjj1s0oys1J+Xmece4U5sTpCE1a
2NdpD93XG70+coXSqKH9YqTn2vhSaQeiScmQH8+u+S9ODPmfJ2A278+JsvxgWDEGqKWdTbyTGck9
MVXnFYFXE+UKgg0Ac2/lwQVl1abELqfDPaixqYT/+PGSLi27Ek8263WwAw69xvo3+GGfoJhMq9ln
yYmZoup8tpgKBpqkbQ0goo9Mpuj1odmo5UnMfeI5ePlBe0x5PxpM2CibtwDI0FNi/06I/Y8anPaL
elsxutdWKtbACVyLPHWe5tMOYdo4WszxDA9UcLHDntAWYRlg6HeAfcgtExnwmKo7ifB5kShZdLZ9
9oObE55KK37X2o8rJh/9qoLQhmfJyDT3e8Iom9Op9zw3jN9PbykiNa8Yx/dLeEO4cnw8+kx83N0y
yUdchE50Wkg78WpiJf95N8D7GijZDhyfIryFkLRCQhZeIyWwrzOJYlFqw0U2bedyaVDsR7RlQiLt
UvglmqWaj4Kedcp0xaSPE0Qs+Q8vOEapfgInNNYP1n5OiNeIPSkkT0aN8CcMR2miwDg/fK/lrbQM
N7RI/MZ+PZ9MQnO6B5K8wmPZCnoTmnnTh7j7k02fN1SIKVybErFT5RT4g7FI9DHTMwYN+jXYK4Ua
qL1WtiB746H1qSNJY0Dlv4EE2PUbPcUUAmClTl65IVYnmnsvpDHSjDxEDUnfds5WxfSffOGZvQdt
LIIymezOQrVeWIJHQtxj9WUVeAhSzv6tkE+aJ5t2vHZl7IU25DmGj71aiHii0nEHoc9nPRq85T7n
+G/d6B1uapCnlhKDTlePybEJCy9TDaqypcu2l/sfCp1lzNMA/9FE5FY9ulREcgiYCp/jwb0ZJobA
TH4iwXH/DPSMcPRPiCrMP13qaEUbdgaXkGCb1VtaJcEJRYi+bddPAoD1gj+5VGrRmPiGCR4L7EVC
jmMwrhOOR/5jP+rzwC9e+Hl4u3eeFK7HUblpUIEXDKPG2eUpmm6ApFWlifc9Rs6pDaA0+p5eU/EF
ZYU+9Y4SRP1JU+dk+nyIoTFQNNMYgIY7eIK7/+La95pNolMaCSOhtUk+UzJsKU/2rTtzeZaXZYmD
HVFT8QBs9E6ftLylBjqdmaE367CtkqIHIXbKlvVn2CNkpKvNvfp7WdrLK2+0ai7hAqA5D/LjCV32
3mKGc3rdn1PZsnv3qGQuMzFT2aTx4H10vn567PNTze5ep5fzAGGphwLJuqBDiPIudJ7MCDfPFB9W
iV+Hs3C4W0hHgyomqIUbOdJA1RO1mj+xuS3Mg6X4EG3GE9dsTL2TkHtZve9rkhiZEZxMm4/JOlbZ
iOcnCgKNGc3wKj/NHnWPrle2WwVpDpQlxEV9KYtktZyGm/jGdmXGWOlyGqsOy3eNns/4E92l6seC
25eNdgc6ScxwAu/bGiNEV0U57JL18uinee+FZxiaoEzb+lalfBrQVTBw72isiFfOngiX3X2geu8c
DY8hDCmQCwqVT2jeHTFRHd/6C+ey1tGGKJSHL++sDktfQOjwiT7oVTib7NBFXGBCEohe/Jy0iti4
oG4edceTz2C4h+SvZ+fObu7tid9LSrvqrX+9wUwb5xps2qEa653wENJa9/01rUT0SzGpsMpStItt
a22tcRuhYJO57Mkl/MG7HBoy86SJf0PreYJUz/j/BpREUh5kFJKE1JnO9zl/YilaQ1r6HdfC3qhL
vEnN1W/RrolbCXyHd8VwXB/VxepZ5puLyI8pSEsLr9SGu93qHcv8AmOoBPplgQbEl+KFbLN0Qxfz
ih4HVTVCy3AkW6bjuuCjo2F73LfzIEHpk0YloVN6CRBgov5by8uAoWOeqc0w5xlpoO7HOpFscv9B
/WxE+Mk+G1Sl4GfuSirBn41Lr9qdkypXxiHuH53peujoQp6k/HDa/f4kYZ6Dxr+Ei0GBbZa90Vid
/oEgHjK3DKLol9IviuLZ1CKdDGU7uQclxMHzVGlNC9InLz+S6TcCdgsJBf3K7LyULGnId8xB2BHC
udYyHEV7mru0fvQsLYDNPB8smodJpeJFE52YJ2HJAdoTZL9lVjXOG44/7V7vau23i3P13NzVuRWQ
1i/ZjFV11P+IlnlHf7VX++tq8Q298S0osjEOoccUGfpR52LPrrfQtBCOUd0q8scVfCLZuQFzL9dL
B5xU8nCu2Vwepxq+dcyxj8RkQSHgdHyenLv/UncG6LTvBpXqUw/A1O4NxM0bsZsfWuXbnIZ/icQj
OSQjfNQtdlhIpSTs7OBoFXG53mxwThSArvJBfMREwSI0fwATPGejSQKSiwFt4aNonbFhL+D0tsn5
Bn9cZs5ob9Uzai1hs57dSDjYdx5Ek1HMvhrQ9OpZy79gZ+iVtDUxwxfCghOPdZsYFtLwnf7wayad
FwvWF+znTkEHgJ66KHBY1DK2mf7yqEiSdu+A6vUzQ2BSumwUr6wAG6cUjopKpyM/NrCBBaZZYuCd
Ojlpauioy4jvKRajNEalO95kR8fEmRrjjWjxkHCAKRms9So0UCHZrH0iZSxmX8Pletn1q+RZKKsW
bUUiM3kjaUcntoT3kaQM1oWap5QXUGO6qkcuLrfE211+SLGYPOhfkCGeGmmDuNbckH9m3AMmsVd2
Wr+KAoYrBGps7z2NDDt7HEqeA5IvNoIoJT5LIbM6+FRSSBAWrkCsXy1hzdhrUUEGzaOMl4ynvwgn
1lGGi39XV0WII5j8WWQsaNBtKsC8atqXKmnwrbHk8Lyz7CaACSgIygoLGQQCmlRJYXl3Yv1Bluk6
4CR0dKEttyjWsluxWuOvFaHq3qa/QJGsQVQ/p/+nJWJaSAWo/2wgXpjtvdVORnQG+gSsmqgfXGY7
HoGKsCeiJi7ifGmAtZ173njGoc93hEhDeMbaxBzysLOCVvPy/yd3AGxRDu7IQjZatj8SC/GLVUzb
xy6t/Wi24sfaQYq1Iw/hQGG7HZ4SAF6wtVcZ6LBSB3IEcoCHtVFchEdSxg6a7CQgb1GI6QtFWsG9
l0/DZaIg7lnW2iM2FmNCdZdjm+Rhk0hq5m3T0Ra17vIzLh3SCw2FJ6RcZ2SwOekNJzE7xTPJ4bHd
BVCTdm8Y7vwBgJskyYESeP0VuBbTBG8Va9Jad1Bw3+loM8A16bm6EAKR2KHw6sQF/4AODbW/G+pY
grhQqddTOLjG/k+2DWspWFEK+/k5WRFs3B3fD//xZvtQIjX6zFs7BYArV/lm8nRFq89D2e3RQ+Qd
bVN1gWMnmWPJu/RYTT3Fqb/7ADLWq1SCoPB+XJNIQ8sXN3tV2Ecuk2+IyRRpwxF2zPYtcVvEhKml
w2MX1J7oi33KUy4/oFQrbaJbZJMYqGMNsXuNWR7cUwKWxg6vXRwG9uRvPvIVebrH7CP8GcpNwz+Q
BlNscIUUulnMB20/75cj0z6cQRmU444jS3uk7jtkMhU5YisnbVVP+zXN7atl1OrFpWzpmE3pWSBh
sWiVoGuj/yaIqX3tKIrMfOEMcRH4sfhNja1Uiu/Nl3TWfEPrmKAZgfzEBDOAvnnHyk/Hq+/s12Xy
9kH3wLOsFAunIyTEL6JG1BySoua5kO1l95NbehVvNF1dEUYp5pfCY0gavXiT/yxBZUhcEYhQlGJI
L0T8+hSp5hO2VM1F24yQxi3KZm7feg7xGT82WWHKDEN8thm9nHHZBiub/NPzxQg1aKUWSrGyrTa+
fWl1dpmxUzNeBE3fDUUYevWufu2DSDvOEc9Oq1iaWbY5hy0YMrADBJN6I6HSbrNWhn9LS85eJG0k
pmXFpGgDEsoxP/viv3E1T8lhdBlToG7rh4flYWCKel0dy4wqNy94gXoRU+xRMguKeDhW1kAPXwRl
HLs1JhmnoGty81Nqum/J7fA9+PSE5snd1TZtTD5mHMss9/I9Od5w+R9wmHt2j7gTplu9wYVsevfL
85u9dxgHUptwE63BVpjBHJL8N6Pz+BcZcNs+cvOm5G8Fvy4r94zfF/GKqTYqFu6Lm344MLpoBMEK
Zq6vkyKE4jWHjujHVHlWquXjWhW7HidDkiPLcZ5/6Bax5I90tY90r0YU/TF2m6mlukc/4OK/p9Ge
U0CT+ilTsFBe6Rd3UY+11OZEsYRUwBVOJXOKEUzuSP6hkLxUe5JaohDRqj0hshVaN8MvyNvKQiqI
JnCZV9czuYri4SiIqtFj2CkT3lTCiXBjSac+wR2dhMkpP1SWPg5sUZuiJuVhicazWwYP6XB9gne1
j9lkpQyTLd7r0p7y0gpXKOL2mfyoDuL6vieIjkzpagr5R3O6Hdbf+sQYaylRIdl9Xd1yL89Cjig4
U0+sJ9UWF3/dGLknNfOrlpztR17ky/y7KW8dPH022lYUgY+Lr6Br/ZZ8htbDpCnjkh2W4pCpANfn
rZzMfnlR0+R1myOg8VClRWPa2Iyt8Mhi6Tt8OkkubfhaxpIAJ8IIRhgyiPoZereyssZ44RwMBM8h
Nsi5EsxIVE+PBRSm1XWa5ju12dgmb94qEQSPUUwHt5Zs0cB/VsLdzgaj2gUoqlyg/2SwBG8KVKGh
EgSR7H/28vG8FnipD79bIWTaDBacEYg2Tz4yITV4TcO83WJMztuwoWPZvHqx/pf+zeIxMZi3T6eY
BWgycK0yFo3fvxDhs2/H4hPwkAm6YN4wST/7FLG3Tb6S62Uy3KDa43hmKHfoXFg9NzBq3sKfHRgE
+yAOqSRfHC6CaAWgi1M/aGhhdR5n8+k3OF2G9ujcAmr/bi4FqtU3S9TSQ8ZfkuFIWg3gahrbpV5Q
Dl2OFI2wmXL5Ml7K/I7lBZZjEfDRUvvBKj22fza5uJWLbEy5wT7l/V4GHCEMrpKLdJspzCJYZy7k
abANhy9fUnkApdpIusMOFs+gyCXIiBUeNvaNiEcU/E36DPHhIfhMKvTmr36aBe9u4EZCAEO39w/K
tyohg1xe+Y5fvm2HU/7yLWf0IpzZ7CESvmOUT8yrR0bXs3RCSTa8fcgz3k9yE+fYl0vMtGCPlESO
uzOA/h0/mCKncVzkROnu9lYBXpghMMOvocDnc3pxje7ewYXOvLHvoY7eA61ssACxF0wwkpTSFu5f
Uwl6eNhRoYkLrmP8VIkfEiOueT68AMwcszAMT07YvJI+3U2sWVUYhjg0ci5/u4tzNk1bl8OM6bcW
QLyPrT5j0NFy1xdxIH2FHxVZf+YWqxtq2uLH2562LwdJbN9hTVf4BBVedsCm+nZqoQYqIdLWNkRP
MSm55bS+/T+oPtNGJ4aqwfibfSGleP0dcl25Zp0bdq5iJHOKoU4WnPFN1I5KmkuYbwMCORB32Js8
t2/ztBELXb3qDn8ZYbScFbOL1SUpGNm/RoGNbHiAVjWtiW+bXwmbtS4if5Qi5R1UpeQF9sjcMGbP
ugH4Qz4J+JGD87eXXWxIfqflQczeEBqHlknR5jpQj37iaAkT6O+tvcVzWVnMICzRnATvg3NBuOQW
XczMpJrvhIxymJY1fVmxLJqyjGKqc7KkMfl499Cn6FpvyBf0dVJujl0AVjy9+ULCJ01vvJTpCbf0
UslGFo/r709175M8oIaUXGdgZWe76Xz+kGAZuT1ePnDf1MakqT2fwrNM87NDMIipL9LEmbtNcpmM
YzTgNMofk9zZqY11C1ZeeEzoSR0gxDU6yM9ftDQHhVtiw3Dgw0NofRJ7sIvJTGMH6A8brp/uMNMh
bQpb665MPzKpznPoTIQQ4Uo4PZvoNn+WfCTAJJ28oGUGfvXsK2uaoZzhFIuJbkkKBo3TNotYm7NV
Sej0aQLMnqFuWMTC4bm+BuLs31/G5/PVEjh3bkNCzdI42CW66iQzFxcSoDoZqHY8eLWBTM8CuIry
JsBb8ennzDptOL+CGWvdLoq9S9zgEkGrMDjfBgRm4F8PJn69Rn/fIsBLWZkipclyyGuWElxMz6eK
LUnsYjH7Ct3IVUyc8aAiTrDNNCe7BBgrjdfoBxjZluTa0hYhFJDCGzAG81flIko1fWBTqJOhMwe/
o4wWlrXzlLI4Q8wAaDCLJWf1GZhdCQqHbJdqZdoTWhhkaxBW4j61noMX8w9nEoLNXgE3BdMftreU
dxb9JU0IKOtW5FFj50UsE2Ufjeu8Hu21oGlKV2NjwFFF+i+P2IxM9CAM3r3JephZ5AxQznrl51tt
EkUzTIrcGx6cqUxf+5CPf5Mrd5qtBuHuAvRiDqbV/0oQ1d5veicMceGtqzjJYkKJQT+7THbfbvnP
wbTNf4FGx+lLDsgIhL+set5qMff7WdpfBpuN59Al5qH1EhTsYJJ2zcLYsqvhZe6dVgyn+gfnkEGb
hlHsyYJb1whlmaV9Zr+wMLHtUiBWUh77H8sSx7E18qXT6iDgliI96vlM2V5O/3TuWcA3OTPHCXue
mfvoOrUKC2TNfM8ILI/vpdYJRsPpTfvFTyW//uH6lqi8iarYbENtolZMmL2+szD9Cz4N/s0aqNeu
W5Jinum4+EHqy5ZAvnz/E/i5EvsDdSmICEFplLX5cJxf0+ic0VF3dHTkkyBMk0nDe/bjx7ikpcdd
k4gUgD13yudhKuowxtKGbfQD31JaR/cFOOmsy1UnBOxmHshMNZZhx+O96V/J7emjO5Y5iBkooAO8
JwH78WLvKLQl9U3aNttVVY+bEC38OM9nMjEGrfodqUY0cozYbN9kTbtPBOvIMV2j2axAsKyAjGdY
m5QdZdaNxjlRHSfgXPnkibz45e1hTT9oEjac8Uz7QA1L/i2oJ7fKHfgYYmaJdLp3j8QeThAkyurP
ZSOF28IF0bOvCKr9Z30hdtsdNba9GQjxyokcFOQk1g0r7OQO6yo3bAxZfWcVCedhKgU1+lB/6ED5
VS5a5ID1IGHiDbbK7/HhIQL1YnyYXWoJ7WIxcEfYCSe25JHvOSYUzc+ihD09lWVLi1B+jP4hgo0E
eZeIsEir0nHdd45aERzcErYdUYaGVusmti2ZSG/Ped4cuhTglfHMbu9W46xZsn/0xTRuuVb72Rst
YxrGcZvLZ+aeQx4woClec4hZjJbwUWmOUWFdAZrRWcmcw4Jf01d0TcVLs7khItjBXdYQb5dHPmV7
vzlzTZ1+yUcHs7WKwLaZBzIfVk16D3VE8LfoCy+BblLFpiZtqDicVZpKQJNGPhzw+jZOJEPSXv7l
ipbxafQ0+a6gN2t7I0jeHC56GTUndVVE/MzkhV9UEzCGxXx3TASU3Mbs9qNXLgdeI2b5IxOCrRYs
msadGjwjX2gu4h6Red0e/ziqb+PDZJO95Lz/XrF2sVpiVYwhdZQxwNopgf0qUScXh4k6rkOZqjLu
UgF4gjl+QQ+4bHvYlgieYXCtmw6rPsS+XalDbY9hVZ4cwpt42ag86UlafVLU+QIFoBn/LCHJQ3rq
RJMpP95glVnwWS4XCU4sM7TmC4a9vl0+4ffk30X0lO2/4K33Jsp3nTJonDlwvyevUweUZqtbansd
NS48VnjvVlGGsjeWJvKqAgZf5HpLmLJ237Lbi17GeYa4KCl3clVOJr6DwnV5LmqGCobAYhHc6NvJ
YYHlUOsZx6iF25LUv695w1i10F9U+nDBqezCRTJBA0rUk4e3odPjvbNNq6VsEwU10UBKvLfxbJ8K
qFEbTaQ3UtXk35EIcIpA/E/xEyL6aFXmjPsIf5JRu5a9bCaAdQfCGZq59/7+HEVt2QHe6RbvD2p4
43lOsSl9vAZC0YQ0LM/IcByTT3mUTMd95JsI85gmOV52LKuGmmcp/cqaSi9Ep8QEyfQrSqiQKqdp
qSbRGV4fr2MTnM8UUvWNcqZxN6e/2wLfMFL702eNyiI0cZtk0Prl54TjM3/hxqP9rlR+hz50dGzG
rQA+RcO9+q6u9prCP9eUDxZ6jXrgjeP4tAsacIq9srVZ3+r1ZcUX8JJN3CPK9MMxjX6EBIf05ErP
/+v3zKGMuZfybyLQXrDaUmDKyIJdqYZ/VxQP881V2nDn4YhPuHXXminR9sup1WUQVdm7/UusWVJJ
syOO+tCUlwIuiv8oXy8QBtN1V3CfI5L1eAw/5QcPMcAVgJldS7TcxXZUhoXO7EuIW35on4m+GT3o
adxSf8ZSjYafeLksH9yq63HGdIbqqd72qkCV3Z9Vl86O1qIdrX4dXMgV7UQcMFHMhbYXaQdRxnja
gbds0+X6vncrDFRC0z9Xyu69fnUnC13OTFWxSDGCCzST40j8EiU91/hC2mLlh7x1IoQw3gZYkxh7
Xg7amuWOvGiC0NlXPEnQhJa1pXbzNUPCUSlvA2SX95opkZzmVnGsqg2j+krzdjgnVMBdFZHEMoe5
XVN/hUEBt65CJJl/nBI8+iddUmebbUiuXLotyPi03KyRrdqa8GEYiucnPMs6cTb37BEWw9CgPKXF
RU0eTqHquDRmW9Itl+HXD9AkXG4pduOSw6ZKAELPnfTqMw/0rsQeBoaBWbdhwWsEGVfaAWN6S8Co
T319jWt27MjEdp1cHdEGJfSLd9pkZDbi+3HgLvuC6H+Zy5XG1eKTFLaZc3SWdkY1CtA9nTOf24p9
6+Yo4Ttr2h8dxnQCr2SjjLyMd21DOfZ+1A38r0KY3uazW1GRD1mFO6XiaH5l+lZRjkXhiDMnI4dS
WIvbUEA5kS6AqynryZ2/NIoWhLjSnCHDqxSHtGovtCZsoRexscGGt9DKequhrBUwnP0407EWX7Jz
b/9xWBuNQKNW28Y2ovK3lwmhUcv4GorO2ChQzeU90rcZrQCw0irp5IQ0mD063Y1IRMixCg/JipQF
EGAenHo7v0ZcRTlgjrKS4SdTI/qQrBjKI5xTC4446JDXKdeFqTjr7H0RHH70Hh7BhJRt4NMfewK4
aW2x8BZZtmRKItnxnpWlatde2TF3hxnfXzyV0Qh2MoJF2h7yuDTbo7CsOO2CQslyE1NvlNMMZdb0
1AM5oP7vbABub3KAv9pY8lnNObttrURc/GJbonVJEZXR7DXazDn1ojjp5C96UCSX94rc13u3XfbI
hUL6HKFDbd6uTUDFa5QfvLcyPgDaaKAVtviYchgm9E4m0uBxbnqhKxONk+Nqv+ZVl5/HFqhT/zAp
gQz2RM8RYtiB4DRupK6QLwkCKPN/TH0ZhsKboXdyK3I9pXr6E5sYtqm7DgAoQz893Zot/U0jzqrB
vUO9DSzgDSg7q8OC0dF7ITJubG5igFT8cvBkWm+dIoXZ9QesRgmbU+jE/dgbIxhy6q4ZFD8bhnpT
ar/bEWeSo9bDYerzeM7E6vqMV3/fOlsnbZ0Kq5pY49ZP8rsb/tcwepEDVOjz1i/kr2PpvPWHywQP
dreN5vTSRGmMASjX95VKMCAlCoP7YyJNmjfRt+BLmKhqD5a4KPS5DMytdJLY11JUO73yz8zMwjid
3zmdHhk+XC0GZiVjRIxTf+YQ1PD7nc2xMjO/77aTOUoN19/vLPs+uNvr3F16PUN41Av8zNHE6VEO
JRnNnkv2uGLyZnzm9eLJufhakNFrDiNiLZYhWgyzw+RfJ0MtG0GYaT2dDSv3m4xwSojeUNnNjXje
dT3EFZDpY4YAlMbCNqmMWg053sXQYCtJB4Unavu49smua/Y5msKfoN8Q9jcrBSwZUPwNJT2xry2K
6c1JKxOLRhVqVVGf1hwbu34Se5iIO5vn0crUJdz+1hF+ThzvDXNt98uEZassZn+X8M3o8lma6EUw
7m2oMYulzUJWm2K3diqKOT3bPh6AMsomJ2Dqmjnxr/Hv3LaTYgm2e6mM3oKlvXRG0A7ostx/WJwg
vc87Llj57qF5ap12iaLLQ6L/t968JoABxBsCDKcIzUTdpR153S3xGVYWZr5gzGVItmDGcYlLsfh5
PLpQ9FjcwdRaTrzLRQoWWWetlT0iMg7rtXp6xNPrnt15GG5V7JHs+L0UJQ1RU6ODmnYRAvO+KSDg
MWLJRF6VhIDVLUPAlk7Iaibbu8Vu+WdFT4A2NaRmaaVoA2CYC30jwySd3LUpUs+ibYTBPxLQn5l5
aUSRib1yUe89rTgZZC5Pygq45yl0s9X7Ib+3O5K999boMS2xF9Faz3cUX6IAxInCSQ5UliRoS7mR
goZ/aWxcoJ3mZ64nMjvFt0MGr0BtwhdiiGtJIKTdExAZk79EDjC8axKLvKE8p+9FnTA/iapdb1Ef
lwiwCFqsZ25sYjSPN4of/MelaAeGl92y4BfFOVosDAVp3wBN2fWLrFCbmc3B/ENlzSSfYNM5rYUb
kEUCk84gTUyaChX8BzcsebZ0bWh6g6/SmHfoD/5sfhjE5sGJnn4PspZn8BVgL83dPamHZ0xEq5H3
O9ndLA+q6GuDJlSOnROIb/izue/4DzIHJxoRW5NV4EHAMOBwUjzvtX8qwSOeoBQBTuRqeh+d+uGi
x074fQU+Hj9V094gkoqfR2HfiSqMGetPoucFRwdrocXS/H60WHhpMaFtolCjHX7GUjZ2frfelWvY
BPa/IXYryVRujpFrl++dD12/KAuVd8pkdiGhEG/ijuXoAdXAH6wvFkCcO9aikll2MIBHFZ6SE5nA
xz7CNwK3MyVaiIudVOPuAt/4EsXZxtoXX9bRkLQBvnUM8rBBaqMJcpiNw0qMsLXL5wljxTe3od3V
RDw0UkrX4Hs2GlPF6bx+YmyncO2Cgd17p4rA0+iY+Wu9GqxaBcSf9pILJQHelLVPL52YOfEeLj+u
zLUrXWDgOQcktbOX1tQ15XRVTNGsRkKL6+ANwlsrSVlOGoHcUaUw39Lvq8ZvWqIjxJFUYFV8M2gz
oHcX+fWSkNiLxeMrtxKsgpx96kgIxnGM9gOLeeJC2ye0RHMcvENxUBx8mzvB3uk3dj9rg+mnUk/6
PXWcMA5Sp7sOIT2czD/h9OdWLTuFFsY6yKhjKF2kDuy2j7DPinGgjs4eSmInf3cnsZRqjjoY0Y9C
/Gf/U8H4J9T8e90TuwIAHCmOYL75UvRAs2L1rUtikgfSsgEEBKdszRwD2UUu1wH6EAWHePaQNiG1
z8L7NSlHC8r8EjUlzLrHF+G64R+dfhx7q7XH+S2UEO5wI9oEM7gIBD70ejcePx68Vx1ldO6JcBnb
xitVvd+titij2BAIh15gJMhZmjVTxDhCd7c45csskbMKded32jh4n+psCYMVmB3prTKxyFKB5zjl
m8sGMEVELeu+sGYQqb3uaUrcjHndfqIAlVIbFLct2C65nDXZ3J2GDubLi8OmIBZjBmP4XcUbFi2g
Q/6RvNZKpPLm/6qYct+92awTnP/SdTQOsPJLAJ1aC4k1EeDlKIuxKmVSu4DkEckMmisBG4HrKydQ
SoLjtUqDV0LC5PAwyRb9ZrhpMVUkgW/UTsWRTY+kK2Iam4dIZ9R0VxAbbIzKKOr2zXX7WGXhElJr
yrOuRC5Xei6NZOsAXdeqJ88ezgQCqKjHf1/BeMqOfgfNa1Q7RaI9pA1xRc1CnYXwjgCLRFqVRvdd
TqsKCEGR02n37jRenaksg1OdKYaqx6nuZttpe8EuHqlA2uXxlYzY2XO0QbI3Dsvht+DDc6nuxaI8
hMvJmC8+NS97Xb4esUj+z07MM1hcEooegE5k4C/ggT/ae3D5uXFWPV1/Wa9koo+r6VE4c8uqr0wC
HtlEK0PJ4sSu/aZP+icfAqYY7EJi5S9bGoBtqqFhRuJnoTD7hTcpaTCJcuS+dXPRgAHv3FG993Vh
Bhj3OQx1okKYDjEYCCIWQUrG2lBMtbq+3QvahOFq8TSjp0jbEVd1zHHPqrURij16hJAlgF1MFdBJ
qyyJv/K1mRRFN+IYazQ8nSU8Pf6a52Jyg+cNp3lIs/lIZ6RrdOLZ8WvSBQSlxzZn8dk7wSMfa6yY
b+JHpCyd/pXHQPPct44WChRVbK+W6Uz6DYaY2SuiGOgFuLeW2dsaabEw/o4NyJVN8e6FhtqvI57x
SRuNEEHYB9wNJIXi+s3LvFoYTiavEXcJOqvYH/nw/SuJ5U363NoZSFoWLTrMbrQjdR5LoP57Gl5/
BP+bbJpUMsrVF4vlF1KUy65SIDSiAY/2vPlIag7FAfaho9rrt8SExUIn+OZWLqef40SpdNib5ix8
XKo2j4ocPXuW0tykaIgvAtqgX9kGAEXrxkZlxZKRMp0yiS4H2d7YZZMPMfFv6Df6emrxWh7MneYq
m7vXXVOM5UYDPynuc3HPDhlUbjEK/tXZJgu3yXSdOH3u3xkd1S56vc4Vd49p8WIUfYQQ1NWCE/PS
aeZK80X8gKBDC0QM1BfrvDY0cvvqrNjKxfGx7Y+E5gtDhRoIqBv1LnMZzYUKE9fTwo7Yy43pvf88
3mamCB9AKG6yc4fGAqnmp/wg01hjLtLuYT3gDBZA7gxoYI4yZjzgN4Sk6MMeqmv40QuxzRTx6KMr
CJ3QBD03XD7C4MqyRks6dtOeypHwGnSh2dSuUxyMTZtjr98ZNVfeAOGICjedSFQty58VwMipK5lR
nUttr0oxhWMN4UTKedWnrl+jik0ZymaDSj5RSsXASuM2m3T3yy4ekk1FUxv5j3/eQsUGILECIZz4
Xj2LrqalSlXq/ezdhOUVRqkjXSCK1cc1YVfd5+eP0bYmJn3tofGUtaGI4VBuobvmUQWO/k0pMiea
B42gUK4iBAWuaZL813XSx8RXAH92TQjTRXafMgLuLFImVZ55a3MH8DgdAM8PSEShVhBOWIBvw2za
QO2JBs48dn+y/DIf+9iRvt7EDy2oht27sR2Hoa6taY6LuR98FNWoseGHT8sM/pGzQTbK4M6h4ph/
ObhcEvicSDkQoL8LS3CAcE4XN+HUPKsx3bPhnnr6z+ifrQm/09VkdziYeFbss8my2yBqJmcexHGp
DmI9hYsnIrHtp5qV0/mKzKyeRCCoa+whjKJBQRJj5f2KNOZH8cF6RSRTiqi17GiXIfdKiJcY85o7
uUY5pAga7JH1C+oiS8rqvGc4fng+2OMQVdMFJYwmOg0R4xbveeDcGC6CuFj5tbrBcEeTRrk8BRtw
j5dAtQRSNC5OJD1phfuJUH8cPiwCnP8amaUXlRMiTiAV5gBhK0QG8QWhOmki0ZkNRJT/pw7zJmKr
iZeU/t0SQMUCcAR8lrMsZNbO8LWu9Ns/XsD//aUWV4ivtNJ5CaRJglCBAl3AgbNVi1SwO7biSnOx
CygMmIlTqT8fc9+axT+lQ7eg/zE/3E+Lh9h5Kjr7kf99Nxv2nu6qHliDI+SzVih4kUqaCmDYWOVr
wNKLnTg3tQiJNL9VOmZhGtHwENiTRGgcG1yoDmIHKtV3FDHsE8cahWy5o6/AuGQVaAw0m+2ceGxt
RVUVpmGO0Qm2GSBZ+VkezAAc42c/d3XT8vKZBVwLuVtqbgFEsoDiS07tWZQ0JNfIs2yLOj71oCRd
5GlxUD6kFrhq1Quhga1/dElfR/JRBUbMLTBeYg7jgdUv9QK+tC41RaA58L/Aoc0HEwEGrHpfcHrg
6MySvzBgrBlmvfod0aJ3Zse8kdLmjaiL7wzTwnF4+4Dd60aQYgdypiaqRHMLjk17+XSVqKTOxcf2
YV713+fkvprqobmud4cisv+Qb73fkOYPccyTr6ejSC/AZ54a11zWc0RxErxQrjrb1aekqMJ8qg/B
oP7AER5k13o2GfWZzUbt9LO4QM5SguVZ3L9OnrV1el7yhkWWdHqKMWTSK4vZMxObtUnYoddeEVRs
opczczq8qFAQOrVc1NOduawiQrp8a2LaQR1cYG60yXmgidqlDA+lhetdH+52Zu/Wah1XzCv4BFBH
SewxGm2Us4tql4iFEePscVpEKQn5NeemSYVYQEcSr1ixEU0Hq4wj2tWqsl2Qdd8bYUStV/GfROjj
/GcvAYQCfFLsCJkL5YD/7yEMVPL1ta4hmAik8wHlpxwCge+RjUePJ37YhAmnD9knp46EjRPcAmeO
T40XPKluIXkMBQ02PnMhEvyyrVON6UfC6HQ1qdI9IIVLSI1cmkcaoxWpSnlyCZYDvOJ0l17K98z8
Pnx5UhNrIu1HI7g58AnbfrDC/XmMGR1Om+fiP4k3K/M+zCiL+n9KDnvEE2AqJ2ccJ7ch1yc28YM6
xMw0YeO/DaNMohC1W67w2reKL2JWyQ7Ue6SmxhJqeLplmxSOXQAVK/Sbruk2TFmpE7Exugzy4z+J
MnNToMtmlGYcYaCLgWNfS02yRNxIfQ44nc3TShhNkNuybmFdacH9uyt5AuxJS/9vw7uKARmLOaGE
jDVoltvObJgObm57SX8Dv6I/MROtcNHMz0CG1JKLgiRL3lKAAb5Zzr645soxkPsOhgn4RCGaJQcW
vAAhf2QbuW5RRH5qGtE1DAhoM4aN91icyhK3lcqoI5xkmT62yr8RX1RSL0z99nq+cxxpbOkZvivp
o8FxNEawndgFiYzYo44RqwLRnFRNZWAOvGB5CPTrpGOB7fEpyq9XK1JuWzwj4yf0UbPJ+8OLpe4x
iZSptz+0yZWKeCIskmPzShLgrrgJebvLQ3m0P8UALdRi9qPLD/Sw+1MWXKZD/KRZC/mlrCC/71b1
BGJighAE+2w6398h3+ZW1j8AZ8mUALbLqnyB+fNzOCNUAmznboagtu4hI0O/1UlZbp9Ow8rtKMN5
0DGnYwsQQ9SVFmGjyRXWlq92A44+kP+zmO5kUUJXqn0n6sgwBjyTpv81LRAf4DBDo+vo3Gs7w+zL
tKSZMolz0XTtGHB94KQTHhC5f+COdeYt5F7XHapk2NuqUGknjjMLL3gT52OR4oUZSG3pxm0wbJ0M
ZohbdxhIbp/dpRE4bwLoINmgIBU2hGZtxRPCDEoxoHKGck5Fl1VfRQ6/YPIRPeDEzJktI1udKCgo
moNft9qb98SuL+rg+h/oOhaAvL3PvZbJQeRXlTq1UW/9Ev3k0CeQMWiUtPmAfTQVYYPXl7qjkPfc
DLiqiDlVAYXXln/6lIxj1Oct/3DUwAYclwtcB1j8Wb3vAidyXz1ll00HG4aRSS3dpFbFOsbryUoS
oONupF7H3h//kfWTx0pT3rxYyn5lPBbh2xCQeQHScEjVgP060Cv/HsxLUUfTwIHfea+MSiy4kHnB
bYDPIieXElyTTgJ2oTixpkl6RVCPUFOqwf8rPebugnNUxHuZVgbLCB/Jr43xqy0EDghQThaHBEYB
k/hwf519t28PQ1w2oUOmpBhUAm9NP7PW/SmTfGVREb1KyfmBT/lpNzYXMQyK5iehZ//rHV83KCLY
A45/qqdyzGXPEB+lF4DqR2geGWXzn2qtnjLk/2+Ng32hNT4gG+oLIspC143GQTdZH02L63YKMzx0
si4k4GRIVz7nR7+zote55HDDeBZhEiGTn7xgA8DNQeOIRohr30EAlDm6mAEYwnC7rX5LutZHQJZ6
byb+m5CE55cpwxrowbcg8nqxoBsxBLJ5btZneMn8vFN0i2lYt5BmvIEpa648quYEKOaYqQlBkFWU
hFdGblPZwM+Pl8ko4skgO3HZkfAtc2geZMepL1z1Fj3dep0u/ILgP0ilxYGkadZah+kAdus1RWPH
VXKhEyVFnasvAcIHpkiDMjBT8DNx2VFxYzQ8MyDcLgxvihcn4/P4fRwEJR2BBaZ+iF5xqGqvd8uW
eJge3/RdKonS0aiWFvloVmD7qSVPDvzYfKls7bmTL8Ca/uVxNyZms2p02YT9E/l59of892UGlkdT
tfLK47UM1i6LnqwOsCzf+LkLoCD2NH0O2uc4pT4kvv8/Sa3wsu+c2ZdAWU1DA1hmYhJQgrA3Vtho
9EsrNK9oLjvCxaOmn+pzsWLiKxpR6g8VmgjsWIUzhLJEJgX43rxuQdGwP6ZkhkFT3c+Lh61PYBCS
iumC0RLStThABklHiB/JY/Ng5modKB+jH5Oo/2yMhbVCF31eJXUARip2II92+eXJfVThciGqB0uI
LO2RV5dd5VdcGsaWy0LByZvU1pWEiV8Hmy+Agdk7EPJtJWBEZd9r2RBUtzAPhdFJBUEM0DI5WWnG
NMXaOYDsU8H/1FKmsd3mkJwk2DJ2M11a1rtda7F3pTIucGWE4F/U8RaLX5GqwPsipUTDseVEjmCQ
9m1Uc2G6HKmM8SYlHAnJqKZ0Ak8gUQB6ZCtZIVOT0nRRzgiN0am0lHPgryq29nSST3N7+xuuO12L
15sJbkTS7K4Zr7dO3Dq14tbb+Om4qRbGy3pzDKSetiZpFwjkomjU9JSli882CvpYs0msTNUNtjo3
k2UCnUJSU90ft04O6ihinj2XsZO4JbOkdGjk6qUUddjhg05ekvtb2vP3dR8pDkhqi3+1hEaC33DS
78BRdb0Ci7GYOihd1lr8oYHqxe5tPyZ5WXmvm4AKkB0mPFbHBXq/6KI2VAONaWOn2h+y3hpYoPyz
r5EeswLO/wlVmN4hCk68tAy3v0Ko2g00/3LNDg4ykmDJVRme/Tp7oRUzXjy2CEg3y5dNApT5jhRT
y7+r9nkqrH3fsdmgcr/uf8B6Q/ksIxPdhvqr6MaUDOI0vBtuaAQLrZ824kiaSfj4ildySXV24RUq
8zbaKbFmyEYyGWPxeaulWoHh816qQQzI7KCqflHBNBjvSozzNvvRqj9R5nxWdzVnLa1WxN0/zF6k
bfn7c+BbWDxf75i2EZz6slEJSylm/19Zab6ETogf9P3fwZSTKoPilwtoQrmo2Hj7UuUAec2MDo9X
4iLUcgXpm1g56isY8hTAJklDWC5JIgyqRW8Mk9e7BRJIZNN2k5fGNxLSlOmSOmowgsbq68JEs1IT
4Jf2UYOJ1GxCMXZgL03fBtQEnPhhOYkSfvJmP2zXEyZw/QDWk9gc3EfSTxLNEYfVk6lXR76biaJs
bbjMiRoug3tBW0um3A4e4QlY5esJ1HlHb3E6x/pJ61FWnYntLm/fUzHZiigMqoG324nkZqCZXl/E
RYwd1s8IVcVOBgg4/54CJdzZ/PwwZII8R9bvEZz3o0EX5dA4zS0ZJ0I1ovO4i4q8URvTw6lghJMV
cWccObOcfWf6CBHFKTwPi6unsT3yEpZ0mjjh/1Lye0TUBecsDtsXAy6JlGeyLZ5086S8olLFVi5L
vLmqlZLzy9idNM8aNb1vMMjXd3kx+4fd+9rSddzZkvgEEdcZZ1CeBdDHdCix8EN4k9oOEy73a5VZ
E4A9wS6+CDQzLNFSnDuD8dkrqjPok6lgHXh9oc+tsQAbkFFUuH7XDR+3Dg73iSkviEUqxOqzXpCS
iFm6jsYyNvXUavfiNrkDmzMFjCzKriIhzmL972qIk1qKJvZiPMSugKe0QWvzI893ZuuG6eY0D0gK
+0IsR5Q4t+v1j8foZV8QtWPbMJvkqkUEOESicUpX20OOIHsRUeS61UswSI2O95oI86ALHm5rXoEW
jEiSNDl5Liu0JE7zRK6UbQjnGeF2kHrYpLGszxT8gmYSbN7wZGvojizH/Xk5En41sDXiYfOCOWVJ
bcuG2UF10p3gb5dk3FKeWv8f6CHnIoltWVcON4SeICDY8UB5p3yBWkH06E6huPQG5eEWrMkBU/gl
9A/mbN4WVpd3AnXwX6+SnBjhFWhuSaLGxXgjCEYkEQdp77ZO7Z81d7i9QT/LibEHPtvSl5jNMZf+
SiW5LovWknI+c0Vl2/hORCkvinYoM5Zd0cBSC775KQyqR72xt3INPuA5u4ycQeP9wE/8xuzDA4AJ
bHLNZIHMxGTGPgxfr9h7ySeevIZOhwdUuxaIvGyMhG+fVXxQjnau0Wy4bO7DrEMCh/dU5QainB5f
o0qVMrdU0ElMaUTrRx4qCE81RMW7o67bd27FZZulfwgb0vmHS6ihkrsRFq8WQsogzLz3GwPUygV2
Pwwflx5uYyKUmZhST2LFhpLrFYhQvdq+6+OkhM3U3AP4k9kakE+yqJcl/jbxMZizYwTEZOn8Pb2F
avr5qQSROCXEcNnT9LOHNr2kKidWf1t07uRWzU0pe4Vxt7yIQcQnMV7EqK4isN/XuF1nVIOek/hs
603bKcDfPKxrFlLSRYeUtWw2PUMQOj+HFzlbFq2WNiYQ1ijwXvsBUsr3MNsRcMlIqUtT6yYwyqcC
/BtVc1o43e4/okHvsMLS0J4KLY8Tog+VhYeULq/ZQReb5UiC8S0YpaSMlBBeJSvD+yQesrWDIv1S
IyNMTpjgbbpWFdN7jhSHLJ12HP+Qrey9kNpNJOJ5TiRakbxbaQD2V/peyvKcZFViiYsLLOib3Ed2
MlyohzH12YX+6jLYf2Q5Cv77kAemkfut/QsNGJyvILRa3fR1ok2VCSD1N8qkjZoY+8P2reUnaVBD
jdsxOUpP6yQigOcEndw+MnLAlldFwL1Faf/CGlLO0jxHB2Zqlj3fD3wYtEZMVT4tqznUp20HzRu0
2Ag5yB5YmWkjsuR7FOjCGBNfQsMvgmhbgqNOHAnb0hh2gh8MrYOodXY94lXjvr0XJKWzMYaOjJAV
X7AN8QnAA43OyA2AopdSXmoDxXN06dfBJvL7L5y8cbjjXSTElLdykh9ELHHqKM3xM6ZugtGZ2xy6
37OTypaU1c5O9lEV53cSpn89Nnig3tTTJ4d3YLxSsZzaHi55WdQ8JE+6L3PXKqyVsYnzOOKptDQP
bm6mPy6YslvliCWCrq6xbyOJX0atPNv7yRcsuxBON6lmBW+j59rCCLOW+W/uEk5IVr+d2c8jSgyA
282Wexrd6GN4GhJ9INscd4J7vS60k399id1NNYK9ZIKyHj67k6lgPQPNU8LzL9PeUb/axwRgTyBy
lxMuZ9fRiGH8oASBxg9QOwQVpzo87bVDf8gmR11WfaDS6NDN4bw8yRYxKfarsGzTV9vF0qCNbyiR
7+yRSRoqtaTmWohwXpNEe/Vw4/2GYebgiAYeocuXErxlgKlbMlcMsMIGi/UMuGGt48qywDJ4ZSDO
A4fJNsFClT4d2wwix2IPSBkONOv+w17bWdAE4Gt5HObQXkhSfGRRJzwuH4hdmLhkihFq/oqMIMME
QNcfwfDdGGgNat//dgKq6n4B+xfTQvXoQz1B94fig5FFgBoaKFtOcYzyezN2GUYhE6NYpjsBWGFA
N/sL1GPl0aqeqwM8FQc8JN2NSrwhJZ9iSszqfra/VUjU0XIXaV3oKKcymS7dMoVuvHl/EwgfyVOm
GrakxtObkGWgqKHeOCJFlJYWbixO9mDL/juxeY4YOJocdaHtyMF87k2KBuGT8B7QR1IbfaDKIfkg
R5fVg7uANhCN17nc/1Bk00UPrqUmBe7sN++MK+hF0NO6vI8H16sZk0Pk1ACchul+ryRAyWJAA+7i
KBAl3FmDM4yPicV2dTBXd2nklTjp0YJjKNDigINzXcd+qqC/UchfzWOrPy+lqXTf6GwDZQ5a9TWb
jfQRD6FNc+Rv+M1pPhKNEEYauO3rXam0mGm6/sKIOWmfZIZ6n7bUAqmayBjiF9oLxJbWIgDyNKBz
crOn4gZwaTcvDmpbNToOVDCe585SJ3qKgpziUu1nJIa1Ls/Q6Jd+k6+AlZLwCccUq6670THfJCTb
300S7LRysN96SOa6HN+DU+nEl1/VaEIo8LkEsMdlDeoUaNfuX1/9zhoAPO4nN1SSQFU2I7/krO0m
Xt0vU6NJpUlnfc+cnlk1KwqPgSLqg7JYAYlGd9oTrse6g9ZpsuWXhNStb9fGnN+hMhCiE+FHaBy2
zu2GC0BMhcSemC1nTdn7bJ1Dy8TXtpx9C/yB23ehRANwoY4AgOhLQZuHiM5G85lHg5lnuiTnvVAK
oprlNiv2puGpMwqm0cjz+AFSGhr38AfrT7w7ci07PK3/NFaAtD3yPvUl1DLF3OcdSc9f4VZJxTru
I5SQC9vaORVmznZNDxThtT8912AKDZOIOelgkQoU5qvmMDtG5lkT9ak4cYbzrMOdo6XzGKNmt5Gl
XQN5sWM4z/ZcZR2uwjI/gLpVbNnbIhILsAEKav00fkvJVhg8OXotNqgDVk7xA8JOIT0eaXle0MuH
rUeDNOUucWoh0kmRDjmKtW0o8TgMUCBMFrY9CfIvScDCTSf1mGt6IlpCrltkRjQfCLxewxg5adlY
gN6T85h4QRoE3Ss6FI3CT+jXccJab8Y9WivPCNz7iGXRbShALa6VD5IxA6Msy+gQzz9zjQsPkXZe
PqZDiS0NqW3rhshkyiBvctn5U/b6BASlLbKPbE5kD1Swc49B4Cqa+jUUlrM1owQW3lxeiWrOwtHR
iRsYsnS8NzEtkwXF4wJczUqf+fD1Y38j6+zenc3dLC0EftTfhyQPddMVAHxyZrIx3dhS9HgP4BV8
GTJ6C33ii2z1gqQzZjWr24c2GEb6jglThD9Ther513im5VzQ0Pf07qrJFQqxGgAhHWYEHW7FHRMv
bgHZR4lt53+MnKPvFsrJLVlH+pPm8XqcrPAR3qWFUecoijzlRUMWoF7EykDcUAmSg8rmEgsjfpzh
pNDEy82Nyaw6V2sebm7Lzf4ELI7AYQHhKe7dyChZhc8MyOMcKGcv9/FUENuB19pVIaPbtOikbZby
7LCYpQb1QWKzrQkA16BioDUdnwHbYQErtIWCO4713GjWFQEV5exuKIYvbC0+6i647qtxh/JaxxG3
Tw1Vwt8uiVnpzRQkZn+JWZJrSxSeEmcVoD81dqd/wCOyUoP+pKuHLbHTr+eTtg6kduf/CpsuzxvM
Na9D5LAuFiJV+sEsLu7EhoEBwJmuSMQEoYY69VpySf8f7LOZHaiuknm1bfMLGgtBXsp5ILVxYtvQ
Oqj9iKGQ3A4nTzMZRf45SIS+MgLAua4IkPpn10/vLpxcOt3ukMLoltOPaCQTnDbNLrdoqb4wfFti
eyeVpVWaRESHi9JEywxkmMI7iALevpbWQuzThVtBVTmQaUv8WtiI3L+i24i4JXnsQhsDCtHfG/XV
cun76f8wDOvLxRyVRskyeCrPZbO6X9wU8/6l+Fcz9UPjwnrX1fV6Ev3DUdGYVnoNcON11qo2QHZy
Q6pyFF5G6jXPrlVEb4XrxJ6lk2zvsn35M8iA+x3KPRnb9vYsHd8ebvVOjenZFZEA784CxoB1SZQM
RRer0iSeMH95Hn6UqEd9u3PeqwFfRYKQcti8u0v4XDPb+kEN4i8erEfpfK2a6y856f/0AMdeK0iA
hH1AsADrX30eTs6kThYjvAHcRQl4/sPHBnt5uFTzbCn6f0t5vg0rDuTc6mCC72oqLMEazKlaGRbD
MEZ076GFD8XBqCcfloLtIK7j8eLYqz7vF1+UuRtF5azuHi6PbEtdefeZvHY1cn+XD+OTZvafmedQ
SW3NjRr/uLGn2WIlvLLSuZTnTM98SVJp4xethcSQ2/Z2aEtiKkJGIjoxdxOXs39n5IU73upYD5KN
YmhMKHFU8BpPEBcTzkx+ZL1TzzEjlYi3Lj0GxvUmbGKvzm527qObXkItWFQkjc43MfMTt1GobygA
2eUvHa5G9F16JAaAqQ+tpks03F2D9s+meV9v0E2bPqsRpiZ9ryQMIvw4D6dLKcHGqn1gz7cvnMKJ
HPddOULUs/W5Xt5W0J+2y48stHtINIyhnYweXEb5DQ+QtjiHNvtX9cW2NyiO9TGI73ONKYqYOrqZ
TTeV6sw8XC4+UgNcmQUYxVfQ3Dl+gb0IhfwC9vtluFC52LzXweWYeqt+DkHPI7YWpgmPHQpcHm17
eFA8JqTFKAuEQPftIZkFNmsjUFUttoUk4OX/phIHiQ/QalVuuMoQ0RFG/RSIGAa5IOO37jFq8Ksy
rtMZqZbOhcIb7MknUtD7Yeqaf6vuvSYsQTqBLII5k5OC4tCz0fmZBcJ61ASHhieDSyOzwtbqxlFu
2hvreI2y18N5sn3yr1CP5we65nAfd1CmnjSzmtrSzTf/zTOIlnthM33v57EUih741oT21Y1NSkQR
jezBoJpNdZJOqSpnFIKDG7mUDR9mmIdKIKkKIBVqY3kfwAzYhUMsfB+zKvipWKD6GVAt2VroaCn8
fcWC/o8cRqRGt0zxGO1DvfUNljUcNozgEkMKvX0ZHIdpna4/lsANkVL9dNFJaYxMxMfSQCHB1ElA
8N0hpYBJOxaigxARXAlX+ar+jeQ1zW4ggAVQ0CN1PyqIC/bZXFho1CJmg+RCcUFrgyCUdnHb8773
LbEBu0EWIFjnuwErX5T+0n3wG4zDtd9wDCfQVJT2LI+s6S283TgyORce4fbTHgKuiZj/bM+xWXle
yOb0gk8U3Ko2ahnMSdV7vKxBgNPKtmTl+7oy8MGQTXAH1hR6fdRL1LuuQgI8Q0zZrS0HvK+DBXGW
5VQW/15wKusAqL+TNn1zr2hOYo14hWiR9yx/jmyMPO3FP9gthacphZEeWWkzfHCGr+UOaJko2drc
8wBgsrsTl2+61R0y7ALnEdar5kAvxZewHz7Aeur06tIHAUD+1OVEItsX7Y9+UCtZzx5BQQldXS4W
XuAhQMfivf8QE05Xqsg2WbGCnqQOtJvUsIXaEdSkWogj9BrMDCsIQJ5tr1cCOSG2gRGhPVGtvUrR
MJwGATsazEz/GHZQ+ubZMMMFRXrUppJEcc5WtylaKSLqJVhxnBd3Fngn87fzDAhg9xnfgp2PI5O2
aeMn2vB3PXEI2OA4GofZeH2e4dypHCQ/NMQ28lTXjfzX5ghALURNoMTOpxOZWP3vOKnMZRg4SU1q
Poo3wgPL1C37H2Pi6xLRoOfp+XUBpESQZgWXoQcykn/bqRUrIWof1uab50rhSLUs37yRvjOFESP3
ZDd57eeI2vkUAWDbXbb+/130P5njU3cpS3D94QldXYJj6KbMUIjnWfptbvqKDaN+qNWEW6NOBPtZ
0YeLVmADK7PvRrszfrM92lvwogYj6YpSR8s2j5WwgiFCz5X0IdV0dh8HIdGnDzABlSlKB1e6rLvA
06/UIzrgwePx5hJ/FULPoubqT/xAYjmLHxHhepJfMygJB+VfUEDmMpX6r+8J7zJQhuwoXla9fzNu
Ygil5yqgy3XKblQOeX6goP0YcuZd45Ooh4/9wBhzPZ6wcQpWlxP5VnW56iKUI8AG0q+VpQmKDi5K
Ga+nILuWFRBFl949GJ/yX2s+tGnQSKOj29WKIyFpWmbimhGvNy0xNRzrnHtO9CJihLzybBbydDNV
HGGEXCx/d+VSWmxKe8YfrfpGD6GBmCWsPqY3x3s9e/cO4etwBQq01W2iP32cG64B97epikKdGvy8
Zo4YG1SWm43mbXfIjPVw/G1MAPC2FS3vCUJqGV9UtyHCTdqZOarLUaA60vW5u/MKZibuds/Qwual
ZzBFn3qO8zVfuxQhKTT8rkynx2ZxXZoLXhrXaALTC8X6DBDSYCXA7tRgrSnbgQLY+P+UafpwbbI/
OdymNl8nDyJjCzkQrhukXcFF7M1+voeGcll7SK2qBCUIjPUHZX8jM1P+V9iUYxrENVV8J/EUPhXy
ctdV4JIg2IvI7d1xXDoMuGAfTT8A+/ImARXiCd7G7iWdxZeM9NVUyRV+DLaJYsyoIZrj1Stx+0HV
9/kGQ7FvS9kykvl0kcdzPG958uCNopgu65ZLrTK0e7LF0C4AJGWucgdp56whze58FartzqEXPXFB
w4KpzHFYDeuaN6yeG8RvQ2P67VgLGsg4EpypP3nFN6onj6Z8P2qMGX1Idwq0gfU6QhJcgRT6RU0d
OH7AAyiG7McEXwMLZ536kvr6XUed1kNG4BN6wuHkNNYJQz4r8c3y615Tme92XA6FWfts/qlOMKJo
CidHdjWkDGSe+5HTdadmdJhbX/pkRx7g8w6YAhjCyf03XsyIRE7Z0NqKxH/RzCGdXkBlbJdBE2uL
/pXe1J717zBjvAqciROryPcNrRIP0j2HIac7BQxFmgVlN/YShnzaCDRIWfTHCx9xkT2H727dZxfC
8wmKncEh+WI1nB4PHBQ9PMOmOEIDbwo+1QBMSSniWcCmbzr65QR7ySAVyiycTWfA8jiT9VLCaUy9
vqYdZ0eoi96cl7fn1gk6H5+jLHrNPlvu3yS702QpQx3GIQWNcmZeprl2sv0NHxz+ojcuCGt6G9fv
ufunwMWg2JawYyrvrZ0dP0PLzeERlRcQxNf/ak1HKW6+Djbnb8c/LEdNd5pfALpu/at71SbQ3lXa
nW72YRzVaUhte2MXia/A4Qrz8LMw8wlx3fysxsnZf6FuRcBkO1hM6eO8cfVYT9qp2S9rbQ86DsV4
jFwjyv/FcNmS/d3qoPEgew9Pl+0+pFf7iK/zDaDuPRJJZ44A4stZHDX+Gt3aiF5hFGU6h2TpAYOh
cpqtYj6aUDSnVxmqMFH3dL6pqhsKYvyJZ14Mrby2sH0kTeXAK37kbbLRul5OEJvTf/cnZ7T//ILo
Hlx/zT7xtwrViorvtvwuAY3ZBamB12AVAqJwW1/ew3qqVXn/Pp5NBFKO5va2MOcl5aSb1pGz+4+R
5/08dZvo8e9lsmLpRtVFR83fJaUQOHZiDPmf3f+DZ6PgPiKZfHPp6IrqiZ+zZmUL3WT26yFcQSNX
Di/aV0aazgOTRg7t9CSggQtjfbsUMFo+47d3A4OVkMvxxHEwa/mENLkFtfk6UGaWn6VIF5J9YXrR
YFOXVw4TVMSUi/W2rzzz8+vj2fdjo6II+0vHWuj7RqF7zJXZcVdji4wGy/7kb91IAQcEnPoQZXbw
2/iS37RJtsc1hajQqBKUvAlLHRgo4+JCDuZr92WFtUDJwYzf6olYadfTW4I6elbeP6Pecm7b3G9C
37ulH+f+62n1yVJZfLwK+XC5pZsnXuBE01065Ms+AF96sHvZxe8HGXXWcNCFAlSMmD8wcxyC5D/f
wwhFZ2gryhmKEOpHrawjqu9yPw4Tc0ChG+lEai/lSzRD6aMQ77nwMk1QV2MSwi5VXI4gJfk3dmaZ
RoYjemPvDbkHBUjKeSqMwnLEqz+NXGFJkQqml5h6sRaqUen9IQsOgJpLcScats/WAVaKKSXRhMm1
gTxSn+CPdKsTghj7mfv6fgpdE2UEcTsBf2qM7Tf6/6LZrNIgavS35087RxDZcp5VdxSJj5BfR5cm
ykntrfL8uTEl3bN+N/kxAmKIyFDcLPjinLty/K74oGXbdC9+FNLoZvOui83/R6l33pjzo8qvISDx
LIXrE86FzYa5fzg8XPKxgkMCgAU6yoVdX7CH5ln0+8NhsOgqZuQCXT0/J08LyYup++Q1uYUOxS15
CPlFFxKNdAOXW6RIxRaNxoIFRl5tDF/82XyuqbVWDpkTRCTZHbf7gHlRv194hsbp2cBObYyNqgX7
f/5+8j/QwLd8ptlzoA5nsWTrTFsVnxFWCQ+x9e7bA2PmwVvnBshUqn7M8Rx6Kn4YO1Y+sF8Eh4M3
huP5fHM1rWHJ7hUkCDjB3zZYorjKP4OaAkvh+hBoLc+2E1RJ/fgH6GJEC5rRYREkf/kC/X9/+kEe
g7OY5+czPqfiWIXp4avMk0vn/DdL/UqZBmwh4Hx9Zzstzj8w57+sylY482KdKBZggjtPm65KV/UA
sMucIsloMgR71lWFC1x6pFxnxIzb1h+A9A/qPh8OGGuCYVrSVO7J1JyTa2pi8tBVl2fSn+1sLsjT
qmAe2/QtH8VzxJn2Cz3W+PVFfY63cw2Oa8/2Ub1db8thmOQkiazfee0zbwwY1FH0K4+ODV1c+gWp
Z/K2Fam2AVP53UaPRmKgDSWGs8weJcaEk6NV7omwnoPOegNAxvwdDfC54nVKqoy1yWreqpAiFFAp
X6h8ooDDfv6t5vYE0nKI4sNiUsLqpeptdustboYv35Gds1iAdLiNpMio1cdiM+GWyOxKKDACtzW+
tjQVvKRe4NVHP2DpnwrVM2WQZAhvS2MhyRLcRtUEctZYjSfO7pppTHamlV/ovu3aM2xm3xXcp8RO
A/i1qUZaXSkX0EO9qfJqSRRLUhmUGr3+NW1R+gdl9ZLgg/8bqJ2fZKxI0XalQxCJJgHL5W3/cUfB
YDavx6w2gkjk5h6WAPZEzstPs1rcmreKUx9XC9GXru/uf04lenQDr2yanzV4IkQouMGKlSa2jXu3
57UrTj09oLhhsn1h7qSM+fqGa83l7y0I2tkg0g/M0T8bUsvD+IDv6EuNERl1j4wXgZjbHD7ngvz2
t9W50jAFlPTxlTMWnW8s7XK2+B4rgojCvc7ho7PFBrEL0R3rVyG72P2eXcMr1w9kJ88yj7Yqr9dl
ot+EuewlI2FtJFYYe5YMZD5R9Gpx0m3oQ1d2TbI9VdpXsiAAI9AVdlgfg+zn4w0q38dcTZ7X6RFn
ZpCZdorqKyArBuVNyLuO3xTyNSfv8U5NMKjlylmRwbH3JaLuvi06B8cTLkXjkof1rjMO7CbW/uey
eMnSISBWnM0o0baweYsuJwP3otj1AWptoafaGgyy8if0HdOxnml7QvYVJU1XlNvurio1/2wkwRcE
+SPKrbz9GkoG66c89MfrV3KbpOzyIf50Igf98RsKZ8zWGtEayszWN4u4AfQmxOTiHvgdx5e63dfQ
mVgnqd21PHB0HA0fye/432L9fyMePkyJ0chWcFv8rEYTlCyMyJPOU9GnDKNxdqW+Pe9D6YcGpZwu
nKK2lL0rmSYlUJrAZub6na+uwzHFzLIWB+ixWCiSt6Kb7EzdTKA5vCRt2ZzSrt+wJ9s91IL7V7Tr
iLrU8n5F5U7w6Osm3Hx5rCClAipsFMzxsmKcG8M9+Mf9KJufAVx6gz8pEDSGu3X6jke71B7x5SL6
3M9tU2G2OkvHcocwb5X3FPvuN6NPegFDXzbYmEp6EZ3ahxov8LJzEHSE0UImlmp0uxEzpZflAufd
u0dxHYsl0KMUvX1hoN62SilX2fObmIU50BgTpN05h7CUHu4aCd3gIf4s221X9hkL/EIgUCrK6YGm
enkFA+srBfDvultOe7DzhOzBJkDlPlkivZViJnQxxpieWpo/Qb8WzD8V7mygew2G5cRtRv2Pi3d/
USplSu6h1bl0KJiVvJSBL19EBxIzj2hxJq2hNVA5j2tN0pMQbviIN0gud9L74ltbE274ZenGvkIR
lCQAU03sWHjN9nuiIr4iI/UuT9tEHrScZ6DM2VyJz6w94+PVatmxmH4FZN6EDSCp5VtbQVgN6GCo
eLaZVneWRS6yGyEYbmZwZC0bQTEpXQTnnnOTeiWjqi33QJbrbeqGvuVrSA31ifF+IQj+sNGmW8XE
DXTtLH8p+OJAaZGpA2o35wKvcxoil2SNxNao54hE3dzQgsuzFkEgWk7afY9NUUndmpXC0U3wR8Q5
dxCtZBsNZcrWVks8Jou/PeD19KMDE18aQix0j7HuPy90x738UiwdD2qQN1N+3ZGAMusfqlP+TTmv
eUSAMPL+S+qbNtqg3/ys8pOVMqxOiIsA8jbBnsuhkmIPcNGav8OY245a7ny2cxAW2npQFT1jnJdo
d1Y/ohMk9nW5kXytNqQEkg9npDUdavhRgIubnpTDZ4968W3b/9aTIi/kFTS/1dEueCrtKZx/FhrJ
2E3p15FEFt+LSQ7xP06gQonjB4YNTF2eQqd2TlhDf+1AuV6h67CRlwGjPMqkLdObXYVXYMbhyRR+
0sCGjuvgYMpNC6k0m0g4RDProfX8Ll7JGRAfpQ37YL0POGN4IvewB6MnX5nnApW/9M28ld1U5SPa
YZio0ZpWlJGqH4XiIYE2pnNc18P3G+ikmxpZ5I3SL3ctU9O6+rYwby2Rz6T8a6Tu4awRWD6TCHAy
MOX4dN6hzmmU/IKoR+Rg2adp0317Hiivtp88AwcYYHTaaUyNC2Hh0wsYzOC3aMKiW81jxsulc2+r
JX0NS9I7RxamYAMxohb6wjfdV+nnv4hx403vpDBtm1ENfb+bo4hilq5OCpib9TziUl7YeTqmX1k3
3/SWVGVEQqE0yKG7VrPupCnZRm6iBJAFr408tb+vK87G/72+++ZOjR3mQWKbd7lTv5Nd8Ck1ILvy
+a5009TMf9qWLnmkuyjfEPv9gmAAyVK2nA8HIEPpadZ+2Wx/PpyV85A4/eiy/vmfF2hkQOusX26c
8V/CQS/qct4Cn05mTV+LsYcx1dXCHt2qgzvQrtK4mlLgA02mrWyBUjmaMlnlrvpaaR4Wvj8FG/Bm
MQUQlyqjV1r0S1lP+ma2un8KosFBDcblxm0bCe1RKVushihGPQ6D/c6AjfWhfROCFBQtTBKOYOgb
AakHmUnEgVO7l4Io2iY8dkcjp/UivGlRbELDj0cMqHRm7zbtryk6jFsYIExD7G9zur15wAVn6wyt
5sCjkQFrLaSAr7ksBV6DG0QsNgJq5m6TAgJ8ES8LAHCsc90QjscXrIXPjUCUKjF88cfIRsVl7zYl
l2Fyq0E0fE78IRRY4rm+pXApkPDLMO+xyS66lGXPzPFlnksl9Bdgu0YJHPfykTSyCZ1iLBT48yy7
Yy82yxpZ4fodKA52FMgHcvFFkAJ+cfzidoXq5P9Wjw1s3LYEmWvKKsvgm1b1awYptEvX0ph8Bq3j
EMkuiM9EGKOtgARfc71ZMs5VrosILSdn2j3ORSgN+ZJADiEcLOJjGw/lI35nQhgCHiiG/dPBqfnA
S3M4sM/+xt172zKOg3s51iIXwGwlaM3rfNOrZFKVg+6W/IOLlONnukU5r78sQtKbAEPVHVIvkwJH
DypBD87sldVkOfxOrbRV9P6hd206SolbcvXoWifJPE+cO6edKn7kphUSCk+0yN6AIMGSdGJx+LCq
wCeRKlif2hUDJgF1/NZciJ/JTeZRgGqbXxLPIkVjdhHpDTVSHniMDcJVYrWSOtD1tgM9Hf7CSR6K
6hsdWNsbnLqAeCC7QTVlEb90bUJJd8GPQUjCTsRWprHGdqU8HGxPj9qQ35xE+oZKNc9jtJOHRnM7
RGkHITMeIHP1JABilzlDkm1U7x8tg2tYlCZnl3syS0jnwzKMiH5GnjQSlzzlmlQ/PrVx0b1CDhim
ljbRJ/fgVdQ7tDkjfBguPmuW/bgVyazaCAA4mLCZTbptnsunUGIG14EwVLD8xJYE8VxfZr/3Tk2x
MCxQxsVy2F8l1X3d6/+JHNc1xYy0AztAZNaytqdjbWu7jXirWtIUg+pjCJkAWxVG0mw8vt9YtZA7
IcOB/qeVm2QWvtt80qsEuER1FQFspCiA7vJVEHX1Turw5Flnka+eVuiQY2Z/BitsGuvM0FwZQY2m
lEHpPAFxLZ3Xm+oc7KSGHtC8DVKkQd2Z4i0M+4xrwkOEBFVcfPoe9IrKWc9afnnVg5of3bldgKNe
Lf24hwJgzUNbGd2wUPlmWzKVPvGTUXMGk7YGXef/H0UA58rNB9XnEeId1gUiSJYIfArWHcgOW/5P
rdZf5Wb4y9TNukYYVc0+brwoNnrd8gsKO6pkQ1K7W0Q1k4kkDz5bK3fnyTvV9rJBcGp9Speykzg7
31+ZHJgH1IR05eLpYBDaD7qyxMl1+xJN0/mYpExhCPukE5Oa4pSaDqYX+vDNeERkE5XncOhlGxw4
fI40yKyTbDTRpzfgC6R8+lfTS22vbtkW0GqM/tUEkjJ7pNTOG2sZb28Ms16hhPUrxtMVxbVBbf15
nrGQVqhKBaim0yxijDHZK1YZD+klnRIHuJ9RcGZOoszHzak9Op647Bf0tXxowY6zINvCCMfZUorY
Nl2MtWx3RaydYmc5/q8HqixrXJoL0hTUwBQ1fjh7ZfJf8HpDAtkZUVEqI6tf7rwDWp2bWCGxnnBj
otv8iR4XmLzzczztBI7UynEM2oSALq93ylHuph+MppM04hVz6D4SYeFCr2qJH+OcPZ3V2qe9ybP9
+bVmOu08S76JgdHr1GHDUtzyHQsZ3SMQDXIXYqH51n99Le6s3lHvczdbEcIex76AiIUVjRrCXcOr
isrIn7JymG1iVsQDdMbknVgy8Pbg4U7opR8kgOAgfcqmtJouEEOwWXRqCPqzZXAnlZTWlb7hmXbC
KHJZ9SlwJhjKk1lG3u9CBkujQcwQ7/yqqANQA+kOaY8I77vOUkYGIuGnR1fCisi3n2ri+tgCgkOB
NRix4Ld3fdLkqCJqpNpRNlfmcVjvq96Hsxiui8C+xgVqGiSVBcLQpKctDrRvD9oMJgd9KJtjmfzX
kKRNpDtTqgkuWe/Socgu/8c/7dhlbm8I6JpMxiAGcHCNqjthc0PHzTUv1kZT1P7S4tyYVizk/Kv7
SKNTJFSOXKfyaGxNGioLpAWPE5eUOo1iNTWGVPt7eDMpvOIuMBAdhG/HfYwP3SdfFDyb//4LVuaj
pG2ILln8AL9asrRo95WgUh4qcyqhVWDe8w+P2oEw9t/LSl+hvjqw6PeCNvvifkOsumQF8e/wVFnx
o3/3tNzAnVz6BSJSmay1rTnzSRLRLwrxSXezwGFOQ4lhVm/1ZDcThgpkBCZu4SjXpSU+Ayc/ynZD
UVBNN6JFMO1Cvu+fXVq0fWhcwSflEcOr7Guo0ydEqpV5JMEIqoFbaDP0GyrUg2pnSqCRkGZ95pkP
I5w/MLoSej2H8ntliy9PM34Cdc0p0b0/XrSxzfJbxTf/ROy5fqNo7F4sB6xyuH5p83984iZvoBQA
yJk+FNxFFkC3/ycPxGP76j9RBF4kEfbyKop3uaUn4Drgts1vWg7fJp1X5v9p0UUEzNfUSDBc+yPo
mpzlf+SWpoVMAtBdm/wk/6UE6hUZwpLwwFAXpXAszkoN1VUTqZJY/xpaq5ptNuXTzpBA9sIRLwNE
sBvFYgnvR8pL6zb9XFYLRjkJLbfFlAUU6H8D4EaWeLjRLf+1bnzawS2OKwyhmoKD85R372SMs25w
RMLpRhRo/zM27UWPP4OxyUtnV5Idm4zMk5cvhDg+UN9V1Fh9X4MS6KJcIYSg5TNYdQzc1dvgtClX
SjVRZhRhJZ8jN2ChzFwLZKbf2pJVBXhsRiX7/yzYhXKnd72tDrTTmjfGMks+cMpCdJ8CzhCSbOP2
/qRIScdz+HPcehDFLofCaHrKHuNgQwxTqcAFwj9GrkhMTn5ILOtY1MmEE/e16XfWiENkrchCyECG
tsKQjCJkJ2t710qcIr6X0mmTk09Bj03KOMbho2RiyKxCTE9hjI1DoifkSXkxBz8SYmQYvGxeJq8K
cR0r1H8CWewbBfqUyogOQqMUs/1aD9z8X/h0SPPttsiRTL1YV6iw+rjJcLu44FIvA5ekhhOGpSO6
Pnv/GLG9eVdoL0EGjo4YvzDRL0IpCbLysJSxLapYEu3M+r8K1puSCGj7xkq/OzMzGF3yOXQMCgp4
goomlq1C8NWM4rvhptguvWTp0IWJ/8TuKTEkXhbz7fQQpXb6FljiN8UUqqlizzS/gqLJZOYHq7tH
cR/m+Q6pOMwAg9gLihCU40a6hAZEJ+kXjvjMSz25wcmFN9FhB1ZDKfZQ1yFoKqSgax36B/LGsDXM
52p7cEQYw/iQXO6z+9iE2Of9DbH5B1dU6KBdAn5/sPbxHOdUcZnJQ55JhM5V3GvAZuqVfJOeUz5g
k3KnlyDBcSmVKaLV/f98piW3C2H884vMdOI2xdc+0wMiOP+vhBjDbFJqg7jcN31MByPgvZIm+ZSk
XHF3Fi/U3PmT7cjoeO4mTi+hLWowoOxrbJY4BXDzKsssXL46aW4oiUmp7NBUkA4gMmvO4tBHZv1W
34sXLZrPLqXoy2FBGzKLvlEyAxe2IhHcwd0aq9FaF0MNc9Uat3kwDEfPwWWzLVQHpyXl1+w+XjW9
OmdAZmwBVhKF5WF/jbENBnq/LNj3/JJmFYxWjpaUvt8c6bl9om7csNEvHW7LKXJlWQ16cTQGwjOY
Ll8hknFyENQCGpN+/ec/5TiH79wmPjPyhrGZTH2wKFgbvVIEv1f6+RUVAXtKSSQEEC7INfWrANmO
EK/ihY7n2U4GvBHE5BPOGNjDvCPnx0QwZCRXIyTn80LVKp3IqxETfnBzGXifQ4ZRnYM25jLDntDD
wCJdEJoo1a3w418YdtcjW7iQ/rX7ZqMCKpe41KYsE2coAYYrS3FTrXzQcJtQmGQgY6KhhBTwe5V+
bWEsBfjQX4CJqwCUs9bn1oW7rGzdCQPL0KdQAxOm8dbm5ogMzcOG7etTT4Cwy4zM5bA/Pp9UnEfB
Dqi5T3DO+O8TcYsC/8iRFQbgGweqXwmMmtlYGztyIxn6J6xqZhiM5oJn6YzI6HsCLQ1mYUyaYSGc
a5/NOdJTrHWvQTGj8neNwsAhx2rsOK2NqlbgikWMttMNdFq9Y9h0E9+4qwytuE6wXM5e3w2Io4TW
dVzXh52G8MHI4n7ZJFfltcBOlU0oTn7caSG5hbX9cAow2TbHTgnET/dHPYTKXsQXSdBPWR5ZvFYA
vWalLTTQW9sjw9pACoxavj++ARG2HbsddKDS4vlcfN1XsXni8sKCy+43QRWI4geUGfMmyZIE/uG0
07/Tjg+i09wh1hS39IBafafj+BaB3aSudPG8Hk+7enoWUtmS9VA0A8SVO21doXflRHO39cdBqaEX
daZSC/a4KC2ncuaG84ASszd+UZ3FfnD1DasgSA2JNgpUdd3R8iNLUM9EgQxxeLr68a1t8XgYcgJQ
+/MT/dtS95MXvHiygO/52i+e8CbFrTR4KpgQo71dWUZd1Weuu31+0b1rOTyLfNMIZ0b9/3eQ5SVc
kCzKBNGfNnGQVpxxpMubAwkVdUeq4eJT6IMagS2NaSwcscqfz+EyR/eI7XMoB8E5hdalJU+azy72
XRaacMPvU6voKEpy1a/rxjvepgay5uWjpbqkbJ2jo9kDJGcn63ZF4QJVw7m1qKeGbEPQLo7402DD
4coM/zOWbbVER6Acv+7xvXfjpNqwHIVnDPozofgXS1JZZqlNy7z40ZBXk5EyEZ+7GEgu6UU99Uvy
1psPiDzl6ToiuglhXP9+DCjpf1QRv+oT+RpJHsy8owze5DbxW6GK73AheADR3K0KtrYSIEZdUs2M
/LwuL23C/MeNW1oUzjM8G86007J4Jm/szXNH/eW0Z7CkKpXy1qHr6kxBoNk1VQUJVCQUbfOaIAJD
g/98J8Sd2wxUxmFGzwPkvCmMzFQuec8H7T9Uid+LJ3LVMgzECpN/ddrKz26sxE+kv+Q4cC/hnqTk
BBlJ2NWgNEAnatvoTjwVSWkDCnSoToZQOWLyqv0eyYX4qq1uXuxc4roIAXpCXLEJ6igukpXO/0vl
i+GhTOqC/SMpdnZfR6eR8ZSMaSMrRBOuDd54r4aSZlrmZMjgChnz34hplU9lIrwyu88Bqw+eRC1t
4tlQC0pKRnWWPFLG+8MFN5XZ0lSYN6I9rZx7kVvubHteTEJ9aA4xcvO4ujcHUn86FVbBA60+lsUb
k8Utzu7e7hlHdOiBStgseRwTXzmmLmRDN2cyVJ7oMMstJLxhtOGWPzLvhnGhEWfqNEzLbnf+E+3T
QWII4/qDhulDM48WawDnM4/YKQqvMu8rrVGClvwY3Pul70ReNNzcGx8l+IE8WVy4L0fUznvuJQDd
6xSQgr0S0FbOwHumNSaoQrwcqwldm3bBZePuEbvbxYwCtZ/cZJBlbnnUBqZsCLnbBJQxFDGxhmmQ
hJzabOCjK7vTlZXXvkLo202+fQ5u0gfzYAU8zZf43uQL6hTFJZNySPeyjfMNE1LYrPAgCwQB5+J1
VH3c/AuirozXwjQDfm2iU1PHvQtS9i/0ATl0waZB3VrC49brCLKWjee2RevNLtZMVfpff92LOG+T
bS4OS+l7DmUkHE7qHmOFpIYpW0tez50u0/cfmjCFqwWE/vg1xHY2PJfnPhSTIFd3SwQBtndjqLR2
cqSlrzvEHQM9Y9/jChQqozLJNf9VGavSE4XYmLsk3AZ9RDw9K76/IJE+UDeeQY0ijZPLOX8i7y5e
lZJweniVtR9xM6DwDhGJapiAFoZ1A0jCybBS46BXiu3W4yxg9t5N9Ewyy5Fxt3rHmgbiBBZE711X
70R9lAuNKWYBj9BNFdEdixStOoxbjkuffzSSYUm4BM7AOZxxH3LdoDVikAnIMsav4pvl8H/5jq7t
BwdTswyXVILQtEDLblY6Xa0zq+wT0ch1Id47bttqDdHh+rkhF995toSPxxVowOFEeansm7egZnOE
WFkHMHo2rKB/8qeul9BSxhX7gFBPi4wuxyYfrHYL42QlJ0jXpN113OMtPA0nTWPX6BVKsSOG23x4
/M210hDYB58H32veloFo1u8+qoE0eRbc4OKsmwntJSrK/CNXowDuh4e3HSvs4O+5ta5luIB7dgDv
cTJg0oy2aDSyQ9huU0gn8fzAQwRL5V88X/wSpmB+hsmowaIniVxKdvlySk3PUUMR3vNnDsUFHiaT
nAKhRjMwm0PgnRQCj7Xu0fZ/4s2bj/EnaHBssqZ6iNQ0kAOQ7T1mqMDjR0Wps3ck3DXjUq/IqbWI
N8ReWVh1bQU4zyhuII+QLFA4W73xnYCVMMWjJrfe0+Ph6AGHzSRU2VDxSk8haArP1V6jUjcGNGvM
wU3sH2zmWUAa6OVVNLkgHPR7NJEPYjw4J5Gj8EPY88oUfLM6w9ioSq2Qk8kHnK4voLsfsLDOikjJ
T8sT7e1V+HhbzDmc4dPhtQwpor+DadBDp7fkXFmuy8oPF64QSCZyKckzvrSrlLDKS2rPViUDSj89
/dIU+EH1pCBSOvWxg8DjEQ7VFLLC3F5WOtD4gK7bA0DZGehLHZNQyRCY3Of2vUtBCK3bJSeQFA1X
r6tjWGNU6SbHi4M0TZqSEoK++pE8CE20v82GBynxT02W0Uzdeh/b2RJ4iJ5t5AH2qfgbVEi5HfiB
v0oz5ZEjEpAcGU5ck6nrsVhKp1gQsOUSIuQDmcOXXTDAFL5SFjA+ro5ULPCAL2fyWpZ+/+CD0b/U
RjlJm8vLs3tUiG5aQQ4tkluOM8aR0BivcvMkWd9a1PR7nqKw2JuZ+zu+aNx775VAoJpqv6Dwm3Zj
sC+0WKS6Y5Qx/ufogcEynYcX2KUs7yZQq3XtLpUZ4jMlKAhtmq2Cq7FXyd/1u8egfcVGtPBm4LP7
i0j9QnCkU5qI6t/hD+ipXkzhtzZq8OuBtMldjmikPZ0ZYRrCAAV0ueQi0dduOM630A8THKtq51ZU
fpbP5BE/15AeY3K0AtdfeuugibIxqyiiQNYbYyQZceL7a4hQ81eMZ/0e3rV2u8VnTV8GAYn23FEa
2QwnE2sElNHrnwFr56ofzHiDJNVSbHui7DXA6p8HaHnKHVexZ5jQ5czrINYctZTIE2UJg5Npq39+
T+mBtjfmAyReN+iXeX1biATRUK0t6J3XoQS2p7mOBx3k0TsoDciMd7TuU/Lw9Ae9e3jDFXtYqsf7
0LiKEd+YXT/1AVPlPe1DkZcSSoyMOhDNkUOiCPLGR4LX5evoF/bB4D351B+Fi0HdEv2ABcupie13
1k9WjIF1oH9IM163k8OdvGj1tV6xtIUZ7H1w7Gyv1nRVNDbfNOF3267kFI4da2ET5uubkvjbBx9N
h4thxltPEuzPd7bkaXtD1QYhwDMqkFVNJruw/OjLp6Zh3JS8ivtQJUR4Z2CEQGvpFhFQGy1KS1Hs
OXUxqvMuQGoJ9HAxCgsvXWW3QdIvN70yfUC3qBQDjxJJZlEkey45mZ+1xnCabQvhHo+5E/m4csKE
KfBaciQy5w8I5TLe6E9XDgzqBPdOfp4i7RcZZti10f4+muxBADybEUfjrQmGAK7FhtdPDq+YcUWR
xqDNx71AlWz0RDceICXXDBOsCjLeMBXCoku5mkds3aDwEyEAYz7zG3SS1smrnZuMh5hwnbllLJE1
hS2b1zwHT3ccIYHwYW+biuWRZ62gSRpRcKb+HQOSObrnOYI1rwY8vTvi/iZVYf2lVt9XJ0FrWYFL
z7mTsE2NGHBHIX+N7V3depvyO279Sk2qxhFTJkpZyzXC2W0UnF2c15TksNEH7VleaZv2QgfPqVPb
oHMyThj3lVwtrXRvRPObeCmTvLPhvohb6TpE5dj88RigkWm72/Upcf1/ZzLUfUXu0aAP3Sd/2Zrc
olpU9L7fkIHRopwCy0KR0pcHJZBwYpRodSE2eFo8XhRa0pfpWLEzJ3CgTKxJurbPXubFjBLGHy63
PtejX0q8BklS8UbH7iWz2Rp/ylFiWY4fqhFQXQPqeBeyUP3tLtBWMjdxgPt5C6qaxnEj4/cgW0ON
Zoh5xpV30p64/Bn/iXKPHg/toXUel6sF3ahrlMfc9TND2XF/0R34Q5hazDEU1uTE+SuKPacjUYx/
vrb54a/5E3j8ERhLwWubh+2ZOFZIQujza0bBHL2cVEi4CxlrO/S/tIJx08b+ROWcOsmW6Xkj0pZr
Zn9Nx+TM39XOF3BxLWqwruIw2r64OTcogJEfb7alXxtQ4bY5iG0mf5wA4bRuuzfzpw8dwh/uPieW
UCGxJ748db9WhoDflbPYF+IiPy/BH6/pDOmLEytmEEuJ36hdlUSuZxExr5Ah3XaiANCEJGUz1tbk
XI1Q4NVr5s7Pa26eVoH5OSLI5vkzjzmPb5Jaiqz2HAvMRd6e4XL4lkimGKcszN9AC1r8aEJGZjfO
yNvxT98ULPNcthIqH5SfcXUmU43JOl2di9RCcewxGkGDdP3qkI1+dakbNwifwkwzcVtYVLhtcouK
N6CPTv+KpQG4sFpO3qkIhDndFdTcOw7tnzAv0bl6otGRofiqbdH8SHVauGttrp8dz1tTqN6PZant
VfWkhNwbLe6zaKTohoL7YkYCobSm9FEG5nOpQ0mD0Yyoi+Kyl2Gd7FkiG/mBJ43ttAa/qjpZOaR7
G9WqXrxUn5qzVWTmR3FKjWYrk55WKK1wJjMc+LcSkbumu8vpQRdfdjX9n/4KI1tEs05HvSwZZ+5N
5HXlOp4hmOahn8rkuy9EVcQzyyH+iG9nEwdrYEQFTNtw5JJQdTyO865ha6065JV9kFGZArGSdGwu
u6gMlxzl6Wt1qk6PMpRIJSV4B2oF7psMxmFlSKjf+erQyA4dcLBAjnxW9DShsJZZVEe7Ze8nO4s2
RhbQt+5tq7zv6+rNt75rWKD3ReGB8Q+Z8jGqtuDBcy3fhgNc1x8TwYWEXcmPq4wFtUuaE0V8Y9XD
1quv/rAyKDY6u6U8vWjFZtz8qgzzhM5lqUqDqd6uzbaIDocCl3apnimQsSfbmeiDHJyEkbO0iZkp
mXuuYy48IxuG9cwYY6F95RFBp3mIzl1M4c3DOcTCVTJf0bdcS0uUHLpTLbhnoRCciAGEsd5qCMw8
9nRMopmCx6UgVakckDa9sxpcIsCTxnrrzzENojRptfD8Pz8jB+RKGg6M5B+WceE8+a8RTKli1l67
0+CIt868Sd8HUrFupMbOEHgPjiUbZ2K1pvpp7/fqB0RArvGpDUw+fojVVL1D8zeefP/SnubCm2Kt
8AcEKgtimd92puZGau/5I7IEMKbUdoYvoBoJfCyxavnzm3ATZm9eG3RgL5pQZa5XMhcHIngrsk+d
4W3VsVpVzuNSYm0uQHVFyZNxd7CJrIRBN5ooFOQvBmp55QSCugICYiKlaf0NbEKLxz/gJnwM3/rI
pFQoru7R6b16K+PXn8M6TqKcHABNaETIMUN2c6OwUKT74Yz8QCVme8VD4MbxoG/t67YLHoyFAMf6
6UJzbzGG1LSmY9ibqp/5860Cq1NuPLQnRv9D8HaZlLLQQySTQ/DddTI+9dSgkrc10oTVxP6FB2ZZ
AWdvLcL9JVBX4gMKY2oFnqT7nHgUMdhtvvyUheQSaqUr8FDiSXgwf1o7oSrHI6gGH3XawEPVfOx/
uHG36fiDphspqYb6CRuZy+zjXPBxAufkMyzXHSlT3YqBCyAUiGsxTF1okQL7/9Kt10/3Jt5IwD+p
MUdOlsJRzUJ7WG2xbF3NZMCn3HNfczjJZGPpCy3iOVlBo0FuoNlaXSSd6qLaCfRNcKY0tMIX/47W
W6khdH/cguMN8yCBOyMMQK80wsjueZgcg1LcwgZmNj47PwpSt3ZTzJLEadnN8QoOYd6LjPjdLvQt
sBie6hMf+P4Ccz/tnbdTVRJhMbeaQ/bif0BqexM0aF5OXtiNwFhwAflMAIL8FaMv9On+4WK3Q5o+
lH1h6+QCGNbYrGV2CgWQM+YOzn1XnqraUtMFshqjOrZnZG+WLbjdWFsECO0jlsprWac7b1QwcBpc
KKw9QwEUzMKRSj3TuNGz5GIUSf+/xioJIRvsxecjfQtpC/Hl5esJqtJMbI4zVlBHjsS0q2mNyWwI
dU7fpM8NlH6dNW0x0Xns5wSm3l24TrM+9HucBs3qUeVxFeSpwZzLbXTlm2vwulPXuikfn+9BcZMh
+g0PRaWQ14O7A1dc0fm3e1YDfFo5mqAYT7HdYeaMBVNtBN5XGBvVRyAODPyxZYSmpemz48V+Hugi
IQoOdhdXCN06NAEpQ8Zil8lbcigLmF8clOmDKJ+z+Gr3nf9rYIgVrDXfXCkG19qwKHZbHplGKHAU
cVPy0BIGa+VU31jdG5CG9O0KQrKL0xhZt0qDz4SQ0tS1JLU/G1obwDtJxitDQIm59BBPAWo+gR+5
clt0zDxADq9EJJ9bc19CqmW+7J4rJsZqCbpJU9V1kAyXmLN+XylZmtIaKux8PZbbhl5k8dXZZN6b
m737sTNuiwrSHhujckQV9eP9+XdL6QtuKoeidROozDj/tARmwysVQbdqsw5P2EawV1VzPSbjhtjw
Z6IP0X18f7pi5rS+l78yXrQMY0MGpILn3Yj//J0tlD9UJ2R0HztB83MWTL7d4hWf9celiy6+pqq2
3UZlyVLBc/46mJqo2YnTfbGInVzb5VaiaQgckyy2b3pxxw/hamqnmAgTW9pk9nR+jI9FTr5u9sQR
9WKVJN5G3Trihdjca6C9rJUjBGwKS6+MnXBHCvgvbUu6G81oFlJgSy6PiSXWyB4WQz6D9yC5Z9Rc
4c5zR69Hwju9URVPlRAuvm9FDwz2XgjhVPpmXXP2WvMwcI3fqZBsFSbDHmXDKnijByft4C7hqO9I
DiJHCYYr0LPWA8e0terr6uBzYS4avyqh//S3KUKBUoleUGJoG79nfjMkfRACtdvAGPwKELyMZKtY
+lT5vb2DEgct//fD2QgxM+zTFQbFD/ITDPc8c4/kA0inyanFlJOLdvrNP4YSM3cwralL8wnImHzo
q8KA0LTfYW8Ekn1VxWTBrVYJ7biOLz0uDOeQK9ygsKFYOAj3KiDVo95buv10gKXt0RLhRx6mLTEV
hErjcb5pmevh4t7DNfw3OfD1vaF5tXHaWlznM0cEbqdQuS0q75fKo9DuAIdejCZkJGf9UYL2opdX
xBBnY24tnM5EB6tlXd+8ukegwA40fzo1XMnwpqL5JUsGs83pkiUY6kv7u7aL9+7BNSUNlsDhCsrA
CcQ18e1uCSTh1w20bD6qfahs4mvB6E5Dq85aM0P31I5AOew4Ex2nqVczWotfvZvUt5PC+isjLhGY
IevJHCBSHB4n1weeK2YaLqvDMQS91wr2sA/QGk10EO0b79gdQFGeydgwn6nYcxWJa0fVrV8S9Q6/
CLAYlSTJ3zTd9cSqC77x130rH/gJK7M/wMe2rQ7whci31rJOM60nQMxyP94DBmkfwiwU2QhIID+u
IYf893m1YkiN9KzfEl/YZQ3khv6BfUuU2uvQXcQdOmVtz7Wla7LccCZ27hdFANT8bTLq9nLnDKhx
0iSVDb2ZcHRF/T0fl6J9Un1na6tj4839LdHDOuALAPfOaWNO06AFzItWYYz0l5KbYcaFyeRH0Fke
QuGCVCL+JosWY67i27mNqtmNjTsHIxy0RJOf0hNG1igYsZri7TEsFRwFs1wIsH5SPfW4X++45p2n
s9DpyYITpnwADqDKLtzMamkJeXxAZ6NMx5mU9BTEnUke4wPrVmuF2tZBpq9RFLQGayqRZl6u25yB
V0FhQRGz2OIAnC8SflHAE7AhhF/BvKH81u0XOab06azrU9HNUCJNMqbqGF2Lk4VGfFLXHnAoTGAs
iedoP3/r4+sUJymQlEtiVcBozvqftrUa8ZerGaA7V6+jLPyI+nRaaPWhAk8veyFSSKWGnoQObM8v
Bx3S1sAhXNDzuEH63rlLDUzTRmb5fYpLGDOiGzJC+R/kREmEezEfzJXX8ySxT65mhplQc6m3zHDi
B8TRLCIFjNxR417C/BIRwfdXvLsy9Flt28g3TupEpGuo0q1HiB0PxRTtWDZl+Aa0JWMqIbYWRQuX
pLm8+oOLnT30HKGF7Skl5AL8GfqWAYbh66mZos+1k2CdJAko8mWJF49n/a81pVG1mWt6RfwrQstu
zUXrfaaPq14k817CfbBsHyC1ev0YsExKWBKk3V25mbvOuI7OOUnNgR2msLz/MhH+fXCHvkXGdh24
aMBB5RmsGNfO6E66yW0QWtvP4OyHr4TuojawEq61MlHMId6f1WUVZl/t8C+dKBDy5GKeX9/d6Bqy
mN4k0lGBJsWztH/oec4jfeVyKM9cNpy1AkaaIiTVR/PORGo2NkO/CfCLR05N36IAXbfX+es7jGRf
izowD3Uv6jb5EH7D5JrTaPBugHamZ1dMwFAxhELUIstI3c+VFclA19JqJNtclDIDZA6F1lrpRRx/
6SyYMSA7tV3mu4UBBguh4HsWgVTtRrad8UPHbHdMCyZGod4/xyEt7Ww1Im/ewHnsJQo6eAvva1Vx
38EOSU/ZSJQZznEKJEp0LN5fLaqzIWT3Kb99kzt+8r6aqV5Sd0ZrUx/p3SHZ6iydsDAZ6gxjmOQ6
WOZ1RLVT5mk10NR2o6rROJAd/o7DOqqZsGCwGguDVILYOB1jHp0rDJETq8iEJ5SlicRiahSbtSVf
Klgo1ZOPUgmUPKyQ3mfwm3BQ/LN4HH3XZvLCpJ7HNPdzyvXKxAwNPxAC2kBao16H2sGZNFDxYZ0J
n05PpLHT5BeDMeZBI4agNmq2iTJXoboI9QIJoTI4pIhm1zF3Y+Z5Q1c61Z8HGjoJBsYk9rvP/fY5
8LW3+B1BjEpDqV1L26UsgTHUtBO1QMtr/KzqH7Kw5/uclGcTJXjznhUTTZCREdpEFRkVpMNaze5N
AQA7OvAlaTBaFfUnvgBXIn2HyrX3XxoNi5ju9WGVy0iULXmOjY85U5xmhvi+hFPUep0N94eeEcN5
0WMv2UbYwU15VTTEm6FnY0RmVUVDWjBDABFh3fXwdBUwqE1S33QHPfEcJ3DJNH5BoxvUIyfMcKmj
FGz7Gnk+N73g5jl0iKUpEQUEix16470NxpFnuiB2zUP4GFOc+KatfCe5wLoCdLWV+pzbS+dwkAmG
13SNSkz270ooD4sFxnXXh6fB8OBUj5Q5pejVp+/I8i/GzxVLmkSpmafgf/womTmcw+BaXstdFOjD
9hYlY/UDjqOYQK2uQBqdSDBvcxLso8cMSgGPlP1s5c6Dy14h/4QIdeRYlZ+tDKn8kDf6iZ6XlCn9
wpWrPO/oDL9Rvmpj95raKHfxpEkBl98ApA8xOOpJTX18ht1j9Y5Ghi8QPguXH9hU9vsENctmD+MK
kCZulYjDjAvF/NRt3AAzkaVvsy+KJj9ObDN0C5F7rCDLy8wo2q8YAwjI9LKaDRi4UZnbxsiCaJIk
bf4oBaTYI+HHecOOO3aR7VBR05OuXnmXRcsuXJWzlCwDUi8Jbs7ItfUnoxuFBCy3tSVVkNf7GDuH
7JFSxwjUr8ijUUKqCFAklMEwso7RA9iPBixI1MuJusKCDjUGs4rB6aKsnh7nJT9K5I8qVzBx6n1C
+vPTpusLTVERhBo3Wh9EWZTvUeEQl1MogQv7K66nz/khxxpgOT8c6sDP0AfuZx/G0tGu1EomPxlh
TgooFiaB+jXs0L87yaNKGkx3g7RYg8w/MprSkYlEQV8pKLCNbRaCOpzM6e9tMoh5YFk7+rOK5+fC
p6HE5LEWLgUMuv0Q/UR4oN1oo5ZMms+rEZHA901+GdJwlWiBAE3nwMMSzc3EmFi+9vDI+OV+rEq4
xWdsICCodTfqIF4gDYElrmzy9xdedh+i0fuPEBN5gr2kmq0M6SDCQL0v+u1X7iDGZPayg3RZjpKW
CsRmiHmGEtcnvUVaTbuyOUv2UpyRigCF7yhDLW+xdqH7AQSvEEeu/pm5G7WZliLd8gwYYi39VWoh
PDcXIJi5ueSA1gRN7FrEByhMqi5pj4NX1HcgYrCoAIFDTvZuvT5CRmS/Hp1TWy+olMHJPSdCbb41
Ks/kw9qNYnZmCbVInpG1uqBw2+HNT2TgPxcstESVefnJqD8dg59gYnM/L3coLC265EzvxYj/ZilB
9X9HLcKUgQWpoUsPi8d+BREEO4xSi/SamXHPL8K96FtbJpy5gIzJNIPxTw5FPv8ELrG9P0evQBbO
mi081jzAzuAq6KRcnwZYdIMPRyAmKqVe5xaGzCE1Nh5xXtKJODB8NX1h6Xw9/N392lVBPdNvbhkt
b7Mjej1ww9kg0uOlulTXD9Uq+OdFS0XBaltgmq2mibjdRuM4ZDcyXJo9gmnj7eNGt+m8hJabLXPx
fWlGMM1YKEURQDx+SnHPG56zoo40/LDhIk7s8S8X8snTK+Yc+CMttK/01WmaJf5Xp9LJ0b0cL+sf
l6y515BD+2wruRo3rlaPYFQaoMoxoGFoFLQytqJCn1QzNFSWaK5u2Bc/F5PP4f8+cBhaRaPjC+C8
lRNpqZJXA2mtB9ELgHFJYBE3nhxf5nFkLf3ke+UZovapfNRdgy6OvgYypw+PEuiHH4C6O3rnbZuN
bDR/r8LCuZUZYN8j9qv1lAaPab+RzCYG/Pe0neUCm8IHLH3cks00UkaSe63vIAt+6TvsCk98nlLT
c6M1v1koeeVxM5X/nkBJikZXT21SHhaIuVDrZygfDVZfz+0rICo1ARNgIlCkArz/7i3mLSplZYRg
rSy3pg7xZiCvGaHtBPcNHzx409xV2VDxOBGiqwV3zv2bG7ArqywQtaGMLdHLjjOgKXDaPw5LYwxQ
a4MIkThqFdqk7rRnYDpGfWuu/9TKAPBAuCc+KuvHfpvAF1Wjn1nU2QyeeS9N9NuT0/k2rnZg1Eax
9We/UiR0hf682B3Y31g/f1kdR//PIjsCy2fjsgdZg236nD3A0WubwgVkNPQNX11DzGhUZjswQ4kA
ryro+/AeCDCB8GUbphZwwUnEmZWt3n2oDXyaalzADcuMtg+BHc5GKWv9Ofp9fkxO65TV+Csksxr5
ltAhV0PLe0SW6dueO5iI7tGlSDQ+T7hKkTETZeHDtNO8CmtCOhEw7YYHD/RTG3goUiTDY5GY0T40
js3U86NKHvZ+sgc/qtf21mIBzSsxiErb/rSYhOgYiQVAbxmMspaZO6Di4mqCs/v+Y5w6YkUqP5eF
17ESdEoyvk+0s/sMed8b7/Sbqqq9qxArmRHEU2Ks2Xd4Y3GJaAAcr/fox1b/FdisoSg6n7XwmNjx
3MW3N6DekT/oftyVNHmGZDmWC2b4lJPbJpov9esMh/tGb5IUyQJ/Tv/KumX/kdCA9rGbYcDaoll0
5RU6XW20FyTbAbH2nM5iTSPVOnyuWxrh98fNYVOnnlflvpUib8ea7eXZwgn+mcH9k40oJJGooofi
AyANQvbyRfvu7ik8GT3pWh6yT0GVHGODR8XvhftcLtq4s7Ju+hZjszCM4stYYpgw/F9neEumlXQ6
zw+SO8qUd+aGj12T4Wut/YLGRL202FswwkW8ZMJPNZ7bDBu0+NCJcPgTUpNbUJVP6LA6JWEEkIZ3
8HjjdbRsKcFNm73/5DqHrHBMV7qQDuJT9v4vsqNtiivltdYAdxgzHFDU8THmY9alpYrCw55isfV/
aIP6GShDGBNDs0Y0nJb4PIoq1TORxlADLXNV15KnbQ/2c8aMZ6UjOVm6EvvQvEE7wkG6hV3osYYb
cZ0xJcPc35oai5F3wc/3KzYTbEdPMttmEvbb6OaGGAETnOc14BoKLfRpwJTekiulcDQ0BpWUmD6K
Xkk9A+lcGyk/7jJoreP4oy0qOx+Uk/zHyqW7EfKLyWKmzSfg9oLP15NmB7EtGJuIrVzA0t2f5hq7
BFvv07TVDX0M6ayB4ECuNz5+JbyWOPUHwLkKDyDEiVcIrYryii4Y25UwH85NFXndUG/5j6p7CTmL
IJPmAyhs5h6wUqhOC2Ra5+WMlBkdkuufBEvfxzDtL8jHVcZIik4VU9CoYPAeAwZjqP8YMIumKUe8
+cZqTyMq7xJ4/ThD1en/Ssiq4C2/hEKMbKAFHpnDKTdVa0pVvAXg07s4U06YswXgg8gsHwHZrOFj
bUEJnTutLm5MQ3R72v04pwn1tRZC9xecnSnOFv3ST/dheOVWElqALhY6m+kxtzLJjzN/6XcWc451
F1aIkZaCtGA5vWUdfok+oHRvGkPOIB3MssuQ+lhbpWsGMBhK6SGAbv766U7bpy7KrXF3uG4WuJJ4
4pq07yh3h0yIFpTgbdvzGb4Wi9Ov6UU+ulwjQBpRPRYG/9G945thtjYmFhuxNEg82+VPvCYId+mR
afxiduViE+vLVo3PBpLKeMRPEd13wmwEMCBPA+mlf2eAvnNJYJe+FhcGcLd5QQZTXnriH66WqO8k
uxgNtOHjIAYtHhDa5s1j8jihuG6pWjKFPa6aIb5G1QXhL/7Dx/Ke7OnqOI3m266ABd2jP2Z0rc1B
iUVIAnJPtZR1RBhTp0PRG87ncsWl8RWRPL9ERyMKwlE78WJtVZEk5S/D0PIcZsyvLedjoDrvxX+g
n+Ht6igvmOzAAKksqV6L4shsq/gcM7CfV5A9Lm5BGH9wa1H0VMm/CGiz4AwqOyhtM8rZSZvWSWhm
2O7EqKBHFLFSixCEBBI07vS716nASUM49RYjB+7IniJFKC3SNMl/C7hnGMYR5e9YuTJwSloQmKA1
XRZnHkD9h8NbrB42pGPts5Zh063Lp8pUYKnspProrqV6iTKyLqlbnwENaytvaeoLk60LWWtEEMki
ZXnfPxyN6dAMKi95x6gp7XL8nc2ndFoZ5G1Pi7CG64mDxeVwrVXD2fhF7cVqLG8dc2HdL5o9OF3h
Fr/pp8pXC4cVaPFEu8w5uMxlucV9P+btU+/CBi2SvPP5Bs0yrmtDC35uI/FRISloT5K/ZmoKxj0L
RFkuSuLPPguFO5tG0qXE2kQBybMrbMNH5WPXx0Pdh1PStew5oCNBhrUQCWBCjHdlz6WIqNu04AJt
f0wlp4CDVAYvapoFE/EEgiwo+s0P98DWpF2zUfvF3nV1qAIYpVKYGE6DEhjaJ/aWMdqY9B6BVCLV
5y/fpDlp1NeisEiT5t2xvGif5jhY26j7DW/njiOAtXET01PvSwL6sHr/EPutKv1SFv+JufEKkvr8
wGUVMHpuneqPuw1b/S6GlcA1QFy8SLRro4O5nd1/HTqZ1m1/D3e0EN84u06o06Sswg+CR3n5wyw7
dj929Oe7catAedxejt74EJK49+raKLE0DAmYM2JefGNyoajRzv9V7J23JvQzcgvcgZLS+/pifLz8
Pgd3QzHOioBV+VxZlMYqfZ8dgfOrSU3BYl6wxB0smQPpaSI8W/reLM3sAUNQCw9R/GnPVtTTw1HH
aaNqPGB2KoZuEPmhVzOXZbeg9E82Ox/zyTRqyQGuO4nlT03Er9SeCnvRvUjr/lAlaSXFG2osbtQL
T/IH9piua2ONqm7Yxvt1TTwv7AQNssD5Wrc+QPhMZhs36jHJ6/5ZZsM7+6v1kllRA+97YPN8ThVe
4iC3cGEJzjnHrQWdwnAdP2V+98ft+WuvF8B0bvGsXuLiOHY/KxGkGaObrQPSXJTA3/xYBuKHsm0U
RYdiORkZhoVZ73J+2puIlAAL/a59xk09ZyDMcEPyoyyJsK1bvEfDnSKm0T3r7nNYt0PpZx5RGh9M
dqY2evZqNicvkXXzfnByFWVkjrBc+zUT6e2Y5KkA2D4l7GS12rvbY4KW2u0sngWgvMSM8HU1mtIH
JgdxzmgqExPBlf1T1XnhLzCLMVrvPY2mWeuiu0f7u6WSqrR/r2nJ8nqvB5MPN8lwejq1js4p0+Eh
CSLuvQfZqfSPkPTPjM5iEtSiR7bCsmABVHFa+ZIYgxZj4VdOujo8Bqy05gBVgbbG/pe1OfzrRTL4
VKGa5YCeBLcge7kN3nH3ml6oZoee4rM8nzE5kAzDrSByCknhgCwGzMakZUpLPrOIJ6nsUbL/8Lwv
5neJxjl2eOrGyaw5HHkfoOj7WGYP3Kiwtpe6M3OA0SMB0SSfg3yPdSe4xM3C3CjP2DNOmN+FuMj8
cLGp8TW/znv/fAKTk0UooYiwTwYdSh40/4xwTuAY+JHRPgYNahjZArFMDFyf0YAYzySy4JDCKFN1
7Mg2+hNpnkNXjyK2NkIiVPQF6tlQxS6AUvGwZpDaFUFEO/RgFuJfYwan7iM5IcUW+RvSYTq85s4D
PFr8TWOcXp6RuUP02TEJUY5t4GXWzzpSQyf8fzkxnwQ4IrSg/XNZQF2YR1Rj+7QmQ5QK2wqwIlTN
TRUBb987JmqBkrhz6tcNTjax+ekpjk4SCYch8EZv6tnEtgs8FcBrBdGlb8fcKvMwdtES+d+us8PF
lh5d1ycu/QAKz0c/GDxHC/jQsdcNSeCnMuPvXaIAof8fTyOuzq+FejdZVeYEfouHl7Pn2nc8avAH
dc7BED6U2DL4YIm0aQCYMSNU4K5XbaXBDOSJseA/3wzHARNakL7AsRFEbAgR2WkIHhU5pkh/+H5J
NQDsh/v2Tiu87gtK6AcB8oSLAqQRrv1EBLhRfbqHgfdLCOuCtF6cqW9RQ89axYUnXiAqJOGcnHAl
xdIsvtm9yWD4qWjIWCnFQc0D96G7mJ44QEn8PzoBUIpCoRx2Q8KzyBkRaio6MoRK5WF3fWKrcCWp
eneohHBlAZHGWTFjAjwgqV3RR+wBORMUvyIFQ2bseVHKVpDb/4FDuCJcTBTdD2pmpXmnuAN4bIlU
uQVwLuupKjOJ35nxhTUCv0/A1JEOi6oAIq+OH9cVR72TlmzeDrBX/9SRhKQ0oh7usp+5j+zFsgfa
h87HKIdQKd4/FI86hCNhRdyl5/4mISFt2lRyhw8fv8Yz37RCoemkrIws24+aPLDo37TezxN/dKuf
EzPw+53cH2WfAG70x4wg8xOwRNAqPqpdOe2MrZQToukS/o5WQq2OKoZE/NVetwaNySCIvCiYcb6D
2x8excFw90lJ8daRgCpQWoO5FIAPql7T9vnlGr0JiARsgfji+IVK9ceHy1Zm2JKE+ukJKCiEEqXQ
Z4JOLiK1Szqa5PUg0meI6zLmLtAiqO6bAf6YW6clbRkUHZ6Aeyp026x7ZnLA00dA1p0aQm+7Jdoe
cEEVS4MGXG7nwP1K09mZOEqNmgaV1tKetmE/v01uXMgoore1nCQCpC+hn1CjvagYPvfOVJo6KafD
gj9p5CJFAasZWv8oIA9XNYdNJLiDU+pHpnNAxoA++lt84Cz3HwSphaKHM2Uw3fCSXcNuDwsfyoqn
qiugfjTZFeXEWLeWaal8Zjf0lpjXKX2g8aNtk2tfX+DSbD+uHvTGLVffJsZkcD1bynaiWlNbhdUb
LFdKoWKmhnXBEqg6ZoWHsSgYfh7i2SQufHW7Xakx8AHc7dk71w/MchzdU1uom2cvsRMKmKNVpo13
1hxOthwC/NiWvn8aszU3ySzvTa1vQJUjHxpch9tGFxKyz32w3Bq3G/qxFMlEfAxo/kYRdyAfm6qx
uRHbDcMkjr9ssxyHDvexWN963+pxa4LgtbNaz8rOPEB90q0yxGOBfa/urYskX2jPuYwKV7LFqEyJ
CVpyhAmP/ezWaEFktyV5UqUVszBRizWKc8e4qBaVXaf3c84fhAChOMcDqzCvBn53adPTRFqjd7VP
rJGkCK7+hrrOZaLAH+EoWUr5BxXvf/TRVSkrXWQAH9V0hFBgsOT7mz036+EcctW/2japZ3VnZJhp
rvT1vTN/L9zYxEkjFie3AAX8yb+87VxiE7m/b8w+H0cFgtYAwBum70qQs60FsGYeZh6UFEc+NfsB
rWyjx6826tQmz7s0TfQAoQNWXWgpWebKI0O3rxF/+PEr6x4xbRrrnRIT7v7it2b1UOqAboG7/BC4
AMbJF5ooW/mY2NFE8lOlJ1rykNU1zx0dvhxsCbR1KJ9MBuL7kQ58oD/IUa9J5JgEOxIHjP1BLKYK
U/4t9i/oWO3W1DR3hSJGkMj1HYzz0ynkb6Qpl/vpH7yijOgaAWayvJk60wGpEKn4KTNogp42qatx
BSBEdmOBi/uTiKu5bS5OK6tDOgC+aK1lgIe+da3udGoe0TUwld+r6RaFBCCvra3cu27QvBPhWTNN
k0kSN8k+m5JjOc/4cb6rJVq0S1SjdRZu9QtwiKJXJT655ohdvqutfPPD6fxef89p45zmwQua9bhu
f+C+ms7WQ0FnNl3W/rfbnzcXVrlq0u7ZD9GSAVTx6iqbpEzo72nSKumICC9ZRj7AewW4DrnkZwy4
N0YobTmrvL0eIIrgFh69YVZ7c+8QvcDIW4XYwuzr/ZsAKFtLHRJDP9xPf3wi8OdmiH248lqBEjio
Xh2K1l7hdHdfsTzEmzxtpm0lLaZ4bUEUcaasFVJDJyb3BnowWpPTREQI6UPisyG22EC9kJohaUMk
nlX1sYnh8cVh+QG6Jylq6qr3b23sQKxaD/VHDCbXNJejS36eXQjo3dZ7ijB1oqMlr3LF5hUr0LP8
cmTDCrooaApizHx+gTizzUucC9TmPrPfP4IndzJDVpfULu7ksmnsDB8d9jBf2SAHgbxm4MdZwB/v
+jIpaT/Py0WdZ+pex93PouWxHCjp+a5WpBtskSHO60jG0O6kaa3gnMGU/andkrhUr2jnfDW10HsI
kTZBdwQkFgMVOMdZwQDnOdnLxxAFhY7j7bNxdmwnsc9hImW0ZuehqlQdENNi03yoKl5lBSYGQ3eA
VY5c0fIp8Tdr48GFVKvuvCZ2M7BqGh9i8YPX/9TH60Khj7YswA90UatV8kEaz1YV0VTSMQjTRiqS
5RIpL+kzGQZgSkD9BQa3hWtZa2dBULolpO28MLLBrbkdifzJY5yMi9lZoUeXG3Isl2N3wD3nhxvQ
+dipgzdZkwDpFsQKshUxFF/k0JmIwXUKzZJQPjMB8mhwTrusbPUq+8Qn2nZoMO8jdHaBiYD9j23N
nRo42YRUK91RCVbscrq5y3J7hkd6ogZ/fbhoD6hrZBegkYcMTvF6gyln8Q+q+g7eKFx6TO0Mxxks
dleutCk4ADe/dnX/3NiMss83B4SuXAWak3j23FX6LNGRDmE1VgJmCBpM6/CPbLoKOhiVwNcc94Hn
ufCNrdeA2js14bgiDBVFXoz3Xh/VV0850I/vk6YyQkQ8Ay5mhyZJ9yJ1qaiZ4wo2KcsZL0J7qu5x
S8Tc8EtGvc05tIsLRnuKM07MH/zcklt1AeBAmTxhfIVxjCw6EU8Tq9UJ2Aabv7yKAjynm1UhOFre
K7vOg1rrwCXyildkv4kJOepuP2elAttXlmVYm4pak5DjBDsdvSA2yDsLtiv4gWRbEabF5KTZ6/kK
FbW+I/MitKoiYwUxp1PTWVqTMkxacHgveu/hm4jKaphV0avh8iNwxAjX/Oq/8ipVjzs4HJarP0Y3
NuUf+hP0LAttJK+U4AYq8Zny9QrSATpO8/pS4PKYtDhnh1iWar35mu6pDp5rAkVc3yUbGe6g/Qp6
PaTMqXKrOh7cgMSLOrBFj40/mTF7zQsY4vR2ggdqPf2PgCCt+SfXrfAfMNh/ZuNmEnHTAtn3bSvn
gbYGReSzMhlo4KY6l6edaNJ/ORDJivkYthWs7hLBJ5lrTvsY4cvlhMdzb2bGp/iX8V4YJ83nBELz
MfjZAuCN5BoAZsvmUMtOK2VQwW3dfaXk28Huq6Na4iVwufkvA8nJPaM1K73VDpHuTaZfwZrpGXub
2dsoZzRfmuGW+gRSadMLx4iUZsTBXnZkZFnz1WNV5OSWf7M8IblhuKHGPVP9lTmal7CF/gXF6Lxq
9CXIktES5xFnpo4hAnT3I11jzvZQueSLcCBTIW14GmNjEohu8PI5Nsbp5Nm/d1FgCb+Uewmbu+bf
YVYin2QdDxjVrF2K7J2fyBMghtG1sDlwG2r5MeLWMC8PkdFudzY2Sjjdx0PuBkzItY+avUakGfJx
apmoJoLA3FXa7QL+y1BT54vUDMTPAV40h0zEDgfPJ1e/Ueqtw/axWFYL982xuBWvfCg9HTh9lfYP
ekZHoEKC+Nf8Kydob7y/SFzGvxxmWwb4WDmRcMli8VCQCO7dgK31GKmR2My9yqjBs6Vf3a/kWo21
SZyLPbUKvWeeyADrnJ0c48WT9pfSmiZH/CSwMYschG20tEnDOuBN1FcsGh/uvZYprDgHqe8G0MGW
iHTwim47TXYkexwu2m8tNxVoCrMRV3fb41vuCAxRn0F3PSur1VGAzlz0vDKCFheN6TcRb3y979pw
LbL6lEAU2jv29Y6i/0cFgByOSa8RXl6sllYzhLntj31qJ9lwMj8kXISk2Aqj9CJ2yD25ZzRqRMYs
+ClAg7G9FL9fJLrszMpsy8C1gocsUnlavzpv1hMalqLP9WS/qBBVtdWsEQ17CwPE4ea9sRStHDdm
fwfvpffE1P/W5AELFo2wlI5L5j16rKEEyiaL2dVeGOVNUINZ51Wai+eOPOmkTTwGz3LcS2nRxzSV
ceH3wQALZk80SymUrWCeI18xn80JHubpWe9dtbJmiJVvM+MXfsMF5jI1h3CKzjKoNVY20rP9fd/H
4RVu7drl9EhuS8tI9d9QxgUeML3qVV6F6W6Kege2+tQ0cb9CpOuVtRwRQZ+tPhzG3NPtXt1f+wTG
fTpwumOD8oVJggcP6UtVLK6dbGZR3yxkIFHpX0txdo7lX6x17rbKFd5iYrneWfa8sOfALLugLYYB
WDAx5Q3itPxBy7yjFXNRRsEWahMBF8NRXl1Y0mRE1pIh3ttB6aori2kFS+jL3M6QPKo3t/n0du4p
kWdU0SoxkEBry0ugXFyijx5Gqc02CEtjvwvJo0pD0bLcCGGxxHT5oRGmqmdVxsaqlEZk/nE8pu8M
lP+JXCggYUGR++myv8k3e26zbkMGWezTQWX7Owp2RrpV/pBsbv6dyDFFBHTlpgLPiM10NdraG0B+
hmzNnvPFqJClSRxGud7ZUWk8QXHWf/4jV9fkvpn1w9eDTKDYy/dQpQf1P5mOCLlgOtTCmqHA4pKe
7PKkRRSBr8JreBbuP6ypx3QTJvZWumYndnvnqfSMn4pm3DHRGMYTZo9m1AlzqUPABlxeeEYAfo58
IclrEU/MrNKcvDPPD70gmGr0csdDUppUw0q6ODqbacxrdoc6Yp88nepxgtWWircqHPp0eWRnHujc
gqrQ295tKwoHyL1r4T7rajWAx/kEcjrLS6hzah2P+FxednzsbDOx4AW/ZKo5OMv8dh1VQ6u+Wtfx
QExlYaivm2QLwM0rWzGOc3RQUMJfAtaoBqpz4OHqM8c9mKrnuj5tZ06Z2f2L5SkUZ/G4vq50QPPl
BdNlV6/vP2GG1qJkoeSs7LYU3HpQjhuaXbmC/ltmKeLKRb360fZxiXCWCLKLdF5990LHQtb6FFwg
hc/rOj95958s4W1nmVMrO2RIe2hj1Mw0I5B6PPTmSDEtVoifjs4zblE69oUgsvyjxoyUedUVnrDQ
Bemx+GNaVvwqlpYRJ6ffzkH6d0tYQ9qGsJn1hh1sXgW7qtIXZbfQDovcxy0C+6w5LTT+0mj28aFQ
rfCE428WhvIPMN4yBQxbu/qeGDSfYGA06P6hFFGiXASi7GFu0WHMZoDEVO/nIYjxJXsZ0wku10KT
BZzeMqJVMvTwhr1frJmFBhpcThs7HRWwMri9y/6/VZ0RJyvI9Zh1bRXqHHaho9X5s612ADFo+rmK
BZ48ePnF98ktzS9bqWiFMSlBy87/bEmqjxHIjY7z7e8lhNvUHkjnhZNd8zbNkWYh9ArgwGBLeK6x
KpqwSRh+rLj+F2QPFm2cr4ltCxUO0Zgt5382oCcO0J0bp9GbgYmPCT7mKo0c2si9NgBftDmjFjvV
DNsVQx07x4ybUJSKVnLaMv4bpe9zNkDGr63XGczqcqebzUxc1DcAFQUm/RPSZHiVzJ+3L//NkQAP
f3caWNNc6iGTrKHzGB7GASSBl9u5OCezNx4lr8jot+lPGcA54eDDadC23Vgg1QKYn3ek1RoUNufB
FV/Y5Om7na8gKqipDj8C901npn6ha9Q1PuHd0PV6jKU9iMzV9dbQ73LB/fg7K152LDDEDgWqUSgF
anflqrI4Nzs9l6ofyptL1WLRuotGL4MxflQvF7z2BPjyps0ezAknGx1reqD/hu8SmuuMCsDEfITj
lMXSaR2CzqpXrPPETH2W1iS41aqmN2aplpzrVykG/Gz+XUd31Yomd1etnaZdhhMdqWqJudcY1Im4
kRdKM9Dz9627SP1LKVUwzz5XloRO7EzW36gXBhJS+LMMHqh8Vb5CIEWSulY5+2QIdHW4hIrDoGL0
wGMWi9latLi2z//jbPHbnipLQnU9MiYKeaFA9BFSJCghonP5EJowniMlLaf2HVJM4VV6AFeMAdRo
X4GeeHx7zit32NQQ6ozlKJHmORqZO8QyldknRuj5wF6iw2QHZ3Us3hwFYAF3blVululjZngpL/Up
ZBV5/nmVOvfeQondnyb1AvLAqk6+4o1j9dHQ3sO8877vB8FLx5N5ohp9r2WwGgK2Q/LTTeRQ/hUf
zM3U2Dt+guOjVr9XfJYTCc1Zxo4jFgeqfk5AfNF9D6whfrvRKfIKFk7imUHq1Yt1HuVVleCuK6L/
2nclFzeZmCP3vJCfhK8ku77H5aQtXVjoBEJGMxDzzBZAxHkdrhLg9thr1RBjkUO2Ddl1qH+W3hz+
bgGqJPPccU2YIwJNi6ZJz6qpd7DXdSxLzH8ozeoODvlmYAuQY0TvrXL+txIxOI+MwqTg+kTPhkEJ
nozVqZz3e44kH0a6gmr/C+YYkN/ocJtujlhVOiEOwEwtIsNutOfz17lhiBLG/BCL9xudAnicuNd7
V/j1QxtH9zcjEajbd8i4IDAIvMyCdoPPbaPnfR917gZHH3cWuU84fEwrC4zu9ESXAUi7+Rd4ciyP
67fri/IaxcVVFpi46PpQfbVwwD6KRU78oS+vHVV6dqolkIE9yuU9PyYe6bgjk4415W7Gd2iIZTY3
6qLgN4GF3IC1/9M1aAwid3DkVNw+YMmDejSsZPrc5AWKLRFwX1NTug1PpNRX8VWSPiwl+T/pJlGy
uEXA9flGjrbgtjHWRbg8OHFQPOvbYMw5gvmSnZIjYDKYIN1AISIktKDtTnNgl+DR22WSXCm98uNB
AtArWrZ8CMeLqc9MZBuvYgR3bH0gyOymeGQD98P8WCng2TxM1X48pMHX6fHVcIabTIu5iXEybFge
h59C0rI50dAZt3SJoUIG9drulHMBZv+ZtPrx1QPwhhHQom6G82/qrczlZPE/1c97XO4UlB5xltyx
rN577ndvup6hLb0Icj1tTlchKLBE0Iov3v5vDin26GQlATxz2pryrijJfvxw5dLNHiZpreC1mgGw
5FPVlJr92StFp44/s748R202hE6Mm0qike7IjnBYD51ZyRVLSsV0oBjyIgVFO7i4Kt8zOg37KAyL
i2H7xay7B85IAUa0sCvC8YEgp+xBs1v7EynpQQHIq4hfHQP5ToyUPBe1Q5RMT6oPoRuZbyIbHT7x
xKNOFlQ1tbG8kQBcb6VX3FvBs+OYpiC6cbqr1HXJEaJUEFGy5hrD9ZC1PL/J2eyETZ97ub9sixPE
B2uyE5z1JKaIDERjkYAsgkmpJeB+JYr03Fy/i2lTKr9z4Yj2m4pSPMHoA3o3s4feO9/2rmb/DShK
eVFo0MUl2GJbTWTP+KCuXwF6J3TjkUQcomgADH9sRtUMWUTxfbwl3JDEZS2lLKluwLiR616UN3Qe
2eXFI5FQDGSfyn3yhDvRcokL5cjd1Or2d3gGukZxiOYEopvts63xcmZoPCJNNRMNizqI9bHKGTgl
/H8T7zvN25wt/jfnvRXi87HgZSFrlVyJj2vD0+USynMk3tC55+p6N5U5sikUKsuOPzRinn3xQsT0
bfO1ZI2m/y4IyDkdogvPywtEDwCQTBxxfjPQ5VL7+iBNFd968ahXjbNqE4/q+/KTh3LQE0z1TjAP
Sshd563yk42puDSzi/Fyz41eMqhXLEqxUsyBjrQdv6jTBPq/BYBgSYGZHMZRE9AnegvZZ66F/qrd
LLmXaWs95FOmvqoLcuZcNf5py2Nhws2617bnXRqafYwEOF4irMmR051tHHzw4t0dZ2UX2yI6SWND
j2v+0DwY//gCXl7Sdv6IPTSFleY4pb28ZAwblX4oKMJZtlCBQnYCYD9uzMZAv6TAo4jZZVjNlOJM
yOl6YHwZU5G6gdE78s93npaDidxIwmhfIAOST1kKyRqhbMEyCDjg29oqJch0fBurSD8aoIs7n3oN
iCChyYp5Ig9LZR4vIUXx5tXACqcReExI9Xyt4ffuzyLows2UmxwxCp4fsAdjZX3RofNSjbUDbIxT
nZ7rtNkjrWbYu1Z+tb0mmtA0/+FBvtrgVGJ7RClz0ypHJvXXNXDH23eELl8bSqLP2whBCihhzjwD
TFmaeKXmfdjr4xBuet38YjIcq0wb00yoo3VPQ7knjdl1oUWvFKngV9U1lq8dEnXPFvN8JL0sHHyD
nnYaA4XcBfV+jI3tviRfcYrAHhnAVrEXOVr1yhwiLSSXHbqNfhCltRLZ/tmXeC+DVGcRTCp83ktf
E7Nc6/BTVze+X2xcVNdsDDpU82HGzHeCRroXMr24uXar466LtPgrh0Zjm4M9rDh8DTysMaTbwppB
QNZyw69x7vsCGnfMab6GF/b9xdLScGj72tSZcPpJpzu19urWIllmVlJS3MTbZU1X3vtA1vUpjPol
2ocMNgAe+lEWqQ6bZQJpIi7ooCm4lUyW66Wpcz9gfgKgOzKm5xlDFnmR3I3cmZXTaYWN3kciMrEn
x4yQ9JlOSZdkwmEFsADqCXhFx4nhWpzSm7FGEpVwGMCrMkadgQBqIGKsXASawvIp7Ak/zxQ2r7OU
TzYyeCnGS/zGtQTXF2TSGsBfBtytJQt6uZ78RTnQNM3w8uTi8ONXAUBNZAyDqjAvg3EdM4LnslXo
IHnWwQBBeo5TRBfF8QS19M4w9tWlpXKTc2h8sVkT04Xt6UsYyc6xxC+kHlcxq3jrsaH3YtHaq0Ny
9n9goEpl81U2HNd2mxOeC+YM9F92ACbHYoHfeMlMLSJrrTU+LvVhJSXv3ysnzeiGH1dtlvxZAyTR
vBBBcb2F+Wa93sr7doC63zRBgzN78hvai4LvID96zQsP3iy14yMXVYx14zjm67M90+uero+nDEHt
sPELGdJ4mnm8SMdiqg04f/s+s08T8lea1MQz4trEzlnGSgLGNyp6cl6YvtcYLhPu9niDI9h5fNDh
bD9qAaiHehdYPwrEQ8+/EhbsyLEotsq1ayLRtWYqz86CGqOwA1juGaEiv8XEucFqMi6gMOephuS0
CbfHZM+uQMeryd7LU7kG9q3Q/dgPskyeqR5RsBvLc5a8sNOpr/JikWSsCH/QuB+A886q14JSQzw2
Nqb53piR6lF2y0SVtRBN49BG5kcimzgdf9CGB7TBpXv2hINEzmDRmgZBG4MfvYFPUA7MoU5a3rap
3e0IUOu1s2Tn0lW4tJeIyNpq8QwWuHsUvR9hSoxPMYZks2o/yEW/Hln8Z+ZzMqsbmcaNrNqZ7fnr
XYdmGlVMA84NUxxJ9ZBjWSNpmJFmKzQC4mm1p08WAzQhqILCw+9GByScBwubHPpSrcFP6pv4KLPW
KdWtUczGnMDHAJhdgHubEML+MDY8HzOh4CKQdxjyC7NtE3K07ePf1E3XoBOcJW2SUSoD2Z6GaBYX
7uFkvPLqPksVJniBjtSG1QbOaosKcgSNDQLEcM6UGwEVIL1QCo/lVJS1K8JU6SH8HbASve1ZRAAy
TbsitdkWeba5Dqar0y/nICDILa+WDtMDVOncpoeSIDftbxQaqq6Nrw12/UR7mgxu865MsQXpXBMe
BJm5LFfebg4aF+ZOJqqvgNRdrcd6nhK32snZmEqu+EiazuKO3s4/nb/Fyo5Giy+2oY5bp2mnmRUk
ev006X5Qm3COWfQTfqBMrggZZ3cH4xvQIbF8wsJsnpQML+d2QfeqUphWnAWLcLjPuIIlgBXIXqDx
1HctYb9+iLuG9csSdKhVIjOwAcs/O059DW8L7Tl3mE2d2Dg781LT8i17AB+2yszn2emkEhLpb9EP
j81Ca8MkOp/WjKYBdR9N6N7L6mAoxa1GRz7swKFXRyhShIyLKBpl+Q16RYTU+yHUB1xFH5ikoH5d
npQEai1eVfV72sy6jYtTEm+1/50W9NERwMojEQ41vxOYg6uo1Flkp26DPZ5MFJr4+zdyGIqOUDle
QBe5jpmhvXN9MAq/uhvZYp7gAHHvruqOxoytTaIEfDhtGbXCgwHsMLoRmqxW06ZDVXXrk7Ifdme8
GCWguaGep1VtrMc2ifmDzp8qEO/8mHhuAG1/TZhATPVFH8Uo+EEoJZtS0Pm0Nlr7MqnKBcWUS51Y
4+PK2LF9wWINSRrK533qiGU06MQQJJ2EvY8F2PGtevVMusYg4HCW22ATkDxgR9WKr5UZyj+UnNSV
e2UFZ+HenogX6NJrldvMgqMlvrZmBnVLmf7Irtu8TcnEyJtBr4j5gAx8BOf7UPINQPe5vWTxMs/N
YCIXbuSXPUZh74LfkNJhkYngUmqQZAO2oFKIOT6G3T13WpjnFbwOCNJpp8+7B6TftQSny9PsHBxh
flVIvi6xuGdXzVJYSwDfMDYGUKx98Kzg6+RZF5kG07PcS1uZvrqeMXyZshlfuBb+tS2qJ1ckKSn5
BFl1ScP5nLCeNTHeeVcXFjt5szCFT2BE62Q4PtohEI6eWRq1LTpb2yTWZVY8lRu957o7Vhrddo9s
72FlJDck+m5ycb9SCS4O6qj39lxzWxvizVUpvmWoijSDxJNYR1P2Feyou2ohV+3PwuM+heI/szxK
BqH6CgtSJU24PY/0v2QdwCpiFezMkiJyLSF64LpFA1P/bOfesBtOFnlIhEU+tgP1FoNmlcocPRJP
VZfmi4K0G4/ML0CkbFMwKGfLJCDe8YTgCOVDmXh7OtrZIdEQU7Msu4S8t87QaYEOSZufg3+UkrtL
SEeHW6WBiq1O5Cyee3bXuLzoc+7KZ7zJsWjTlNYjKM4Rd+RZ8EhdCWIr/m7JayL4IzL/biDR3Imb
IvUzAqErDbwxbEaIc+yFHhasygIWvD+MiuBFs2/EMRZbAEEp9mg7mukEgYPnhdNv8K6D3KYGgMjl
VIl9ErOGw3bSHwRBTT1SXT0xmOrzAwBON6R9vviDMHP04kd1Ns6KKeN6MXgb0DRCeTUExTh4EUQw
JnrPXofuRc8XH5v9sL1KFNIpE2PS44g99Zr/+h8f8xRo9uTRfoDVl6K9KVJdD0FKFo0SmwUoxKiF
UHqs0iMOofpQefd9aY4QpF0bnj8InxjYcQn4Ns7KvLeOvvlzEG7JMet0FHVEsUfPNUnojhSSSoup
FHjJCHlQ4fLEvTnLchjZgXnLh01xppems+lU33UDCcMOaRgUveIK6RM58oCamUlOjBHnFnfKsxrW
waBl20k4yGaKpHOJlworoODAK0/VBX4B734R5CLzdOmyxbKnY4TJQr+HgPggCxgn1heXoUtmtDPA
KU+KpHkyA35onowB21X/l+UNnW2ulEnj+wSZcNzBNoRCKGe5pEg2pFyxrBJrKYL6dvY7mUabKWea
XDxJoW+m5V1y0kcVk//y7MtaIXpNDsu1iGchZ94bjlcP5PBkWY45JxuxRajT6LKLU3aV8zcZ6y9a
f9VaFdVfaPzPFG1UC7L+73HkLn08wwkyiQQoJG0aNPNPKrK1IZ68YreHbek3DXBPZVlMn9Yhnllq
k3xsTRVIVrHR1jMPdfcFHM2AZawFfhrPphP7pD3GpV7+psGLXsSlVr875BDlJdAnPaoSPNrVPj5X
oCzi1aA6cnV74xwn6Zu75soez8WCQiFk0JZ1Y9eQDl96VuPTLwAs7kfNBBQDTC+kK3ue2/Jfjjhm
wzYNfTVqq1N19eirt9Cg6igbDkbVgWOb+b3SeFf9TOStnrLkczCLVDJR0ce8oT5gcHLCSzOigNrw
HooyuqfHGx7qR3A/LY08NIUiEelLG35tmw7tvXeHG1f1qfVDgXK9HpkGnC3gAuC1KbXCdGEwS4BC
SLtj4TQRAfQNTEEh0cXe1GydUJt2ylAuUeTVgenWTPK14HWJl+bdjspVaSaMfnG7PMeRJZRnCK+k
3xLpVUXBryttJq4KBvqAHKPCfMruKAqZPHBn0seR9s6foyRgTQxjrh5yI2Dcki7dxVBZ8DI1JRgL
B5/YU1OCtv9sbeFy+dnvx9L4g/9n5ORKMrD0MNVyJ9ibTsGd3PJqbZa84apy7uY8L1TRCcTTBOI4
KexyWRKfxpESgHNvFKhKGlpPwM0u97GpEL0ii/mshbpute73OJdgwB5Hu6DiYjGnbbhOui8LzZsa
g8OLV9FklX3wxKOCNIlmNROCuIK3+tIbnB4OY78pNshFw1cGMV8mzi+/HpuFi6KAY0WpubFLmXnN
ciZ9Z9R9fSN5WaRzFXNQ73yCGpN/I3Lm5KzgQ6MG61F3mTMz1Iv5qXzyhiA/QffAHj+UdZpoTpzn
G49yT/Mz42o0yEfuEfd+NQPqmx5+o0PopfA9DvKx90aNPH1ljJPE858sfZxfRrl9NhMouLmJedA2
wZQd5pR7KZl0qpUuhnMOkUC4PupK+LFMxI0bpd+N3IgX2MC3OOPwmhT7QG2U+wjAgaHCQwKJ2QBh
yI8ynod1IYxN4jLOF7BYcnoVhJMCan2VSKDifDjVBDE9z2Ldk0DYv5s8enS4ZzxcMs0onRQ1kZxp
KxBS5OFm7cubyxBJQhMNklVBsvbrmX7U/k99DqeUkM8g75CrV9IYvOOSj0ZHPKl3qKfO6DrLnRQz
38Qrx/lSWE6BxOIqqOFM9UoxyW+mnYEMbnCff06lljtaOtXj0GbSjq2S0ROZ4pjKemRX1I145iLz
HxBXfegSASBUGPRxkhIZ0F/JZw4QhS1djtqb7oTVA9zVeUAeuQ5F3WD6J5cOLnQ9/t4MFlQGUIE2
nV/VLqY/YoTbmEeP28FUlLn6tJskzf1R9E2qr+FyzzkLxrkDUVp9EHZ/bErlN78Kzo/JmpfIiq4R
xFr0+H9yF6CSgg7Uv4B/OD2D7kffKyNQzD7prnfhoXblV8xoGS0hGu8sm3Jy+DI/K5gW7K5RWzni
thxAA7B1egltk24mgDmxHjeyQDrUGrZyZ4EGlv90e/h/NsLhJAxx91znqQSw7jF9GyOALNLmBWZz
zbpMRymP2v+4CvLSx8WFu9Bk+mIP4Ac1zmfKrxX6D/KnkOc2LaibU0Fpv6MStghRYZ5DHN0gDB6w
fKU9p8gcJot0pBwu6LX3gHipj2sjcrFiw3jGVpY7ZsJvCAMyOsVWDHQqDFNdt3IWn4E5CcrauUpq
uVaNcbwqZ2pIIN98kyDuGH5g9eXNAjCl35mseMftsuk50T9ISccqjUUIV8YzFhVfVYaG9VPM5ekX
/1RUL9UtKWrqAIajO0iGoxBYFGswRFDGm0qgnKwAtt7TOjDJIUUrzm8yQI5ssA8aE1edQUBoYuoD
Ng/+rsTeU05Ahyj0IfixHGrdA++anaqqEZ442CSWpvF0fosRFQiiBMlqcEAqh0n+KJHqFsvH+JWj
x785LH7/ymODz4/zUGjoOoHkMJlvYyAvKngB5Ak8vVLTBEEx+xbO9mlv45JYMbc65D68M0rn2mVx
iaPGXsglxr+A5QCHXeA4ktK5/MmwumB7qaEI3DfffbwLvN0xyPXx5+4qVDZoIuumplRWegHSNcOE
YWOsFp3PFZjlpVo2rD9H/RXq2WRGP0//jIAWYdTy6pLusd7dv8miDQXC3YZc6ptQ7c2hMN4V8aXP
J9zokh+FOA2/QBPseVuDOKZYvMl8AKNZuW48CWhPvHen0BkUcsMXtCb5SAMfjbr0f61vtWbRXm64
elu5noehC6zn/K4+tBKiOxei1kc2Voh6sjQG/LbYhkMd36IMJ2qJ/pgQZ+3oxmepHhbkgIHgpBcU
9ghh7QlXU27pXj+s9P8JORfPmw+negOW0vyrRFQAApSuJArmcALjC/jmDHLKA4EV9b/itcPXYWbf
XLaklYev0nMkMBw/6/Buv8Poya//7I0guXLbYS9GqjL8hoMcZDgZHc9XL3JW3kTKn7SegGiMz7G3
P4cEF2SIZDdigeyRaNw8F75sJruVxJLs9NprURm274a3tAkrF+lxrujaNhR/Fi9isDZu7ACQ4WPE
AgR8cuUTAKl4E8rcoR0SGan4boOsMmtKGfxU4QTtnyRnfVBotFg+Dz9hJzHkiTWaHXgunoIKd6UA
Rlr2RzR5YflZFC3HsZ8+FJLeCsj97X7pH7aJA606NzBg3hDHvi9x85A2jbxQEpaB+iEPXyB8Pzmi
OjDny318rtxzPqvqYnMJwyVvvia5F5Lg7DoWdJIAn/GOGtjTPfHwpfqQY6NdvFUswOW6MHBZF/Ld
6ZZL3KRfr77o/40viNorCaNg5IB4tJ3zULefp5OK+0P03qraX0Nn1D3QXi+rWmYvscjS0lNR5OT0
ULMyjBx/38u+1zwLXLtnENQzBIxK7p+0ZddGe0gPuzEhqv6RVtIX3tzYyA/rNjxGptM0FXmixavh
M6sEjpFtZEkJzVSnsniWGauEIwES91bIqKNsDeciXIBYVI0VuLL3UvQ1vQ7qa0qlD/nX7G/bvs0G
azD52azMPxVLhm005vX2D/HyrZEjzjBAF5bCRp3lcr+KecLpWd9x1CZ9noQciaBDNsw1m3vp9a+5
k1xwk1jdjS2tU8DP6IWFq3wklSaboquf9xMzORA/VrhmJeoKoqq/WeRIbyzwoUCwneCemjWUlQ0R
OG+bHNPWK2mHfoH892muLiiWl3GG1T7EmYzp5RlgoQgXF19tWpiTgasYyNbcwqeOn5dmUfSvyTiv
HuPY7PpCp48L+amqPLbqLsoOCPD01hKaxn4n4LleDh434R5b9hZzPCz03CVt+uTl79i3IutRc7Bk
SB5VcDBLmij89qVtg2gVFojeVRtYvtpe3M9hamicFNgohBsifEMlCP7pvjXMJrLgaLuVTIkeYm1G
bGJ0lDwzlra7AuOy88ZAPhMsXAPYUMTxkRpyb+SALRDXCYFKtdAbecnsmba4lteOT6RPTXs/2LIl
t1/+gSVXDqmVZXKec0XKvRl62OP75AMc//9vaA7Epn3v30BLi6XxjlRs5+iHgtAB3qMeVliYw102
yNia/Tb6IcU++ySSVCqRffxsykuCZ6g2a/TjL8QAAxq9eZPTdX7rcvFdyiZgeghtUjY7adusuu4R
ooRWm6dNH8wzTCWxhMvRB09WMLzLyFk3W/FN5sCjgtSx782EfqCJVv7+6a3ahgK5qpgoNOiPPcui
N3AzyzqTAgc94WeBkQaoRzSXU6HS+jCH9LQCpfDFMnrXO8+VIyiQWcbX9Hz698nDfp/YEu1BQ+Du
+WY5+2yPvwfLj6lHCskcH60B/naM3IDZJcUVNPXHF/mXpRqzlEQ1tTm4EMxyvm2HDZP8yEeHS0Bz
ACvlG2RoifT5eLIE14tjjXD56ZswG0RtwRwdOnb60yah8ukniNE71DsvpLXnuu/MEMZh0FSNBfuz
tsYgCWpSmum0/GtRdVk24pEHl9eMoFr5ZGsP2tUWLggNBFr1qi+k+UqADI9HRt7Aw9CwjJnPHN9k
Ah4aXnxjjTW0baKYhCvsoHteeQB50+s0mw/IT7oBeksdayr+g9SZvEnhrqQdLY+0n6RzwHXaFqcN
i/3jOHZbbgGjV8Xs8VYfocRC5+2IqmwRS3T6B08h9+Emp0duC1OyyvaKRyXl5mdfttOhhcanbJdG
13E4ojGO3KR8WCJa2YPsaBmKWxusdETr3ntVvHfj0L2pT7K78dSmBzIqRjAdfuGGfwsdGDkILc7V
Es9yAu66KO/hOBMlNynd1ecnin8Ig/Cu7Zge9z5PNPn9ZLkbc8HlJT3p/H+7sOTjqGbEe4RUPeAB
vd0n778htv42F8TeF8flv8vmUDM2mAb4xrufJzehs9mGbIxjn2COd/AVItf9O6bYRyPOy9NmYRkt
2H2nfOoHRtWyZU24FqSAUaKkqO3azGuI8vDjn4ZeMBNU2/3n1+7bbz+QnGR/+GvOVLjMKmM6OTwi
EbGU99m1pESV+FKMIzcFpVESvHb3yPA3CpNhfvlXxdgSnDEXGLPWZtCkZvIl9Pm9NKDLH++c8ksZ
/a6QCB6NoGVJu0DLpzFy7MSQQWxuWZKdwzMkyqqbKXSF1rs/LDueh3p4G8Mt25027CrR8bTDBllf
scCr3ZsOzqGXdN2/x0TkiDUk6C9FKH8Y2JhhEKrex3ia3bivXjT74K83lTSuzBWY1JDxSPqyhDSH
HzkM6lZ7G7Yr/Gir2Q9Kgi6KSLe55Yn6L5Yhj6DniBHKeY23HEw7hx4QwoDM2Y1iqp+mSV1EbXY5
4t3O/6ATGwTlX42uTved3BL1JE6gIA7Q4ATklGJJqqBUjN4Qvf9TuF5UzJysaH3k+q/o+55U2cEv
0Eqe+qsG19BVvRyCQmEalSrI25kccssJ+l69hROiePZSE+86dh4rXUl7GHY4MxfoKKfX6M578Im9
YnDfO6R3l8PNy6n0y8zkZ0D+7W2XXB7I6xALjQASRO2KCwuGuq6iPUeZzeP1Qm8cpFBtylCh6tKT
AwQANThgwiEdEQ1dq65cSY25zrtKLz78hVR7PV3XtmfwmrLzHjd4bBE5potPiAQqmBXQERRppY47
pvSwYHPeiVVaqtKkb/0TBd6FrERagBGfkoK7JIBeNNQokiwQudTjQnpkjjbFSZid6H8yzVVhe1Zg
C7FaX/B2lJ/P8DstJlStMF5Q6DQ1IyK7A6G0zF2RIvjPWWJaDD6dceY/azJlI49dwbVdMEcypzgY
EPckZLC+VtcLM/CmCYlhQWd9Y2MMC3oLR77RR0R0Ou7YLy/l239+0xFFoO4gShAcpfPAafXefjZ4
6cJXIRsd9QKy9aJ2sxjfIAk2INuPXTyZyHebQC81hKkdEu9MD23CzaomnctRnskzvKCzEMSkOAX8
kzubaohHfmD3skpdXhB11mqUiVhXZAV7ccgoU7+C6rn6XfQ3Q31ir48/Agp3WcOTY0B/4GoHOHAk
EWp/DHm2gbI88BCe6iSKlNUSdoJCI0IFYC3mU+tt0heccQpK/1zRsjlWL6qKLU9o9USsUfycmPmf
jvpgZa8XTDNJNWWivzSh38TkBOUUEY8wP2IqpbbUKmCkT5B+B/GLP6u9qIozR92YEBrc7rfuvZ++
uEliZFGjMJN7mpjXbWCA9WVEh0XXI9NG9KcpKN+G0Ex7/YMAu2PnABB1EnRvqAkQ3aT85Ehzkwgs
ih1YM7TToiqz1AZAHhRa8mobWy1nQ/fhmoTDgtmT3IEVZtPya/N9biAkrIgBRatyvTPD6SBOSUPx
LCCjhmmpzHckf9gPyLU7y0oeRTyNzvP3QO8FUrlo2EFAZMI6EpggGqVWjOAV6LV6cqlIQdwkfRZx
MmCb7kglsbDcJR0An1vwy+dxxXVmZy2XG+MW+I11IQCs1mF2kxEVRuCxZtahBxseeLOo06YphfJE
61ZkmvOdDSTUPRn6hm/EmtUBVGyfv6LRc7ARZAm3b1LIE/StnZjpWkrjThhCNdLJRCur5oldCp09
AiECKuSKMIjkt5eOL9z73mLQTDBiDHhVx2bFyUvbHsPRVxpQ4Y6fVxFu/9ZZ0IaKcbQm4PW/hmBe
Q5A2HbWtQ5HlpUPwyIFyr9GH4vSr2tN/ZKRHDxOKeNH1FLTDx0kg5xxTzz71EWRMrB4jvUbXoooe
s028CeWUBlE19IvG+1joKdhKBpZow83XiGaXdb1NmcCzDy5PwnKFQV9um0eCTt+F/61dVH7woWNe
QL8jqWopV0s9nRogcoYmKKKNLJAQy1WwP9Ctre0ihbYYYaOwsZbaTejq3UTjlbWZUEfUtVfpQ1i3
sWqDYkeQylCNPcV/9I/4puGyXWxVbD0L3ihdWYQkKPyBxGLN6kz4q6sksN7Yljxpo5tApVnZdeyv
jJeQ6jpbSnPnDv8IfUj1phhSyy+EjRDGeZkNIM/dklw9eMpagOReNZRZ+vqdtTQmhCJt6odvkAVY
vDA5G129b+TWgizuaufsD/n2IpQ7+ymGjx92ZbvVEcASU3BOLyvZcvqSgwLWBR9eqMu1YRB8rbqY
Kf6MNuYPJ1B32eji9+WABldPqcjBcYjf32IdgTACUgSgnWI9ZWCOnXxxEzJ3DdAGnPBQe17EkPQm
qxDNgSsU/i9NqSjrUkvERO4J0CTpg8R7hPZ/h8qg024o4XsEH9z5YV2EEB1eLDwiyrbGcFfpAsR1
kWtnuvZf6Hemgm8zKXIVgNYYck8TIJ13gob+3aAg1pbPffXMZSZBska4rg9vqr4e4TU7qy7Vfs9X
tk/wfy9M57lXUJSs8qDWqkifRWhFB9pgeXjObD3TUzlQlqyj5kXlbbrD9FYeUbnZcam/nb3tOzYE
BACki1tXFcUjus0iRRvpgGOfjHFrcvFhaef1R17LuBoD5keYDgIDgbkPJCN1Ri4TG3g8uwSQW83U
FjcRbE7DoIjL/0FqG/33koHqjJVtYO79ep0m+5bSkvT/LoO/5tYnQ/w3YjQlzpEYu2oa1kzX7taq
vuGmFrtfOW0g9PnO3tIaVlwa7Y5Vx0NiHznZLeJHyfrOC5Q9Fpe6l8sI0udB+0vsMcqByqOfnqju
bD8d5mPzVzT+k6dCKRnpvPHL1y59NNn+hbdE5T6mfY0vWnw5rEavMJZ8mBLyNfqQbIdPAWiAhHVo
VURVhbK9EOaswAMd53WZ4Lp7XKAIhunLok8zalJOHAnT04KxFGgcVoYMw6GrhLep9uExFwGWoGh4
yODmFRlOVC3nbhLunPgDHfGk5Km1b57vBO3lGnOV8xC0r/2WKFZUfIx37JLeflgEn6K3bpbHvBR3
U+mPmvhHvEzCRN/16BD/zyN46szpUp7R4n6SSv32dnXam1PL+722CleZTo+4tTnUwxDgpgqDK+an
3Ra3s5UmeDxbQih8S8ehFPl8gRn6/MhQuIebfg993vpMZTxMQ/UXmOkwyvD6SgCMqjutbg5VEnKC
VJFloK4eoQ9E+WLntOOtqj3YZ3oD9yKzVbkPxVxmPyULXC5OuJUtqJotWNVEQSmR3BPZVofY2lI8
GT3xwvZoJBSEzuxHdxUFfAei5pEJOUp7f9Nxx8dPSPjIV8d5xcIBv6eoSnlqN0WKummqBy1Vpq64
y6MlTt61I4MzAwl1F8y9bjLlR8CmbfEDuxFEEdLZxBTzGg4yWV7KCF8EW0SLMTukggZvYr5Gk+2I
Fqo3Bg49WhyyPAI20COOKXcWNEhxLvuU2u/FAeewKvj3AmOHD2HdDo4s/FyaLRulpTtnb0XcrWe7
xA7fHXfA/D2M+Bnp7y7Z6meVybHBxPq03lvZm4LDYMAkMc4z2rI1ZUXRafAyFgPAGg3dsYQ19/LX
YPF4um/9ilx7Vdxc9lPmD8vyhknAGXukLAXi2j2/dlGKmb0UvqiW+hhl/LRO97WMQ+MhYDn/UsUl
oau1arLAs6xSUqNLoasRKqWs/GkWIvMu3mzeAGoGXdtvDO0O3Yzd0ekJm3aJYwKvAYcxfz+7aiff
9diEHwcuAx03XmcmlE7ZXocdn3UIy9Eai8ScNOMGx74JsM/XIT0uQ27X7G9fzHybjdW7G1g7dwrx
ELuhr4Gfz7HS0QPc+GEVVrGwTZQda3zBlmaY24H90cHEIKar++ieD3rXTxDzlhCkT8XC1QUk/0jF
+h7IP1AvQeTO8hSKSVG+iCkW0NfMqMsIHqnPfCRp++MyY9ponSRRs4vnOvcpIRIkjmxBx4k8ad3q
We5uohtmewCJSF0CGkI0lsPrTDsjwh8MQ2P2Nq8W0QxJwiCe8GaRzr4Ud3XCh+nGovgQShvpaTur
Uvey0jswI6vct1tSwIYvD3+OXOCsHEfb8v2tlTD3xnbZ0rpI+oF58rRXcYlSIFZ67Nd4pd6tWWuY
RhlyrlRv7HrPJ+vffKjZ4T7bWnIqpYwE6YLaaLq/L4NIkxSUYVYlS3QCmpHpnWXpHMXVsEkNkdyX
GBCmfxZ4UhCEFbtUsuBhgTwfQ0EHJAySZd/ghx3qal8+49/2ygoS2oIwnJJlMARwBOqfT6WfeIw9
t0R4oN9X7dOgW8iKsdsEc4PAbNI3Al30Z/iV9ukIYqSlHrXRrUDaBroqSKDJOJuru8ZxP2KDoYsu
NGNCGfUnANV5DVv1jPBfX8f9MJ9E6TLjc4j+L4PosRkIlJmW6/QN6PogafLofa9LOGIEzVUsuqw2
F/gSoVywDgwKniOfvrW872MLHtlOeU2pmBlWYD7XNphpSPyPrOyA3rXsTp6ITTdvI/E2V0wgCx3l
1Q+wEbPg9OELu2BGa7KZynSgyMSorymDKTVNYljKMPSIx5O8Vqp9uKNGfGPARbfPXlwCS5E9H/ZD
jWnXzdlQ4CGCsbiZUiRAdk+Lu1impyTsoym6kWPCRZFWEhjAXX03HaKMbFpyl2UXMzduUkooitr7
9NYcjym/43btMq34rEyv8XTLJs+pePMzpmVC3T9I4Qvhd1wb1ktVN29dbG7AexYMRtEyAavrZ6hZ
VIt7NjliFKMR92+GunsyMIIqFpPFlFdl+xlYGgYl9Mww6Uu0SpYoE/fAw+H76ZJlMbZbjOlmlba9
fetK3cdFXL3BWSYXBbZHsq0alqnfHkrf63OrRlBRNELttPUo1yd+aSXT1XvTlNcIZFsm9TyvMqPD
F4slpLPHtQAkj1DmqV8nJFFe7MDTa/2onskFhL8HGS6sFgQjknVc8SdWtXvYC77EM1YGfn5SFSgk
9Ukm0UpvHTXqog8xDRFV0UCdvTkvWfVxG/NrhFmylAJWKFTIwgGyIwKjGEhTBXZA9tLuGHisSHKx
I4wD6WQKCkaor8WBR9T5Bs7SyToD9HrCgofI75jPSjql86GJ1YLUbf4gZEuphHagzyBGxB3oBJFE
IFd9i1MbkQC0UZlUDIPknu83ZxP7dCjWgBMsPd7APJ1Yjp6HbvygHsWCoUs9PXtZw+kNOiB65Ayl
ujCSdLh9puM4FQt3OLea+O5+K9lGzcHtdJSyQ26JNTedepx++mv/cR3tXSeh1izN2JMoB3PbNRKN
N+r0iXw2q8njDxEWnjfGGa5hjSQ6xtZ3g22fWtohGpcT94xSKPSJELMif3jJM0Pn2pKj0ZiqOCHV
zuhQvXkzebRkV1fqqeiZbP70MBuPjWTJpTafcxJ4KHinPQruvuL6TXqsBQ8gcfS0pJ0nSzbq13NV
/uzyAJYTNOGxrhZDo32egA6w545D8Di/LO0ALrae5MtN7dnm857mrjLoVlGrIW61FicZ40usstLB
To7j5SnOk4bp2J+UGMrqWsq6f6mV8jB0GqW7x5vi6n63Zv+Aa35dvMpt6uwWEaWFlP/oCBL6clac
0w8gK5nOAxiqc6pCMd00BYyGWu3TI9UuyKF60q1Q1aeZYexwvPykpFEhdJL4jJsNzTM7vYJur+Lu
6Wklxz6wDQfTmOp/g/IR5rUl2CeJfBeF6AbwT8PUfYVaqEoaf4X1y0Yxnok5ls14m3jhfsPsGrcK
8IHZZMsEiDN4xc9Hxcrm5lhY2wD56+MAt/HJnaus2DRGjZLwDGLfpfHzOGGiNTMf3P0sdh9g/fOA
YIXyDgJ993N9iDOmWma+w5JA34vfgdlHOJ8YWokJqOqVOsg7gd+LPZTM1jJhIz32WhE5r1pZmv30
DxW1K2HgxAI5qHjSaisT71qqyQm+YAGPs02jtCRqtrNXq0OEg9aizMZARloy9H8zsgBylByXelBj
QdvBuvO63v9UagR3txykow277VBcsMeZhoHAzMcvnHRtPHL++zCspYyyrIigiWmT3rLJF/54FIG1
dsur+COV4ekP2Wdx4/dSwllLGUnKXKbHu9iW+r4ZUW/yMQSs2YCJDu0BIHAWalRjKSzdLOQRLkgZ
Cb2a7dRS37iUmZfG9VFFL8GJbKLFBK6MWklvWLCwKpERixWPUtlyzNFsw7sEaEyfg1GJDXYREA5S
nYoTcw9xWz14X99qL2dQIa1Jp0RsjE9TbJ3cvTEzrFLZyebWsY4pBCi3vAeNTAPRQWsBl388r3hC
nqM9sSDq8/3gxui8Clf4atsSHT2U8Vqcfr3oTHcXkhAzImq/JtFB6xMe8WehyXcLeaP6SJNue5nm
x8nv9/BhK5jgmiGVwXXyMEkFXR3H5svoF1G8JjolzxxRQSpQEulJP/fSYnKdqdzx35YT3Ze2d/BO
TdGDZBVytefbOQLXYtFbUXBd/gy4BGD/sCZJprF+9BiMasWoRKubDNeiirvSvVHIyffWcAPzadYe
mlGAz1GiqIEjbY6RR4ddPHqCk4TaeJScRS8VBoJ8FY419BMhQhOgz9G6BObYIcCif5alJQ9T1YNy
9wqHnoc79Zfy/Vvmp1tj30Vv8Y8Yn3VyexOn6FnPvlGznwIdy5OzZrdLJisAKEQMETnGrv+cEBoY
9GiQL651XRe9jbmjmsam3eJXGA0/ZXpiZZHgBMwIO2/dwrl0UVkNTtdAZ/oPeBZ5EgWY7m3tDuFH
+jOs8XIIFHv0r39GojiLVG1mSFC+uEe/uAx8HIhUBH1FS2Tq7/GvPNFcI8OFBhkjZui6I/m7WGsX
yB/5p6CfTy7Lfib/Xl/t/Jha/7RtLkyjoaXRh5+kohw3NIEaJZVsN+mfg+h+0OC8KXPC1oozHwxz
YIGmdRwQjzczTfSBvOKDvhw+rrJ0kFkDCeizn0wf5nsRtOe2JHTRtNZh5u2gYRR6hiZCRMG5F9of
DQD3h7P971gkCLZDil9omRcWs6QSuVvb/grzt0J9W5fBRbLov3gATALzxJaLFoaqrwVwldP6B//5
4/8nXE3xwrERhy7bI9dVF3D4z0RAmSyzRYqpCVi+LnnoHPSK2qQzlnVInNzUWQUmyyOWhfYtI2Cz
fJvdQkK5UeyJMhNcBm2oZWynXYpnz9gi4zD9hoz5VlO+v6P3XGiYBmWeBZtAyKJLJ5Z8DQdoZrUS
FL+1+43Pj6CUl0Aq7BE3TWEL8ExhjuHdaosW7F3AVYc7xaZq3Iz4QuQw72XmbFcCHLjxuMjGeMFw
qrES0aftJEjUg2AdjVyKMu5Rg9z8zG72wfovD0excdL3Vlv8oRYa8rwBmVTYTYDqJAUyMqqOP0YC
BvvRLzJYphJLKndcw69B2CQ5mK+boxLAtByXpwU9sRKdONfph5FlGqQ5t4TR/zvGFJgRAOsL9QFE
574V7uNZSAuTXkTP8QrkVOqT/5DUaMFgGg6Fqlntm/eebDf+UuwH2yyfEHHS97JhYGD9WTeBgkYf
zWGwcMfws6ox66xh+QMDU+sdUeZCTM9tO0Mu3n5kxm6H3kR9ujmG5UUrGnYXnKsVDbHqMl6TPxuA
++ODmXHTz1fHJrmlxQhkLVPTYimU9bWTsmZGuaEhT68wwcIlxgXUalKrVAiwuviDt0A7dZzH4b/z
0QmkfjV5oRkPPbc8pCjs4DvsWmrhjyJRy/1iOcdHBJo6fRN9cGWrtLhHvBMC62XAZTm9f+t6MhsP
ls3NnRSDMEnl/ViMDFJEMg0HMu2daDaKQZtdCRbW8ZToNjdbIPXS3LvHYbM8KwLk2R+lvVYO0R2g
rvFTY+RfRmQUZZqWKR0YG4A+T/05vdwhIEfwvE7IkGCigI82K7nSG98yF3OCTBoIgcLzn41yuesG
5CxxtVUYYp5uYhbHD2kz3MX6XnXmHRJ851GC9gal54GVvzUbcG5O75/eUPgucr6tE1XjHddksPjs
9NNmbWT2jGRwNQF2/Zz9w9CbnVl/ob0/a8xSQXd+Bfzy1bPXIkNnQpmvZjuzrbZzl+9KVJgGjRmW
Us8AenczGYq9NQZhcj+WhncwiKdXiq6MyKshLn4vJ8vtfJhGn2G0RiznZjJ2Yn6PY5plxzlamusH
Ppz/+DuGhEcpT6XNhTYdZalhHOJ8sraoWffIEIzwVM5oaE0b2xLvcV/i6Me1IkdQu56wxboGoKO0
YKjPgIMuYL+hKdF9R5sV8UOxrJPkpx8g7fDTv9msQTnsOD6/siQ9pi/8YPLD+57s4H2F0qfyy6TN
e0PZEEkAThnFYfhyj1LhcAEAYQyr6WPBcXN79McPHChrq61X5ktGDQjmyT9zc+nzknk+TOrIM1hc
uv32/V3AK83OXNQu7d4rI3kOwjL3UNdNXv7cUUspym41ye+i55cOS+sjw+ayksPIFHgehi9pg3HM
Ckp08hqJBedUuDYRw6a2CVYZVL6yNA+IcGbqRka3i3YrxA5YYXCoIyM9YqqoRunh9wzUdZpSeeF6
/CC4E933U7r6VuehB0wTiKoHuAIC9pg1mj15QHudcbtSKBIpvdE4al3kHtQltl2l02iQt49E2C8T
6B2L4Fr6Ui4dVzRayJiC1CsmakAeBoD83kMOJ9HDUO6OOxUTNJECz52nuJ0GvX062fSZv5lkqSoZ
MbFqnDkX8QXShgis/lz22l73WYKdhzSy6DiIQK119N0fhLAhxizxv0sDTPCpn84DcV/zwQtf8ccz
xEDgXefS8S164/qWuvdgH8pVrcZVU8cRyI9QcTYAKZvktj9gv/KW8bhNHjnwD/G1olJAC490IszL
qbsjsYTKV1fC2zmiJyMei8lpqOCDzS0o1g2GNsJ3giPjTb5LVmoaj90XVzrzxD+maG/IK3Vddzsv
SaCLQJo+C6lKiq6KXkgMQiWz2sAVk3ge1+iK4wAyR8rd1RHghU14p/hT2eGUk2jKVHG40nzozKlz
uFwFRExEEiHIBbqEX9taqUM+NFQA/zWOxlMQkK1BiL2tZzNoYo0ORVh8zBkCYAUlO1SuQKxV0qyl
eLg+c2yINmeusXxEuDphCC+4K+fRa38kjHRagP9A8vajLQ0RWjq1snh/BNyHPWVDszOzFiVXf88a
Wb4fTStRJWnlxcmhJyM6a9VGp6JPT7IZHeiWyJ6cad0/PAhvrpYNbK3qqxgj5JdhKeHqDz/Ed4F4
M+GCQUs/watHP1cBcwtSV570LuiqSI/jxlZgzW43IJBDCYHB67CLhYza943euU6rMRmU3bTd2Qm9
fuivA/ZgG6U6pXSrIUXGmmtkTZAh1DexgugDNR1L8/pQt5uXeAVlF/yIgVNcNJrGzUxW6lFe6fET
QWMdIqgDV8KkXB5cJAiVsuhS81hqXXQNOxhcKRipgG3BGhpz05bPRhD3sIuNUWud19oSmfEx1wfC
ymcmDVvkjRCwIQr5ad13EMKJHnfOPJCmxhkujNbrShnNHWrhO2+BJfsf414C0ceOpnpGm/Pa+xF+
Zgd6fUZTH2lw/wujDg8G7RKxbbo++2wUh9y7BxW6ICtkX5xpOlYhi5YGdZezQKLXXItKu3DQ4ll8
84xsKauJ7+/RXyG/bYbpX9pC4yuff9zwa4lomT4F6A5YYw/Sw9XBgIS/Qn2BtsvPGlBhjUlPea+E
QEwzHcKI419HLo9kcjPSRLqvbhXpnao3pbThLNUK/F+Gwzm0ZWRhTld3BCrVIKSeouBnTsDBvJi7
eRjEfj2tUjN+Uw5q5+eO7vyzlLrT/qc1YxHmAlMm6ctry82nRggmkjIWaL6mGSPvsIlMfaKWMBfd
aM911x60fCDscqtp/qGbFhU5pY5DSfwRa3B3WGQUvTp1dzlGH8S9pM+oeffFJUznasIKUjXiX6RZ
Ph7Y3cQXReFYxKk8X5YBIYVsULW1zcole/etQBlzqGI4jAwPmn0/N6bwDB5SalQ7eWZv7uSVns1P
utHdFMLh4p67bidzFDPVmEZbbShrXMsBYfS651j/WcQtG2jalCZEI3ozR/eQe0NrzirhMhGu6psL
+4hVCBb/23ajOre7z4Fm6FqNLWfXIQvmSEvk1MFvWC4MUtFfnM/fF8IpU4e4FXgLoW4zDutD4X3T
Nfmr3zh6ZChL1AIWY1XHtEaubRFk8KWhF6ib0Xdj+SzlTdroNHIsPGvPwKGOD2BP3EU8C3xY6omK
YSnJ+dfpTxY51ma9wxpY4IxjBlkGGEfJZ2n5jnWKwimiQinzLpmTEhS1nd5vZ8Oc/7j9cQS/MEPP
Dt4RxjAJ3fvpILLIY91K5UZByloGMqM+QszqgAikoGddMqS5euthQHGIVjmEJQ2xhaeTcY/JiKNo
9oKOlYvOJuA/Qlqu8tSWPe3GbimE6nQpHpscZQdbKYaFuYxXtdena2jgEgo1iq33dl5EcKmnjn06
/jiezjJdLhjHbpVuscauNUUCdWTqaMMdkx7wl80y3bBDE2nFaNO52xMiHVsu8l1/kZjf+4MmLRzP
Ntj6Lwj8p8RMDHQB/Sy7Vtm02yzI+kh6y3eNdj8VwLHHPcbwabf+G7LSIyfz5TUFaY2HBPKhj76D
xLl8DDvKw5Y/AsbSAna5XjUYvSYdscNthJSECdXrxEgoaVGr8ZWE6nhO9TuvqqPmeV2q2tS0qQgX
U4iPEhmXn7kU02pb3mmweP0gi31BaR0cqmNBIADspMDonyW+VQOFbE9kBauNBqdNRPTztHZ4Rrst
a9VEEz5UlUnb2rE2n2wX+M99C/tqnZ0s6rFw64xuVm+JXHVOEcWVYU+exGQ7rHa5TmDm2bxU5BLp
G9bxP1dsPj5BsjLSWZdJbP0qIlrMyERqt7vshMhImOT+oOD0HSKpKy/suMyuKog8UTkRiyP19r3i
Hiomxx1z8viPvF9gI7tj0WzThY+mu5bE/mHTtHpTrQu6m7BRYqJel9T4sVU1OOG4Lmjk4eOrh2Zr
+AyuUsdA3sz1w6vM5AQ376mJcz6aGsKC1W6736/GRnTRT8dpmwQtQYeq0vSTXCMZXFZuB+smC5tc
DVD+yGqEuITplkExHpnxSXciLxN9NqK18sj9BNnDlr1JyoJYYGzUiflOIjcCurzmiHQBIZ9gDMoe
34D8H2th3NgxCyBzceOP5V3NANZjXo80UebOg4sBtmF3pHyak/vfSNtfRhAC+isIeQt2ZaxNUWnX
grKrTFtMmkpvjuwnJwWP2lzxpSibpFHX+o1JZqT/0dz7GduAMLYT9mGHUfhHBbtSAFCX4LyXBIwg
PC4PLIH43AUV8Y7GuVPv7G+xBCL7oo+Y2e8lZ/Pqd/Dc2wmSy850buyBXrTWJJyqCKJWjvTl4ET/
Q7cOsV1r/LfC+JVIvY0WbkbH15wXgepxaRhOpM4BX8BahkYGK3OiewsfJkSJS4cVtYKUYKH8FJQD
2CxiilC92ZSQCjzU8XFg0R2zzVMLubKNN4imNCelw3ZUpvJRZgtdgj1EcpK6XYQrLO5M7sWqLr4E
K0tp4XniPzhrOwWWIqtBFvBFE6mHxFFbDyvueiN6EkmzG7OnJamU1pBlSyp/v3kLVejpQVoY/dgf
eanWA5ncJnHmae9CD0Iv/Gh0Wx1Zp6xfIDbq1cF9kr1czA+fgBpiu2XLaZG0wuTDlEavboHCeDk8
v3rP5wX+qIkxNRP8B4+GnEZQmJwIhgKNeUDnieEVXAIAvn2RjA6jdNC+c+OGuEyvsCmmaTXn3idc
PKJHBTLgBGPZ/bpOWPTLLRVOeV58YKJNXlhs0RbwUhQLy3D7QlcvZHoDs3QERPG0f9A5A7WvZGWb
etRK7MqID+5UhzRdThpm4i/Qfdi1h/HE6nz+6i8G0qydM8WOPDavw2iQPPmrsY8xQAeYymWpAkSJ
A8lk8F2EmwmHr87KLYYgz30K47cqz7uRACLHrMRTKwGTxp8/U+bh3W9coS/aiguPqIJLp/3n6p4l
NNNkKoZ8yCIGMmnYR7IxYQ9Cxb1TNDhF0mf5sWgzbUxPsBmPOKJ+9xEmCswM7l9+DZ+c2vP0UYC6
eie21VeFnW7CieZ8ZEqit2J6ocYXwPniD5gOWK2ccambI6bpgUZOxC/thaLlXq61eW/RcIJzYJKY
vVCxKpc9HIOp90ifbTK5BjKcq3s0g9D6/raV5k3VtOfBswaIy3cqC3orRFHCDVtHPoeqQBEEJI1W
eT5PnSJS8HPoxQdc4/+yYOS3fxtognpQbl3FD1vX9TR/nGKEtYi6PJ6igwFa1vEJivaVZoXzy7Qn
BZOj6yXskhCXKNfa4QcgPx4mYfNddhsq7sDgPGzUXre7yrdpOjKFsBD5NI9v40MSg/s9ZSpMCOO3
ZUURum3l/KuE0mwVSrINZDcv0XRT8wE8ab+1bA1TAuqDN/1QBUs4OmltQjA/HVczIWRlWpUaP1KV
QDjkziuh+pF+4HSGKZ4CqYX02DsT5ea6VOv9slCZUaRtsw7lQ2+VvXHjYaYYlMu3952vCnW5uWA8
aVdn5TmDlqolAPr1cHZQ/z7933a9hd/Fx+QXSk6ad/NIgq7vIs6XdAEDYzpluRzrUx02XfUOQ9SD
Lg7ffXO6UasJpzYMAB0CU28HKPIpDMEaj2bR239WACVrGuNeyXI+FC+LnKpjMt2KqMH3fhiUbQ2C
XeNyPh0A52o55dS7OtEzq4SAAfnbB199+eXjc8/F2W2Msqexdz/Y9tZJCjymL3EUiq8krLxH/Nfs
IwKix/XO5i9RhmNUR/9Z7l8bGoQPtNTPeYgtz3wLorJf583gwc81jET4WxUG0ORZExyyr7cVnTfl
anGtXUblL4nhXtFyWp/QMKu21/xxpAUuijqbB6z16ldGdNiJQ9Or9v62DVxUgbHeF/KSPZcHV9Yw
vbiiMovg3eXHGoosWPvihaDwlI79QNCKW3afZo9KGyJFGBsWf9b7zkCUeQjoDjJkAAy3nJMQYGwp
04EE9ukiWVMDJE7TexTByqlXzyon7KFYkxQBmQmQy8HwMctZLf8YO3UasElufB+SlWDdgo/VA/ZM
Ayee3hwNF2BGCEQ6RcwD4I+YbxHcbqmSm+Ir2p0iX/THss47ttKRe+NhcDzKhjm5bRBsGG5aVhfF
V4MOQ7diAPvvsAfzEY15B32yQryq5se3v2u4wp5lMeTHZM2ys+GMnXG0e8Lfo2wdHWS+b6Qgmmgf
nNwHlkpieChDlXMgCCWxgKYiQlFzxnMKR4XhG44XMC5I2bm15o8rBbu3OqjQesrBuUmJhJAJ1zw3
sUcPCX/sFdYfUNJ0DKzc5NF6qmi+zUUlNNeg9AT/bhNbxVu2UII0mMC02Dte9d343+dQss1X+GbO
J0F2RI4q9ec1Ccx5fm6Sr7uXosLjlRa0rC9NxsDhYIU+IK4eHiM2M+9q/ROWFi0FAfGlTWGJhHzV
EqYGDWKosPcU5UpsvkDXMZZu4is/mwnyDYwetCCO6OAzu1oW9pZ8EmeGdB6pAx0btc7/6Ua8LSec
PFvGImHXmJz+LJZHk9WWRGWdry3DRVdAfPPhkLbBWkz1jT+okZ8tTVhTLnPsUk6ZstJqxmGUzZzb
hQslTso5ZjSzheCk7OGLkjezZvxVNFugANxOnh8J1jWYnzzjVdIGE5U+ToyNSMoohO9qIPEyEiD8
4bqj1i/oyUkAz9zk3ey/jm5W73jt2AatvSFOU1TZUHGRYxCLCjydKyGEDhJ72FBtBGoJOG6EVdWZ
1Ia5GZhqmfekzPdtWo6fzFb3qMgS2rb3SNsQ+ymp6sV0sr3LRpG/hiaVoT1BTmAYVl9V+b0ItX0U
Lw9TeXQE+lvVYqQAj6pajv5Lo6T5Wn/fhBXf85Mvn3pbKz5fkds1a5NAhfoPSkJAmbh6offHFNSj
EM05GM99M7iYBMvejcR8lUFOAmSZgo6rC6x2WD0G2W2yIw6tWfNgu8MZjIW4JYF65wlgXqoc0SQ5
UC2e+muwVT48sN8e1k+n0/PYgoM6t3ZgdbmlOJnPsME6zEG4IUbdpfhEBegavYh75aEi9YldrgeH
ZY9t9g38lD3hktYev/JUIJKk7X0pt9DzdgvYq4AzkNm/H32FDVNDjFSqpz+nHG3dd/ZMLD5Q8Vtd
W2qoJtJJISuIQ70fJkSAa2MJulY6QLaA0QGSpSdjCbvtrgJYeJnThQim1PYEG8LK8MgRxTArVkdf
BhhFu541fRwwa/N4vuwrbeJvquo8jRUi3d+RHf60dAdFeUE7zqsHfMvvgtGl4sSgpE68DbuHXcS+
I7GvHLPKj7AqGrdsnu61VmkwlA0yoYWxvjYKk4lFcqZPDuOl59EZIfCR4/UHdVUEvKYD9D5dZbvZ
hombygikaa4gtuFZ3B9C/sz26wlMrjwvaBHWt5udXrrFjeEix1wIoFkMSlK7EfdCsW52huk/UHwn
8obK6JAmZIhtSWZmEbbZd6DWdd4lO3MXP6bF1GP7+dFHG6fzN/uSdESFoAOJP+bmHQZIRHfwoqdF
rrRn3nCOjVUgBthn8Z3pnuR7vWm91/cK09wiTDdxBbefFuDAi1awPjgdLj+xmKF2jVOThegpP+lC
Oxn9qtwrJhaABqIXxLt0QtE4kV8b/7Lo+wOpjEJy/LMXApEgvTPAortCVr2g/5773Cuh9BnYpyr7
oPJUQUz3HSycUbEUCRqEIAg5IMjn2e82rfEIIHO9pxEc7//K1FuPuCeixBoubhbG71YAhdlUb7Ld
m4FpOeftRNIqJV+sDnFJCFHzCL1v4gTYKeJ32dseV0hFBuEx/GAuG7sqwiX/LREh7WQ/2Sbktkw2
uDl8isWCJpdYgmDowiC/SOlOpU35fWQ2yYjAUBCTs3QtJTdAs4MPSJNeLpLeW8zCoyN8/5j2Skv8
ql9te3zJXLKw6Won8u7zjv62sF/IBnlZRNDTmwNR4sPvL8/omWuPedwG43XHs2sEoPrZ7Ow6obt0
69SgIpuPDlU5WLUcw7cPDxg5AUZS+AoaYgOcDqtMfblciFQEgxJuIvhlYe62IOKCx9OP0TQd2ue/
ZhG7UM8iAUmNhsvyzBNLuUDvmfuQiXCJL62o6Twi3VvJ4lBXp1aDhaN2walSPOUOBaQd5jMhktiJ
vpMS2lB8gHn5L5ovppmU/mpaIsaYEb7f1GRO1lIPPSMhIfe4zLbNCt1TwXWoQ23bS3Enk8rCiZQC
+OFuOoQWH5mHYL7zyp/o65PItEREYxsqV5AUSaxhvq2yuC1RADmXx6x7PirA+FhlQiE018dzDg8J
rHArjsYDsYe2Rv/IDcM/ml63Dl38XCcyHCGgNsh8xaXfQ6q/bIHbSbCrwxvBhNfFJIXziKAru/Y+
bWTmG8spow9XN6Q6lFFJggyjwmFDIEN6XXb4ysEcavN6EdGwIh6hWkxqFAU6k1D2iLg2duUUZMFP
VnCajVNZC8Tz1Ny0kWAI+QUv6+/to789grKr8QrcSS/Me+KaSiYEKc1Q/Zqj9M9MQ1uVCB/USLOj
oHOXDUZKl5aajY3dmthR42ewajXTu4dFNTJAgzC0DM5XkzYtKhRI8/UNiRPb7dcz/TaO7jbvGRFM
zrpaQIcdLx7rKWFEIe22kUwH+x6VVjPFoPqN+FhvLZrpTETZFxp3D9kD2XcGVMk+6K40xpNoovEG
9IHyZ0fASH749ucn+cSp1Ubx36dgkFR+eq6GQALkMFVYuWlezUqij6Qa5uTKa6/D2ZKk0eYD5iAQ
tzmyqzMXzfpTJcBoUfCm1p0EtsJaDRQ3glmmwQ/azCdDdaIFh+S/XUuVv8ZFheK70v45IfWlGS01
N7lV2wLUYnIguVHyRtQEIMMbZvpht+MS/Mqxv4EHRNGSlfbCBKUJX3gHk3Aud+neM31b0VLQeSmx
gzCl9yNzLiNx22eBMcDPYmMGgpSZGewxdgsySrnItcfCxVNxKDiwRr1fo9P5uQA6RvytU7TbBsdx
wDtrD8xKG1e/07xIs/zt07v3NxsCmcmriw6TAYIEzpfbESa8BL53XxZZVj8glYTyAskxYHbE0tPK
xCVbM8PMpL0Besa5R1JwWE2f+mTUM99jLst7iOZHGpDZBuK1glfO299rgNtdNj72m45ZbtDCqXYv
4yRKI0qDb4myiPk7hQqdk3wgDnU8lBaPWCbBdTCUA1DVYTJip/Ex85htCl3CGXl+HEnnKAAx7Krk
qBnZmdq8NhrY+fXyD2p+/4VKyo9tS1hBNhC1oWVTEeIJvHR9WCNervOykFzSi41H3L1GQ3yJ6lXt
Pql0LNPMhI/AFFe91XiNiBcA+ZokLcYP1sRg4Kzn5FCTli5O1vqoV8Ye4I8HCmL6Gjh84A/x5Tgj
JUuIgvsGB5aUVSFfzJ8Iwqy6kSkr37GCCNr0CEO2BaykNh77dEUfuNEglb5lkB1sixueLP3koagN
nTcQJmxVHjnO6mLuZxwmqag1eZ2w7NRZlaNBRAbUgX8VsjhnR8idO571bSis8VIMhECO9bmdAsKI
v0/NeJUYvtpYo3tVCGSTYhYco9PZkgGME5Cs3ykIiL4JrVpqHmwarCXDeGciSHypKz+QUv5LZxqs
FsOqHELg19Ej8TLHq7d8QUXogUUDz21a3W685cf+YMc1WkmskyqZDFCXzL4tewc6AdyKyCJ29l9x
TZfjK/M9/Bkg5h8LKru3+4mZLOOUm6KJQF+tPJadLQQrsIp8/GdepgoqEvdBbuOzBxUTyv0zTx8Z
ede+p8YIHFqQ7XGSGyrDbWH7vPWJt7wIIUWMRt9utt8p6u2w0lpN/0VBEhi4tysh9gLgGascQ1mM
xHsniHrhLcuXy85tjyvdQaxpHVIXT/xv5zIq2IGUIvP959H8wIJBDBcsrmkkOPjSRppnNggXeWel
i5AA+/SImG+iS0r3ZIsrQJYEipVgRjw6our3x+s87OZbUytuZGRIRXmIphhNK814yqujWkv+/c+x
jIU97iYJJQJGpjdrgVQvyQISD8jB+aHxeuvIlmYI5Z5Vz3rGrLtR4zhaW62KJnEyQeHL85PcsjKh
kHVCc7LKUrW8AFcsKYAeYVio+l0Lk3AwAyRO3/Zj9fqcKFpKjy8t/X/p9xHoBeQv5JPMvMyjVJUO
99eeDGTC1rL9PusZYBUiti0FlGGFV3Q+O7PI5GuI4svCD3OKJlpZZBZUKbQKDPs5iv1YgM9wO9PH
/ctp9Y6Eub9S5bigEeavkhiA9DagxhsTLBIRracHwJXNvB9n3W/htp0EqP6Va6nj2FKB4StuXvHK
7cAzzu5q93RJwTjbrClgQtZ5QqZCx4uktogH53ExqeAlDZk8nAZcTT5frLl/k1IJk7wYl5iEB0mv
id3IEbY6JYBli2wWVYyOQ2oUw8nNE3I70hJGg/C6x66qjeXtwvmMDLePAvUYzQ3wJeDVqimpPrEn
DN0iLhl76SbuKr/1eZHTG+tvH5oUlcaBYiOI0Zf+gdxi7ciTcjHFwR9gXClUU0nf5nULj6GXxDIg
qxvWTFymKuwkt2wWS9PujI20GFkMCK5mi17rs/eY9IozY7eB26Qox0Sr/f8cOU3oaXTvAmkQUmht
sxe/50Bem7rTwlSe7fCZTpKRvaH5Pmwf8DkWlqcbiCXaFl015cLMTb7ySWHQVAFfmi/vt1E/pDYp
VcYUX1UVhWTmqDKXlRZct3XF1opk5hRfmWzVdxaAE0sKbYbRgC1VVF1TWGCbH/28K/8jTIpru0aD
rfaHPqbLt26NniVi9oLIr8PSz9RL8jCpTTY6qhePZVz/YNzbYuQHpMxpZPA2zwnorP0z5p1pmqCL
TNA516DY7AadaCeTDtCZGFaqHmD0Jls/OA+W9uJKq6NViApEnsgSYUwLFPxFNJFOpFmorywg9Ho7
QYofyjF21YC+5vvlx+HddiKB9F4awm9yl+//Hmpp6mSOsVKcKL3gzyyN0eHmz+yiXyLQwM9mba32
rkEBLmJDgUxSs77IC9g0qVkG1wDdsg7Faniz1Na7ct2P6UkkhHSJmJiwGQhrgV779awhN0f+kL/S
8a1B3hwcnjJ/o//AhNOdAtlLSnwZlk9K34kdO0K5jfCKiHRWa1uLt9kKvp7kC4mL52PpZudrz+Sr
2bzhyj1EdRYJFY3vfYYor2KVKUnR5CaWvYu92Z92LZFnWJsEggINjBam5N7sQVaCUK89xppuHl5X
bt+ZLtt0TeiFmmA4DphMpKcgSYkDO8Fq1hsNtbhh9wF1H6xdSuHy5Q2iYhH9AoIHZcsIS/Yjc0Ac
vPUhA+Goj3ATDQ0+DCHudB3DOMJmXKp/Rjijg64yjNfsoLLM4EQ35GndTF7wqMXWED8u9wlsvqaY
ono00tw2PipBq/dF5JS0Mh0A2xvdkwIQSORTM+R8+O6tQdfcBzlbs8mHhWyeOmxVO+4/j0rIeEzA
Mv8xtmj14uty48rpxLlS7nRjECvz10+H85hoEjScXXE3J3O3RJkwv9kdDS1ekG8yg/j7a1LiA/Jk
8+5Na5qE8mQZalE/KT4utaGd16rE/eo4OScRPw3EyldcQGRpX8HVrreYEhwZ1MU7d5sy5p4ub4Dq
sQPTTkj33378LK8gfOA4SliTNwhR24H5yjANe5XPFGJsxCuvb407QmmoamlyySnU7gxsLKjye7aO
Vq1jZNC6TMIauRP6+kAGyJNP48rwcUF6hgdoaZYPK1lcDIPgcmg7HCcRQJVcW8+77nSXjImLHrdf
MVE1WnkNf0r4NlQfT4kzRJ/ygrvyZNT2gl67y2B064HX/+WVwWZUl+EyWKx9imYu49cg91V2woDc
7UYXQEf7wuRgdrD/yUIEO9/Z3YUzn8qXGiTpKwqmiZoxyEaTO0ZVecZanUerUycjPY0Jp09HQdYu
qSZOBiXoP6QoRARkUrVELxPjTozYpPGSps7+PtuHc0t7rZEkSPp5ArjCrBqJrLrie+kNRHL/Z1DF
iy2vADBOrrPukAH51cTfI2+fI6iZq3MOdmvrI5nwRTjHndyzciYD9QN7xjYUEkyOF1R0FVYNsMdK
kM+/BXxRImWZg/h9uC5v0VLPW+sXmEF28pVCtDet4mFBnhKcWZofLqJhiztHT38BjtCobz+KAUq7
3faAc4Pn63MU/iQqZOvuVcU+NTgy18wHGzh606uP556JrtmrAuJpj1HRPBJ6a1Dgp6Sxsod2+o2J
gSF0vJrfpaHLVgI22OC2jpgB6FFgwYLjMUM5lijfF0Lx6V08NLpuIzH+ys3CSWd5mf2SoQZRMh2Y
YDr82OU6BnpZ7Ak1ZtRazWDQCByJ/KKWf6fL5oyjXmpnjAR1Yy4DWIxYACiMLJLnISjjslhgYiwM
uqC+dNy3aQpVrScZk4CPYuM4Bp4VQjzDcsPOxW7ZU+X6mQCaSi8WIDqMP9AdjUUTWAXognIGt3W8
vqvLAziyvQ8083dVC//KDOHNddjq51Ka/ihLEOl+sdF9SaifvieFEyOMDT3PHG2Bh1QnI7WPfuHZ
DYVrfpjSIugN6jEooJ0Ac9EdMSfvH3HRAndkSeKy9D++8jD37s4YnilWfTSekRPqLo4kl3I2/Y7n
dj8r2a8wOwePGpPIeU1NbyPIMYfCjp8k6uE+cuOMCi2uH0U2IW5m624rYbyaudXI71WSTBC5ovJ2
qyOmnmmw05FhPboWJSteaVm7MeHPcenShlseuleFKds1PwuqncfgkBTl+SPmb3tXXxgPc/Q5PwOJ
y5CdTg8By7gDHhy0B3+hUqQVuTnWfojBMvUWd9DBs5dCT2X/lzU+0MYo3g3JJl/VAQ+2tt2nGS5i
bhDP0s11CLPje8DEIad+1cDqMQ01wOWYGJNtXgozTCFv3bIjAZzig74hWloRAwCau8K84h6M11aK
DqEr3Ub+e863CPdiJWySs4wPp+JLzDrxLIX3CEAQ4fcVPza+Be+81jrK0e4p69XSdUaf1l4oPrrR
azCDp2XN7r84Vtn2gC5pSSI6fIDtu5MDaMoYBADmoPGlJ9wSj2VEgScNN9Sr6wBS7fGJtzE1ORq7
9aD+LXKW+34Tsq8CV7JoVfjA2mim2eDv/1Z8zuyybDeZ8zf3OiyhFsKXe4td0iyNdndH5aqks4oV
hjRbyjqBCYdzL7AlvdZVm5ANHuhwkFkvIfJZ1404nA+CkhSL01wHwRAi1zyXUMkJcwNdcmTYcrGM
x+o4zuEjI5d3L3+wIJ1QNgHYsB13YcB69WPyzfHD6qoWo7uxzyws2WuI+GQa1KYynDzDk3fZD71H
9R1VY9Vign/bu5wFYj+KUuAPqt6I9sZi0A5Ka5DeqhWlrcG9sePN+K/U+XeM8mQyzlZvCQWLhDjQ
2bbKjiX2/zVS5X6gaLJSOgDwPnJJiFbxu46AzpNAFZSb017eS6JRHLldPhJ+9vOLMRVVYeMyYy3t
/m4IKc8ZYlaubGI5vqxmJ8ijjT3mW+4a0rotSCPGde+7wMHk4DQhFvsfDWiEGVGAPBsk0WacuyI1
rRPCGOOzj/bOV/S+Xr+nQnBEnva/geWKrJJz0zKp2UQmbBGyeX8R8afX/I0INP1Sb5POPyb/QwNv
vKRIqUvs65I70xENgHm5b+qKqtWmoH+BBtT9v9I3/ra8mA/MU7uRZenYcqKA28Z3VNXU08vpi0lR
QEqV+JEpMyTvCjh2LHE05RDe6Y5Z92ojXn8Gq6aCVTaDwOvml+Q7zpPD6Kvaw4cD99nLMW9Qdzpx
MCTYqSe1AKztbDgY6MsaFghqNIS1vCCUMzGyIvcyuxoNU9DO1ZYdRB7VlKvslzViW2QImTOPVMga
KfQSMKOka6N5TijXViTQIH7E/CtJ843ATjE3BtEhOuBA3WDuihYn/sHVnBxVFq0PE1F/1m54Ab9x
sfTrtv6WdpZbXAqh6x8oCFTHlA57jpB6istBjlcD7/3oK6zTPlSSA09tMbeq7l6tpQt0dRSDKpFm
YYvKxJmUvrpjSUIfv9Fe/aUZVeLwc0nC84/oiLvZLdZgd0GRZZXcMF52oWDVEc16wAEq5uVu1Mu/
h54hqcHZ1KhHJRoD78u4r130QATPXq4lV0hiad12ZXl2/RwkRtgyKXbEmVGqOD4R379bswnW5G76
3nngxRWBin2QbP3KlEy2NbRzISZIvhYyPOCQdYDwCBkvdy3BGu1OYifUpzmmO+kwN+C/9J4rZitY
ot4OUqlLXceSWrMp06fBIvc4UMWxyPq5O6lcRe82TCeIkPnimA88WkAvisREeBpsLE+t2HqqM3H+
fkCJoqbO+1h/r/84U8qaaQPnppKjvdrfGy6ZzdhuGjKRSUIXeXpaBR+8jYerad4lmG6uOCm9Bmcj
7CQeZ9Xo+L2uf4PmxCrCjuNND1J2EQDAXVTuSBufVEHZ4q3bBA2wQHXqtIub6+y0XtgivAtwyT27
oNHd+d46CK/uakY+87Qx/nrylalPeYnH+9OlkDJXhyTHjUyP81zaQGPHC1zbHeq6xXnZMA8RkV7F
2EeewO7QL7yV4mM3DVnon+DC1gZgKYS6E7fW3vY21ypLGnINDZ0omqhGz9lhOfJ7gd2l0cAAeX9C
IuCZNgP0pCBukvsywKqDouCSkPhZM7aQ8NB/bP4GSgjmwJtFFccnNMq0RRzpZVb7IljuFNTKnj8I
V1BQ2tIV+vKWFyxDcUHEVRcgS9oy4J6JS9mV5tFoVCGSKOjvObvr7XaoxZeKe3fuCRh/QwrNrA7B
9rYVtY5zj7ytpJzGdc3nZOkMbQ2XN4NaxiV/xmxTWrKa7eUAke97ICVPtvLNYV12Q/Vi8nXUXKXq
zwJekIqjRBgkipjkiIoxu4qdqJFGUY4hMat36RM1bEXNUIS8gFf78/Xpdo5aMesWvxmThSqlFT25
UUZ0DcGET4EQqtUH3fOK08RSY9PNaQZ0PPjyQuJxsWtExEZARLqzhh0PBS4Xf/K0eD6RJnMOHxSQ
gqkZxO5wt/EBMRmvmHH8E2YvEyuKT0v+zFrVZfsEz4xVDu6CIH52UgJ03NShU0IEoFe/64Kq3+5+
HFGfZIqsNZf3+qDhzCopv+Y5BD4k/yvToD0mPF2IrIA9Q8rQ7ksTEpS/Hdi3GvoMtuM3OIrhTFBO
c1gEdS6Mb6GmvlPxPE2f28yFmJJwR4bawlWlYaokRXXDym7eQhz8ZEvCJ1n3hOWc/hD+/pRFe4Tl
dZBvUMSoVov7nYhO2MKrijwEbed+z89aOaT61Ob5l6gOSJLcGMW1VEguVATIbW/93ZaF6qOrPwpF
0D+PFmJJNtXTRo0Y/PbRKp5qAW9FRnxHSp26535mdZCir+Lanh8SDO+zQs+Y57EKB3Zoju43hxmt
VCNOPGy5zv1cGu7Bcl71cGiHr5p+7ZcCjtvJpCQM6bCAlXY2VFAyYr3NSc36CIPiFcasM05o2+rv
R7iWSNPHGIwwSU4cESPKlIZa0FO3DCG0Yz8tafvFJXooirOQ9WaJQeNBXVwJ3FVgXpV7TXlDuDKX
4skOzPmB+5o6Jv6R6NTR/M6bi3f+6YGaYqrPPrvagyUaEY2WYqGQMkU3S6sdfjuDG8rs/Zed7bec
f8gv0alhxvHXOkAVvhUUy4zVERJeoURWu+1tJHZE2GcKyj8XM2nsLTFUKIVsVA6L1FTWNJE3hYYP
XTeS9vTaPjW5pS8EvwXJStriS3dc75ikS1oBqqzjpEYkK/UiVGNRm1rTBtQeg2xMR4obtaXk5WaZ
DuQlCQgzU3/SEC4GbKHD8qiE+LewjlPFywTW/L2/7Y7MiMpEQBCebdsEphErZHIb3gYeWwiIDC+Y
ndh5WgUPNCe/jZvfnrui03Zx6hEvxdNpoBGIaWCTNKYl8dQKAmt36GDnGchX1tyNEYNLpb8z2ebK
uBxrBJihm2vpnKlS4VtpGpwObOcdkG6Sw4Lyi56jjw90zI+TD0vDTwGBvPbhF076AXUyb3CCo0I4
gXPNUsn6IdC9s1XKS/1dwW6pPD0CUvMzGKnSWBQIu4FrgB1AlJxdlIaJTyMKBRLnALp/ni/Pbfpt
B+0GGSIJcuocBenPF7S3OQ21fJDMYoJS04ngRbm3aiEVLcZcnEBkNnS+ez0GP2jhKHvywe23Y6tR
3UNPI+WphYejSLixbIbK0v4gdPe1J17LFq2eNvgRr2T1FwadGTc+A4HM6J5I2PtsJoPbZPFgNGow
DzbJFeVhXqfx/kMdMIg9tMyGLXNlb5FxPP4NHdL6oIvPC9qxBzgzfM/7IHZ4s0gmCeanEhSs5u7r
tT9/WZ0im+COED9bBkYQ6Jol/45FDZr83GnZRQShyg3C7NTZbiH8irUxG6a4NR3IuobVs3AbGuN0
bfAUwQs0yzvDMrNkczwqDghcBLuIz9lQV0Mvz6Df5nKoSqPJtWl5FNYCKMyfKBys0FBhdTXnMsuw
AcO/zVaaCHGvKLLsSt3rUpE9gfWrRGIFv6j+942c01Ek2MMvgB5278fPz20gecsXIrHhvDZH7Pzm
gh9k7k8ojoRkB8yAZr8ts0iRg2GzIAQkqasaa9ucmX0H/Da8jdC3Qnvga/BD1t3pojtuoS0FttFw
fkRwU4opKJeIWA4SWshokBGUf8PFgbUscDkObAKwI6QDinv56GkmS4JUkThYVr4IeB/1mFDwYuWZ
wPFOv4xdUhOJVbFHD930iKNsTqb2WzKHnXSbnG89Xo761Q5zwzNw4uW5+RuLHEWpWZ1oDASpTEzf
vLuZoEyy0mXyTf7iBwW+3EAx+1ZHjgFUDK+1fCQUXa1xcngQN/+OyCyK6ZR0lpX02x53Ej8XRysb
TuQUH/jrtuS2ouwIKdRas6s2OqCzJ9+YFyttijeGgoG6hJvVBQH11kerlHmPw0BEN2aeb2yRNqQk
MmayJH7Ki5gf+chMrZW8ELBW+II/qtgmSLhBLiF1RKQsgvAp1y8qf5fxIAuSkvXRX2Qsp+z1FtvP
RBSRyhucm9pG4L/MrJGlyxhKwSNDeWobcY7VjHqmCg7Co4t/wEWDolgB2DoOinCRvh824jw8GaaR
cVogN7cHdxOJrNGywKXt+7Z4UwSWO9Y3ZXz1tFY5kb95VfvCC5nwwdjeOZwXGlLmx4mfyi7e80e0
tvZkhrAAidVB+AA3jj+46SpmP6fBOmY9s0V2jlNhw3wGCU8k1hHvPREgdt35swAYJ4Ia8JIX7Lwu
Wet0ZSdB3FYY57icG0l3D+qgkNtS1Xh+fpWTWD+PSEeluM0+qZbomCa7eK4u4DNnL8I+rS7Gj359
4cQfYNrQkkhX6Gv+3bvpJDubJ2qsRc0g63bxC4OnX9tNQONcrWowJZE2q2z8GIZ3HCkho39CxG+X
6HyoHeM/fTQOBaJSDEc8BVaKpHWVRcqTDdXa79QkJGxyz0Fk6zXq/bOliluagwU+09G0hY+e1d4k
HKSQTXfHKtH6atY6wHZyG/+4iQA/qTkZA3bZQSClVHbQiLxtQmLwZWrC3uAH6OGEp4AgdesMrmYl
FmZxfWKzWYB3LJaWtkuxg3sHTuFv+am5hsuHPdR9zOqULsySHvk9UdUDZrmRoCcvCguEQuDe4IAA
s018g1WpLp977Sw/5LUEVYqlEvZBFMsOMY4frSeP13yFBuMI4PkPM+95XBClkiEfEhVIJQM979hF
j9Ly4KMIvIi0xvwUUBCgM8MdShj/BhFtwAP9Xppv/4itXSXNS6cUZO/N7101E91B+iOML/CbWCwg
nYEgMUcmYfS+wHLoHFV5xz+maLA7EeOME9QNWA+jaVbQKOV0i2BAFwM7q2aUcWPi4fXIsfWDbxzu
Tncybsofu88wM1o18KzYAurisdOA80uWXOQGSGRhvNANlNhstt2R0Fvc4aaG8EUlzQPXuCZVylNt
4IKVS7jrQyzWQfM8HFWp3SFNCKIbzc1X4pMoxtedrfubxAkdNVTiopPUD581uVo9v7fEs5eMpyoD
tsI9QbJkrN/OY5K0Yewyw9/X7N5UNqvN3BkBj2PyzNkPpXm5uQO0wkpeWJB5BotpBYuj1BQy2loE
4uUoWivgv44464+yzswSeR34vK/HVu1+uwd3t5TDK0BiihsZYXlkWkr5r1lxRfUYNtUANupe3XYD
apEPRNPOd2rk11P2o8KBQVl9kq464pvu8Ck5i1NYMgP9ALh7u/6rj3R5tSAkxsOiM7oHA3+W2g+O
wbvftnnzRQv6wbAl3MmvRKV1WcRGer/BBqWsrSkLciR9JlG/2ccmJbuFEOFgZZp7aN5LLtfRmxI9
DOqOwqy6xfN6niD8rbJoX87Q4ZUnFQR9sqJrWO85WTskF4RrB0TjqMGkltr+D/yedG4xUZLEt9+l
4Emw8azP2LBKyxbFNYxa3N4SJuXVmO+Vcm4FOAIBwl5iXdTO3fYY0nKE2eoP+LMEcIKw2CofMvrC
LZ/2Kk8KLd+lWhMjEcgY/SuYTz0udJt3JyhmwmbTjb+XOjiFy5vmKH5ypmnEse0oJNDvx87c3Qex
TkNbd5KgWz2MGeXnAsFZIlRxuLWMPDM3F4BU56na6LFiVH9l51FMVZaPKQvmJH90K4PQfjIKhFbY
5xKgn7dXgXGgA0TEy1lAzcx7FXIh0EwNPkxfxemswaBx60op1k5hGaeyVvoeKGFwm+dcAnmOkQbq
RuryGtr7YXWDe/NUO1Lzis8rxbkUnuwlcPBJYRgq+0cxY/hoe9foejMQezsQUbmH9JyPlIinwDxI
74CDLSTZatCx0KrXjwp14cQMr9iB/anYOuNS3aWrpt/PEjmEE8rCC8wVM2svSrRCYQSVX26hfV5t
gF3YW6i5kB5fITkiWSokawwzsMTn4E8WdgMBUcBicM5678DPe7nOgL3FcWoiKduIgtfeVDTws1x0
fFKQlSR1M3lJckLe9f9kFO7cyuHqsnuU2xBXlkgXyM/bH8SxVuQBQISaMDMJ/Tv4zZlgFd7WPe4P
8XOKw889iCttlvpUCPc05avxPxBF5NIwTpxh3uPdqAQ3oH5kFCZp6RmgX58o5+Yk0B/Z58lG+2Gj
8tkFYF7nyhLSv1tJ1Nl1Z9GPUoY46cXP9/zzVaVBj4YLqlfMAQT0Isd1pu5GfgEwKMrw5amnFEAV
yhfgHxXBKazkfhS4SwbSTxc7M2PmK+jT/S0kc2cu7NaC3aXk/lf7N402+6k7zjsVmjliRw4AopKs
PY2DkKkzDGekOsY7Qn5q+zlxiiuqZQOCrq/UeVaysBnrnRgkWC/ed1I+d3XF45uLRYM/3KEcdvNo
fVMOx3fzzhYPkLSpaYwUitPRspfGEv4qU5OSJw1Ztgb6Cy2rayHYS5vLrXrZC9XFDYndHd+pcacP
DS1v+3nLeOnBQtSGYAgXRmAjdjgy94l0LwAtl+rD6rkGMVcEzq7UOsuMD1A4TM1NlPt0LrofHf1E
xgzKsR3kHt+zC9yCg17XnNHuKGeEWa8YQxmRAB1RGeBBGSsUvCSDc4IXW0t7lioEJc+2MMNjJtx3
26Osn3mpjfeyGPavQqEP68aW+PFbQ4Lrv4WqMbmeOkAR7lRIf4oO/5uVA3apOTmsC6sMO/cpSZcr
d8pXeIq8/Ci4aKEU6B9AD4eMROU2NB2m27zBjw2t40tumuR+vle32g4MOluFZNf4k/CaufZYV9+8
GfrEIhEKFldccOO8f0M6TH1Jv1J4sg49lorpsltuk5pjhBaG725U2KMfm7+dA8r5Fr3chSEGa/D+
MQ8chD0wMTaTEkRMO6yzdUkycU3v6OhkEnH8fjw6QVlzu1IRI6E6J6PRWl1l+k3ip5Kt4RTqHdpN
Vo4OambR8KzpilzKrCbI7+0dXvii8JRMV59dD24lCSK4Sd1dc14Vc/sGDNj444Ff7/uH5o+LEtIB
QUcR+XSQVrtYTp1K6hGTJ7tAiZVJESqpgPpiyOvNeiepzhNLRWtj3KJ0FQeKjb6DKUuOWVHAbqmG
fq/RU3kCqfK6BVOcDrsIGKIJBv4d+nC4JxYggZs1Zz7qBEb4Daq4tDdQdVgvZH5jUt18SCWFSXT1
Rxgj7hV/kozqWzBHmxw7G6Ct6VM+mIJpYKPs55HCtwe65vE5YsEuU30UeWEv9Q9lloMfhlB5xodn
d/sk+6pm8sI+8aOPKlgjb3VbqSj5/e8hxQlw1XD6mVLagTIsKGgkzjDQ4claWuAigLAEVs2CBykd
I3sJK4BWRLsVTL5GsvWjDo9KLRHI6yPhOiZc5AkN2mNim6ynIB2/gspCEiWHcT5jotXyMvgj1zkT
BRi1eyYF+qtlO9GuPlg6ciHcwev5srl8hf/4nm22Dv8nsoFBPa5iLUlGyhXERItmy8x7A2s3qQbU
F8cxgflEtB5nRfUDBatooAfg0vL2kYa//Qg+gXmZrLOe7Rhjz21emTdhbRmUCMQOOn94qTm8T06m
iTO3Fn75hJOqcGZGkUWLFDTA00g4iNx0mQIUVxBqCc2dsx7tcmazgPCh6bXR5+6ST9XpBZVPGMxH
RofJzoMc9NZ1O2RXNOJPP2ZOsZ0VLjsaXupN+2vGkSKUd/F82B+sAzCMikY377ezgk4+Izs0NL1Q
PD5SlH+zxgpEQ47O0cgeeVUanSHtSQqXLn9kLMqda3p5u+/HaLw/J93SwJZRP5UEyq5LNFefnzUv
/dkc+ntOMKM6VAvAw/hgvt2YCfxP3bR7fCXjtJeOfkZl2jASpnnBeA/IrZ8pwQ3n5CDKQnfeqynN
e02nSJ6oVrjjuwgOsTLD27TESYn3BRNelx5tsrfEGYc1JFwTu2sEo45bnIbHoyPw+AdAqlCbhzvN
Z5+2lAW7OGPEbM5tmkVjDWvyW9aEyREvIVe0EJv1+1N9dxnuKGuvq45xfCKCDmz5a+dxo/RQ4JOX
Q96TN5AMxT7RpfJC2b6CTNniJ/dC6Aj7nVoB86pj7ejiGkaECQBzJuxEFi4pI2alORqKLMdzxAhR
58HmmOS8FlR0AcxXLFlx1YbGH5t6FSEfBuFinRkOJ+XH+nyli/WVzHU1S+I/2nUrPMGSbaxTIOmQ
97lLwGWd8qutN1JbE22aaM8nNuVxeroJagGaq/kK3jBtCpb7aEQsf6Irl1KrgXkdHPFZrVpxGdKz
gRibqs9IMul9WZ+485f4cMKk9rEl6S9OKh81PtsvUlcAvEUNygAPF/UIidAd5HXzUCCvcy7fxDUF
BZSdvKIDK0QQXgA/orTNZkSOg9/Z7RwkF9AqsOk1hKqpSrckF1sQ0/VvdI3jYKFZL81wtzxdNVm3
+etMABSPHyhfcUYmkbo3DVrNvqi96lnCPmZj7u9wRQCjJblSU/xZqre9RYif7U1XGad68AK+Mj7F
oe6b1Gkbm9Nd0ic/vWVhilSvCGh0oYTRl1nx2i7EDB300jdcPDU1NM400lTesBGSiZTjgIzhZxGH
MK3BhMOGw4zUsFPKFO8JI49NIqdSaE4UMsplVTwNu7AyEXWPARL3EQG1+YtJxGtbyebALPKWid1N
VffkQ/kZUeydzS3OGSpbkN0eGAHVVMu1aErysF+JHlrgLRgmZQTNg/SUck8ffCoWMlXtj0jpwF9n
WEqSXdf2t4ocAA74L4VuSoV8xTYnXNCk4/tng5cSfrGzvX2wLldNWTx1clRSmNAoyfpaGp1bZC1e
EDhQuSOENcm0J4kygVJzb9DY+ToSyvXZMPyRogaM1d7DEAUDZogJ9UDshs1YWR4AZUGq5eWetium
MPaBRMqJEVpvsSYRJS1ifk7GHNS3R4rQBYV8LFiNLBzy8Tb3bSNi9fOQEN2j0y6kPOPejH+On9TA
al85U0ElnxBs6aVxTguhhoHZ0yRzlsxZHRFu0uK0i5VCr4tQhcI+IvrDTRmdJ0HiyeLQxRejb72x
C59IzbqFpIo+FwTtJydbMeHXY3/tuJlWf4dmgjOMBiInkFjdApMFar5FT7U609eagRwzL5eDqDoJ
mVVf64yJU8GcLOwQayq8iUCWaCm7SaP8hJogYwX2VZp7hXHS4cWSRaDafwYAaA1XgBdNcxADrWPX
18u78nUA8G2+pi5FFFpwpsqRNWqKkKK4OeUKaoc7+nw33+BuhoD9IGMucUk55E5EHMV+sHCBO0Ke
cAgTholfF4x885hiO/GD3hGpWQ+U7qreHErvodne5TxWUHtsxG+UOSrXpbKjGt5yhq05rDpBQiiy
IpquTvve80vOFKVje/QpFGsE+eRNbQfuRPEccMqJsTKnibdynxbTQulaOR8VZH+FFqblHADMvdiq
ff239LPyvb/P0T3HWYJ4NAfJp3k5b/jzj1xwwjdkDNiyRCF4xQt7Y1WWPijKdvJqQJRJeSY7d0ao
uwmLYG519rYFej4uvNjYOvYGSpBQbzR2Y5yCxSgqUEK5wavYUUeWUjAq0gO3Y4KfGeiTkQ+BMmFr
DXvB9wbcYb4DoH8SvQshagVzhqntmEGBYFWihHP3pR3KEXTNueTgGQgSK/1MpQ/UtoDeEhOwdpO7
p2Pp0iBWS2MllbjNm1xz0gei8+mBOKgr1BnGQcVFbG9Nu3sgnU1geHQr5AS/7VGGvvYus8Rrf1xm
5ifXiGsQF3yC1NZtWOnAGwUwFbl3Jp1I3fE+0fxTPVGYl9+kM8aDB/PwGo/UqIsUIHfxpieSCpdH
5zGBqNxi1+a7NFArx/KSFUECLZATyAG/eMVBFYBqlx7ILhQhjdlO1pJB8MWPp7cbOTlPf32aLm4F
6tes1fLESBmF0LXYfGK7O5mLRDNA8sDPrL11xH9bYmmniMT5+CGDeyhq4ID2hjqQaki6f/Ju6P/4
b76Enc8Jl1SVQPdGonDJC6HP6VoM9L08DWHFBOWoPgrsf5r1VSJGhIzZlR9yvaq34hVO5M3fQ/7v
agG8CUi56M3VtQgbeSUOgNBmoaE4URAO3nvDttbPANDCfkllOVVAy2SPpJ/mgkf4NF/zznhul6OS
qkdjCdfJXhcNrhJStyc8mWJxfFvK9yYAsLrE2GMlxAPHGZBl9EqQai+IQRyp4+R2lPNiUsNGuETP
XIdNCCF/ySwR6JFm5Q46mGr51bbe5uIkbwdNammlLsOKXxZFDv8wYGcmRPxD37eRlVU5yf8zCKCs
ADyjbjqIXfZGXRMAAxx+JUr3Wmmnc52MeNp57K6QJ+HeMEHPUKHDmTvICzxildhPgRJWAeWqGOl5
iQiobAI+Qt4YlYH7m5q54ecgWMN7O6i3FQxnc4olNg1aFYsHCle0LkrTifNmeyAYAOIYBQx9OO8Q
xheiD099ICMlMBvpl8tjyBWPKLxVq2tJEYZSA/6tSr5h7QlhBOvIM7oeuGYwTvnOI5quGDL9Gway
/JjXAOhzktpt7HCVbnEFX/zrARDDwn+H22YtK3MqDHI9Hq5kPSUkW7iRbH9a2paYbdTCMswvL6Qq
sx9J7kW0gOuhNTzxqmSCOlFqhvHr9VsgUjFOS4dVumW1XJCIn/DRUXK7MOL+e31rjz5aW2gv2e6X
Z2WYnRHO9zyPSbNsgjvWuOU1Zc3X22MABH6KjrEgjlmvxzan01s2cpOkqEVchdIBxawJdVaB6mdp
+83iFMCK35FsuKaQTQbDWtml/hbZn4SFND8nZ/yZkEjvC4SDAFuvQp7FBkk21Iy4ImwMFCw22faP
sDxmZj5nqcIPTYkbGduwMfQnFFycf2T/9GGpi3zuk1SueyaHu2+iJ3i/zI/f4s0MiNWuKgxO+OUY
mQ0d36VgIdOJ91Gy/f4+0nixFrKMNHd5o+lO7bSPFJ2Yugsix2+WVV1WpIl8B1hsfHuZzrTgqrjL
9EPZy2Q7RgI3RnlQvzVdGatL5Lk7Ms+HXn+iYvYBe2nIncEUfWInS5x63byVJldBvm0L0xZSYB8I
o7+7nJerHLjzTpvWm+rPqXsslJk9zDG/ZIccXo3anMSr3yYhSlXKXDanbdJA9HHL0jrMNyTlygN8
hNvT5r35FUwmO3AZRL6qnJl3f9DFs7QBOY2kXdK8l3g/CBYQMaPzlIVimJ/RggsQcyxJlpByTx0h
bZktMj9USreLAbJA2FWuoUsqqP/IfzWFMqa/f3jczXdBC9jom21sJSPyIA72IUBQwSy7DyH5Xof3
iwVdggag0oyRv0Zim2jApRmcX350CZhqaJ3U8nQTD8ud9x6hyOj4en8ZB16QHL5NZJKM7UhZiW2r
CUfbjC5xranoWjtqmhT8LZVy8ebYXcYnBC3aTBXKW2jfgDQP7fz52PO6ksR8/TvQ9CW9zALOLGfE
RhJ3IU0AJ8hQiBzqnVK2tRqATg0BaAfkmmen76EoUNgcHlGxxrlq3l3QCznnBdlhJ39voousvuxS
tenPbush+W5WbUKny/EVonYeVsq9mcOZ6ll7AJ3Ib+/LbMBrHaqjONATL48HWS7nKHB+Vqqkrj+V
3m/KOajpztS00UULwAxHrDjVAZP8OgAcbzom67rX9tJnQ4WMP0bfZSdtovfP7PHFwVA+SqQwNFoD
5uQeiL+Ufde4fQZ4nkvJfDKwLryaVBA6COwvxUDntTpLfiMFqydDA9gfKUkZvU/fodfXSiiwNLiM
h2RvM4/BYq+v68u9VsyxEv+akY4wvYx7v/GpURscrPcr8zgs5XiACsh50Nq+RGhJP6wWowrcJe/m
a3+I1Ncm7ysSzhMSmoo/+9+1BQIFjNSAZODrxVmk+Ch6PWLFLe/wspY0SXX9XceH3u2Dd3iLlOEg
Oe86JexvwF9amf6/EQHFVZ2+UBNp8E2ldgCLQsgydz2nS0YY49WHaKMYC0nN/WJwBtUQ5Za3kBSO
XlUgG0MoLFv9arisHu4xEKJeH9PP/YtC4fWu7S5a3hHta31jDVyIswpQaAjtoiFJtmJXNuuLv7bR
xOo0P4YSQCZaQltqmiNJssLf1k+LrI9ujlpXDJEHMxb4cCrQtbXS58xTiG57ZAt3bMBB3WlaT9rX
HDRvRLs7L23tVSZ1gJgUOLNVXVUdXwmD8w8BQ/kA6HyMAkcUenljH9AyDqufOnddRxJQORlhBX9i
Gn/5yzwQqw1cQ1IY0Id9rhqCKIzWwsJKjjCgUjWQHf5n0K9lYMdLY/S0Sm6VDvpQvAIVngTeP359
VIrzK1g4QrVgbknugdPaHlubriTnDW/hIX7zRFtrtdKTw87bduqyfMpBcA3MKgk1U25PNivrolQA
hneoH+y8XhKilEZeYkchczQO49FYB0V5NsD+8HL7NiBjSfl/97ubRbHKB4WhUMfIFYBnRFeXXFFi
x7X9cU7iq3TCipuJEeCfuwXu3/tYa0M6qCKzhOWG8zapnmR1sE8pISdpGPZA5EfOIeeNy4yoeALE
IMZqfLcWv/pqZDxrIBlJp7yGPm4ZKt2wR7KJmQbIt8ahqiSa/1IlWT8vu7UPLo7sMD0LWloz2AJr
tuaKqeer68qyrX6J6Pxa7f3qPCgfrNAnfKLaYi+Oj7zQogSd0YJFaztmD7vdYuq9/JuAXeRWCNz+
yII/Nx9uT8bLtCtD8c2FXkNt/rrFwNdOu6/Ns8vp5wM6BElwzHxkfYxJNICSWbdq1S3xkBSd9YiD
LUf2Zxtc98mv8m6gQ32Pilmf046kSApsoWeMEJtZ13szWVX5SZOMYcCj59Qw6N1t541CidAn6I0J
psa9WrVCrb6bKY2F3PjGx+TtMBM7P5gpZqnGQ4eZRoK4mBoBqvBKMO82kajCvT0nWGpLWfr8aVRR
32mXzdPCQrvzAbmvLW4PvVtnOA6P9sr7udYsWwUMasVUzIDqUQCdzfG47J0t4Bz+1Ocwwp8dbZy7
EMRGZKjeHU/JkD3NJELBbz1Awn6Kk6V8sEN76+Dr57HjLEzbngUa09NrGXe3ksNf2ccUF8qkXPcL
GkiJIXKakGh9R3K8q4lbPPJrvpmBRgW8FS0JxL/GmL/3nNl+ZFZZpvSRyAi1i8Lxjb2buttjJl8G
CanrgYkdEpQUGDrYbIE7hSIvepCSkmAZPz+fuj5QI2bQIXvXunVrV1fGy45VDTWt1GA/nrImbqay
DZbJr1iWuDqoonKGm9ilA3MrV1qXyOtoMRh0VIZgELG2VkMfsZNGr4V4b4gPguYwZDZOuHpeqk1/
cEN373PdxpMoGdljBUxlmdPVk39HPs3BIZpV6XvfAhZ25pp2Lnq499s19zCk6Fv5ubsXf/NsXVQZ
qCaWGKX/oQBx+532Qp1cClocsC9bF+DdnUSzQcI6TjLd53/dBskrdOfKO8Sn90Th7a/HYHjffjMi
vjSrHc4VQHb1OsDbujK7ksC1HTm383nvcoI5K9ZZYQleRd9NbIKg6AZLrIsZMJs2FfIaXpk0ohjK
Zjs5AoDDHeM5BphCRm6GndSXfLAIzBCkRcpgmTNlww1n49FPlasicehwZivzJP6qgYVh8qoJsRPf
XUMAzSM2EF8m1/SxVCrT2ZX2rRYkSuJxnotjBwM3PccpBNi43FFKqMOzqu1A8TqON8PcXAsYwkmz
QGByjIISXpQyFlwF3aybsRNKwwO291tKqEfPUGW/ButnEecAkp+mtxokuN1oubjjzGc7uyMGELlx
QCgrjWZ27R488C5OnrUvrWfUpWG9x2XrXV2A4L63nX6NFA832pMZi6KgSyOwUr/ZO4qkXkkHFlPz
+RJncSfXsBH7vb3esc5yIxXUNoTVTJHUdXfSFvaMTsncMXGf9DRldi3FUy+euHJSHqVMMFO1qABi
Co8ZgmqSb8Y+JIZ44usm0To8vfCMqSZk1kErj0P2umYrD6yeZ1bPkZiG/fqtsKvfLJv3Xf9juhb3
eeOH76NMP872EkEdsvkFnzfUssWoXvPHVEGiTYyl4DAlL5pEH+Lf68xwoW2ug1Mo4QvZZtDrAq1h
l8JfeIgT684o32PvpTfhfegwc9uz9QsCRSP2IqNY4ysmhFtkdysdd4DEnKJyi54pZBrDGhXUSkoL
M0WtVeuMxxUa5dmtP94Ab3tICkAmk4wV4q4fKzQoGgrKXtF5k8ID2SZGewYIxkJBh45PdfjOgleo
d3mzGljcpN6WaUujALk910e++On0/DcPwUj8PEZl1NJICBXLJA8jiNGLU0LIiuDWWWCgru6M8Dix
D9eUibim6wjn83XL5b6zds5H4N6L8KDi7AHryRtVFlkdbYnH3l+KbaM56XpsBWPyyUufpUz45C6w
F3rRFfWIMwKF9yjp43d66h5zzHPWpvqRKnawKQHIic2Zxd7uYD5W+bSSsGxHUsuilEKrDWJv5KFi
5qdVt3BZdTbYwnDaBss05/3fl/GCxmc5v2omjvK2WwS99Qi/gZIg+rsJ3qRFig81TmGo150+W+Ff
iDMNELB/L+7QOUnaxxjnAUn2Z4xfYTXgBRO1xJqgAta91zlpj7tqcKDGsbWaFpoWg7sg5A/uZTl0
we21uLIwwUgTjZetvIdymV2JUX2CDsJwJ332MRcQdG9sBQS0cu0ZxpscZkm6ZriS4nSNIbZitRrE
eBFzOi53uBA2nZLhw9s6z/4Jepv53l7A1k9e+4jVQZznX7rmigRC20fueq2uQAz5uGD/cwDY13le
5qnn6fgOlxc1QHgTOmPLBGWfO+VXojm+BV6almaKW2rh+f+WeHPgEdLYiyjP7SFSy3g18Jc1TBMa
fbGdsSlGM/TUR8J1ixewm3fkDzgd9EjYxl8FzLjpN5vLsJJo2V4sISFEtjp7TMTc5OL7HBsYpCdG
KF0y3QsY7FqmtHzpSkXy4+XpRehof2/vamPt4hYg4E6vBJYuayfx7Kg/kd87agUWXZFGYQf9WxZ/
S97ICFZuMJsOJD+7gYU+A2lpfVZYXbtA74Xt2X3r3pfCOnhtt/uETY8hZJzn9HiIKnnjm9Ygs4so
9vNf7h+OdVpr3TbS9OnhZ8NJSJ/WwwzfIWPe+oHzzrgu0IgwLuVTzNtj65SinN8KGEOBDIpR6hdG
5dF75qi8grybuvJ8j6ZEbel8kKPIiyjKb6WiRyYLtkQkeAWrSQ9IL8G7lXRCLY6mqe3M6d3JjDQa
ZCOEFOXtusMjymv2ynP8BrSfJJZ6lMkFCyMCNUmNoLymPISnmOvi6f0G91XFjXR/VVGoUBD2Mm5P
eU0ryJVYBjFVc2Q/ZD2HLAm2dxb1xisFFiqD/eUmC6Uoxt4XXB/Fe6UqNcmWFNUAa7Phn50m4PeA
8UW7sRnZsY4VEZrIKXQ7cntUArUTwoWtx3e7ITRdYZWiWpDBWLRcvN/2n+Qvw8BggmicIETTfZRe
B80PWVWE4NpFg6i/nSp3gahDiuAcaJ+6fCE0qcgA/Z0cU7pu5EBnMCqhIRvBUxXooKOaxIu86RH2
nXvfFiGeHGAX56Px/a70exc+akSI3RSgJJwambBsKaVXqqZ+JcffbIG49vTAyBtsh1Ieokxd4Idn
VY3AKPals28M1OoW2S+BpO9HwrNZes1v4ocwk9aBMYWqpy+659NNr0N1c3GZge73SXeQdnvUmoRJ
w4P/23JewUpPRAwqyqBN0UOJtC13Kn4bVHq4/fwBTEBLdUwFbS34xFDL//99IG0qF1KWWo68Sn+o
H+eIdsARrlNM88pofCYpOF18vWveejPMAZ0hw4uw/23U1JtDY/bDAv/YrE3XaDoZkw5vcVnkR13h
b1BygJNPvGw/kD0VV4UuS6JECTpOHHpsIFDhBQUaFOXAuEG0vBPE/MDYGYs6rbmarNOKNe+uFoBu
ZFYzv0DZQZBZlw44zQyjyEakeG96gme7n41n7X0WoWU5HFjcmRmkBaZVbdTX9TlI4Gona2dS7Z1j
sf90ZXS1cvlP8QNAbekHlQcIJyWY9Qo1feAXSxAXntFmbZ5WDnoRqdfRu2r8BqDucO0xXeSDIe3m
LF4X8aZY+4HaRFypdZV9oKaFKp+W127i8O8GvCE0WPMOov+4jBByMGKj61A0WWE+7/tS5NJpOG25
V+54K0/J4/3Q3Rsyr1lbo2aCb+G4x5kgQkS3rYOmfD5SM4Ur8SGT+oMb/08wh4hRr/az1ESbUbpa
0FCznwEc47r1P2J7ku5Y/NFCHIB4JTPIZV3yvIox4ccuwqTuWdaUCCh8gWC93bD3ItG+6VZQDWNF
mW6BM27ypLdKIOx09zJ7gP9rLW+exO2reeFTrB1rsw320nnBYgxWzU29ONTjbY03guMJh9sFpmeJ
50fDKWS6x6WL2+85QIg59CjWayL2qdJI399HRBI+rhb6QtftfiX1806TEM3Nr2ozyv9qUsWroqui
80Nh+Z2QP+jr/iDjhy+65cQ+gMHp+F/Cr/Mi4ow+WOta/CajFxeEd0fJVtkYFNs88Gnlj8KPHgTS
3I+HtHr48SG3CKDD87GzBGIFnqrDnx0t1ZGnSOzDmJs4pdFtQBPlyLTtWMd3fyAtCuJQDxCiKhVv
4jzARYEEqeQwitEnkcOgbFxEwVAlVTQg80ET7SmJOsDiDpg6FhPls/GfxnlLmgbCX25Fl0DHE5kH
uZjmUr/AxylNvkwAS2yafI0izIJKOWim6+8eo8agSgedtevJdyJ4HdhCMqSTD+6P8cmt7rJDClxu
mlDhHiffFYkw3QvgMTNAqPGGj/kTwkJsFRrcMcwdJb0OEHOfq/X5AWWONuHnMJqJVjOboYxhbccZ
DWgTXRHFRi0KqICvEdY+QgbmZwYGhTmXykAygg7VPG2w9hStwve8/uEFdiX4TgLxd+zepuSqXg80
+eu7+PWmESIUJLQHHI10KvZPKJAOddlH7LVMleqhJx5+hCMdICwGiKt5Nur3FvmMabhaWFUroyaw
p8mWcTM8BVu3Vw9fLN4wOifEMzLOlgLt6eS1XMRlkoFoWHd5z5O8esNkWyGdQhI/wWj05nSNxu5E
wj7+grrGfv3bnqzFWa7FiaDFxm+2Ex1o3R2G0Y5Pv1HM3ihGBFa15Dw/uw1aHk4PJtgonPUWkseQ
piyj1/7kGQLSLFPjfQBx9SkjY+tMregtxLNwYGdQtD1oHj0kv8seobw4H9aelMdYmNweYL/k7gMv
8QB42P9wo9anbAdDkt0Si6lUs3bX1r18o10pBZHbJMaWsITXKkk5bn9dfaeEPWiXKbroHmygZik4
2KhGNcM+72ljdY6kJSMR8FaTzT9RVQHXExcKTlvt7tJNz9r2UrFMD4kiuiv2wfreeZhHrUG/Kkod
8VUKomNEh1ljsGN+b5jWP8A3blBq+9Bf3RnnyDQrX0vc03VLZqaDTtMmV3l6FafbPeJ6vXMALWlK
Ty3T+G20bizotp4B/2TcPoIPkeXfHS8MkefZMN2yWGC3yRciYqh4W9aLA2jq5dlzJjvaeJ6jHyEP
WBlPZez/qBQ8s/3+9A0m54upWqXHifqtI79tjpFpyKuRhocuvjKdLliGycLoFBb+5y5q/5sk0R8d
DA/x94nJXF6i6j1BE87cgmmSBoTkhVQ/shp1ehNLvrocI2m1ffLA9lUWqN1ljPKCZ2WUAKDB5Jpd
OvflRSl9gV3BlJtI2MYK1zLYcypeOql0II/xQNHD9r2FB9GmqbBnj01zImmAsrPqcbem2R9GbsN4
MJ+m8Ui9aVuCA659emQNp9VYKEu+7jbOtAUVM7ndyqMmBOo3DZuahFeJe61umWNt7zhmJer4AH5D
TBDcBtZ2Ifl7l8TMWVdvTWH3bbs4gW0tVbSchvl8ivjaxgtbpOSPYMHC+Nq5c//kNkvyDLaKI8M9
8u0lKWu7b+vazfX2L2kcRS5+vH7IpzSKt/CV0/E86a5xSv86ewtdrt1SWeUO01xkTmsivdXOOL2i
qJ/dpQ0Adbdf1B6/PFO9u61u+rufg2628VVTgwm666iuPeszcC4VnORDI4dVqOYJoTOaAseGXVdv
TlyJlCXZ7jSXSMbQqC60dxlfUMLSxArzmkhEGUjXhDbQe/h0VlQSVHzbMFSd8Z82VvTNIyptWp1C
18ckezRqQGAe88HEU0ngQqXD7h4HVKJRZ2yNUdekvOmLEVp6L4btnGvdoZ4+yZV5SStKqPM9dhOp
bN7luaHD0cTEp24lAUVd4Ga2ffQ/TRXE+7fNMmR03tVwfZ4xZACdLuXOnaQXVs5CLznr6QpdpIE6
p0jUoTxZZfrNEQVx8SNY0aug3EkQNefk9IsO/ggr8EpNwaTrGHPL6IzK7QhhwV3gIi7i+hqL8VKS
ej8x+20KBjKnfS1PVxasp7TMj4DAHTiIf89zfyd9Lkr/t+9xmvf10px6D7BPVJ2qsKKW9I+IOlz7
qYxTb+8xRbCXC3N22ClVp4IJ0Hmbtijwfg4kKDmTOeKKubVIiCfnTKjrIcgl2Y7ciBlRY9dTsbzY
3gHdnLGcoQF5IFG9RmwLFzlnyCCVgAEchj4KXKMNbf11uDMl0kJFAFAbIMkS0flPfXDGlXrInEKV
H36jcLFYR4W7SEc/w206U7JHS/n/eondVLPDlVppwxRlmhOq14Zeu3g/OqnUHUXNn4t8geDSzkf9
3S8PaMEgRj5LZkN+IB6k+llzn4IijjH+iqtAE8v1dQ6lNMF7NpHw8dnBY7Zu/PitqrBJqwkW4s9o
8v0a17faGssE3dz0ztgD3mHOiMvI01O2tsraVeeOyN33ljOkpk0VC0WYwBSlExR+fks5oP0usklo
0aLAJYJjHZ5UM/gTzZm+jLUpeHYex9Wja0+vsgHHT4B7ayOVRdM6g97IdAV82Cs8QVamUQt+PYMJ
EM3zmqZSodcVhy+gz651z6euS8tTGEkzEKnLubnr9OLdm0YJCc2nwVyB7KYeFSXPjf89rbbK2PyE
03zH58A+2hhTzkEdgSY2QS640loS8DJqDQKdd4ZJ4Ijp1sbeqTMpoRHphNqt6oCAD49+Bqw6/Nk5
APTPly0bYKgrfGGae+/mfQh8M62CaA0eHWqaF5VEsgwW7zC5mWZVkcM8wvztVFdKISSvqQe8l7JI
/NBF29aUsWSvRnQuovMMe+038cICu7r1MigfZXGEHDpdyIgRU37F1933JBIqZzGS5E5szSKJGa1V
V8DWxWtKu+HfkpzKZFDaLYnWwGjrFlvX9dEugOd1lACIbrZndZ59CB04YKRa19G9SEBmod/OIf8C
P8RZlbmun8S5G/7MxPQfZv9Wy5+/FymqqMize30Z4VYRnDmFqkNVjPsuLmD2O9Qs21eWnR50cdxs
OTPcF6XKrxTFt0Es7GLJlwXaedhRjTTmy2d3Ypy4BCuTEZ5dySiN573fvNmNbizQcFGx54lYWhDT
sIx+X2PLmFd4vGXgv+7CWTxutae/DQ34O/lpXfBMy2Ld2eTa7Dq+33WcymNvwq5TcdlfSaD3krVX
iuVlaJ6ppVLvgBC0eqTHxU0F9+XsrttUY8SwFdtcLrNks2Jz7HwfeYWVjkN01RJcCTyg4QFS8FHJ
ecn3ONKmqYQxBoOajzowLAsyYeufLh8tvEfN4wuRMDbam4uRK6087jRfTG0bqyEbcYA7ECvxpgDK
YJR/+hh7esOO8l/2PGbvFAeBJdpi2wsvzhYSpLCNF/WFGulJBe6S5joO5qFyj3ELPcOXec17Nhv2
HBNg5lzIj4/RfcbAFOx1e2p+dCV3fTima7hVx8HEMXfDeRp3tO5i439Gc8adCmVz13QcirI9eVfy
tqu7l1KECu8ws6DyYvSeisQxzcIvRybff5J1bq7sQ9TkxTZLrLpGQ1oD7tn4Ab3+wEf4SLSCzNQs
IozY8PkE8zEuyzthYB+rNYHB9DJFWpdPu/AW7krubI6FRsLxe4RA2jUa7qqK7S56hUHSBp2ZgG7R
0hmVIh1tX0p0hXL3IxNfjRGoOQBEcWFAPtpBgAOzsy8YI/a8WrIvRgeG9WrQtzDmZ8uxC/b4ogmy
ZFyU+LiGdnBtaV4ZZ2lSzQeS3+v3FmN5N7JOY/UmasvFnB2jkSXCupexo3+QumbKB7noIQQeGV3v
3xhlA/7Ykid/ax+PBca9mxSWky0Hp6H4hRun0cYEzFK0cSy1DOwrLdPbW8plv+fLgTEUzJwyjXyk
es2UXAg7dWO6AbGSHQ/98vGRjVnmjwrBfgUwvKTqIs2/OPpLXzwEDPK/4XCf4MGdpVzeq5YPBfDf
11fQr0KIvpjHMP6Y+C6X9pe6iU+4iHe2ddZuYrxeUjClt2wQs0W5F2turRLF+RKauqRcEJmu5Mi5
sMM6hV9emLCb/QuatRpczt8UgM704O5UrRVh/goYVbs1iUJ7fXK0gy3f9MIINqhOtnl1wJMxAaR+
AgQ2v6cY9WAgcohQ36QdIckIGUIGF/XVbZt4lJsMpt7sXVXuKb9a55HaIcs/6Tm62Q6nuc8OmurZ
8vFFlehjwAkBU7JWP+udThZqr+Ct0TFzJFM3q/JYv2mkz078Gzt4jMCVWF8Lxxe9hjJe1XaIzgxn
ZhUvrNWlBu9Ga2+wONq4eAqFLAYHpDsiqyKj+pxVPh/6ZVfJgT7xYX2iYyq3ZB1udbSdMoQFCB1M
R6h3DH7b3Z0BIGgcW+mFCnu34umhlsLL9QUIWu9YKI0iA1eGu0ObZkPm0+3wy6Fxl2jBDAJkzKcb
OGsxelJrBKXBdu0WzuM5opAwTw/Nr/Pv3LZqSsyvExqH23UlRGa0KEmrv2W3Qi1kA9yiQ0+w1btV
hBxZuiPYz/c/ghc33+7s0E1GECzOxWpZlGZD9lIf6nMwxP1qnqXLJaX6enViABXIISw26MsC69xW
wAtI7TgQUtdg6ZXGSkVwJTCLzlPmkcDHH5qUYUDjbddW4Xf5tHau+Ie9raF1DHim8bJKBDGIXNCn
Yv3DvMGU7xD0shvIbsLBs5bT3Wow7viHKREgokJpEj0we8wKoAsFGNRd4f4y8+YHPXkxigklBgw8
YHefLlVauvXbSJneGhZAAICgMW4xI9D/DPD9iVoRRH4WyFIy0r6E/kDVDZRVd+3jdk0H3NXCeHQT
dUGeX4lnDQ7tz0LjIbbBJP+RoiQuy6SlMMdK8KHTba20559Dh/an4qvaaLzoBJI3Zzx1L11PrSDz
JSf5yOu56wmfuW0Dt+AhSEfz1jemB94EVKB1CRN1ZRm+7zxoKQK1S7d5CDF/MErYHz8/jXSfZio5
QeydG/NoIbL86A+Dd2xmGHxnFGRxV+bapoRhn/TEI6SJPpgVWBdZN9tcFKc6UCj/lpNz6YRG8y3V
034e9SM8uIkUIq8Hs2wjWscr0Pp9S2wuZ8WNFKx2BK1QnHRBHt/WwFE5U/gTHwLYCsBDy5SRSixl
OfrPUrFZlEQYY2LvhTvXKyF3QBVdnw1H0a5HHwLHzyhjB+5Ejg3uVu8EHgH3ewNSQJRgbX3Q+aKJ
+MF63tWA5H4L2zFckb8jXOFvB2V4Z/xBA6j8z9IF8bApfFftAteZuaVOWOjl//l21OY3cKCrUguL
fuy1dKOD0BxQDc1KWJabsPQXk+LfcrWCcj+pol2LI9oY1de5xolH/oAi7tAm4dTVR3gcOXkhycgO
s3NZvQ2fEohixhOk0GLSftZiOYp3jQdZWboUpA0u+PgYONmwlQazlmm/Tg9jvvgd9oYGrvYeRoQz
Knesv3IQD+AHdO1Who3Tn6c/yI00cOXIWtMzcJAWiFbQMp/KC5kq46bnSQohbqSM0AY8YnRTta4V
hbW32wHT/vPUzU8Wihhg4ZDAXt9rrqhGRpDr83u1UBPeuWViFzMYdKgsOlH47FjufO37bGCBSjg0
IPW0p6PJHSRqhNcGqctcsd895DUz/BHRE4s/bmTjIAB50RjEP7VX5QHUXORlPnbx96i/LIhlzUy/
kd3ZaFRhYZaCtU1rHhrLk3jsBP2qy5OvZ/mZHtzn8N1duCF//mHsWRlP4ing7KsWfHoNs0pYn/os
JdwO4KBD3+ATVIHk6CXAtFp/HtVi6xrntV8YNfX/IBkSINN39QBDxdycHSjthYCXVgUrwnqMwZVI
exmaPbQcVcUggKLsrDdL9liIzXDdBEKwHldCd77D1AB0tNzOJqENPb5VBDE/BCHZR8NT3P8UG09Z
LS9O8T7Ol/ybDYquuzP/RVZsBYDcECpSpyKAhsalyTEr0keVXWwg5/rqcL9BzHhxcmxPuANMN7HX
LHmVavkMkwzkmyxbmY4qUkA1VmC+TXL6rLSWN2IJ8usdodhJwvRZpDQu4/nt4h7mY1e7FcNGG3Rl
8EM4ZtpWOdaz6mir2Xg9AzogJBi3XQySUfnA0/2RVhQprqqJDr+KL/nmWbMBDXDaUMLTampyt//g
hRCqNB7/EJE7BkhDR/aJbFs0TmsdRAXN183a+7CEEIdoAIMWR9AXe0dkIMagWo/QNvLuT/XVibI8
8nM9VXYjSGUUpNajLYcp3+Ug+LXQPQssMHAbcFiN+SP5bUM8QfHUijriRZoawqrHjyVlGFCUkEID
oju2KdqSKrdOf3230YZY8nkGZEn5fVu0/aR0tNV4LnXH+BlnENquNDbmf0y5TlNdv0+iAzHpX8YY
QGwVGR6P9vX2U5CVsBBd10IWkLAJLgLwjEmiDfqFc5RPom/huP+U0ysm73u38fJ0w1qISKL+FXwN
r3U3izlQSXVcxk8gEtMZkri8baEEFWgdy0H9wSLk9yjEkTawYFPslqVnCGvV+xg61gJS+11IbENl
24lwDYtwp3aGGSi4rOkywM6dtb5uYHnTx93NthSYA86vXwGiohDKFzTIdz3XLtXs9sIQUocxnsYr
RG0TbFEJVWUaX4HzlV4UJfdEytb0lVsQp/X4iVxeR50A2n2DaN9WqQkrLXFCyCu3ftWO4DlR+Nzs
U9YODvYeW3K6vP3rOjMWLS7sRqF5naHePFehrNOhi6G6ehgIVDOJ5JalQCHZo+YCmye+awKYm/Bc
AUiy8kapAN6IuhSnYVg733+rA5FcqjWG5+otHnjR3zP+CEHxDoBI6vRGXXM2bZPiRVzS2BVaXmAO
EayGpytSP/0X0jBYdTqjKuPXN+VIwTd+rS8TSRTk/OZEt547LxBeYDMmj6VQT7OOL/xb9gYTBz5C
g2k6E7c5hJz01ot2PtcROVLBSF4zijZ+4cWToEFOJLqISk1M2ysDzlBM6TeWgPWK6u9nDqffWAO2
g9IyIxVs5OHtLp0P9HWqOv8ZFU8I503pH98A83prbhh1LJ27StodSb5ETNgk8/dcyLXtuX2Gyyp2
TUGGvt4exn+d0rmEuSqcvVzc7K5LH7RvHb/+AKCHZ00RxhgCs5C6jQGsxgrgKseHAN3bzDLCO66m
IGpELLN19VeHqnqtf1ShWnvijcZ+g8XQxlXZN/+btHxyoNEx0LvU9xmR0bAESdmIPjpCprXkptOf
a2HPa1hvMkTAABkMrfPcaTNSh/fJgnMzR28jZS1Y8s3XOcACmIt+pQMN6mHztSHEfMs6IJDLvDS0
HHtkz5gbSyOeuHMXByRXQki41sSxnx+XH0Q4qWWDHh0RKTsGM5ztd9loyB662QOlK8PS1EPEQFq0
eiUVf/65p8ChUP9M5e8FdS++xmYdNTYVZ80/X7YhFWjiNuicSdvhpLv2JAbogBVLOnI/KAvsUTHN
uUDh1qS/AnuDa193nIiio36Sg3QYAqMizF1xAQhADbENqsyFK0ajHBaCaJRMqq37tbLXb70nGh9W
qDmfQ1D1eJwWRL8c1Pp0w+zyUkh7g+y0EXd0R2wXHzR3ASSN/gfwHf52UtlOqwcSc7rwkuXf7s7S
HrlTfMs2BmdV2vsReyRlZfkyDXU9pTUppG/R8hcqBb/VocMIRsHqvc1E1tZYoeHPkhSaxSVIN+6x
3c09H/jM5NTRkeJb6KZsXjptlRS3Ki3HyTPt72yZ9DwZNzqMnYvh55mr2fv5yjPN6gvlhycfLnRE
KlTwmk7v7xKbW9gLsu4UpIseEkjCh/ZYnYxq2bGPn3yzh/Hmrs6QHCYPijofvpqemaDLY1KuIDBT
xpt25zFyMU2Ou74wJu5DlYpPeL825DqeKpcvIpz8U+19EVD/Djyp1YZ4jhPFV8coo6+UoKFMYa6L
MlwaG4iGACE459LjsNXUwAZ9P4C0WeVJGnXy8QUwvAjUoHQCbJJ0FDuxqEIQRdfhq1DLH1mZmyBC
pE8EyJU32M/nWkOM5hrI4cc20GvaVx6tf2VjSFbNKKIPmAjaZz1QnYrtL8wokFU3uWPOOU+pn33a
dSMuY5XZR4I3oBzhskT26n0Afe0/GHrU2fpxuLIhqnX6zT7ua7d6YZo9ozrgUYh+nFs/nFzo5RiW
hjXlCCvXB3koGaYXTEOTvatUlakNrSCrVRfzb1DCSGiIuOa9tDxTaLpszkCEogOEvlfFD/CDl1Fx
UQogtPEvSAHcbLEI+EpztHU5WUOvSQtVoqvwrL10V+9dqeQLQm4tMF6Mu7BLoeqDwKRtRROd313I
Y3wOmkyua4dO9P7EPDHGjaSfYgHHvXBig4S16npYN24KMCxMLR3VKSu96WAX/1lFt4bmjzMeVmND
3QkeZA2hP1ew0wQqEEJrwTNkSeJ2tpmbfeUi7O4OEUUKCBM6SDdpJO1kg0BOjhw9qTBf/Lj9DTnv
ElH30R3c1V0fEaXUJM2ln0B8uP/eT0KpLHGU0O5rXN+NhoJQKijiLjh4PnG2HyWu/s++2dSEu/Mq
AvPW1NnRipi+Fq7U95DAhKXE3lPRFFqea0kwwsXt3vMfWeBYzOTIvPUO0NWHFPmEjVTSbvMXANSD
OVpnnX/Wq36D/L/s+5yQ1F2FtwQ3IqFtLO89KlFS8gTGI37sB/vrbhkXRo0sw1Sy2qd7O+wABBAC
HGQNgblaJAnWPg5Ann2j88lO0Sr687SY7iU+bCuPccL7ZFP4Tln8JuItsWdJCHtaN5WeizGFLLiv
+s2Qn/H04DmuUnkJiyVVncCvY2dwbQPSxq+ZwyK37scCjedDPfYn2OhmSDz3k1LyOVMHAohvwcSt
qdfvJDxdnANG2TL9Q1SsFlmKJLE4qCycbPpn5vCoHcDiJ5YK+/4+Z2K0SPYI2D/GAMWA2+vcqXd2
DuSVJiuWENZdWqU4O/3uUxVKM+Cak/L7akzjuGa5r8McSyNvU1C0Itd5tN9kV9q1jrDVtgy6gEDx
w5uSIn+KLKSkmxn/E4DYVSPDP9NZUlxCZdroisEpL1IprnomB9PXpgRrIdqEEBbDV2PsMHp2XfkC
LumDXMk4F0yk1TPpmCPdGmm6DtSjv8m3n/yTv+nawLfch1TGo+l7+9c2vs17b38DLBcPgdWdr3Tq
BOhALcNlKXQn7vw0FbTXgzioRcfl1GtHsdZdOnifNEavnl0gypk0lr3mvCLu1r47AmA8HRf9uxQb
QjY0gfB23U43q1LbXQsaKJhhoxeOB0llgyy7DNZSr+1ZQa5uTHJmcT/2xE1rv1yhPAkueHsegQBp
PLcChGJPxuFqGi02eLxSVhYvjvqStR9LVtOr4EW/iHmgDErgFjVGzqgHVb3mKNd4ermLG1Je0BmT
UKJDWg/V1JroEiKBu9Za/3PfhqCXKgkb87Swiwiaj/3TcKkFW5cFU4RvziW3i9A8COOA7tgOh9eB
PPHzq+lq9sYDa+WevIn4VcnMr5nWUZMpLLUxI54XJYnqlp2r7cHLsDDYXkZlcgVW4LIGeFViP5G/
xp4Qs5XHozRzmUlm/7VNSoWjGnXpMI97eufbm5g0TV3AhLDlhWA+o7iUIkJjIdE+KqffPPc3Yqmv
od9WZ5BblDE5QiJQBBvdNCvkI6/3pwWTznRPVvRLYtp0MO2bNojjgiNXhq+XOgNsrg1PuCFkH9sP
O/4cz1xaLLLJUPujJ9NVwPueMnugEpCWItrA6QSNk7wxPgxzLOe4oWZS4ppYqf9/wcW3HTnfierJ
APCnY3MPxRPEg+6sSOU71vPh9VOxCvAx7gEDqbKfT/L/FRnLdE26XGJxTz1PoOPC0EsaUrkRvC7/
hUjOqqQLECNHVSPDqm3MYKoaEXPVIz92ojorZ3D2vP5u4ElRDusB9+6UdEfluWQh9mG8XZQ/WxuT
HO7VxqwDnCI+2uHqcqLhLdupnQQpyCljU0vfhBNF54Jhfwao8BwMlVNrXkm8z7z+cSo6CmFq4h2D
MMzB7CFkTr+vIQrCWs3Y6+fjY8W/JRh/sLfTc7b/7Tuq3Id5h/PQJTL+fNo1RrqRkpEkFLoEfU+q
Izi/oj+k119JHd+2dyRASHF86VoLayjDMuUNjKF0e4ZTx9OBq8YXrw9cugq/emDhhgtPRKS4b5fL
bk0ynyMyg0idSUHe2VX3MdICT7szBpS80DndxxDxPyoe9r/aGpd0dBF4mR+1xqIPAVyp6V0OWgU4
7WKt1wcaiN/BCeJXKE8xGrsHn0PpCw9AGxPxIFOnT7k+bIYLWNKPP3VqBr0gcL0jgE8uuYPAqT/O
MIVYPqfj3CIca0FG+m+oxokPah0vURoZ/SarhZZisFx4LvgxXGt4jTyXKwlDv8wQvIPjvz8C5AMr
+6E2vVS+wjuGFnSGCtO4waVm0qLIped3NsRRCgDtCcZiIZlRXqwhdd5UKZVOpqeQKY+pWm1lUT53
6zVyGgatfcMfBpU064kQkUR6TUEpYcO9BvfUMLZal6RX8znqmNZ1T6WfWkgZzHcn8BnwdYf47iFh
zMe56i0myjEGxZd7cr83U6IGZ6MbnHx2xrRLqt4GV+E/eU1CLHe0LHa2qIQgUKFzJi+tBbnGHv5G
Hyh6L+9GhFrdzp142V+3innn94GnUREFsTPm6TAPV4CvjKTg0Q1Vht9r8B/ANzSN6b+rmDpWuuJi
WaZEPKDq7uW7FTpm2MU5EIcU4cSVANIVQbcWltUx+MnfRAbk4LbMf/YGwrr6IIGZIXuaY5biPVvk
V2SmAS3oEie6JsGUWFJlVLrwYoj5mC0WNnJ4albfrNRUwenlwDLigKAXqrV9hBeA7TcqY9nVV2cT
eJ8ltHn2cleudGYQKZ/wOre6limJGxAXHVfcrrY9erVJTUJZMmOwF4q883nE/9MxRk6gtSfjrtRj
GzFyxmI7jwm9Z+B1a1482Lt8GAsm3STSroFGvPiKf23GoYFrzjUZievLHs6ygt9ND+ysrPb8A/4Z
E/pTPAjgcl3hRvKKkWylal8FXsXFeyCmvLd+dOuVKbPox4lxZL8geQiLEYlJlrlwuFQVFa4eotgc
/ARhTof6oMJelcbueMuP096X6gLAYv5nk+GyT8O7kWmLGG20W3YZxz3zwr2pwLRzp+96FI9DNb+S
7bzdF9lcByIv5eqJxGXSkZDFY4yQZQfFQNxkmKmikivHJ5ttfqrzKRGojjz/L3ESjRpFE7/9Osy5
aQuKpWxEQYUvIBaMJwzRpd5Xe93RQT7YyMl7tIhU00aQFYzbLqB8ZQlvyUUoSYII55B00p+Z+Yte
aUVTaTevhZOO6flXKjSuQRCjtzSnEaGgkU0nIfCTZ3A05oDMp6014RZW5pNvpgK3R9z3zYODYxsC
Z8hbJT3s4egEyBqyGsXzK3K3zEXLVk+RTigHzA9vmHB4ZBjrKjhJGMRIsiue9uzeQhophSjON2wO
e+4mbiE0hGKC+xFP7rZk/zmkQRfXLvlOiU1pIRW/E3m7elKbuew/xmpmSJft5QYYzHWfxEOu3Bu6
VGoYAw+ojF+t4PSTvKs1ghdo0IVeBD8XSQ7ayDsOYeZDVYWt2201a9oyNFEjEO8mwOGk68ECnVm4
QGWTFXcvowwHXvArHToVKP1hEvP1Wlk24iSoxlFSyM2rUOk50YeOmM3Ov4urNUQjQYBQeSW2Dq13
GNmxBILP0Een+GfawojPUAIAZOtNdOzXpghlv3Gbwpng4qqntF+zwZr9UHUPIzlHVisXJldy1EzB
6psofbWtAuAxwxJsYyEb0hZkmLLNWqqCOPWhfCYlyvvcT+KRAzvKjY7sYk7MEPwaEVljdEUdo+gs
Cx4WiBJgM6B/UKGsEK6KieQy5NlaBfupvPFswspZmzbr6brQA4qejaKVxPMxqucGX5qz05wd7JkN
JEyfI5aQL+28U1OYNIMi7s5TJQ4mMi+yaJ51Amv93oeSW7eKr+Hkbi+MAQIO8IXmy4DeBKz7NuVN
rwgO4an11tYQAe2iBEpZLcCyzBTjohJFrODSmIAcE77gNjVKF/DnL9nLcLEIwBiMakPQB+WpZWu3
kcfoLx7AUFtfYmjuVdXmfo2YtUXM3PYRPKEe5W+6/OirNNA7zZ8Mr/7KXcWLBG6zleXj/kSIjMHU
VOggvbUWRrC4wfDXLoiG+3i5eEO/LTUOphXMVtjRCS81+o2XX9IJNkHm8O9DVZhvUsXWmGIwg4p7
ySznq3hJUKUGxGxsCiSEgplxe+JibXDCH6igFIrqo59nC0OSXICwTbSwFOLa9+VY6YCQYBRgS37Y
amhTEZwlLxANbFmglHu3fr3fply1H0DLFxNem2dTNMhuZqzGoCLgYKWzf39LQA00VZeRC3WghZqH
RCiPjxZXTlgewiERVkC3nAO2cvABcF+dIH5kr0owCPTLNmYnLklD6E3VvU7N+BycpkVHvu72F9Cx
FjnMOMtw1ExTazGIxke3GHcADsVrfnP5p/UUgiw2K3DjDqLqcs/4zZzynP881PAhgzKU93P6lOvW
dD5Vaj/Ep/AfGGOlekNMoPsi9wcMne7s2BfdIlnP3YbYbyg0RcWDoDROps6yk2NsE0m5nuohHBGc
ggRyJXN7DODrmrccrz5QrjJV4CZBm7yxpxyX3XzB5n8FLMqkgX2wn3zpoOzt7X8PDxVqPs4ptS4Q
Rwch5sZwnG6MKAC2Qqy5QZKj89cA00fh94oKUam+qhMlGJGEtv9nuI03JYJ21s//VwKUvo3k8StW
R+neeIANDtmtQJryhM6/83wYOC14YzPjMVGIJqwZhISEA6qYa7Np3EZgX5Dm5tBgDvhOaPooqux3
UVd1wRbfGnp7U3JVkqvoYGLsejwDmo9dX/3+4JJ0Jn8xG1VkAGolSM2024sURJ90Ag9JK/CVEO49
OiqvLywfi9+x5gmdFdllhqqnbInMxsH0wPSWziBCBDjfTolblp39Y7id+W/oRionrriBIQQEPKll
qiJGq47KOQyp5VU3WJZ8lxnP+okNXqc1neEC5Fkh9iYhD/uiFBS1zDnpUc+rnmKGHJ0DgRjUTka5
OgiiFHbyXRzVKXEDmHiCRUsZfEXgBtVFXV5yW8Qf23AfnIjjMIIRUGjOxMzbnBDMo1XVYu+XUDoQ
2pk4ofi1UgnWFGc+3TE3XldkkjULuTS2HvSIweWYfbSEG0+jDzkukDYj4nsEk1At5clpe1f3Wl+Y
3ygpfAXHkSbAZwdmDd2SP/ISmWeihdt09WTU1WxfNn1tZ1S2zUm/WS7n+4TwKPK857gws8XpwxID
miHYq3rZjKxGyQsFQSeAbkJgWpCjJhVFpJJEw6ujEHIrvWEBtspZ6hCIlZaOZqfp/rj0z6p45r7a
8HNSg0pmk2RDwQAjwM4Qa2cKzClS64NmJDz0n/ymYI5LTqm/8tl69TMFitcH8tE/1oEXUkNigMdp
hHwqJ5KhmtQvqKGIlfaJF3jtfLZ25VmE+Qbbwkc7WlG6vSXz82+CgCz3BQuG4oLcM09tJ6cTBsdN
g3wFLkVLOOx8fMPimcnat8Y1Gh6UwybHwtmzOot7ac7BRF4QQxHKKEB4x09jqOXkC/yMVWzJ+GRc
ADLk46TYJgw8p73EaiqHDpSzHubNFhTXy2a9wu1R+VwLhgeclPOVAbWl6PGqHk00L0yswqvStmJ7
TVyBvHyl4ykACCZ/7UORvp9jj814kTGhvt+IO8++3RIso/GNtoroogfvJYI8412rL799Z3jjAVoT
ORXX+HN1sXrZNXcCFhUx/wRds87Rn/asabxm/FQnQv6KCYrMR0Ugt6PNdMTBWfXZbZhXYajzTzA0
CxqgYIkxGCkWNUfRzRyz421la/We4n3NctDWMcqpWnCX+K4bkaY9K7YqBIyCY61F4AeSk7+SGJVD
f5eG2Z+PbtBNA3gCzoDnClGBNc0+injfXvYlyr94ZGjpNInANG1r0cWNgusnJ7V74HC9mI2C6V+A
DimdVH8vRwPnhRC683JVtRM9FYkhxyQsmPM97oudlC/kU6hEy24V6DF9VrZC4yB8iJOtUOqln0mA
eRPwnPK4s5+MM/E32fGyf8RXWI+bRI5U9H2WWHgTAOYu/855nzdErIVUYGCDMBKQFwNgSdRfJYof
+srU9bceJ5zAfgneVlaJmtH/ufnNotwkNTG5bSngdievf7rXB7yk6Xqjin+g+Rt7Fe93p5jk99d5
x4abFfjUGBVvc2nEfnJXWxdyCuZ2JC0OvP6KNEeRrJ7NIKLfgpf/vUGhHWbbK4ZIBQJHigKYRKPl
ULSno/hRuf6ZMNSqiD7vCnh087OQbXjcCeqsCosfAOSqLcWXWuty7AGR+S9ePcszDtfjOkjhYxqQ
mvKxRDWfU5Sf7Co1US9tUYmmxKwpOE+2MrC/HeUhAKW4+XnH6ac6Lx0ybhZIOwmlzmNWvLDPj4Cv
s/TWxhI213Cko31GsxV25qnbrp84vYtkrrhdTQzZtzCNcws2HmPhNt9KI0xpEcGLJrDJeUJqY36f
oqwVGqRlHTpND6jtV4XUXsr0oSjJ/U+hKbbdfMRqMRgeyA/DZhO94v7LP3sujokjrPs2HhZGzBol
EbjyVbgri7knoUC79Qrd2lyP3UQe/q0gnRdihefIwQ27WVQV/rABgoG/HJ1fBes//7MhQAQHMW1J
PJK2dTY/gUP10JPrBXEeyU/dcH7MX9jKi+O9K6VYcW3vQ9m9syjgC4VwYcbIJInKt8YJSmcwLq3h
Tuay3qk4EGjkvg7QHARRqvliRao+IkFwFEYdnd8sRJ7VFr/PgyzhBLwj+57G1W2YUsAbzL8ah3tl
yfI25TLIPqHfEs9GsyU/azjIuG8E5qxOKSi5Ky6GYgj4xeVGhYBqcJSKGxMRzHNKCISI8B8m24Y3
qoNUa9zVD8XOglps7zQDwGh+OdWY5rwjgDaBkHWKHq82ruBNhxAhKQHfIemUSnJbzI7wAK9hUa4A
5daKJXTMa45n/LdCoNr2kZRRC11WxXu63wa4LtvAw7AEPMqKdm0yR92nB7Dn6Lraw2BpsGxFYBJN
8d5nDR6jNzOEtoSrvGRI8Y2oT2YRBFqOb7rlVVdT7squXP1JuZleh2fyu/tc8r3HUYfX6S+aof63
Gpe0FBt5h0smQ6qM54w3HRhFrzu4Wp/v2CmCdT4vuzwVmzijf/QY8ueleYnBLJHsdFqeqK+XuQ6m
6sn5XkPloJU9V6j4wZsvvThXV4r0+U2xlGRA4/GTliXvTRolpb67e3YSuksbWUSBKpDYOm11nWyy
+LvfpMm5moMrJWE1P0Hk36eNSAzrVmm2F4gK4CIcPBLIBF1wb4n7vUGZk+PP8hUp7BU5KKa9TFkY
Fk99wv30jfpkMtbUpuJ3p4d9g+eeigSYjqA+ZQ/8KcxJ5ntoIsqpWCyxPshQQ7U+2k8LQIzcdt4i
5nYfBohS58HqbJaKf5UtcVBM/7BT6O+v2Md7R5oDsGN1+k5126dLHhxdTesmDAqZHdpCPlEAcbNE
lhCKX+Eki55vei8HlVFNhjhoxa1Ust51hLhdBi6yminIYAd1owRlOO2M/0Kx6QC79wZw6Khm6LaU
6ODnepIZ3omZ/XEsAfA5p9QUehu4XDDuPcrzvHdqtwp08wAa+uqhQb3dY6L7nj9e/9AuTLxzFYn5
bK4w56Voc9sUn+urmBBs/MVGWr1lL1h2kP/qYWf96vYMfye7HKSlRlg0xc5gEGMPMVtUBhUZ+xMA
2o2FD6hLDopJSaPIortn1/a1hNM7tW+4dGc7/dzUaN30tYdDRrlEz+sx/B5jECMRHnMkSohy7d2I
MJvk/yv32C2f8gve6YpdXph/H1KbYMJJieLIZ53NDXC7S/nkKvVLor4nepGS18HrDEFN+yGz11u3
g1//6NANZlASnUl4bpkDPLBf2HVITE5L0apmUzeGOvuH6N4woNRz5XCHOL+VG6O7dfXCEurPWgcT
2ZSQp9rHSXO8ibuaEQyhyUv/oJfWu9DmIiGZCkEN0yKIL8m591y7pTEuI14Q43Bust6jHa75GZnh
Gbhm03J8sMxTfUQ1zobHyMnHB9E3SITMuIuhTAyx/tCrkz1oIT3w2FcVKdDIPheszTSNmf6YG35/
443dI6R0eo+MuNwg3EWNhjfdvgEHSNRC2Rc8qZpleVLQl7GzSivvVt+WKszNibs7eEvhoHpYL2YU
6F4Okl3xDdj34h8sCnmQSYBElqunLTcGunbOt7anTUATadDGdFrfy8IjzFsI/Wzk8oOREuMaQB4h
DlYBrF+x3KVclB6aJagGrFHkrDwSlcCNXC6vEaikfgjab2h4QfrcKorBHh3n1g0uCmX8VrePFLyJ
3XFUsrX1MUhnmv2ct6fdPS+I+Rn6qZIRjgoqhFmL48aVvQqGMcZ85ZRsssUdd3q47GUms05yfY8S
a6YvgGl36c2KEzMylGOPP67Yj36bUUedN4T187KhK/ulvWxxj/Byys4z7ivJRMFX6JRKrcSltrQF
RU9JW29Uel/ZjG43a9MPuffITAt1FB8pULgnKkc+aBl9mOrL9lTWZG1Vf40opg4foOtuOwA2LliW
BbKmZy/57oK2nr3OEQbfwqZMNeswdzb1IJ5RFHZhvppfZEafmP7Ml1zDMOAgASQE27RI2B1kslD/
gt2Jxb5FIolAaayBvcWE2dv66xK1mpHKlXTOEWLXSRs4+gMG+kAmko60gvgC1eIB0CzQrlkcXuSQ
gBLtiX4xHwEqUp6jnNtvcWE+xv5byrHXBwShjLqduT2yWEinMC4KNnjk3u7x2P4rqRDfYztLuXKi
7Zj7Y10Rz0I7Jvlom7sDpPz3K11EO+RI1B9FjO4I9ybneugPvfclRmY00gE9zob2m+emr1C+zDDI
ufs3L9H3Sfn9un07mwqBeDCaGWiZNHsUztaaC0wmaFg6PFtP/raj0zLSK73CS5lU8cRhvDpIFUdf
mvhZvQMBePVDTeGI4jKBl+IxOOWQHiD37NlpUcpMluBIuaMITJpQP06CN+ViOdqTww/th3Wcvpej
PkVbUyakggJqH1458/lzlr/Vc4OuY1SVfpIUG6aEduBfCIWAwdR9bcEB08PNSNuPt37rizXKZG4B
KwVQSzR9AQDA+wVgkR7r2QubSnkYIPz32WgglqqiwDoaEtr/cJm+qYdNN4EOsN9OcSFRXINB8JjU
NdN3TLdR0q+8VbZcuwM/8AX4ShQifFdo3XnAk4p9d0zifRi/JUNbUYo6++mN88dR3l+1ubKKS2Ww
gQYLH4OcHS+Eg5Qn5wmSFDf8mGLa5pYSiaXfXAOlL4uyeIwAr+PxHSlOPTDXCEdqJC4SIxgdLB2O
Cnco7uMuuTUVzNOxLCPi5yhN0iYaJgeS5si9yPazzQe8UGONt6luYtOgefObNoLo/4SXNQyck/iP
bKC9sto9y4GX/6tj+akfcsRFfQa9YPmyueyRxm6BNSsFB1iTnBzvx2m4Z5mVu65Iz4h5bZDnz0bC
w9mXStRHCJyGIg90ZYUdJcDBPSdlUug49kxzkVDtjmaLxfLiVgvzqLzkGkE1OdW3kvGyXtgoZiJK
9GZpKslmgmSVkGb3cv6cF7JmVsnSEsrv6YEgB2e0x22kQgtlEFYR5juwbyig380THY+qjgwr3nLM
qOuopv9on80dVlKhhp5R+HdGbRX2+q9GuREW0s9oicSYt57gjNGtzeorfDYfMlJKkacQ6PE30xRJ
vqVDkqfnR66J9080+O4kntYSJHtMusdxBr4ySVXDQtaX9/C/u3ompsH7m21u043nElJW5pzgb6tQ
BcN9XcOsfCE9hcskTCTJS56Ia38L0UfAdvGWHeTnEMVpWfxyw0UBnKCwL0uvq49AEfw2sWLNuULP
o43dlRSj5uCA1AzjZ2IvYa/qJG0Lb38WRtoFNYrAgUn7mOVUT3HmLr9Rtlq6y4rbQ1BRHjA8kLh5
4ppdQpe273vDLJlACL2dygU8YiCuOtJwmQPwQK6pdkg4Us6MB5VsGQ4mPgZF8Q8mSy2BKskcnxVT
xv1dNqvk9u09icUVZzXdZkNA2TYyvY6MON5MRRV18HB0x5R7ZZtmFkFRFE1uNfGmNgDCmj0adOfU
GqQSQilGST95UsSllKKNHYzRoIDNhIpdRGifc6Tfaxga6gmy4AGvyx9VlkiwmqpD5SYWx4hf8iKo
4+9vPC42I3fA0KXIlwhEYmiMJHVdwQaXEhOSFAF8iUDV0FspAxVHUvcLlmAuaObn6UVGiyg0/M5x
Ok/BrVjvVL/pMX1fm4xXqlebAt6E7PUqWaoQdGof/3km0XREM2iieqjn2p1m5WbkYjdiXLGL2Oyd
/NIdbucFK5E6yFUlaZkz77uSARsvOwoqd8ool8gI50C/I+cp2O+AMxtBkp4L7QDrhTOeOXUcugOo
tEI717YGsePVpVQu3Dp7xO2yEibvfJhXFseFS13YM9071sL9a0mdqtAjT4hvCYWypcARIrfxwvnp
49NKCPE0lCwf+r80IS9J7DCko0cvHxZmJVybVHpyWKh6jxf0N0C6MMXJVfTWvLP3A11dnHdMvIW3
Tph+pzZISC2hrtXteFGRBR8ajOPQGh9gFWUkvZf/+beqNqIrpSXUK+ek6QZKHSbvJVM4ebvRdr1r
fNTHKuDw9NQ27GgLrTrUSBUfw7y8QeasHuIMUNbGuJ2IxzDW6RH7BO6h9iddOq3j1a6IXMLuzrie
H2ocMhpxfLNFDwdESOEIqDD9nCXH81v6Mlaf6vTnUBrRGO5z0fy1afy7t78dKpd+YLO6ovMY7FlT
Y9USvF2yGNM9FaBPiH3shKY5XsSlJYqENTVTrSriNOa6vokMdZH9jNibxO1FaXgdKZ4kmWu+9SQA
j1Rh3F+RhIMimeRqR9EYVI/6eHzyRF41TjhZGohqssRJj0STOm3YjUHJlUBlTpRMnW9mLievjd3/
5KTwbNJ1G68vspLoKeK774t1GPL7HQJoodHvSNXqpX5AcOyJ98+yyXTLWu/8s7558XHEndWLSZ8H
xN9V2na6+6fDAqDqIomQajbLZxiT2m1jpxbgC5guyQvOA+MDILVKl49gxMqFJdfHoCRk3sqSNhOX
EJoqoQRohSvPncoxiV1BMblaHq5GMMxUtcra2Q+X6UKhSazXEwswTG3OED6EE9WaSgO9dplE+83e
LNbgnL9J1fP16fNrAMLM39W0D6llDs8B2h8zqseVAryOjt772eDEtAws8BaQzyUgdufpFYwjw8tf
NWkkLzbKNsqX+XpUFTJroorRKWVXSkk2FprsSQnk6aBkhtH1U/N3iIG5llHedtXBdozRrMlLHerC
tqK4s7npallkvoaRHfvzqyd5IbhWQFGnCM4aRL9U14njKPippxgKf+u1/mUzB6qoPi9hI1jg+4a3
H3F15fWeuoIx+wC0xw0udo5nES9/1VS8D8UVeeakF0ZphAKfbw7lkg1bmRR1GybKmZHU2VV25zL6
BgZsKO+/sgBBbDKGchSuPAqqiAt910HFAt/XIQpm/L1qsncdwhsIzBDDRcPbR62dhMvpNc8Ex57I
anU5xf+GcUjzDuMVmz22o0Oypaqouw6/1GrxBuZkkhiNG48LXjpUz4xgxgzST2BVDJ5qXX5BphoA
IgjFRlU3AjnBDn3p8t/Z/61PRbd7vd7QRZCq5gRmFXaFU2rGe1fNxirzF7A35moo+vNLyqnClFCi
7YSWtTXNd1z+SFQIwVyQxwbaLeAEV+XCeYTvASfjnzALG2eZa+BpThGq2rqYYzPfD63dICMUxWYn
QJAGkaw6G5CWKg+z9ga1Yn6GwwoqMhsmF+f0JVKJIQRUZKCZ30Tlv3+zuppYi/ZiMHjoxwhcdYg+
CCniKR4wtge9eT1HRmG5GBH9fwrMmTWqVwtHY2OgmJSQkIss25ZKyKsPPNKmZVa5wjH+QMS+DKtc
X8WrQR/bdOJuOKd/a2LsgxjQD7i52uqQcGFaafRoKZ4JUgX6ou1jvuFejOifoP0nbE9FMW3dCGmd
8ZOxyB7Cqn0jcmMd4Nh2BmD1IHHau5fW6i9iSRp9vEbMDNDes/JuMpxfWDBqX2kNm2ejaM23H94f
1BrnekoST8q3lFBxUumcdtcnotnABrL7umBPQlpBNkuSopcmR5qeEOJhF3YjzfjEQTGCNGy34Vhk
Hqs/ft8W9wFgggBevgF5j5ABZb6unR/xNIThK1fbogNGFeKsKB9vCq0VM7L7T/fWmbkMiPe9LSv0
dn9Os8TTOYNqXfhw87j2Gx8UhUzOJSFWwKgH4VCObQvTJfE+T6CV5sByFNZMKGPK5ms+lVrBX6JW
dKeiX7lfvk7o/bQvo1YEcKHRE3c6k+gq1ghjUNwyxcHZDpnq65z00B1VRQjULuFi6WbjZ35SXJ2q
EraGfK45LpyYs3/PEZkLq5R0XiL1OikPYEyKED1dsTOBacxHkFOA09dBoeXLRKA2elL+C8VGixCL
EsWGUsGlWwh5T3QfHueqhVDVo84g8zOqKeXulb0qU784QWm2VroVNZL0R1Q8QAk2V2no2dMJEWRd
0qZ+rzZstUktB/X7sz68E9PM8Tm6SBj5wi8D5PI41a1okU4WqkC07McOBYN41Pn/CuHHqlZe2Lq9
6F3cBWWoBTbRNwAMwWMEusUJHnJR8lEHPxsOLedDLYUF1lzU2Ke4blcMmzy9Lr8U7iB6Ydozeocr
XN7q+/a4MpltO6NxF5RMJ4wm66SI/0L1ERdjknemMDOhqxzPLCcMVjy4UKoMN3FAVX8c7K2alq1K
V7FzOVyR/UnDqQAB63x2jO1dnluLHc+5fuN8F0PsqbB0QoUIXb+S/OLW+CdccR6N7wb7imRgyGg6
5wwU2GfAw5spJ5neAMgeqUT5R2sWZTjgPxUfFDS6oyqG5q41QznAxn4bTFn2GDz/ES3RAEB2V9BB
+t+T0kB4sam5tNr3Ows0PgFm5QqMCovQPogVqyyi/ob/xWwy3KY6s5fUAjtVLFsM6yneKsu0Ed08
bvG8gcpcrDRgMbYQ1e9wk0jCl3UmG0Zo6r5ipvbveauLzCg35gkGTHO5OFFHzd+AHvb2L6GTzUVv
MkcYvz7c+jRPuNPnpG7wzEzzbCGFcaYswOuGOrldD/lfIDb0PRu0x8jkOnoxc9cC8XaS32P29jVm
Pm4sasoYkVJMEd+7k7vEHrNjXFA+XhSZ410u9IHUJ6zPXpZZBmAbgQ77ANjHxgOXw4n3NMOmSdhT
sjcAqDbPVZyEQIQXovlFw/xf65/YMjFcM38monzXG6cIXuK57oGMLQdKwluYtNmvJul4PPFxlyBu
jcRECKBo+GhH9HAtI4teLF1HThHyoSyoTRHDGEXS7IxtHwBG/Mfw0AfAGRXr8tsst668/q6BwdQB
mSKhZkBizzP74FNLrmh6ApzE/WIl8XSUlWOvg4A5f5cQyMF2L3BMNLWZTK2sCgW5YfSU+zHl67NT
9TDy4E5BzLJqnGsoD+s76Y6GNcA8XpKsL9hzizpvf+Jt8qrUStiox6oiec1F8S8kF2fBiB2BT2cS
nGy5oS9oKU8ocJMS0mU0Sjo4rRgrV2FNrJQX8+PQ69xav10BMG2vPkD3kV2UeLRn7AphDNu+Mp/X
rPEcTYtOG2xkMDTqhKikCQWJ0/HAsrg203EmEJ3XOhOsOEwE8XLasnjUIwDIe4AtTWYpnKTj1IGy
4lelzjpoU3Hm6ameehT8lOrzb/ZOz+r12HiPAwHXw7/DIpGojhN6c2Dlg6m0T72GeIMAuRfq379B
fZi8mYQGdDulIuQ8+fLeEcr0gPpFV9iEQ9MhvkFAq+TsgOhoBb45ctK/x3QasOLlcRxRLjpNVidF
etswNMae/DngP4aRsZF4g6zw/xBFVWaaJtSZCUMdCBVT9xjowfXtKBbTz6eDwgdddPqbsVlAuxzt
6piJAN1MsXn4ZFcyRYCcWikuDXEt62/IzvDKQHHb95vu8HsK18FCiKgJPylAONGiVcGqa+mJMohp
oOFq2gA2Z5ur0sbZAk6+u8pbyLTHdIFzmT06zNnNfkLDzL6Bo64NG/qN9FeWMgE6Y7xZlEUJIRvT
W5EAUnxI8CI68/fghZ9rGo1i2w81jF906rTbfDD85eetfprZAJKMWWhNGlOjpv3Y7Gnr2yxo4BmC
6tvSDsNr/8fhA0nQ4RDbBAHP88VVpSVwMfrS116NbKDHAHybB6cpIXaixccKHIJH/TIa/btd7LeG
NuI9vF1XXZN2rXDsDgr6mU6X3Dxrr2Z9fwKn2wvDELkv67ET7GUpdXUHCAny5KakRKYWcpjsnTFf
DQI6W+UD4DLZTsIyMFIDK4mKNMizmFBO51J78IOECGKfuq9SSXEITAUHdH3JL0EvMgwHatK8f8Cj
dqIvNhsy/dsNINZon28CZoeABUs66OuvWicaYS2RORqUoHFTyEXxn7L9eqlIHWpK9Mm0bb52tqMY
+sg6v+B+ulLumIiXiDoAjEpxFQZG3y2IP5A/7pgqgTEJ3QpLlWBponGv6iHtobn90mRKSd5/CagO
nZa/PaO9jdZBPjfHLYf5gQtUWNyMaQFE2SGIYbDXDCGb4GutgJS/WErC3JQwWGyiaVUvg4isdPhX
5QBumEVZCyvyyA8UzsQeX3h0jeA7tqn2bcRLQKcX84CIaE6SvfHBKjlMegqfFI4x5W6HLVwZy33E
q4fc764GRGjuk6qgfU4oI2RBz+stNmubAKameJHovK9UQZrXxIxw49fsJZSLClQ4WCiW8KzgoEKl
nlJg3bi4eQg6V5IzNTysnWaBeboPQfOLp0XeRs7uVKOzVoNWeXwTPNIXyBIlZnf4EqlRAOZ2m7rS
MTYjwIrHAEZyRNdLU20ZuqxFd86Xd8gklauC35n86PyhfxDi7WBQ2E60dZ8d9vwwwp/CWuds479E
msVm58/buuT93OUyGY8d6KMoikwKP2HdNvk5o84eLYa5MNprm8po2+5ccq5WxzHpKIG6UILPBG8O
/HbOe0NJzJ6/62smUCfjQMA5IBB611azjhzXGo9rbdSyhH/U1lYTp/yb+aUDVYtatgdI2dfA29AZ
ajYGGVeH/cFfaOs7ln1ezZTdAfHqG59MVuZbt1T3l1sdgyZp2DeJHtRqaM09hEJ1s09Z8Z2N5NkU
38RvRUGb4Z+olwv43gPbiVHbgaj3BYA/SJK4B4blXlIuus3K+TA2AsS3IIifp88cd2wf+9/sQhCa
iqAC+MlYscBbErsQqoH/McHxSww4e5aqwX4T1iu0/v4kVhkd3b7IezOiJl282awU2EyUp+I2Ivw8
1zOa8YIWPZi2Z6zVawYKSOeRLEXHSJKJybTqBRmfWXEsZp13eh4gf2Rl9srQ6g3ckgmgC2gTPrim
5M5TKfytcLKwOMcQA4u7JxdIa4BNCTAV068AHpwNWmuw/A1D6SFcgYzvnQD9ExRuHs/OugwYkzfY
tPiecxFhIBpdtF4orhGH9OGzQkolSijm+xC1JEqbio6FA7y5v/Ds76kgKX4XP8irdMjr3eBDIeLg
oIkIprqlJ0jhw2FCQ7TnCk1bjZO2wXjr0DqgRJRL09FFn+82fk7+KNZxFZQgfmfT3GE2Y20m4AOA
UvRv7PahckixjYi32qSxh9Z73MzRl+F3KzTn9IbSAccX8qPx9WW6jWX7snsbwXgvjCFql0zzyW4B
k9TUDG4g/8CEFGRoI2SoD0M+LpefTgmtrNrjhR76w4Ier5tChc8Tv03DEDfVV82OYIVzl/3fL3I5
ZQh94wbVwFOEEv9cReQoMvPfevGdBfVCdBqAUDz75+EfLwZdUeFQRplaPbYA/HL+HNcbmVs8Tx9R
ERsCk28GPsHR8ZGRyPL6606k888IZVC2k5+j2bxKWK7GlwwtOvJfxfp/p0R/fz4XEtQBCuYlnaDb
gFRQuBo+fz3CNrgwOgwPqonsmYyk3MiY2KY9j5vSL0i8VFOuh6djfL2NW0fJz/7Je/xxrS77dma7
YyPoLSCZ8io1ItV6XREjoddDCzFU2sUGkcwtSTtbB2yOYk+BMxWCEJr3hPjxl8P8T7xJgKq1WtrT
akwaB37Nt2uk+rONVl+nKNBvdsqcFNfF97yvngR/aeYmiIIr0ZpsNMZwFv1ltY9F/5uUMPUDhmDR
OXlokakD4jcP6gZhjdCGHltKqrl0LE7CoKNxFM0TnlHiWxOh7nfdup8C/H1GWGbdoLaniCNFeDOd
NhxjhbB6xaWwqKO6lkzOwsiiogbwnrRo3horZkXpvpEAumfBm7cScF+iyppSwDI9h+W1bJDl8WM6
XwXhJ69BmDWly8t3z9bSkDnE/RgxFFL6t+heftxZr8seeCQqF3xfsJIiq6QwMPo4818Hrsb0wZLF
G3slOWnW629BiLAA+oq76ONfspKGc+zg6EM7aWmjmvjt9e4fuOyUAbIGZc2PnlrD0Qhu9D+81rB3
deqNKQMQNDBnEsRDweCuz0EDUrKAwpV9GEdQAZMweu6W+TxQZKHgAGRnhz51G5PqddGtXn6KjtGF
Wfauw3fZ47xNgSlvniw7DFLK1nqAljchvu5leIS9OQ12gi+VgLZLyYQumsxbj+LGSlf+xBkF8Ioi
NFa1YO4iZ7QqygkemFOWsWdl9hl0vTDf9uq3DDN56Wts3fw3Jk9FlhCccfuRdMc0LSGE25qoBesb
hOgNU3owWOBH6A+BjHJHTuudadea4YGBxPVQ9M+Ojfio3AjFVq0GSXouuDTL52h4KU9VdgoXOrbf
0BIoq5Y2w+ouiAtB7tg3I0/A0RV/fpIvtqppMONF0PJYdHHvmqq+XTPLQcVwDKneYjKoYqp5qvfq
+B2RqmFIeg3es0tt7HFHLNB53Lm6MZtamM2khdy/1qGioQ5DXWicLFOeqiDb16d4wZC4l7UbzeeJ
9g/t8UkgBwiFi8NcfFk8zqIvDnV+DIwRovEw+UBlYCZZscjL57w9gFjkvi2XUAOSV+r0OSMJeBpe
mINYqamkyCtTJJGzcBKZT1awgKaSqS4JzlbZaKWf8I9sxxzs+J4Q7zAQKlWCksg6yRn6XNmhVeE+
z+RjJI897lbXI0JwoCN+gtelcnEUENQIntfjy4c4SiIEPepb6AdD+/KmSaG/6w01xtQZtLKp1AOe
01I9GOhXPfQR24ozbsNPAo+4T5K/ZzPMxTroGBBb4XzfXsOn5xiLlL8XCZhMypLd2WVSupj/ZGir
akE46hYJiIWgkXFISoLywxx/awF7E2DqNwnks/GFetmae8b5ZaJm24mFCOEhpW0Q2PWRU3yTKiC1
2BuBqJEJKsRHkitGgq1w8kmGKBH4fcBrIg2X1GMzbaEMIRmlu7kplW3JVrOWDfol+zLLPrLvWxec
D5cLTPqdOsWAd5aF7X3j/8npI6UPwk2F/9Eu+LHJkz6aJ3C89D4Yci4woYgUO0DN6G0YINj1xFTN
bxsLT87rlk34SYWW8ERUArgd7eTLWURE3FK34gvroqjKAHz7ElciTzEHhPh3woHocRzjdrpsNBzD
PInUED2HBVZHpXE1G4AswZ44REelT5h1PxG9YApU4jen+dQeBHWpnydIVuV2Pr0zrWxZHJjh5Kxm
6w5ghZyGAnMsb9l2iAoACSxctUbbnEezqlCn+iflC7ac8GZ5rz68dHjYeidIkyO4PPOVa6AQI9Ng
yzTuuivj8T28YEdBfEkF+nh0X+5QqCTDMkevqs+8+dOxNCQbLregMg45vkyl6s/myNV+cqaCoxmb
qKF7X9eIIP5KLqN1ozoA2Bt6tXTcnN/c4G0Asm5CbKKpeZGSJQLvPFR5B3IOi02pU8oSHTAazPEc
jsO1kavL1GG2tUkVuhrlJJXNP2owYMpAU/Yd7vE0fI1p/pmoViBIXQwvirRpLC6UsKvYUy78bOn5
5UujAVRFVlRNErPuBwktS7YM6m6ufaoUfyT5Z4mM7JmgGUVhYgbknNBWcDw2m65lDnUXnPGYdOb3
rQhRn/2+0POofzz0XQLsw1V9+Jyi6qXERqdqQyuSqScN66av7nuV/siDSrQMSAQkCPsCJQIccHGJ
LEV/srZj1xOFavRQUYhFbWgF6Zs4q4CYVDpTXjhbzT7NG4hDJeLpP0/rx9PGNTFTGTMzTxdc1lT2
NmNv3Jotve16YQFvXENS9tBWrusDqVn8PQpybgY7owe9TgsYlz4Yay9DXsOT8X4p6ZmtiUJOgHa4
AkJ+ApHZfI3oAxmQRPDfoxa0j7EEalqqEt+h0aLJkJCeo2jA/zNlkj2HQqzXU9UkvxHlqPUzQAkp
vVS0IRw5TD4p3poFPfhTtWaIv5jgf8CqvOyrJiTl0RX/4/9ceQo/rf+A5KenU8VW4cRRe9g+JdkN
QlHMdV01na7LTLMfC+Bkvl+bi9mWeQZrk0uY4vLIJrSb+MD87mGhDLn/3mwxgyo9Xz4DBcl9Qe5/
EU+ev3/A/OUV2coNfzH5XMXLiWwr4uXB4pKSIXtIuexqOP4Gft2BWRvJBBo9IZDuNjr9AsYj7rPw
HV4AhmEUBEqVrJcI1NI8iyms/UR8oX/5FbiL95hZiawLvoPIGA3gtCLdc++vmXwTCIFYAWi4icXr
AFUbY1zCF9lMnuZVKRXmyjiQOks+bNjkfKi41WpXwKYZ0GC0bsGl6f1byLm1LmBdvSMkHaK9fHLt
8Ph52QR9ETzm5NdspqD5N6x/T/3XiQT7O7/FyoTIHZPcGkUiBIgtvL8yzAz78y6apSj53h4H0QAC
nS4hjH8uOedMfs4b1NF9wo81f99dfkd7HWZw//K5rc3b+GRJmDx6SRe9yMEsrtsTPXxgEKAQbNam
AKuHPqkVzulhF37bXAdPKhUrXr3HP24fjk9ZCeJPlMSImPaHhZlFBbm/bhmgR0T+WCDPOyHDLo2k
7gRFqK+5cg6mHuFbCGk1BEYIztnSm9RFShAaAl402IKu/bW8fzcqal/UTRXHFNFOpC3AjzRzRyVh
DuHh9EWegGFrEI9bIoTDQtgdmRGUVWvlXyyksCd6VAYkdusHlxKviQH2CUj/cvOQ8dmyaSSdLmWa
H0bPZPNJuQmuZz+WpuVngSI6+lom0UO/trIDMUztRF/jT4tyltze/EoscDU40tlO1uzkTfs5n773
CUDn1DtZn9IaiYHw75R1ISOmBVMPVzzRe4NG/7XTbiKfasfMWpUl5ze0K5T/D6zvbCCx4bdD5WEZ
N36HouqKd6M8rEMs/Q0Ejkc75xNNpStD6tY7gNNgEjoq3nkXx9eDs9zNtFAl8hKBtR4WMJZpTc2P
Y5th1h9vasc2bo54xeozU1txlB8e0cWc0Q+Us7dqKjRUqKKkSjBdNOdTtE4MaGEeauNz7x0DDKNv
tMiYjJKk3ckpoNQ44aGim4XkXCXVeDc9/LjDHlcXN+nfC1svG7ZWhNFqudVZh53ZsbDjh9evsi4J
C5S7Bqp+QjBi5AfVCuglGDLBfdOb6Lu7All1EfWuNqXRPjQ7eQFn6YKw5QneSiyf332t4BUrkzgk
IzxLK9YzxbOJXuCSBBXcIuK8D8Kp7zvVjv5ld2OBhfCZ1zBdJs0w7d0WKimHHRfO2cPYnL8v9Kb2
q00vFH5R5pcJOzloJ6mofNd6efIJrY/80zBlph6CJbgEm34gffOK2UvVYM1gfVBLktReLRullCJZ
Gp7HMSRKdEbxLLLvFA4KOh2F+YEX5SNIgfTyV2iuE4ufH51js9376Uh3TCChPB6UqsAoLdxJz81h
LtB7sJP2pFdpyFuav+N4ec8XiOaaBc5RChM/U2Oa+IEvCJcOnYfUQUgJyco7dOgjOa5LRguUtHZP
VDspGsgZKPWE5I5XghdY4KfmSZIG5Cr2ABGQecNll/dh8pX+IAfZgDkIJCbGR7RyAvhLuDE87KL+
fp/Du5pCsP1TN9ACReXkCQyx2WQ2veb8zEsOFV+O6sLqeG6dfKliLQBOg7I9FTRalaB2NPnHU08Y
Hxh5HSRdBUVo9Ywy6Z5U2pFLPBgri3/Hmliwdrp30VVVSKQLviyulqd1a4YBtBThE1RyEvDmD1CM
YYRkno4oSrOZPJgtVRG/dWZ9j3NIJU3oLag9xpobtWjTZeuMtH/SPx8sP8a4Vni/dxgtRv3vVlIs
SYssgn5qpCYAAm/cVXneUal+2jewgkxKep8F1VTeJMqzpniiu95UW1j+0QvW7ZsYZF19ESlx8bNm
yKQ8Cjf8+HOotgeYJ9miFHh3fS+U1JKyR0jf7wUbdsJoF7RtCNNGGdC5+Jvzsw8M8Sa+kLL9IvyG
TugAsP+B51WGrLXaXvbLPxmoeU8gw1m7zy5J26osjbJ4R6lzSXzDoUHZZX5BeIh5r7rkizJKhQeG
CPqSBQVgWhPqhtBZmCR5Zoa1Kp7ABS43jYBDTTESzPxRPlMNCKyXJaZr9OTFUIEB+Nvkz2QVxlcv
y1lxaCBfZ8lcUyhrW93o0HIgAjK4BaNUI8Y++c+LqZ37nBrjiF45iEJSwx2qe78x0YadeX/kqBRF
A582KZUezNKNguhuJnk5bsmZcN5bU8KIDOUUVrQwmhcC6+JGnht9bVX+yYIh5/8AalVzxeP1ZWRK
30Jx1uKv2b4II+HaAfC/YRiDfRXY+rEu9g/UbPxA4rIjKwUyuqHEdX7oRIXF+uFAuOpt28KaR6gA
1juIIof0nqYE9yDHHs+6adBuvC8cEyoETdP6QCApW1l12gMnjSy7YxUzAK6Z0xTVScnPNzwya3T4
aB78/Gc8Rm7TGzXze2i4Li2SRMoGz6O2yO6MnebPWHmSyJHbD3wNzXgj3HdZpfWYQYLqCxfN62Xn
XAkA+l3cZUMoQxjE/ebkcH9yvazNGFpN1z7QYhk7kqN2uaiAeQPndEX5dzgqofxGHajv12irFXp+
AqGoK+XJX0gw/Hv7xFtPFJRb1GffxISd9T2Mb4adiCkDMGTHaiIF8vmKjI1MHu8Ja2/wb4P5HdFv
R+2GdtMFVb5fWxmrH3X4VkFwIDF4eErlxujpva2jmlfg5QlQAwAyIMuz6OpreCtkwMbYkFXmvUck
CvI14aswr+2Ek30tkMe0EXkvahTiJph1POQ6PzMdnQAzfeig6YC6p84pJo5uI39DuxFOGI8Q9xDN
AQYY/BrCLJz5Z1tejWA7N3Xbaa+8I1fjIR7B9wrRGz+1slIh0LZbN6HxRNfCsyJZzvILQy3iAtlI
Ub5fqZ7aF00xQsesDyniUe3FK1zEAyju+qMdLYBfKxFS4ZPj7CJL1bJBm1MzYvBepZeXkK5ABo0N
Zo4lG6PnyTSpkhl+FKvfYOqdKUN90szq79WVBuIftExjsKOhit6FwxnLX5CchIEnzS2W+wfDV3GF
mjZdvsgeyM16o9Rky9LmaWkWiA1ODkkPz7Kr0MtpoxQI3jcMhf5EGuBvnZhvG4fULtISf2b7MIh4
FgwTY3OV+sd3GKQRc8glEiR25NHYTmaHv6Wah9yTUJ6WZIxKiQtdQrDhFMvavw9p2RUI8CaNES3p
67RAnaqtegAASRRem4AGnVoBkwWm9iAk+HytdPIfMV2wsQPXdx5wKFmoylHAF88VOIyvbwOfPfR8
qLIOj0hFZ8jHiaqvBJ8+yscnTgKrRxgogd77AFGeGsqRxzVDdXZZ01CWeJthVO7hiFHmK/edkvo0
N3wFCd1Wa7UMFXW0JYRx+JJ6vd+UBsu0KpfzwxtlQEy8u2gr1jYiYQa0GABtpEbQHYLc7/2IJrMf
G28MIlzOHJDbKDIxJtAgiSZTBF80Rno1774CaqrCsHDjZUlEKtEEhARS1Z5lxYLaIEOn6W+/BIJJ
YxJDcq54Cu2dejjJU4N1hgRBrGXe3IVhVtD3+A9LO4cq24OMZvgwDsMY3uuf7A5QoYTSaFay+Jw4
vLgQb0DlCMK2pZQvN+G3U/6lP92+JvnlDkFTakFfXW8cxqi0kybM700LzItEJwaGzq2WiggfDr3H
TDR7bjsmLtn9j/TNvwdLXn8AWtT1JKeUdOfUrWE3L/BbiTmXaY2uhDbIWGP2PDNkmnrJTxnbxti3
iIoqR2lMNwwASTo27Wxvb0IeAcXDVetssZufpwp0YFr0WRlxhH3bhA74jYOiXwoGg5HATn6ZsjfG
9TC8d0oFIfVD23BpFZkT7S/ORqgvTRiCAIzoSw2O9BtgYjWJu6kGg0grilfAZ+zCyYVevBx62lMi
MeHlAEMEfub5jQevcpHYvNTKNKwBFK0NtasoSAGfW4s3Zle3npBJVE5OxX9fnjj3uGmXiz+Tzw5+
cSnZycHcc9Umxi3VmWwSdDDzZJ5hYCXgQsr5mTLIJv1PAByOMpdYri86rueFsIGPMiE5hznSZml+
FI0LjyZbjORHuFkxD/7KkpwZfLPWi0+u/Udk7YM2pmUQjCvjWDDQXop5E0/AXb/zH6db6krWCtgD
4fxMTzopAufZbFUmvpcZcy8S665QJghdGCCaACZ9wqu63FIgnrU+sJe4w8sdXrxceabZrOV+mbKJ
RrCSnI5ujYaJpvFieBArDi0bs8jyk+OTKM1mjCPN3kRiwKY8sNb0SrlSI5pl16tLMv5eeTJ/lKr6
5Jb/XSn0u3VrVoiDSdjiSxSsu2bj5Set5qO/OVqcvb0tsMuL50k/pxGY61cMB8uv7pies2YYTnI8
4albTkLWeFkxRAWDqFBmKRb5ItKcgWhv8uJsuUATXTVrXcwNVYztAeZ20kMkREDyu3dkGpVdf4Xr
rcTXxAnngXYwY/60Px6ZGiSTwqzESFyAZ6u5qRtqkpZjLfPXGWJEgictWsxhcj65fEzuZIt+DiaB
t5Uh102xNGaeJSC2qIILYK9axv8vuqU/3ZxPXiGG7eSod9bXN6cOpFHTAY9JVYaE7/Pc/8JLqs8a
s+ZBeX4r7QtKepnalyeQnudPAJbCv/NbVns4TwIQcczU3t/IPyzzqBtfMHPGGbgl0X5pCE0U17O8
DWpo33ZVm9QazPiOsKl42t/f3xB2Sqy8vPSCxdTt+nMelw9ULVakZv1XS6x+xoy7YP10dUKeLUoS
s6favHDWB9h2MtyMptZij6EQwX3vzW8Qm3xCzJ7k3mvInfhOwmGHimeAibv0M7yVcXQr98mipufC
Wbc0aI/Fp8Lj/teWoFHXI5hL3qOopzcnX57ure40FUdmyX1KN7LdL5lc0wnhImoZlvGboqwrQJQU
pn5vYFX3oVhoocEfLGzOqH6dUziLj0YWp5hfFAd5SpyMWGCzAuiMmKITkIB9/frwoQJukdN2nLBM
dtp/P4oAvk8nrB9hpiBXcJU7IdOk5rjb+miLIwSHlI9P/PzXDMN2ASkX/3qWF2AlqiMBYx3QrPbT
MCYku8vYmzyGEcDTTtQ0LGq/a3ElfV1iDoA8B4S7zTaL5FqrO1yqBIf1r7EMEQrP5tkv8DKMMxyO
DwRVtX3li0UxgIe7DxjBXQPrpVqpq2fByEXddc1yo4sGOyOvZ7pKhJaIUz005mPDfdqwOA+QYdgf
9lzokRIXQvIDtC2iNJRCuYHwN2xUSJxi9x0UxwcMGr2EVfXB8dTHufIVbavIMBg8UJwKpHvWOGFJ
QEqq3cdwOfb51P5+CTMWTxXzX/2JiNzqIyCYYukFfKdvhikdHycDkZ2WSdDJg5noToucMTpQZ7Uq
Ox8+co2DYLfpTmRfGzNqruysbZxsx9mQdJJTWhu8KVtDr47HMFZhmwk92ce2vO8MSwOAncBk6ztc
2/+MxiyDOey3pWPId6Ul5kHydwf+yQfIY+C8l/Nx/ajOne0kwsyR/xf/LVQlP2at910/zd6eKlur
XgFV7K61uy8uocDt9JoDVSNUhinZ2mRrc6hFKLbotbDCNnCfVqZB4/Bf9AaJYhm/MkWIb2pjVtq8
sHYh2vMJVATSvAal00MqOZ2TWjp5HI6tn4p7dEoy9a35DKUVs+WK+Faxh8E9Mkw3luL080ffmsyw
CW4zasrJAAt4TBdOjUZJmVv8ZmVjWHrLr9sY/FOhnqgvD4ec4xwM0+LlrGN8EUgbc8Bb8+cciy//
Bucz7IS/dB9jVMTJ6rhkk16pnI6HgLP0kfHUJP3BVMxSco42VTNb80PyapBDrmWky24GaaXGSWYH
y9So+v1dqARrFB02zyPx2SwrDdaQyRnVfARid4PVaI/19SL9ZShJu1HqVI6bg2afNqOr+PJ9KzyT
4B0jHvv/2YbQvTjV+5FSNrX77MZ0v29FaEEHS5VjsV3R3QjccY2JSvxmF/omvy9zNzJVSCiR4bYO
AYVS6o9/DWRg9lawIsRDOhW6ZSLc1z8BRESi7VwSRmDB2HfF8vgKDzDXBUq8NpY18zLZo0nyS+E2
GZlewDnVkFjgaJvg5RerteZBMtz8KHcg9EP8aigr5og36NbQOWzu0y8UECUZ9y2Oc9KqhPyjz7iX
3ISPi43w+8f0zKvRvyGpRbeVIoXmZR0U2qwmjZELNFH0/vAUhBsE38oJ2b9I217XvuNUktdXCQhd
+/zak9pFJsnSE9zllpJM3L89ET3wROf61IOAE7uj2Vf+gZCxcgOyNSx7IE3TXwTSjDPSDANKN8e+
sjRPsEXBIBxi8gKV6Fyjc0ZtbTYTocFKYE8XqdNplimWVMwORoIMfdWlo/A9MOXCcAiw/C7b6sYf
F24NhNfgnOgR023Rye7UFeoYAXHdRV3QZiyTWkkdbcbavJ2imxijPOCtrX5lceaQfmafC66x8Ix2
HUzG3TST5qNk9mV9HkIbIeABoxZg85fud43qIkq76hIyWCHJpm6gq8mKQng7KEI7zsxBiZEeD/Xy
Yg8rOyy/eQymP7M86shv619QN+lEvUSySPBbEgx4xtThL0tebMl0BmlwVoTOH2oaUcno2hfLHA9s
LLv5LN9Ngf0xlBgtHbbSlEuH3lj2tf3+XaBwjNPJemwZM1r322MrNb3dYQ9gyN29UL7+6t1Y+sQ8
zoDx0FrCxxRZyK0dUSAb28WKgTIFUV2/sIwdk5PV2FPt4jB8WENpg2FEH+Eyf3Ug5aUcNFSJ49im
8yH8vx7NwWSy42or43Npl/ed7bNQhK3YcS4PpV9lzNGzhbZEpesifH8iLfccWryRhlTwwySNafXE
eMWId7JBmvAKKkLEsB9i5OXu4+oZjJkNuP3lySSGBabsd2KpanOHrzUc+9P3yVs9QYQZXuI29TjS
EKnjOodp8YST3OSzwvttANrMe/RwKK9lYXTYKVwBKqmiZWBN06AL+gwXd0dJK/a3z2zG9rMVk5/e
WXusAi2kSrkMZ3oHScP0BuisYzV5u6SE85Lb4u/k1x8u5InqZIkzricjKhOse9WkEvzyiL93YD08
L2LqKVjagYJFdkdWv/aTaQyLe33Of2h1NgMrM3hmK2eLh5Npnl07lwokxM5yLban6MpQ0BhP3q3J
LuNPFdfcLmSRddz/ck5S2ED58CzAvc28/Ztzutr4MfMxSZYoNqVyyAVFXOLfwMiD3vHiXn1dnc/y
uO3YZ9KeHaWsIpObSF7ckQfyp0eyUDBXDidez+6s3Ndx3rh1YewfgnkNj1aLtd0H2RAw0Ejm6pFs
ipqCMdsXWcTVnULkBP23qGWJMipyYN02oD58FowLUU6JcuCIc367cWBxLBsuHmmTzOKkh+2tRCdy
pcA+IgCqTewJQ1QkxISrQrBSXbeuSrgmtlnU0Pfk7q4m+Vwx8/zRIy0sp7Fq3xGKvyTypTV5M+p5
GRyF6kPXrAmuN7n6UaHYX8jmGyFl2qXJrxtRMJhsRvP7hYzgsMPG8slP42S+dUK8ihrcJl1MBcFk
stUUNYz8DfyN4X0F9VPkt34bqNRyDgP2/v2T+j183nWGL5NirmdqPVe10x55OrMDl9cyxRHq1dbo
doLk3fCjwb/BLVSqFw73Pz5579Tn45Dmw52043RhPfG8xWurHaEutB/Eqiu+9NyxxZh+rsyO4y7h
glfe9CTy8VKPhUfl2f/tLDGfPCfWTBfxzdOR9wXZ4FYprlhTL3grw0EqfTEg730985MS8oUBfz49
STB7dp+ZlHKRcoFMFxEyGtnNIf7VIDy/uCsMNgfZXTZzPEtnrj3Lyfgq1jKk7nRpDs/mV0XoLpDc
RiCoJs2o5BbNbkI7ryiXiM699vR5CNwaRUcAFOtKHpWUpaIcPM4kjecZXKzm33Qyc5dxXOXEc+aD
nm8V2OuESmc+WN6mXsf4obbJlfixRgffvS8xh4BRG3nOYUiOn016FLsB4r+qIyE9tcsHCNo8E06I
9W6tOfPW4+cXvCyzoc33v2Y0PkXiexBECu8onVCDvdgemeXt7dYa+cIEqFS6QGi8BFn0ocCGyLZB
ZRr90EMl2gySh4vNaivfETNGki8lnXyz7RMsuxSP08dLHoQaIXTpoUjwcZ1ZkXaLhbhBVag6crNK
ir5uwOo9lF2D4blagPh+VBB/PWRfnHDontjvjcMwzxF8DdlFXaJeMYVEOwlAxtenDuNEM+sQS2AV
VtT7oLpt22zLtg2dMBFlmL0G52aDWFP7lRQjX7AOIMYyodcuYa64OLbFNP7UdTIFmkAQnp2DSgiZ
pO+KZugKPkDA6++MD6hCOmk4uEiWw2WspgYgAsopoo/3+elc+h1amjBkxoYltOXq7xg4VRFGJFAk
pCBNYuLIdHQRe4sWulqhJD72Sf/hmdOH81PX+NIQpt0q4wrY5wvVRStY3ag+DiGQ8lsK4thpBNqX
j6wC/Kk3hbk1C3B8BDN7GHhdiNCQJoRr1dWunBs2z+AHZnflNbBtr7XwnRUDfTBUSj7FYn1TgkJd
rsXHzwpeF0iN0mzkQkyfzzJx1TIbaRl8mHr9bGkvD1yx8p4SPuf8SFTnER0hZTfOSs7TPBgVj1iH
fnuF6ewBgJHQbo8Do1L60gRvwCbmB9wlmAxUxwQJzyI37ut5bzb+Nfkl3qehTi4eyaJvMVbkw+3f
o5o/9SprzqqDLeZ/qnK3ud6ow/46IQZoiAhmyjJI1RMjpSoUGSdBKdwrJBfW/eT3X6J1P5AOF9CV
CjuMA+JAqFMEPFnwKjnbY6o6wJwn0z7ZZpqNSrEhPjtCx1Py1+tUsIcfvyf2/w5IBS6GisZ5m3+p
DneNtfhpLM0vPWx4/15jv8aCMJwpv6BjH6wHj0mme2tQQMekFC6dc2P6LiE6Ndvg/1HmpagMetQ/
J91/1bTbSnU8EYye+LYgpgW0StC32LNCw1+ValZf4bqn1QEG/M1ubRABdbXhbrhrfVCWoWIby0xL
TFnSn5wPJSK3xJ+iy9gxvWJLvMzJMX2e5l3/t7ic8a6/3Dlnlf2lhN5T6bOWABM8B1sp8cN1XPZU
S3RwAnWGopz3t8rQhNSlmk0/NsZAfyGuNw5p/iyYxdpac8Hf5TBlgGnEp8qEOIB+Nqb2ywA3DAf7
wsh7M/binO4n5PztBxyTAGqUebEeSvbIZBvONgSKsA8JqvfXlMSRoFau64lPaS/3Kj7iCXT5/1AA
+a/KzgMBYG+07O7dLhU7/OgHVL6eB+7CcmsazSirv8uUZuXOxEsomLuhygiQ251Ps2tYi4FS77Xm
+K8k+NF+BcfFt1Q8xRYtVpFp32s6KAkKKKUjIhSrnh8RpzsOrpQ+LfC1OryBfs1bFhrAkmbcd42G
jZW9e7R+p1myRrjOLp2mJgIcohvqroviOiZ6Puajo8cErIcrQ3YG5ECZA/YkfzbdN5AE1NlNi063
WMVxGHIwrd1llQaoXU67VXG0U9EJqPQHFBSS1DVFFT7iLK8RKn3UvWZ/FSRGFtNR2IbrtLRSd1JB
uOttuJ6MS8CZ/5LnW33RkK0vGVQXy9QeOwIiPdWUEPSz2mEvHYrkZYLjIixS/GZru/z9Heubr7lk
BQOkYiqhY4VoQ3tC0NkuR+jP9GsQdepG+azCfTQxWdfxBWiMrPyGwc7rLpA+T+nCWfpesIwxiZpm
WNVyIHU3leyvR7HYYw5elMePu/M4E3vvasRgoEWg8gKR6GKNWE6NCN/GcHp1s9V/6sQLelvxfbs0
+vxU4QfN7GFGIAN0z9B2SIYLqEACs5Y1oZdpS0wtDyBCfpQCSYlpKxanbb//XXyMJRWuHizeiqkF
5WtvvH1stsxDCGQj4oKEqqoJcTNk2jJ9uAwd4YX3AlubZX+PORqn/MDKyWYdLDotDpGazqW9Xy9h
GSXJvnFWBTphIXEsNnaIJ6KsxZyLWdvwD3JjqwDHXpAJIa8Gpnfg72oMiMIKvqeeurMnP1CybYDs
EUfZfEZVwR2jNfQBnrQxJ8xVX4EcHrEZZ8c8eMrk5H/HKcao6Fob1fxTYqawVwcMH5NGKroac3qC
C/8v5UwAX+UXKtcTnr5x76EbKPT3woX+kwrvJjr/yEbO9QxJO65Gp8qSRpTaEmHUZcjZk4cGpywB
QSiH10fd8YRmQa3uit9W731Zdz1WaX4Kz9utwiNjKPCwmX6plBQEewfKAKySFSQTyXAQOUV6lvDP
QtkbJKAjOyr66FOGKBlKhn8sO1AFWNJy3jHvbyBnKj3Kuc1PZmoUg3dtbq8R4024qWYhV7JJwfkL
lKPBLKHqFVtmYX7hNjPw1NbJg3L4XcWFmJr6EarDLKZUpVIVXUewgnkbP54o7AS7DJcf03mzNSXk
6uneRAB5zdaEfOvHg7prpAe1biH8pEjSGAQTAttIOp/KYf4dHdU577Vkv59ruD98WhgBgf/C1Gts
4fEkxgE4y7ooZcBiP7HwNsoLELQPz0S2iRb7oeF8ul6X8XBYd+T1c3BmiE3q4B/CtdgfW5FOOHCE
iFakY789Rqt6LrGCwL6Qjzhg0qnXkwMCTPmoGtJJgkS9rGSmF7rkQs8Q4PYgAnIDoF1Dzw926o1w
5DnkxyMCXs0AHnQM8GfR8J2tYUbyQKky6hM172nHj3KialRYaPWdkyNAmkjf0EvMrx1V/+ftpiXi
PpBS0cwkPYMKPj2IHXkw9LTLJDBzokz0u0wVEwhdZDRQu4G3UCWsZWDHlavMp0xqhlG4yLKsXEtr
kM0IdzbH62qCucM0yGHibWwVJYi1w0cG2YiQbFGuF2fRf8OUK/aFLOaASnH5H3sZaUjoM/hvdpYr
1qMjuAG7sDd1dTtGokxmrkeBGroYQEsrqnCDg8PGhKPqceKme4FidKI9mUl7jlz4JJitNZjOLvwl
thSSeN8j30Ew0P/u7Mymtvoa2mcqhY0u243g7Qp4Cp4ry6CjhvrW3lm4bsN5JtLBHWem0RJ7YiPz
dpidaDEH74n8972yLerogctKKg8ZInLityfxSsjQYCVOxOf3vyAQYmOhWXz9LYl8xVBkUi8Me3/K
y0T1oQw9mRdghpCtyboCoqGoIR1IaOjnYg2O2qiLysmB4hwAkMkGJWSJX8LOkEA15GGwRyS7Yw6Z
k7eYCJJuVuObDHrJdcFKEMlxl54mYMasTPW41+mtT1BjaI5fmRDZKxB3wmkbD2thnZDp6V5rNhe8
Uw/GPCMgW3r5Q+yuJqcQwZQHOo4LtUTmkQfHqpnUafEdyrgD9R/EkjyDBQHn/35ESt5T0Pob99/r
gXEf+QWECYzkMxLXqKMvdnFRb0bW335URuajxTN0dhKaN5CQ6ibhHJfAKrKYnDyb6ZF3FhA8SNzj
iXyZAwRM4qT52EazvI3QebODOYyIwn8qdreGefrXjBKOaU8H6QmsYMHGdGpT3Z2milmaTR8glc+z
IfYC12bURht54G75B/7ddcbt08A9r+jKHPU+AUj1BqVcM73+BxO8ISEQ0p6A1mNXSNEBT6d/IQrl
eCS85dmhXSh+CNsfkeQ75gBv2UYuDM1ZaUk7cdeZOjwzfE2Pi76IRu2ykLvBq86aI3SaObTAZ2Pn
Xst3Ab2eh33+75dYRXICyAK3rLHutZxGsWAeHF24fhjxAMmcwXsmTWjGDtMbDL1pC2YIIhCe0XFQ
k5vPucZMIUrd6mBlWLe9B1eaSGyBOtACx6at3XLsMsVaCZ2Dd+3sWIHeHhMeJ6m3/h0usHSN8X+F
zdNGFpWdNyNFAw9Uq7uAPIFPKPC1Zp2zyJWHXdRT4xuvw6kFGhbCdLjOr4EgqUd8odNHkZovaise
yaii6oc2plpPU6hnOoE8OMi6z+za2oGJ8JP46u8bAcNr/ONl+YYCgIHX++R3injyHrusbeeCjQQy
fKef6nM3z3G4U3/iTUOAaFSnrRwoQ4lAmbtjvlmiWvnjy4o25kIKw5XgJ1fXd25ISEoznIw5oRzc
/V7JKgWTdVShkxlUSy9nZSBvs3HvOUTl7WdyaoX90PdLOzfCaGWAr5x2GITtmiIUGoKmxG/TqHFu
/A0UudIsAVllckg+ohwP0L7DTRczzWvuoJQNlUuuRviqMVrqnD9ushEHCF2OueakxOY4V14zCIl2
iGbVBUqKVHtsLOzUHS45hmKF3qBLf4VARahQUFouBjJ+pbxC4jueiHkWIdkSE0ncfOEdF8j3NXpJ
EFMaq/OkvBcLIoxXpAmQEVZJbXVg0eE4ZoRQsmL9wvVbcL7NxSCfu/n4Ixv07sl8CGEXNypHhAxe
LCVykOxnp5vRaV7EPMymbQgDzIB8Rsy6HOyJnb/iAe2O1ozuqGrJ2kKqstLWE/m/VSiIgWceGeBU
RpSWIkJCKFn78Z72KiQYXjZEZtou30RYab38urqQDPRrNmeR9spaOqHuCSOG3Lcvu9aa9dEUu3kH
wHV09pEYOiEaY30wP9SPZGMPafxyGu+x0pMuohiIBG1u3cu8hPPlqtLfUS8HLew8wTBmMv6ZxzU3
AoRnUl2mT02zGitsIoDtemgVMiJcnPr9lxZBNWht7pZKIgdVLtlgOBLT/qZ/vtDSQv7nhDecq4pO
MGSTq5unLwH0gMrWzvDzZAApNXQn0sulVa5iD1dAdbNKrGsBp7Clfr85SmGmBP+Vreq8lFKTjkla
AaRzQEUoFKLNqEONga4ftTmQjcFlyTezg5TQ+vqSxtScisZWC3j5Sv2BTctn1F9w/LfHYubEY4Tu
pnfOTElighdA4n61oyga9GWYQfGqvtZ59a67Qs7i/8hSUyEJ1Y+eYroSg0ow7Nbe/W4FHJyuJDH2
gojlmqSz6wAKfsXBbwvBKie+Q46ppZL4y34aEeOMYJm0eO19QjRpZvpTde5OzEpf0meHdfLJnnVN
dZuSXxpnoD2T7lcKEwL1T/z0pM/QMaTftoEVLMIedPxmxW7JzbcfEnyrWhjAUVR3Li3Nkiyfb/8a
iZ2R9REnUOikGh+ucPssbq+azz5oJXrxi1piEBjtShKzYTY1rX8ayl/C9sapBqq6EZp86fSnTh7E
nafhgNQxMYTPT3vPvvt2x/CsLPw9y5RL9hGfIGlAoGAiBzT6w82qTqury84YxigiQvswoqrs9JpX
6k1vZySz5Z22ATNZ4TzhN5VfdRdoZlHJ2aggB9JvNsYwc7/dH2OpKKlV4MCda2Ryj8R9hHu27zml
ycRYcrxPpiiqnfdVSr+CG76pTSCMFOuh02ESscetO36taKSfRruao7PKzvpucVS+Bn8Y7VGmLOI7
LbbTXW5P+UBVBYp2mlI/9bgmCy+LLFt6A6ROsVZqqvaO2yllfC9yLgBFZ7jubgP+Xpc6ckCn8uY5
ICkA/bRI0f9+wugdUY7mf5eRQM+65RFCLD2nVGsSgZ/0abouq2fRpnzJustkeAyE9QPGQls2YFNU
JX2xgguEkGSagrtdfdXMoKjgshZIoSlT8COfpbFLeghzCPW9l6cb+BxNUgzXCKgBqqs0MpY9EB9x
IUskBYzfWkKeusq/BjNcdAbGQ3ZDP9Lylo1ra6s7w8zylzfbFe5C5kMzyzIfoKuQyam4zCTEkeJg
3jTaIIPcOB2NTYLA37Hti189tzFTb+I52nWHbPnMR3RLucQ36xA5vBZ1uLNOacdJg3xatcEcN5lT
fsy0ja7ZW9AFdhNQdxeVU38FfiWPH7XHJcf9mPQXLGo3Lzu9VtRKqhovGyQfj33vX6DotRLyTvA7
s3mlAKzTSAnx0OyODk4GQDg3S7xPuJwV2APTegXCm8nTpDJoahjt5/Xm5pl6hynGi+Q3mxG9ebEs
kCQvXKg+E4LMuwTX8xHMwLyGKTvG2f/38gcxxiQWYkLD4QmuG+spfeuHUkrOe3Y+dFmH1MhMs7vk
FuW/o765cK3EZCPS66gHFO+jXCOfeCT4dtpv5ve16XJT8I/xS6xsTJasvFooSodMMqv0mrJKvPvW
5/PGHMYocGUAqopx/m373U+yjkIXNYwzijXb+h5aUEwfv6KBLgHnoV9nwdcOvVRQdZ5RlY+KtNe0
nq7PDpBBKEvx6I1CgfLayi728odocLa4dkotq80seP9dr7NyRGBxqAYQuy1mdl93u9uDzglcPEVl
s6BN+AVgKYWo+qZsWdkZ55zvNb+cyvenk1UhzxtfpnPL0V5HmoOSHWRuhqK0ltVgZSlZ1BG8gcKQ
kTv0KrH4s1d6oRw4Z49TRCbaOmo6Pq9L2rN6+wt4/ZhS8bKcPxB2K+HCiWy1TU2jI6fH50fGzMBq
g16CZpv4X5CuBX9ieGVPPD6HpP6iXDFxI3g76NDyVh0/9mKfU6Pv5SPlgGAQ3IKHzddc04fBaOCw
/UnctXx25be2vg5g5gp0r6F2hG+ZwB+FiLyO7aBsQ1lZccaryuvBVFhEBjEuYQeCuYyFN8u8EbfY
wntzs1fU2IwNfaPAvwPow1SwJivacNvv/Ysx36f1CtkR/youajKgDxBCLZD3YK2KTSZj8eZ5Yt52
wIWpv7ESoKLibN8AnK9EyARji4VCO6lFDleIFKIeminFjqcDRT5oMusEI96facgerixn8R5q2gz5
6VOEhFpWJLp/HhvlU15u/xt6pPzxaHf4ty+pE/240x5qcydOP7u85JR8JiWGP1FvFzJEJG+ltqrE
phm3OnwKhyc82JBm+Ij6K7bX6w6oVIwM00LXvxEN8UOctmkrzFSq66jUJ+uiIG5qeV2AA5E/ORki
KpWXKuS/UXwIqu99tWbUk8XD80iwo4KC8bX4ccHtD4hqlxXmmM1Ygmx/SOuOZIU6x9lwKjUhcY4C
baRTDkrrUhomPWiy8s3Prfsu9evEQtQHOWkxhWMJXP9UH0w80g0JCyYHCH0tcWk3Ki4TwpO3NC/G
Z0IQHVRZuH67Cd01oBAMOwYSsifChdbjgppCVp8rlLaTEHMMkDGr9umAWr1h0bnDTh1wkxpoMhM3
ED14y5q2WjA3M0hUkHHcmUfU0+zjGMmoeLntT5lOGU655+mpm93p1derPr1BMuEdT2uRDaPfVivv
m0KWF0cboiukHUoKZ3EXIDZf5psGXmzGYFgWjgQek+GKcKccSlz2sk70pg7yF+raL36xRWAirrVK
aRV+Vx3jycYAXPDwsF2S1Jn/bhhUA51eEydIlpt7uT7oi/gF49BrDjtHmsk9q1l7Xh2VFzk5DVB/
4CwDuBc3AbfHuTTlyHkx23UBVypejASeduLuIFDoRh+UrRUUkUpclxG/lNeSVwTCbJMqVhpB8Xjy
k4gLYX0G4QGgZWoI7vAlDyqsYAPtu9wt7HorfJ2iKr4zS92VRO5+SiMO/p5xqbvVUD9tcwlPv2WM
DFErTM1iDY8teadXF286BUijco3vrqmSiyxaKZu2Sh8E7tHzqUGbIGzEF7/Ps1WbDKzNBxl0izjs
ZU279XoT2n2IHvuF6tWXlYt+4mSf7ULRP6GLqKLrZaba28aA4H+ZUvQaxUUUXPsf2/AhNXeDytTa
H8Tx67XZinCR9Lwlsjp5zbHLb57gFM1+php3lwpIAM6VTIh3sZ3DCdbcXwfvB9Vw2/B9kyta+nwj
FvVRijZd9bZONImUsL0xVM9ns6XflEwLQFAeCP2fq+//WBCv5iLDsC7gXV4AAs0cPFdRFp66iENh
6JqO2JGYX1wk90HK3U0BkliddZIqXvDM+94oMYvEDIGvqUSq2aIrrjDbbTEaksLaDoAal1PKZXPT
KgFY4cUN9pVLuYr6qUFMb4oD7ech9BDQIsz1Fj3JyEM6triTxguYxBpJhMyssKiwNV4Vu+cRO1RW
NlfbQkJMJtVk0a9X5AucBKldjUB4UO3qq1QJU1HG5BI+V7UCHz4WI2B7dCYNRxhW6VEzKvMlaNNA
mNjiT/v9smh8LjYg7C3HrYh2oLeRFR27Lw7L6avKnrJrFLF6kxsvOulESjcZJhu31dd9IW0Z8DoJ
0iVDEYwIF/vJ75MhJBy7280lOG2y1WHnwZ6TOu/aIT4P/HCh6DCvhJPC3fYFzfIahn7SkYTRZirj
lQdOVemESkTt+wQ1Mdk4DePJi1GQo1BlBYnKm0Y+L7wyAiVmahcXXjdfv1V1WjZIf/TW3QuJEgQO
u7tBQ5YU5O8m/xRRkUdfAClmRqykQFcnCHSZIiaDGcn/XHUInVjccRvcqRFRub+Rab80d0sQ/vuQ
mQWzjyU0ek3GVHZOlmQL+slaUAurUTFluzR66Bv+aJenW2wESICfsSzutvLISOeXdIAfYYPpufd6
tBNNuCfR0sYWiKSEzG0dV3X4MSlZYpSdfXuWs8fZ6xy4HOpCul0ZfskyYAHDd2LaKG7NvTErn71l
m4N7Az5BbWjtDkYky5+ut/6iJ2QgYkpoGu1i3TohkSl0saotf5Ei0AULZ+gPM9yfnLG4gPbNRT0/
ODkPy3sWEJgb3Nci6OwjydAsStfw/Wx00V0D7MOjh1Ora1X9VLnxyule6FLWBDPt5H++p8N5nMoz
DuS74zL9GrhhidS6Eq7PnzFYC9jg77OSz98tJumE4YJ5FMYyzOVd9WPvfli8buF6Bch4EN8pP97t
//mzEGvBYe8PZLJ1v+z+tQYqdZ87TLOYYOBys1/UXPj+GFlnRlt1AXGv/Avz98yWVtK5WhP4d4Mw
psw/fBCUqLo9qSYzkTOY0wSaSEdE6KUXV7zymF65qX9npa9GutCauScJ4acWjVgY/JBWASbiXDiJ
VDc7pX+4bKYkRIm0uBnw8N01EbItW0Udy1Zpp4rp4l4ErVqeV6qZQOcTydxmo+/hTu9zMNg4UVdp
a9d7+68zA8ZZBFjSptg2yGyf/GLgqWJWX6uscamwWcoCgpzJOwIVTZOr3sjtFCKTy1nLxUuZgezM
qW5ilJ0APc0piLOQeDv20lqrBkypxvXtWhyKLDLrVokAS5w5jdBCFaCJr3Ct0thfiQbzjkjkkzX5
MNiOHcbZMgc4ldaZbibgCST4hLcoic52+0Ecj14Uz2Z5DSqJcxtHh0Q2d5CfdfmFiRF88wZlKWz4
HfAXiB2oYadS+cfEP5qv0FL6pamL6kcWQLFgj2h2//u3Wq7AzLPdVQo8i213HiR4dSlmVUyEJXrQ
mUajeTMi9U5SiIsjDkTRrSuhU5HCSE1iCJ+XCQXyUHQSA2sj9/bez2PBU64GTKIZm8xbb74PrBg4
1G0dAQCC+DqHQ0SWL8lcZoEEw7BJOYtW0npBUvYIm9RgphZGHCF8Mtumsdgrb3DOw0Xi2+kAazq8
rKwXJcqbQOSPEL+ReOrhrQVj41vOkYng5Nh+g9Pn5o7hOQB1E0bgx67zo5v5JmhipZDFIWNh19bd
hTmqW5eWfs3oZYM8z0CNgNFm/rAXMhFjLL9kXkgaocAQ6srfrYZCv0lr2o+38XaGZkGMzTDqcvh7
A2YDvXdUksUpuJKkHFLpjAMj2cOKZP5rTJxRHxjl5BMXn1aJLjNQS3sb5S4v+gSaboH+vM4koEhR
6G1w4l8RLOz7Rf6cA4BxNoNTTbi5a+QpF+jeU+XAV5y4KyPBRF9BOlTdXoJm/0W5FRGwDwO5PImR
39/uBqezirtASERn/SWxviy9FdoEQbMWY2q//uJR0ubAh8LAUKJtnK/X5btOqytxVloMuv6Z2pwt
DZx+KsC9eXOhF18cGAx68ZtFOmBvFjtbmrqC5FZcLNQfeJLO5+yJvyDEGzjSA1vY74nf1Ujy0y3e
HVMbEaGgWraXp/vgOf64bnkEq+kUy0cQi1nTJYwIwzArlbdt8lOHQAVZIKkrweLoAzWsPUOxWvk6
qMbMqpxmPHS1yJ88MKUT3R0gbw395ZhSXC/f4i/ABDzR6CeRGFFu7c0Yp78Pwrh3NVu0evudr22N
8dfMId6i7yAHejVR2+k1DLUcx2o8n4wGYTks6WyPYgjNzH8gvrnmBcxXnXGQaHHMV77zg4zg1AmG
7RTg9JkhZ/iXnzbgr9lXySA6mSi6F1r8S9CaTBq0arZDQWLMYikZzLwQ98PUq6w91i/wdC4UEJ8e
99QHI7sKl2pzrdzp7RXVqD3BL6Eb9Lid31p/8KHCESg2ew6588Z7WouoIXz04AIWsTfdHGugbyhu
kR2HroSLOtVRrHzTdmlEsBteN47IChZQcVSo4YVhdzag2p1I5gSI+LqJ3hlGoDkpg8mGkBOXKnyC
00XqvHiiogG+NbOwWAGb7agZr/jK434Vn8EaG7zjfqzxY0aSPYb/KhSfR2NPeNjl9jZEAksP5E6Y
76e31gf8QRHSALOK+Wczcfr2mnw2GX0ZwvcSlcvD88IM4PFSAgIauaTphPZ8gfhZGVyMWJz0gGdm
yiD2CI9opYPZZqNEN9VCLC5dWfZdk8VDAdR6Ak3EiLWVqxwHlqR2UL6yPQLA12hWyYKASaJoi+BI
GRr3Eta5dLf0jSpqQOtZhaoLopBGBkPilwJkP5iyEtl7gFiq5KtFu1c2Ke74TBAr9nq5QgM5Ho5a
6PqOm/0ngVBIm+aH66499L+GPT4cxCOb2ITRQ44T+MIAD2V3jKYvMKzbsxWap+gEXITL5wEYlx3i
gVelKDdLv/yOC9oMZnpK1AwxIb08aP3DvUOwg6XNdI6N7HSolwbVIbcbcKy0Ykan+kQ8DcdPDwxv
dOOU2dGhWeYaDl23T8gS92H+zmzKokBQuJv+e0KH7vmzDIJ3pBS5F5OsZj3LVIwjhieObDEhFWCI
sz+lqnv0Q7CKh938x5HIWQiKv02CKqSN/T1HQHVASrExAZmBG13tF0dm165ngTftz19uaj0BBRQd
LAkwxTxNeiPgvrClKsi/8TUW4Alp7TvzEMbd4AQmS74i/9BQgdo0nFcEe+znMVKy3ShsYZpoqtL8
tccqHgkxAxg3OzQ54nKsGNttRIrwa+DXwZpdNatN+H+Rc96V9d1kOuvvKK7j+I1U43EF2aeBx9py
dSXavoY5g4np0tbdEqDV5PoLZcR35Xa8wupJudeLk/VFm9RhRxuFPHJ2RoqbQDF37i0llXhl6riP
g59RrSa/SVnN+QhCbXxqmrsP91wmgAVpG5AB6Xy69efX8TbMlLXNC2K4qLg92SxBvzaJWqauqJcN
eeQ0zgV82fI1CQg49Wsgv4kiEJ+EEsg6gGbTLqQYeY/GIkw+NPSGzyxP4Vjuhtdu/3NMXQiSZowr
q+2oIEe0O8f1qjW+2PBiufHIUvMgCZPCUdmDpmmjEfbB6FZVE39E3nybHTGvVLcwfjUVMgMixwma
BIi2cimiqc3+wSnx6w2MzlkoL8v/SkQBRdemEr+6O2ywRVrJEnydlsvlsafqOiMjNoQATTgVe575
FnFFYGUCwRUSSoKOoD8zqDftXpf2Zxc7/oWVM/NfAGdKnEgzpp3fKCIL2DXqF+CwgNewvlBvzDZA
PYf00nvv8bd+6/9QOJJoQbqjb609L+wavqT1AZLgbvR3vFMrGuLurCGCr3Cep3Z3NakkkvgP0Hej
bRfy7/73gI8u12gx/3aeOap2F1ERqoqNOEEEx5/0VkGNFf2Mku8utHE/6FfpikOCF1S7Y0M2svNr
smDLGka/X84lhJXQqLYlacqwQX5MqfhttAkPhtgStbwpdq52Hxih4nqlczPsTFUx/juhXM09PseC
FfPg8hvYGWGPKyl2ogu2AuF/W47KBt1l4N0eSHctaiOQj6o1NNuMTZZFnHI5NJDKBuWtg++hHDRv
LZei2o14VNpIN4NTaS/BLKRxxg7rJ0P/dsm9G2JrMJieZT7XdWcNh4PK6wPy7URdb8QJpwbDNYx5
c4pLFOgfA7vfFm8hS+UMXpmhwwpFI+1sHQ3Pj6wTGq7o88s+4ip9eWGKdgb6Syvpk1hFXyezkA5V
mYK6KMJq1bt0NiV/84kt47DrekzjGBNbM4wxcWitnanUB+v/K8tli2iBiOU8B/ATZ4qNt7J/FBjV
2lnyWF9uUwqmdYZqotpwkwuvs+UdRdfun3oAqpiI5J4xVFjO/HOyanzgcOZCmf30bGXORla0SI8N
mfTfEGhSdK8Vu2zLru/9rYYs+udTDzvqNcIVm6BAGk0RlRGHLC9wPdQt//UgDrQ+OoY/t2sfOzjV
yzfDGsH7mFroKI8UNFGFYkL5LjSfV4jw/XrFMQ0I4ywjRjllVCjc8uCnVTyxLDNVvkuFqePT2cik
f9pw29M/7AlemKRuxsQSUY3Ivje7ClH+PwPDgDR6/KTzA3UlRzsF7UzY3EDwwZBput21n6QM3YFz
pp4mScfZVyJ1HxQODFr88QN1zm0a83VfmrulCn+jOY47h9LUiUb6aNEnZHgYVOnOa/whLgBxOstg
yLvmpOiyzhXZRPcUmUtnB7kbEXbUhzITbXutn1WDROXUMJVuc9HTnzyCllcPW2+i8juTNeF/AV9Y
6qGmAIObHO6G4vW96pcd/M4+Ijt+cgkach36UUmCmFYHUprcHf72KORbOooGFy4YrVDVDGxhhOrY
Yj+hUrodyY2zNtsULqKTNhUMBF6ZQQjs0rWRj233I0a8MTkA+PfA+DcpqENs5iK1KAz8AQkLeIV6
ez6oIcM028SqOUx4N52kHNdfwN1Ws6Rt8yEjumjZUw3z1myJiv6TsD0JrG7FVfXk+G8zsjmtZJKj
rW4v2sf/d40ZVBe2U2gOd1Bg/RQCvEiTl964f5FwwmaAOEZZRk2HIo+0DoaeJCX5FC79GeUA5fe+
m/yMDbJE865xwG5oWkuJXQIt+1VkmjytNOYxqid5VFgXEzqQPnN83F+KtDIrY0wDa0Kf0WGQ9SjM
xm+fra9jA6y5B6pJ6iLqJXqEdkiPVJF/ycvGXOqyTFcU6jEbuwD0hitCW8qXinX5UFWU1SDyuvaQ
3OR2G+mzWnDX2X412coZyQ5k1p9aBjBsX7QvWzKfBIL4fRu1ua+KOmyFG3/Rmgp/m2ZI6ALDl+Xq
ldRRJEp97GoBLrmW0GjJLzqDYJUe/EIT1VIZIuYdojrv33WHYJwoYPgeiLK0MLniLtKZx5njLSxO
Gk+kwJDEgMpABj4imXlBHy0DTziJzqB7snqyheLYGf6bspbZ2tP68g/1whac9HpiPDPGGMYHXnnZ
GxSUFDWJqS4nYX9XvjWpwRBKctNUI8PlZl9bkNpD9MpfQ1QlvIT1tzLXIURcL5mV9995rEGjmEJJ
2DyXQXxR3S0kmwVh0A8NHST7dbex93lFFJ28cydZIs3rARaNgJIQnPPSaEeT3g53UEQ/MC3dVNz0
KsrQvxD7s5I24RqBnuq6PnbY7B00dNcDothz0SsNS64M3kKKZ5RJiu2CasTaw16aIdoCrIiJ6qkv
3MeLL8tvuLsasxx/KHG6hlsf47r04S3pLB5keBz5FqZZWwBvePzXu7wVzfIbN8xUx5IwLHLp4buP
Jr0pcF556s9qcwM4yzur6oLyDlA4HepRBXIqgr1tSIV7XUnOBUu6BSzthvJbClyZEhVYcHNFsJXn
RChxVsZKnEV2SMrGk0cIPw3IEMrL/YMCdsQI8PwUGOimJf1X5KyWIBSuaRKhIT8jG+h8Of2T7aK/
p1HE2LXvUv+pRK1tFRmb7VjwRQfTkPmX4PAxfq/DtAjnD0jnfQm2uR8FsSFQABIS72hKcEcOqP2i
cJWkddcRblNoR/+jHLdj85VOZvqN6PVRrBbG84CbQkMvbmdehnrYch31yDF1Uu4w5O8QlJINSxWM
uUs0VhlDRPVdHM+ns4ANhKlFjtxxoRGHKS96dz5GdO5bxhnRVixZ1y7E4rf2WItF8NoEy/5AmDzm
C0QLASPDD3ErYlPAABsiegPuQYyysyt0awwwIBb3iH4uzWBNteK8p2JAacXJ31bHsknKEqcFs5w+
usgRrOKOlLFpHC5gdua2A5kW7cwB9DFfo9mzR2lhBazu/Xtu3Zww+z3DZBnQcxGKYTKybmVMY4jh
7XXOnZd1K091vznn4uLJPs2f/Ux0mfyN+eg+iShIoLu8lGwU6jWS7OrhT+SrNBSzGqOio3dvMq1c
iIGbMRATB0jovi3lOLFWuf7H5iI3ZsVyDK8iCLyOLa+YnLEBz9oGccQuLyAG+Wtwh0RfToUOF4eh
SToy1f8C+yQAWFzmusLXoshSuMLZWMYXTvbo7EM3d9SEUeYGEwJopmnw2W3ulMpmoudDhIYJkBq7
Jb3SFhtp6/JWwRChXz3CEckOqf2B3AkFHRGqiCY/X9Uulwyt0eIxdd7PqOD39A7DpqlXQ6iwc/IV
lMOgGnEdm8LoC7eWSfO2zCmPFdudYS1X0FJyEyM2mEBCS35BkQWWMeOgTr349LgKVM2GuKp692Og
6KU9LkcPL78GJBcjADzyKKYtPhf1t23i2FyCCxvM2wjFPOjhXMtW409+9NxWCBDp2ZJX54UihW2P
7d7YUM7vo+Nxy9xfGRztkrsrpMIyFPtbk+jwJpIr1e3oF69mhFkH/MVz0pybR7vM2t7/LxrSAJyD
NZbPnnN0c6iWjk1h5iNV6povrf/G0CHsxhyt5fAJy+j1HBXka/ey0Nuk0KHDIqRzFoR328P9nSQj
R0wAQvF5lVYbmixeunau8+z35r+cGSTpYaerCJaJdDH4mEjPO1y8ayfBQ9JZT/kzF+t9WPKKWb6Q
YErzbDATJNru44+8Su15JifszG0OAJhHaEpGDI33WZ3k92UVebBbBWd4s38Z5Pf1w2o0vQIAHWiO
U25UpRAzkkY9yV5gu3gv/e8lzbs03vKeITY6rK+wF+Neia3O5yjrF+iS7vRZ3a1VIq1URSRwpHL3
OHT6025Unflk99vTd9m4lbszxjsPvtf6Azp+TbdShmkV6HVCKgrC4tZTDT0mXaC8/PP3orFVcdx2
9l6kf6iCpUiDnvlrtci/89wDsyPgPUIlivNLIPUKPfd/f6HwaH2nHQ2wTWcQyLaMrqjoNfp6kWcN
vczP3sKSuzjAx0pDIk8x94i+h8dNH6OAl36KS6ZL3lLWxrTU6chr425B+y4OBX1h2Ztd/KYuJqxe
rRY0Pt70ZnSGZ3ldfKiUyRmbQcUIP1p3AS3HMpV0fjIwi3DiW5aYjm8MROsGd25JyLRf7kZW+TbC
U3vVfz8EH6sLtBSbSJVtaRQFV/xMDDKCIOh/7eQBJ3RkwgeLYHQ3QJ9mzqFOM/rGmn8oQXOhxL8H
k26YTZ8DKL3wENm0Gp2AohcWXMoGv/AEFRJv6/o+sZp6sN4ODWVgBGnM01XsGKlmZIWU0TlPmaA1
4vrNq8yljEGmnWk11ovOpGaHhbAGFwwVfAHtGVnwGxE6SlUxQ1P4aZD9BwIJME7Zwrf1K2alYGex
MdQTfmASZE8ZSdOF9VU7dbHG0b75jrBlQzyLQJX7K6wk4FfBeJZLWeh6i7uRNj67GNmXTKGUdgul
t8u5M1xNK/voVq1zn3NuiD5II7oaz4XzdydQDMWfmJ2BnTZ26wdks2j7DFAneSwurzt2FMpLmF4g
ctdmHzZ90qrShN5lylWSR2hX1NrH2zREXj0MBExZE8t5NRBlLqIZlfY5Sal7UW83dIp2q6opuXzk
wDXFhXdAZbFZXboS1bqAxeUeEQ9qgfNdEZPL0BaXWxm1cN/86M02Ken7R4kzk4BHgWL4CJ0eIIqm
xkBp6Tl75QhAtgbEtCrnwP8OF0WO62EcirFbYhUOE/8oHRbR0874c4SCz4biQZNtCIunjpvl4sJG
zhptBLK2BDf9OlD/DGcNfYSicow5eF91ehjKiIQZHAncmK1uw3ek0fI+ffDjap4xXLA/eNLuWuzC
W7WOli8HHnLojIeu6XxMRpMnpySVwOEGkz4Rla3xxNNu7RvBnY46QFquJYDEQpg2cldW6Izuabz6
p7b/8ym9COj8pf0vmXVZ93Jt3Y10CDv42qg0ECpYjHUcmKLH7FvuoAhad1zxNyai3Rek4+1xDLyo
k7bUMgHYmvtlfEURGq+z1eD40bqJSJuNrhN3hHCIpTa9uC/o27HLgB8fBWluws8Vdy/fb5BLMLrx
nJIwDo/5T+MsLv/1cNrGAa2l+spQH2iShwECX6ZG7REazQrzY7RV+kZ0mP3FgGfer4G2LGSGAvYb
a5ZmSA2SrFHh2nngUXlX7N2yVqKo7CDZ7TnYzLO8hRMLs8IZXkZp2Wcf8T4XVsngtcEFo35EQWUn
lH4NoE4UBEXx6B5/xhyZk+jETNm2bWltUYHoAejFKgY+5aJVBAnTF88lLcyeo0vNj6jJh+o6RNL8
j53gF3PLwsPmDnfq9fDOhpXXFcVUgUYIcmnfA1n4uNTmQx/rhbKN1tX0wlI6PjXQo8SFVLTRlOtB
U72XeEoFQsvpVGyqtfIIeoGE3Ily77d326ubnb1aAcnqAJKuZeLf1TDzLvr+KhA+ScDdIqz2LjJC
Of52bXx8Uu/mf0/sf+eCfF29Nwz3ktHQNJmLN8LNMTTxxgN+WsvdaRa5r1QRM8GMzLZHJFc28NNi
8CixP6lQdCG3AR4O4AYdmrHCa+uyDBjG/npXDlaAJLhnSdA7rcic7Me0nDCzYOoSl9m0i1GZWVfQ
YhUwTwwngWLnssIQDoK2O0hkWM5vyStT+Mc/FVMsOGFx3vwrepnBYd+yBKQ3HYKySusuSiEsdo8K
cBTadva5AOP1QwBW1dXc7inLA9DbIkH1Ypa3BBRkbjnfLc8WQ92VOhdxUjjlFTA8D1T/W0ZNBatO
0bEoy2lwS6k63UuzPcgV4aILhj830aTW1kDdqqTKWYIKAtdK+gApoKcE7l7J9pOapLmmnjZmEgoQ
gs0hGGyI73j2a8X3lg8VvpGzbXttsrPAxy0AQnV2p3qt3TIc+zvby1OWy6a0GE83DGzefG9gzgNW
1P9hRFzEgKUQ8NQPmG4YBBqlG3pALceWxJVHUV04rMtICiM/bw49AhXwrAWQ01AXFonXXTwIHfyi
oa3kDcP/ylP0fyFrAK68XCG9KkVE/K37qTIPboQBsMCKiqFRKofaPXE+VvZtxqnUU0kFt7KTrCRF
hQniJzeDsfIjeYM1JNpCRK+Nxut5RAc2PgxlVuMb8QcfZdr4vjNfVOHX24R0DGt+4Zbx9cO1H+vs
VgOtWZ8cm7VGpsnS5N1BBE1K68NsQaK1Mxt4YdvPHJpp9k0nFW4HDjkT+i4PcdwDYlUZV2gCDED4
X5o1gLpnYHaOCcaJRHbS8hvooc5pQAYiv/9dTIrFSnSiXgYqR/utjhxVfStjZlYcW2dH0PbXa+OM
ba3HAJJPiQ8OG9XMwUOONm47u+h3vs8rgkatCa4Fa3yWn+cmhLpC5p4dmuLKshfkkalpYHNJIr/b
CjqbUpDDmxpO04xYljEqjFdKj6QzrkJsUcR9sVKGIcymCx6N3vxTkuLha/ZzESWNpB6MHJAk7Ixb
gQWALTOPUGQ8OAgE3XpMefquJg/zFFPitT8XjAStegE2mmzrGdnK2OLiiP8mgnu9prsARrfZqGnR
9vLhUU9TXcs1tFvvYW2zH93E9SO0TVLnOKUFsS9DM4zeYoqVUzcQMAcvYWMH9G3ZuUAdiVaGyCgv
G7poQl/NYlZV7nyJ1ByS7bycUSqcuu8sf4hcKbjDPg2x1btkr+DQ37WcVNDEeAhVGyVw5z5HB3d/
byD2hWJGoNlcm+CPrxIhKiH7v8wM/t2ev8LU0SwXC2pSyBgP82pb+nW96+0vUbK5BB2NqSQWyyu+
3H7LuV5YN0D80A9JG/bPpyQlHxcq8UKKROyvqtMf1j36UqKhxvRpOy+RbFNzlCwiJ052JPVUMC7W
emxPBENe+TkvSCL/ntx2pfirjo3LCYPPYjVe0X0jVRcV5ldvtfvjy0iaOyzsM8sXUr9c5PIxOEBq
Ftff72mWA2jcmtYXvHidUy0OHopOMVsMF4jVW0L9xsFcLTltCN3ict8a7MkUMPD7BSYe2RKEc2D7
2RQpJgaR5vf3qWb6eRMSs8F5DSreBxNl5j5NqNvX+GdxF1o9r735GYDbNDJPv/HSIhJ0XJowfui9
Xi7/v6XKD9vWDrNmLEURIzzCil01y6ljYUs8cv2mw2F2nD3jbdkumr4M2XkYcK7RQpXyp0G3cdnB
3ijWsv0qx3/xvKZ2oVIzjn9tLoVEnVHZwIJnTmduRfAfkXfkrk9aBP0Wrgml5xjEruOVbqE+ms/Q
ExXwzhiM4gb5IZF+mTrMadTARSk84d+WCBSKf6rpqUt4SmmjMgOYvvqJVKO7NU08ZJJK5jxzDy+Y
vD6JisfZgus6M052Exn3Yp9Mnix/+q+XQGDpZNBBYet73LwETcy+r8s+JhTVl400d9de6NVJkrrj
HYE1m69hgw+rj8VPKtcbotPc2RwUluC3oPyAKByLOHRQ1dzmz3jlGbtbc0lx9wqTT4x2rSoe6ZXY
YBNqlDU8/M7m4/bXWnjmiCoQsdoVakzMZjnjBhGtCXmTaH01Fx+RuOI/VfLIvOqVfYXo19YDn08j
7rVat4VsiB66KuF171uSkdr6Yn8yOtzb21RE87fHxDVwRAKPbJcVuv0KJ27BPL0v1i396RURVFh7
AvI5llGFJFcsfP68w2liLp9TgaoWhA8PP5tZvYTDwXd6TJQudrVzmG9Aq7Q44MnMTNLPxnSV6Z4T
SPqZxO2CvoXqibrhobNVjTu506vfYqg3jJ7OXAAngblkzusM6GmW7qcss/mdwI7Av8n/smTHeLSI
uMlhhynLaPZkJWxyDBsBUKDLUZviXX5J1gOie8J2xJjFR9sisYXXeurtp7JBQqsIOIabAyvAiWQV
wpumTW1pf0cb1eWMbfTA/m347yoHDe2VRpr4rpnkUeS/UfETUk3CW0cdpUhnz8/8/2fi5hY5rVLC
hXQZKX0KlFLa5ayt/QszkuMLr3fdGG3Clb/WLCGDVIMD9uGuEoz37CCZwZcmT7LPdltSKO74Gd2S
emSCvQjbXRTujokNsOC+cPJf/fERVbQ8LkrCFnJIX8IdsyaZLwgvn7yRO9N2SjqKR1TPJ+ydKTr1
/1fwkZHWyKix3lqQrO4B+r2eBS27WL3dqTuuOR5Ss7Pa2Q2jDQAj7V4yfvlDy8OgIW4eJ5OqMz3k
CVhvCA0FxsA4i41pYlHYvc5tboVJslaeTFAxDj1aryR+0FmGGy4t0cvZKiWMO+7vyFlfopwSywkp
bDWfm7CRgFgy+GBGbyr+cOWtHRs9xF74eGkTU9e+K8T8EGlSup350+B9VR+Sk1AQjXZuo/9lBEHG
qfJuXJMlCQMpt+hDyNXoOWqDFGqg1FdPjb4kZqfbuG5TVz9KK+k//5MwfEAUtYG+fCCK7AyupU81
lONpejGBm/aXD4aPDtP4SVZDkjq5njmbZsK0h2weqKmcxm6T0pKa+tH6frknpNTbjWcDOXspPk/a
nA4ExPrZ/13ssjRvgPyFgaPC14yFj7sw2DrSPw1BjV9+GkQoPtknAHyv4TF6qUgK5as0PU6kYvr+
msqkd6nj1c/ZCcLm6icLcr3Rn01Ji/yDx6PCm6wXF5l0JEx0DIUMXvOf6ushaZcd7a9ljBNyxvUF
aKw0sRG+gzqcVaOP1V0avCULoHEJrtTuVTRCBOFAse4LwYPZHJz1Xt5O7MlDz4diD8vya4tyfUWg
j6BwEeGRgAnF+jAODrlGdUd6ooEfeyiXspM9DIEACuQ6lyRssVGvRBudy5qB6rqA8h+t4egzL9yZ
78nBjC/cjChQ8R1EIJ/VCeGxLFxzSfYsOZi1yCOI2PNrwAUfzeJ2JhHzNiuQR1abOYzUq1R6zKPi
SdVAi/XwsjtOa1Vqlo+1Ft5sRo01gUBp3NBEE636P4Mg7yog2b4dqwwdOn54W81YQVt6zcS6KxXC
udEQRLUJZyl6AIulYKZTmdpRSrVgwjmGW3SowbqtVVU9vh+x6tKXKhFdNHeAUZ48iey0W4TiolHN
AmmA2RC/M7eHmiI8QvvOyEDNy2UePxwIQRZMz3NJ5ttEjOLW2nB8/4/44kdR9PNzO8PXENoGRjMZ
ss4+tzWiKAJMGuqjMUWb09Hd8NhuCF0iwludnvL673jAOB/qb2Hu3OqLM+0QtjUKWVzznpjAg8eI
UQpoGIm0AUFxexjza6+fNOoe2x5lRxPrtIeYXvk8PNpxWplulyf/KyfVqnXZHizJTscq7pr+sH7b
tuQ1LkhoKn43VJ1d9NAFt1tGT4VzRSjXbWdmKv92c7+b1gc3gYNTE/FwTs42hN3Gx4ULSkb9YhA9
DLREzwDuWFjou1eAXwp9LKqOzNxhdwFjslkxYntOcOgNfmwOpGdHP2JdLhYCTe3CFTrpQaMarq7U
9UC7oCNswt+QyOekl3RAQ/klBE3uArC0mk8iUiTNnSzFYGTd7vY6pR0r8RJIFO3q7OqLzkq3mdM3
swBu4/E7dQj7/FaD6LLlUw1ZEM4mDU0clyc8IbvCUd/7bFzydJHvOKCaMvK0xbD+gbMGacOR7VZR
54hAc+bXlCeXOgI/GxcEnVRCD2+J0CLWr059oEYdKj8N52Z0Jww8EhFQKMvvSTT3YuDbkcv+aymK
0crQm3CM8/JJUSypED9I6W9t8y1IeH9zToBdsXzYvYuAvT39i7QeUP75V7IMZ31rCIDIqUCkr7+5
H8Rn7AKXY1gk3Woh81KkCf3dWzmiGYYrUXTRo9Rv6K6fu3hFbEkLZGundVrFuuJBd+Uh86Hsjx3C
jwnSXBiXbxjKdmzTVqVeywNpnOTvelXAoBqd6F+igNxbrXW37ijcXvIy6xGjWrm7RMc7hHysJXDe
28k3rrzgNTMeUP+aT4/Gba0aJoo5EXZpIW2u4Xtzyf2lrZdcrvSCVH6DakTavlWUPrssqcbDG+qm
GzslEZ/KBsX8lauivDe9Qsb8DgQMEG6hAr/KeU/gbs6TUk3JMHf8gi9e3Zl+G7kdErky8WGVwa3Z
/YwYv+TfIqW2Q0gZJJw+1vRonLj4wGguri2JxOfnt/ZGtM3iZzJQLSRv83ILRAT1eO5eAIHIZq4T
HEXD/ACnLgItnz9UQt4ZYbWxIw6+u17r5v9c9fvz97n3tbqEStJueg60LDyGYHZ4Y9UdEFmuFYkb
vKZ9LUuitf2fkzkeK8cWTBcundXPHFiFW0bgtGG2vhl6ihBjFqiie800YKWXqlWNmykIu6NnMLG1
L5LxnZl6n0RmDPA39phz6ZI7SU9wTlUOzGhhLkyKXddVW4ymAACiLYT86porn4P7gkMtwRF6BZj6
G5OIl+peRZ4cLiyd5yA4rRRZgb258dz2iT8ZAJKs2Oal3SE9ReV8UKBnvBt4cQXbNRmW0gZRMMCH
788auW1Lf5Iw38qvE0iS3LE+grhc5uR4VhRJFER1nD3NmFSaxo7y7w6AdxweuSVqdVuwJCZYDEfA
D6qTvTv3XLIAcPUXQ7IXJgD0pX0vbsG8dhUgxJNfW5k2gtE9DcBjLGJzYKqareHG3uhzZPSt/q+t
UpxbRohR6q6V2fiEL7D8enqsN3tyAUP8UMS6WpL6jQZhZvKMmctXsqieazey4Cxay34a9H3y/Mau
twH0NlyTjFm+bC2J5DVqU+HxRPW8LwnOrMtfXo1/C4bg7OloyXFL4VEIIaav6NHyrgleCBHJh4Vm
6KrhclSNwQi1lsDaNuWUP1cQNP2iF0dnutJMmEaxlNhF3Ok2E2nR5+RvmXD8cB8080HnRpFVH1oU
7k8AvV7KwDK7ga9AbM/cWJqNSO8BIhLBMRAHZh0UnhcUJrr+Vl+8WRRKUOV1d6hawoUDNsiG/yvY
ET7EkP2KakN80rbPWWLyczNHsAUBxa7XQFgbw4XZ1hOJCmHfPU/YFe44oFFlB8VTNYQLyCsGEgRA
zlhcDw0WTsgOtKu5JNMLirCRif07v2/TzV8Zo9HoZf0eKdLBcah2yOTmO9XLYoiMOsPb9dU0kWUn
hdjE2m3tRg9KXbv08NGdbaLwQJFnncbCcMVT/FodgalnmzEDZLrUYvcbXhOZF87LKepTUjswfxEL
NlWipEBeeea6AcQOowlRqoXnXdYhkVlIhttc4gKqM0VMZ3nte/44Wf+0N/ex2a2lFlyBfiVlpbNB
qgNug6atjDWu0Xtpn5wAgWkMmmi6yT7DoPOL4Ix7hOIPIdfDpYhDP6uxkvI6kMI3BYaCY6EhDzj4
FGrOA82wIvQybVvJb1XWrTndGDUyPk2jo5FRwO7bibeALLpW4f55ia4Y8VYG0FmaJ5g93ZXVdq2f
v4t4mKCpHKjpGKA5BTYUkUs0eS4lURGyhBKY8X/j1jJFXbr3JeIipp6eTYRGAT3E3+VwMi722ph5
f4KNDI5O9kNmUgh+Ma4sH9I6D76p2XzUAMUCYgaJK0gpOLq2090w8vTker2aSFQCtYyMHDd2gDyB
ZLZ6riMnpJlTScUOiwo+kH8yo+7zM6yEzZpxS+72WegBlEDSc89Dp5vA/5E+LNnsA4XpUXIUmBlt
rWDWrNB6Az8zuVy7zfYcNb+vDNAHspXYSAsuLxfCDfYN6XSqeHM902xqr4gUMdybBE73XCMjnJ1E
UnCBJWVJp14xuH94H5KYKPyj7IdhofdgoKh/8Fg3+RgfcWudQhAM8kNKnZ2Ct32+xOF+H7VZmh7w
RwIugxf5GG11j1cekw/CC+VZBzanm95SmIcUVygNiAms0nP4wjX5Xtuf9SO7L4uqgoirMjJCvqHI
DOfALGzI7bLnlCQ01ukThWNv19ZacZ7YTL28UMB7j5WZHmwwHmnysKgr0MJB4BViJq4rkak6DdQH
uwT2pWOcdaY0oL/DVaVM3MpsY1MbgdNOBYssH1GNlLtRP9Jk2b+j73M+h8CTtMeiN5dcQ5YQmGDI
WXNgY9RpPmhN2QmG37n3tV1/xf4ygsJvyz9aQI3EJg+GQegsygZZ/BhRVWvvUupVN8jmcejMnV18
N2a8UK5meCFKFiSleMQToSHLr4KXGt9u3tkw9cFKhOFpnzX+6IdsZQKZvAWTvlRxg2DROIoNCs+i
ubSUrf0+eRK6rPHjDPgsB63htmIkzW13lQg0Z6NS4V+FxAbWh6+RT19nwiUAszdcs42mVQ7vLjQr
xyaCnQjT6zl4m0Fl8HNrBuvZTVUELXH3DHTDRB+ItydlbyyMBbZBO/mOKheKBKNNpfzww9CytIqJ
Bp/sxTxBPZhvRhiXRyXOhWPr56ZJnlAjRBxh9LFiMj9n68U7/66rEUiVQsoKx0mhpiUZVgdWjIK5
jP//tnoJkgp1imltDRj+vNo9+P0/Xo2Uc2I1K4gnDxoUOJCFHfhhrTyE9JYhjnxom9LjQy+TOcCI
PLVrU879VUNIwTqVsf0AzG12s66WzV9pA1D+CF8CBNRK/Xwbc6uLxgvfQICuGrBHtoHQ2xxxpUX/
jqY3/f92LgL9WL+s5y8T7uGiGgRDI3Dz2b2lHbr/7+QHjw17jTzG3IGvLC2EqIw9eebYGgxUMOq5
AqqUOMwYDVbbkB6M8vwtekbypgBiWaWELfbfJDE331Q+Ccmu2zusSihvFUVWa6KmbGyIQ2emxRzH
S1qw+78bBwvq5tubE7piv1pfWCOWUOwrRk8WCXCD/y91l65AUupXMG1ppkAA+mePPEoFOOdkouwJ
Xs8f13k+oGbJYx9YlmyZKXvkPphLoxdljTUSkTkuPXrcvQNdPmae2XKYv5zxvIwoWiTdjHeFreyq
rLsXmbj1PCoo+B4kPme2bePqSGXEXwmgbqOJOtwxzi/00RucMHsINUwniTqGk0n0E0mzPubGT5N5
420L0XUf27Iwbatwl29BkJ2L+uBDp1ybsciQE3H0KcRs+5TVEzQrZBirhb6I9GrIXdcCz8DXA3lr
aoyscigM9Amz9UROWx3fHj5D75iEYQ/Dpx8pbZLN7RD2Qf4WCUXI64kATha+6C/vneE+4POQU3PO
hXBVNxdPRrFLmhSU7wAaIVJxlS/UBe2j5T3uQ/ePGW3T7p7RKPmw8D3ozgXHJVpm+940+L1xJfbr
ec23zzOmw7m19hQWDJo9F8iifVUpZRU9ts372xWCaFmgS0n/R5/OpR2R7y5ar57TZCwgrqH+3MF3
NCQ9FXNQKsMNH/wm2T+8wB0n9FOPuE/vGlvpuc5DVBuR3x8sT05DQBHJk4gr2+3ILlNzaof1r1H7
t95p6Jm5KYe/9s7TQDn0cu+nSaca4OWQrskM7WONLK3AlZW5NUfs8XJZDKseI1CWJnua+7EfFD0K
L93tmqkoOT5FI5phphJ8kH4hh17LMaAVPnJb/14H674Juzre4nV+yEBCkZFim+nNeqsrsyz/1Nyr
jnmYfxz/Qq0HAqgeF5PLt939Fe7i2hSqXHpuAnZqCxmQRA+Zgkk/Ur8qzuEaUOHkofwyXBzuV8hG
LGEa0P3Woc3ubGiFrIdtYFKhu6YkylPwI2W6KTao8nZOyTAN/8wR2xsrP2WXSfnv0GguW6T0VJgt
jo+MDghsOKFK1Iaa9Yk41Tf94iGA1xn2bNtdII0kzoTM5xbTnPRXTw8leAR+P/p37bhrYPatZGbo
kq2SxATBg/mJQ+2VDRclA9naAFHnYKY80qa7yjBKohwKYqFbxKPSBPRGfjn5IUn3CsklkpaJb7Wm
wXpFAsne+/72u8yaeVAfV3B3Zk7549U9WKpNuhizoZXV/jCLpO66txejTBGoTyxknDbKHSmq3YDj
9l0VW7WRt/k3tmha909VNvmlPTNy44qBX7GzvtJELq5WX0YtH3ubEvVNcparc1iaLbhT9vuG/Au3
DEahwpE/IcXvXjhVWBAHym4E2Gdr3F96fYqHK4LWgPeCVorIdP7c/tEDN7CWIANLWnHVzuJnhVkp
EEtYa8TVWT9hRlAOAbJedf6QNHzaCvQ9rW/lFGyuD+YSEDsgPYQgrgm+8utbJ8dMs7yYlnQcFpUu
zoFt8nmdn5sOMsavnysZ9+KqFG5o8KE8bcJiQF0QckTJ/uk0j94s+Fsf+6lYMLlNt64oI17nsuz4
0Ti8E0iXIVSPWvZM0Fy3XH7aS4LzRV60iXLP222eNX0QgXal1n31VtuKUqxRgJ/E0A71AySqBERs
+BscibpaFNKHQ7JMB56Ll43ukZStT66zk8rtR9kx0b0bRu/jj611Hy9OvTs95h1jUrYsNTsmHkvm
rZ9LT0YZ/OUIWoQrk9wMNZ/FOmeSxYMqV4EfT+ekGLfnmgytNAPbM1dmNN3mD4RvSjxVbtb918Z5
KrDRM+hat78+DZQfG39iGf/vn1NaRX4P3w0rHQq+JvFosF+zldJM3lzHj8WsEGF8NSdoi23cVpqc
khqXKoJeNYr92PvVgPb6rZ1uhdiOmo+K4PHwNOhkUEPtwIqvSUwH4RSN2nSXxET9TKiTHA8Qng2J
xuWlGwO+VvNmezPbydVHRp6Ha3ocgtMyrogQqzjiGRKy5wnJtROl8azJH0nX9vWUsXGEFFd6u9TX
ucZHajLGiXbSPcZfsV6ij8bsJs+xxzrm774MLHkrTHuwQ5uOr5EMnaVaHlaan56lgA+50F09PMPU
nu4rtSqxEmRDaAeAzY10maUTMhehuOw7reVD4qbLXrZSB7VBKuM+nn/ImDC9KAwrhhp43lTqppRb
FTpeEbHxub5RhzvAyhkxpQaCNLJhJekEgyvDCDXSffmCIFxh45ci5g4Rho+aSHv20koLpCXmSdkE
FR3g3aQTKgspWt6wyoJmrlgmvUIkAxjiU+Jhutuu2IastLkJ3zaLtolCwC99xs9XeSpm1TTKYB6J
JKiBDg4i/0CghG9jXuUbzwADO4RvdATWgmzcku4SQlQC2/qVjE+YMFbZ95RDejapVNyGGSklbqzl
4DvtKVBY7G2kfOurxXmyid9VRSWh+9MZgplxQvWTWbGtuWhtanl6TDFhm+jOAw1Vah7UadwX0KI/
9hw/OM+jcAA0FYfnSvXoCeLJZctyCOnuLTT7omoEMyJUmAsM2IhIVhQNose9FQDc14k10Rf4ojtZ
ME6tHn0Rggvft7c+rpuNR7/kw7KkfTANuzED2iF15PKf/kNyq/EnFh6Z64igErXbkTBhK/2hVJrp
tZWuxWr0B5tzEY5PJvnTrSUBa8wdC8iQUYUumacOlMraXwP+AKvjYMwm6Ar9EG5dJ8Yd+KIVnV2V
JncOikX/dKVc1t4pzN6ifd4p7/V68kK3qQoIb87ADTs3dPB1tjK4WSVys5MfIF/r5QioDyggoTBT
/V4Hy5yP+pJFhdRSLuCELiEJxuRlCbKOMoVJIBIRWGRdCTqxp+or4itIgBY0awVZEEOtmj6Mz4hV
TlwMlNXWaywnsDVOFQntZsLvRpl+4tqEW4+YUIZezC25isZcM2saWp90EesLCKMaYeXWHPH7jmBB
bAaCKSxU5OagOtjZ4Wu6vLaYqL00HgtRq1arLpi/18kzIe4f3gG1YjLhs6w+yoQ9ayIdfqlLpAI8
As83X75qEXTztODSEjfcmBpM3FvLwbwgxMM+kFNjZcrYTYFTNRA38WL7E2mvg6WuxAmKr3ceJT9J
0xy95fO4LNQxq4hZ7YgwHsu/Zfb48qjJngCjFJvDOIryNEoxRteJn4Q27aQid+7nZhtUT2O6LziP
2sCgzzyTIJa0J9ixOC8di0AiVIltzY3pI5j4etLKDiu11ywCwDUcBJFws2prRXDjN+ynH9MMggQy
1uERdjn6E0HMfFV+hqMJuCwLRrjWdUY4pVAer64RpXcPYfKKMxefjei07j3/XLeaNiY0JImKPMx/
WH8nbH650GgDSs6zz5FnbEYVAaJBCGlfKU3woRo7f9gZdEHBqdAcoccg/y04S+I/gUsqCXrheJph
JRvJOOkYNdiJOT6yZXHaGWmxGTqbIkzn3DkY+8Ooe9zJHAIaCK7YYOpY2YniX/M9nbUAD6qKDjSF
V18VPRd9ilyKmUdiCPdzalZZTrYSdOIH1AkTi+oq0fX+bPeIOrV6Co8WuoC6sKLtixja8e9eP/YX
vb+ecjj7JTQP13gZ5A6h+46zWUJ5EwVHDuASFGWVloLxGEMus5/hiIa+Xj5brn0tkTdNGukYstVu
J9/14927KlwiP8djS2c444iGp+GV7qv+0QWUkhC/zwZtF9XvYeDHVeZ4/Ulp/5Hpx6OFV0cys8Oj
OP7yMuJbYNBCnlNUhsCMqIFAE1368kmpDXJ/AFQbKVvgdH0baauLyTBNSHKdgMAN+L+IJAniXC9p
e33HLfgszBDc0DCK3SmMuAj4O1+KztxQiJOib/sKSx79dOG/x0bqKiapUCboXHUDbJOyOFTYN1zE
yKvKPCJdCyKcc4wMcZRqnNaIK/qEGuCdDdtZY55f3ZCA03s+4XfzpGRU7mhe3GXdE4rxbL9W5JuR
Zc0oa1Zt3DN365s5gBp4q5hbd8UeS36A0J+6MxAxUJcGhEIfhlk0M72m6XmMGmRK2b/A1gEGQD8g
72mmc6iDtixGwtpwXJQMvoiKlzqLMZaaIuP4tF5UWORVuEHBDMsX2rm31ZYdXT3X0QeXvobal9ue
XoHa4DtbxyxXp4cByJQheOHG8TTDv3z7vz/1JzzpZ6iURN2vMudwLk9ATZOA7OjOkbdyw8cc0i8P
9ljGNOlDrSC/zjCg8GNhAcLZZ104Y9rXy4QHqc8rZG52Qr21HL5S4I3wNN9CynGbe6o6SMFzCokd
+6hXBtkXtEAfYwJQMfC5R15MOd3gIhQM6SqkKR7FERdV6VWtwCjhngPsINuYKCrUzqK87IPZpdG2
eRiiA/BCB3e46rYboCBIAvynGSWzaJ6F0wdWoxFC3nBFNfLVt/QEBn+Gej3GlgfOv9fgtYLHf5HV
1lZkW1A+UysgmztHa82PsDYDXvUcl/SIaoXjY7Hutkqwx5WRmM8tiDRn6E7gEE6prgzk/B5fAAz4
d2mrBW/WCY47MtZN2xCY7PlCKlfB4PDvwS7ums7CqFCg4NpG8BrXAV7ADByRk6XWsHQ5XjP9MPcr
c3T1eDQf0sEYVBYwD5RpBPXng+2gfVpd2bYE5aOyXbYpknf+hX0vK4MmliuG+30/+n++yxKwhnMB
5/niP2PawQerm7f86JGyi76sqGg7V7Mgu+8oPK4lcy4+tblVcd2hb8H+NpL4bJUJ3J75ixCkoowM
EyRvGJTwYoVipVrTdqIPxx60pcvDMaWrftlC3MjSD8AYiCwXKgf3yXbKlXlhi4PpcwZ0cQnVLY74
Yhdikrw8iASswTj6r6YDdZk74w8j3qtgqR/kyoBxpK8RDUBvVAMXZnCxje6IqrXgwFrOt8e/sr/I
7b7d5bY/jgml1gC+UCaegP5Ukjq0vouY93spN8O9YKbeqGxxGPdJu00yRHr7AZh7NQnHihgDqjLh
Kinfa50Jevot04Oyx4Lo944V5LbcTc58DBRn93HAw7ORiMBIjp/e+3VNALu5cyAfVtclY3T0bSo/
DQulWldpoSWcTakoBaI4BZnzPFMB/EXJf8Km2/NWCigdH0QFbwpBXAMo7o2H7RD0d6P1f8TLfbMG
bsi5UMEvSJ+PLzlfeqRSbWr+rT1ztzrhpwhKe5YY/EW2S7Fwq2/YfOAPeSeSklSdJla+l5BJsdpi
Ks/w9x9OejQzPDWsi6LQAWi7kFGQgkCGTh0qvolj14gnQTCvRcclCD27vVr2jcMQizjvTN8+iVB+
oiEZMku8rL1E8X0ZIQyeOiLCeJGsXb5xgF/n+cwIujOADN1YPs9tIRCWpKn0OBGiK5rdHWS6mFko
lf66nYZndoibcFFsGv0bMIKB1CqVCCaaUQYYQCYl1ZrNeJxBj0yanv3OTcV5vPNZy+0EQxgeGRi7
eb7qJhcEc9DJyCc03LhuOBgndvBVReCA90JOfDumYTOW7k26RgLyEsr+GOmenY5EVH0XsO47ri9a
n4twlNIzRAaYkt90DfxOYucjeYhy9VRV/EBrBGmEDtE3GTbKOYIz0X5r+xAuG/onYIJAxyNvfdB6
7P6IW6R9jzv//7wwLrlob8GOzkPg8BlfmK/t0sp4WCpCKe57lrCsVMc3T0KrpWFt84Tfph/6Pgvq
a/Eori/ucOItUVLByLjn7yJLEs1XF00KLwO1I1tNK0mL+PHnmcHq15wn5iISvmGNlG1vld6YydaN
px7CqoXYzn14k5Na2SIfAbobg3V7knDwJ+S6joKC3Xy9N4tzvrcqKss/1FX270dCRf0FhjnT+YL2
/Awl9Q41bf7ySnsfH3lVohbeD46Ik9Iza2RZVkgbPwiWVZd+HViwllHtocnayMjZDTTCsXWJrGCH
HyCusyGcBCL0XrxLght86oGPAwnzNs//JpDa4Fg48d+bZvzCl/Bwh8X8jFMxNDANRPFM4dQ9HxER
bLNzxSMQddQg497TyObGePZ5EaunF0d8ug85f4ZjuEgp6Jme4RypBwO6O7eTCR1Wchql+pfliOCj
HRzPrOv+sM+u3l0TD8II5jEkgWwhNN6dqaVmZvAmRE2tx6AYcKoVyOKG+v17QoEMr2p8FhMzJkpn
VK5NnPDlpFiyAsp+Ad50DHweWpzWw9RHDaN5u9Tq0yZL1eBAaNzqOX+BFPifBVK83mC1Go0igE8N
HfdzergQVyzE5HxgEFLwYyCfs1SJNVIGpKv3ZL93wH7Qme0jNYvszU7jONLDJIPwlL/YFyFBBEwi
swV0/RBtn+zltLHheF/JMjQ+/7Vb9/+oEjwwijaJ+rY6Lt8sYzthW6HT+OcA7mVWcBm2nj2dIPyk
YIj1onjeSt70v35wLpN7X+sKY3aw2LJ9tA5vwN7wJ4nBIDZiPWGr/k0YmqbdBBvAthVcH2l5UmJ/
14Z2IXEWfixt0FN/mS+OOh2p3e/9JqNo3gOanAmyCI/wPOUMLzbVmjDC/v3bgWkN/mz/Y7mOzV3v
hCZxevSU8k4KQpAU51iGCIZft8z1Xd/dYZTG/OQGUt2wY0YVKacCbcuSVoJD4twoRBya3KnmHXw+
1gzJhTOXiEG2jE34UtgigTjMtleU4Aemc9SenSHHPVuLkD09BCu4CSPvHZ0TztNX5LK9U7/8oC0e
e4vlr62WcZwhJvt8V6PtKMAqPcA6v6fmMTYpxat/Ebq/5ZzpQp25ViewwNBqsYmPzI+wUF0NjAa8
q02YRfq6tnCHKz9Ou1DxQT3XLbKqdvKx/ErEkSXBrDWrGZouDE709+W1KfpMQ8IMFfkwuSa8jfM9
zYqBEXjBV6omL3Zn9rpWtVcMZEsGrk1W6N67TVr75rtE8Ey2Fz7UYmD+UJyrF8edIq7rdViivC1g
9DPPabEuvBo/OW2jfh+zZvJTx+KS0MSPNWG+y/ePwIbA9HYulhAvegCq5uvKa7BkeidN9ih7nNkO
sJsnT5cDAJM3vhqTgutiIa1HAqJBwaUwtr///L3tXX3WkhbkCAIRCSvQ54Ua7D9W+cvBcsr4x13g
+gK9Y5qThiZ0k77M4m0NAUqULNIMt0C0mql3dm2a+LSI/i4v9rvV0ZVElWITs8GORguzKD3br1EI
wfngE9thZngxzWJvuZnyjxXmyag/b1z8xhPMEhX6ZPqAZl0Titn43Vi2IUpw/BOzLJfcY8r8wywP
xZlm4LhagapvLP5pK8WEHL0tiD/DTT04csgV+ASv6lAduGHseZzlyF9AyP3jqbnp4tZnWL60o8Aq
tzjULzw12zD6UD6+dcTesBfpddEdSk48IJS6wXMwXMeZBk6KiIvxYfhb14dMvxCW7tAz+Ew7TTES
rs1THI9NWB9A6Ro+sn9Pbax6iKhVw8W+XC7NVzOy+BkGpMudjTq1ELaPxNpYjibFlo8nzcpUoPWX
c2ebVPqXVOO+2FiI8aGs6GQ0t0ckkXGou9Abha8xEuS0Ng5H37CjZe1ZvFY+nDyT0Jf4nQ9cIL3E
eibN0yTdOqeDvAiGw53QIheqaLNZNtDJUcXas0Nyzaz9cjxfLAiSZmel4T75+PdlIeTjF0R1zKdk
S6KbwVGtl4+j3tRmzGhKfZZrKJXBlepRzqKRwnJh7uoT6OSHWLtQoe+7MxkvUZcu5NdYxX9doJJQ
oc3rI6Mv+iccfbbtZ5QXv7zc5ShbdeO9LSS4bYqNkEjXVdkxKE15I7uBxbNOgEzA4GdDjgjSpkWd
ik/HZlnu3cRRAXz5gmA4v5obppU1WwdBspmm/v0qAwTw/pY4Fcz7U3wbE9zv+H27+rtWczuJzjc2
RCMvHhYEQAT/h5dY6yZVd6SMoDLjv0P/uQ7Vmr23coHcQ5nO9L8tZPbsZKfKQdN/mxPRNqy54N7A
SHuIruP+5GD20hFgMFS9NX7yWxQg1rWabfSg0wvadEKShndGlWp/vHn1wGcnUZZEjRVDKPODZXNU
8fV0QytH/tyItxhAIyw9YonGbEk6Hurd1eY8NkgMBzdz3rPJGfiLsrltashsUBJvUTpaGjGiFdtL
qrz6xGVfrlBAd496kRlBiHY885SSAd6+UZle6PgyRf1esZZNAjti7cGxZIl2QOwUbHVYGUWk+19E
cXRuSzYLSVvjyn7eOAZP95mgxILyxvClqhHYPwhOgJCeP19yGH/jPL14m2RQCDOHzRBdyBfaTP2O
7uHkHiI0VokEo35UgjaX7a9Bxz9sEk9onxTezsUuhCLz5EKzaon/ipP2RUDwOuLzo52HMAdZSpQu
lyxdpQQdJBxdhvxXGZhS+moNz9d7dBjeaSE1eqPVPFtyxy89IFh9BvWYOn0mRhbEOQEWoEXNijUH
X8dVjsTe7fcr4jwi0BQ8OFbImoQXkSaV3qEpkpr1aHZUE4ypD9UKCgj7C5gB+AiuQcpzLYSwF/ZW
JtevM7jhbh7BSLVTj6/hP0vFb0otW4ht7uQngpILCE9UF6hhs4YoE+swHztzmWF9bISujmbBR99+
e2MzjGAi9C6fmK969ZQyTw8UOduAyW0KhA+RWvAfvwXws2Kvtdk4V8ge5lnpFHiAgPCfaQbU3d/e
gD/xgpaLqkwGYTOa5rrWVTz1cL2iW7utDnQvE957WUsnLfxbM4TCrpEQvxb1uXNHN/fZh0re1OhN
qxlPoM8snW/iDbuoNan+KBT13iaBkuDyMNP0phZJfM56/CkK7TPyjgMnWn8guYzf0CDktgoqO9Gs
TRLtfx3IcvzyMz1xHvlq6fmFo/aN7PGrwXrRkgVqtxPsJfXfp5X0gF6Gbp6/5EWJRWSpzfy0jYXl
T9iNTfZKK47dMfcWW2Jln0SFV6YJXKbqsyQg2UnDa0QKDTtTASE/cviY3ayyJhLyMimOnerosUZp
kKs+e3qo9Vw3lluur4v/N87s+vdboq65hPjM7B7Od54zFVPqjpu5NgeE63+qXF4A72eMHupWwD9W
p7PQFqHGbl1RrNcvTbyPz3UJzsMGyIVyipni0w5nvfWnnjrsh4yxMhX7ANSxnWivLqbZ5zkoHiNy
WQn1VHeIQkY3pRZdswJ39rSrT1mCzzKdWGiTWf33NWv1aTr9Vl3eO1pk1YqpJWyDjqbKGrez4aSV
ewX4R9FEp9ro+uTi7EbijtMgVXvPRNG2L5+l369qtsV9w7wSJoOVd/eOfUP0FhRAKFunLwO5WBpv
Mz0WXVJatnBLrB3rzuJ6l4LwsA7ewO+SW+FymDKbU35aV/enw/0MJmOuEjJqYCwSDYFnyDy6jGm9
1zJxXBnzucAg19jWtuQJIPFEQ3Pqd2tjw1tay7R1yMv687iBG+se4OT/ykWkvFxJKDjl8/zfriZ9
WhR/3YAwRXtied5QCccwHbnFAKnGKK/5cw0V//rN1+GcRzWcjj+XUgjBbiPn2jy1OS0spV5CH7OZ
GjEzICPwTckQCiLZJnJGMbJH16dgD0M2d+ds+M+rYtdCvvIW2WADuirpSI1s1R/uMBdU82nkNcDa
9T2h0axqJvbS6pDEcy8/LT41qzsGeMr5aEh2271w5vP4P+gP7RuCaiGjMqO1duhm4XUTKLRNuk1p
iVFSakiZmy51NXc0SJjg7hIGPZBc+HSA6W5zB5axnsJu2D/Kw9DPyOJ3COyA+ApIH0ABc0b67TKN
QM9NMbPnaBNGz/5kzDzbO/IXfmEHPkFIY35ZjXcg/B7TmkBsnvoxr4q36oC5HOuu17/AtdUI5YBM
6HKTd8RMQ5HwJU/SAkTT9fm0w+nhiRf7mOvUSdI+I2UUGFNSRJGHJk+jB0xJfOZ3GX6H4eNJvWaz
5/tW9xyr6bcS8aF49jA7xpPqKVyzK3xizTHsm3Q7UMPPqkzBF8fpqYPe1lVBolGAJz20BwtNOfX6
12oBAYsnSjLHrNyYtb+fdrAQXn8v5yimLEF2IB+N75vMKTIgu73bYIjY8Pa1nco6LKcSrNxRzutG
8P71yx2q7gWXclFVXn1llqzSgFaIgPFnssAoY4xTTeTMFhj71akj5lTTWE9Vk4d9ogXEfaCE8aGp
hZlrJko12sjTkiH2IHJzj7LgST6LAetzCnJoSz3H5+Du2wVKR30PFQGaoCiVpe827mMtfaD5U2Vs
N0qnl8xUAoyEVkMR9NLCJ+jezJzVuieebPdl4APy39IdZbAVQwrxxUV/zxVdvTo87a7UN3c0iUJg
oVKbBJk/VroksxXBdVl+8t/s57GSiwpY+OW2cleGeJX97ptRjgtuGcu1k51xbJMdJtQGllOdIpDb
PAFNrVIyj62RArraidojb8g1nCmEWA6S2vBHKh9yAMaCjC4OOOdXBivMphYJi1k2JC12MPeutSlm
ypl4e1QhZb4470YQQtee6Y8/PBLZujek47SPZrWNmojnBl9u354jCQcyGyq6gidanyyHBivN06ZD
nP0WJpIoBcrhgdW991ofatTuBxsvspFWb7ZJAVXWMzwAUCvRF3D7uOGN4GcEryBhETzR9AJ+retg
61SM2FETFvZWnXS8/vC2bjPawVZIOUqNNzYxtX62KdVGwBpcIa12t1OVTFRDP8TGM6uISL+5yHxX
jdI7wDk5r9dnw+5+4zN/hrSpRcoIT2VkpZ6YevuCVHiRcJ7dyQr84ILta/oslbMqB8Pm9Ff3jfrA
9N/t4ndGMp/V90mQvHq0FoXk5wEG8nOD/x0LxQHeX9iHh23MIa2Kk0saGhUISL8SRYVdbywyIkaT
eMcxmC0XNiurLqzQ2jVeFetFz54zdP6WEipqzkRnZGhHzTz0+laug4OdEr73yMPJLjQmGtjI10qI
23wrSCtBCzDpvG3sOCNeo0pShbLb267vF5/hOx6bY6fF1eE+YIXcuHmmCYInPOcOM/pBnpH/dac2
ydI9je1eL7qYLMo7+q5nffOwctxxLgSHOpndZoMEOnJkMMrHaLoT190dKXr4WnhlJqxC8gE9l1yV
IvXZzGY1xpR8iSaZi81LdhVo0hDvQEtKNrCW5bu7Z4AKekS/TsNubaC4phT0eW79SUHgnLyIT0ET
dnzT/NmR96YWoaRu5Dddf2XCb96SvyUU0csT1AU1u5PLPr1V5IAkz5A5NGKqSMHBH/Ox1anH4fd/
2aJZTQonG9d1jJ3iNrxu/Bcje/8Uf7pZaEoH8mvx+f/X8UOweN0odFatUMB4w0Gmgt/NSEouEytN
sQGX6FsN/TiQ06kk98VaMkmwII6ZHgiVbuhOQZVsd0rfH9Z51gEIlFYdLX6ve536ZkvEDeP5q3+C
2brd/4BxuUhYOSTkSYcaZFSCSme5oocKLGBcqxHKyN/jtAYsmC1Ht2P+30+/vv/l4qlOSr5GY6qo
FyPyyR8bswmwm3H54CHO2QqxoKRnBZCQtx95/MnMJwHy4jHBBRUhJf0dthMfRbzE4x3+C+vJMhiK
2D9oj0MHHM9uAE2fHa+l+qgshKemo6+0c4H41GoRWiKU8Phj9JnYMXSWgpcnikAcEjdoK7I83ycF
adQ9FsouiGIvr6l+Al6Nk3qDkGXyQDOa032Js6cV1GU2KUPJD4al9nVSDqc4ZE5a69rUv5LgP19D
j7LlvWSmjACybaHMsCnUbmXBswXJTOTcO+jqDJlbhIB+BVgV0i9RpR2WVxoCUULf/f9CV3DRlwob
ZPsdgvsmYK5sqMncpHGs5EOREemqV93vQztUZWNTg6qXOXid81u+y8+LswsS+ovDty5TkGgOvSH7
2Z1bT9x89jhCH9qe1NVTR286NNWk3IX9Q0QSCOx8+FygQpFlIFBRBO0XpboAONZ3dRvX60x7g+r0
7wreh5NIhnrkS7p4arzPTIfgKkDRwEvOIY+Ngfim2B462C84oZkDqF0dGi1RIlhqDtI3S4f5z6Ad
XXY1hqmBxZoKi72NTxhRHMGPgyNy4U60TsHcMmFIjh9RAvcba+xML8i3rI+KPlnFB8Hs8TH163Mz
TYKWZXiFOQc2fWkeShqm2ojNod3uHh81WUx8mukByxVr6FQTWzelnS0kTyQd8WitU5DK9MuYeL/p
DcuQwoJ9F45GHPlBEGfgXfVlA5vyM5URqccz1qaCcGSfMsscE4Th1hOlt+3MC+ltQk4FoCprcgyL
N6yeGrxP+5h4FuNodZocx8NX1Vo03UB7h9S6dz7aoBSDhtLRT7Wr+XOCABdRXT6XiflgWL1cf3oU
8c7BxwiOY8/Ou4ryGhafmoeceb5hTmPYMtMPJv1sAOf1kbr/X5OW12M6KG8SPfeq60a2/ieSBxTE
mWylG2OsbBsdfePZW77oP8780SwM3XIrQsZyzIRKDy+8H7R91adJa9pM0b/rarZf7QhEkggLpDub
cRFL/xHSRwefIo4klQ6KmmH4JPm+Vjkk/FAb9wAaj83H0oMu44TrXhyFPHn+J4wmgCoFzGJbUBw7
rqsoYkQ2pJkEUpuYijJSFrzZSlA1DYOtS4QgJo+U6ybOioT41E5lX2fKwfzTAOYArcBsBwihZmxV
lFSYYjv1Qd4okZnfE6e7Xbmmja9dDbUON0zWQYYWmeJ7YHoGaYyaBC2CtVx5ex77oQ2lZORE6x8r
R6WxcRy+ouWYjtPL1wMwGV/BSbFuFQrMfXM4qIGC6wU6SiS0GpLcSz7pCd3lUkIu7KieAcBstucI
2zbbCBAGuSgxl05aH8gYrXMGiC3MQe/DB+pAoImBrHkVxEQ+kv7q0GE3Cf5r7EdG/UH63q2rUQ3m
BvpLJiiJEpH1mzz9S5zBTUpnfaHESgMgKT8aObYwPFlJENmC0Afsii3iTEJRz5oVvMLxk5HKVEeQ
vYk0neBrq+nVTrMbPjhb0edtffe6uzY8jv+E1zW/1YoqltdPU+afvZCJkQp5+JlzrQ2gQxwQyOBu
gEs0eYrui5XhfEjyW6Mg9Hr5eyXBfg0YhqVB2pJKD69fnXPW/xR/y6MYiMBt1W2U7WE817k9Dy7r
bcu7aXjTmZP+JrTMGeA3DBabCP6MC0OfYYy1RD/S0s9/Inr1hSSEzrbh+dy0XqQpsJuwOe/qDwXT
xwwjgMPxX44NEZ32se8BZ2dee7A2X19UGRqNHy/1/XHqw6XyYXH3mhpjWJAUosOLOo8xRLlr3tPG
TnrfmrZcxqjCtZT53VParSWU1oSdU1evS66/JzVV4QgKY/XRwqa6LgEWF3HL/G436QY2awLnfWxa
FhLWnNYs8bM/o/rYSMx/mb0GCmhBAvjDCmjM3et0BM7SEPnt682mT+VuC8nyA5q3WGiXE264/rwZ
CAT29nYk4xnSY+9idD8DMH011UKiAvEBZrS+OMeC4cv+ghpwcnySvgkCzn6VJVrSYmsZFOwrRWJf
ay05RgzVkXOCd88Sbc1LPhzeUl0FO5lUVvJ+DCVvWuQoh+04zd39AlGYIcoCXQgMSY3TAkUMkO1n
FToNMP5gU3h6Xart4YoGJVEhOPDrHp67NQDrzlryQUbzxR9Qd0ilbbG8fPlt3ey3fHaB5thHvFq9
mHrIk6bUaYUY0HOtpbS1x353YAiTzpIGhR6Xc6BVGjuR9dpuGB2Ta+nYFBUkdM69GMO9aqOT2Hcy
CT/onWgL1Wo+wmmtyqVlUc0WxqsxKm6W2eANDPXhbqtrNn8aC5vklURMc3p3l5RRNaVt2C88rI35
nIU9hp+jo149hKi67ZZyX6DzrgM9GgTQ3StnQy/NDNjpD5Sf0AA7K8x0k3DqPXyJdjzoID6dhHAH
ntZNM6Vxbh8JKElV+S4JkbHHcwfaDjV9IvMNCjRRvCBwJpL28Yf6eFAIlK03w4tTwV9Gg2PyaC5E
J2E0kdHfLeH5pdxkRmLHAPSfOKh9ryqhi1zszVJF32nP3QpsQ4laW3m6V2E/oG1sY/6iamvtOj4e
CM/JHo0rT7L3uCA6u9Ol8sxeXqdCKnJLu4VfyzAYT3Ux8CHKRb/oKztrhli1uWBLtpvfllNdGcTJ
0ONvwjMXbdVMntQ6ctpYGLc/1yiwAnkv3jMGnrFd8JJwX82wykhZREqgUH2BuX+SBIRVS7YimzYf
6ZiFW3hUlCaepse3fpRk+nniRGEFJRG+7H6+/naJYhDLkkSWLSmtjukvUYumSCDP/UDkCQX5wolm
haY0boYuevdWXE/x2iNlZUENuBJH2HCCvCdN7tns+gNqx9bXFwvycmWRz2+Kzvq380tfut4na1fy
Z/0ItGg/mkH1QvfzTMQ68aO/BuVZfuyWBCG13WMh/Kk+3ahixciUVEyGda1pGdO9z/RGSkMSR+eW
8aXL35WxeX+9CoN/iM/hxDggqzFIfetqC+85lUKOyHT7vTlZHzVrw3YgMNGsOnHjTReTkUerGDZv
KjeA5+rp/zHNeL2nVOkkuWH1w/Kw1mf66Ow1KII3cgeD9JWOb6gudjaQtjeoQ1VAbXqE/2pOh96J
RUio5k0H8pr/koxw2/m+RjLXtGzZhuPwT+xtS/N99dPTnm528Z1jsHxLo+8V/9dCtiim+kEF/Bcf
CkppIB4g6kWe6N3JGhQ/VKdQFKee1lO1+d2pZ1X/ABEX50U13DHFd3hM1iueQHeyGUxZI4qT1rh+
wcSmpxMQ7DqKZxU5odXC8kIopZ4somCN/4CTnOZJ54kI4OuiRDF8bg+nNIHePHWEOGH29Okby0cl
Ukc0Tn2hImAbLzE6KPonk4bll0zPdjQMubStFvqwgIcoJRzJM2f3c4Z0JsK8HtOegmGD3ekkO079
AFqJRK2KnoWhrjNYeDCClD0uyBGtGFoBteNHFVe0lfkL+PbTEga6cZf+ZSDsqd+6LI7B7Dieedf2
p+akd+XDp0bZyBOyXdI3bwhqQ2piy5RCUnQN5Sbiv3/WuBMMwrn9MjWc8dJJCuKwjMpJ9I3r5ymj
acxt4A82IbFUR1wXDo3j4Vdv81dPWqOpg8TodD+JBnGlzp5MMQAr6Mfljni8RKNpYQiKQAmEQwL7
clcxZ9Hatx/wiJtldYDHyr7MBIbMYkD6ZjFABiynAzkjmNXGr06HUBqKJuG99SUVI8cana1xv67U
DAUQgh+Lg4Zf84p/HW4kl4Rp3GhRXMicpUArhAcX5YdFZcfTFisf7T5aNNEMjtOJSMEiVF+Y8djl
2PngHUlKg6zDk54SUzo5T0wS07z+ZhpXr/WT1IThcncCvqfxVjCj1TNTYHU1COt0K0m8xEzf4ej9
i3PuzeW9PNgIzu5ywvqqzVkqpsxvNXt97zqzRyWz51wOM0kC9HbOTETD8d6maFETbdN6Gp8AmOPy
rJ8zEEdekEW6yvhqmEMIQAJz0A05GTUTusHsDhczWNujhMDnS3GdoChTV+hMLAfLrIkcYJHD99XG
YrQPbgnCElW8PqL6Qptmbdq6C+9SsqetBMq1oXpPFTmRliIthJ9f/4FyBYLj9blHf0VNaIVyoaSO
Ix93Dk/P4kC3YJ6bPZVI5nzFGqLjwZbCtw/ZwJ5TcEqOUJr4jetpZQAWyPfnIv7iPWosciK4cpHQ
HaLMfn6ATfuSBIm+ym4reQ6qjBacm/tQ5ZgJs8K/NipZzJ3JvKza8oH8veKqmQml6EoogLqpLZQM
U71wagNUlVxVGTzwxevi97my7RK+jkrz9CEsKAW7ubOf0vXu8FRwaJd+8jukyoPfEQWBIPSstj2B
hsqmXl5ghOWAapqtBk9yoLlOOQP8W7dKQR7tVrnujMAuAPOLza7xcvvXMKQvmRijmOHW8mp37uWa
7zIupgt9vAeAGhHXw5ZYJhInu/qIrSNC8NSctTWTIQ5U0VsYmmMWwoqYD4Dm5XFrYQRGOzGO1hAD
D3PnRp2TlOL2hW14rP4Fe0Tiq4UntCAg1MNig4q5P+5ojuBwNzpXPycgifdVXmQpoP2mFGETVbEO
WkxpdnEzuLiakity/csqo5vxkqT/j+OoxADlSLuWYq8tVvc/kTkHqlf1upmUyepTviOSLhVOuPw2
MMMtRff9eZn56rUutoiyPmog3+QIJqOBqR2+f/NMuea5S0HGq98JinizuiZir4K6nCwEBk2fLRyy
+4tFraN0kKI7iwUFecRhzoQBG1uZjqha2/n49M+pvaluapOsbFX/u7e583pW6xVP3kVB8WPks67E
1NZ2WIc2jt9oxjQXgieVT38EXTgJytXbHC4ncySFZ6zoxnus8ssuZvg6w8IG8Vr9kD/5X35Z+Xff
wmTCt6I0VEW+ugXJ8Lcx46srdu5hPUCjFd+3hKotNedmlwON7Gj3Qma5PKwhXNhx2NOhJHd61DdY
Oce1kLwinMPoa5luS3KotBTyinGYnKxTlMM83djt7OkNmSt6sXwnb25cp3K3DpJ5lpk4ESJ7v4P9
ptmksstL3PQePFYPPrWCghYqYRNGR8tkyfB2z4eXYJANPtR6DBthxQsWiQnCQgeUESB66Y4Me0bG
K9FYoM6PitOJ/ZuqWoy9Cn6Ez9WBDM0KNlIp/nPGVJfV01n+JO1X4Qd2HOGIok5m+5/HTgojfV9g
G2k1oBg4q1Wc7R+mQ05Kn2avBOG+dwsWqYqRrjoqNhBggxWptNLymNKWQbg9QMOb/szKXviI+vBq
36x2RMsxMTvGkpSWyC2E6Mxa30djSwoHGsbpEGsfom8x7Pssd8IDwgp16M6wRD4MlWq5DsFhyWXY
rsmvAwrHQ1Z3rSM6BnG1caLORAKv0AhGMCWAPzBcJKKfCczbD8+pQjLA25KkISySh3Y9bpwCrSu3
DrkCIZiLiDerUADJfPSuiy/jDd13oaaIucymgj09cYKw3FcGWVNY12tlyogO6+EVhX01Gi5SJ0QW
dBrHQWzO5qBKD0c4ON7IUZPCOmm6cgHr4CWL+UGSIiP09POQUNJdUieOSKJ4GTSFjnOE+4Pw3sl4
H2CBM8D/YPrUFYpEk8sVWiOK3QpvpZ+jiYmQp/gE/H7EGC5evDGFObCrVli7dHemOR8Vp8nQDiwF
5LKEFQO6IZ7dcFXlMuC6a5pb6wz4xyq6wrAnR25mEaNZ1iQnKckNKJnMO3WspGOABDbNuOKedEPg
BzlgViNZnR646N286zT25gF5MKsXhHIVjAjOqNhg+7fSRZiYrsoyRV2hW/NvcY33YqSgK6eSue2S
LVe2dU7F52Nlpc1NfndmVdNiitm3V9DwTv5QR6UN65e+6UZUxORgdYKR6GZZaktHc+hV6WsYdH+8
6cg7Iev6AY9lrgFpqgQwTeJvzO6Ocr4kCf0OxEDyxKH/pfUQfwak/95GElt9FyyhB3BXYRDEr2XP
2PDSofC8vJEuKcNOWO+I43v9KqpTQmjhNRuQ16OqGpmMvSFeUnpA7pkwnKkWohJYQvW2L9a7PyVI
RSb1sWO2ojpkoMRY+md+qVWZ6jAzCLaQikUmUgfVEm4ZNH2Hzc+KbcUs/XYayTRW1jTp50Jhm+nu
LRrv6CdguFYf1fi0uvsN6jEu5v2EyBKIgXUx91giLWiIttB5hd5+Ynha71vG+kCZsPikR45gSLQ2
6hgkMtxdqlkrwSOC8lGClLOqWbbNmvt60o8bNXof1hBY7G90+S0Jg6noHMwgDryevGmUDQf66p+Z
qYvJT11yRTFdSyrxAzANo4sgEP0bQUstQ9vMy7RT47iq6jZh08tNegVEGWRWKtxoh4gs4USCNCOa
VOq3FSGyUwuHQaKffPN+v1DiQ38VlO0p13slKiqjq4ElAf1x1dyCDahxUkPgGkRKgrebXtklEqXE
77QxV8FnnxOt5tVzpBZCQmb+I4avQPUas0PYp579j0/RDVp+dJ4vuS+Ty0nGxR0tJ9cIxFNeBKNB
z7FTEZd0yWZoxijj48f89swhb6r6YunXBmOdz6wBQO7KecJ43/5DM2g9x80k2+HsE5ksltXszJzA
ELn8JzHn4Z7ddAnAE/tPkW/jjHXOVVbBs6viT/bQRCi4VUWvXYEjtJnCuUp/5182BlJau7ztWfVp
T9p7r1f3dTQiVovo56eXRGp27URoMVBD6R4J9zwwXaCwQzJJlaMnIQiROXRsX5MvEHDYknezl7qL
UBOuwNtG9hcd2v2EGFkFTqcd9vSYX/Q3h0ZkIXHAFnXxrh3hA1dttTZ/jaD5aULtbLNDo+BqOeyt
v2zhZYpd3jar9N7q0rPx7iKFRYW4BsmYrn8laQvQVdR0cPqwOTyVJ9ZBQxatXtj/3xBZJJSYdmzp
oQwkkHDCmpRSECmEZ3/gs30DmdVlMg0I4lswQHPcCc50fyrpkKCTc2ddw5uePZipWeM+mcTB+tPx
MBz0E1zYAvEriZDnk4vExB1V/HaRFPifk/z5dnmQ5MhcKhOclGwmbRQIkDeIMZ+8jtnt0cmrlscp
t0Kk0ITPVE9A86KRsa4dmaJrGOBEayiRsIw7WOxi9u6OVzF9n5zJuKBZbJ+LC2LU16MV3GyOLCd8
OfhE6D3hqnS3OCaM4W6FnmPXq/Qc+7yGGMo36AI5Zazwcv/hcsKhwaEP12a1eRZYu0eakvw+3p3a
E3C6fOfa/M9iNqMtSmIxRt5GCrgUWV6eimFgw2rYDTBX7IRsWlidNqm2JGIUQNynS/FomRQq86Bs
Tewy7j+Z+/tQTIPcGeqI+EgIo8SQcxQkzpDMFx9li1/FVF6DZD+gF+qa7A/31M3P3CuRp0Ustpnz
GDbXuhXmb4rHcREwZ7HoO1jo6MDhjNgjibBlXxXnDGD8ynKU6FgWsdU8BsxH00MvR/FDaw6SNtXa
40OX/0cTCvp+dz9jzAvnM6LR0GnDWiVUx6ciFuu1TKxk0p3DGuWrpcM93z6fS9SEwNLT4sU5xZmn
+V8BaxyY6XAf6PNoSEKp7Ruedq+5if3f4q11dU3oLwBlY1mRMAfDCdCcAMU/d9a5sUGi1bpXqg1Y
Teu7H8c4GiyioRpocjeVGtq97mWK9TK7vDb3fr+9OT9JciFL5qcjBAL8WUw7OCFkgALRqmkZFyOi
aYzcf7xkonRb19xRETePjsjOQHt7sK/KUiUawlJ6sQgSPu1givLSY1pQttUYEwHIXOBvDYJifLMd
VqmmlZu6pBW4sq+MauYyZduaiqxTzbp+AmZMn7vKxIXYm8GzhTn0VGLWJqvqwkTHR5aB2ITnDhXK
HcpkMtP4AGu+KIdx5CfLqOFG2qCzqjLzTT8InJ/qLWu+chuhccK0DXOFgGK6Be5osHh0XDePIgpr
NR2qY8z9xk3EYAg/ujB7b0kJwqSPNQeOdNAvEmp5JWyacjw3XGf1j4QZzmJwB2e7BFxg3VvSYMtZ
IuyUsgg11ije+K2uZ0130DToVUp91YICiRQIEl8D2QjrAC3D4bTRyhizb9OpsPqZxv6onDJs4cQq
ngyj/pmXkkNyFvoQDJKQHCHjuzbz1e/VZd8YOk6WSk0vAqlrYUlzNmMao3UBiXalCkOKN8dsYnVS
yRR54c24ksdewK7acf6tNMRMs5KZimUovHL9t6mYlWcUTEX/ApZhFt1JW5lDEWu9ZGztBylJ400s
7r+Mri84ZksFcuACG1HpPN/5iEZa3ImYrPKwf8vxb+ta26FuhllJ9y+IZYp26f/9JZhimCMPGK3S
1p/5LWsUGQW2BG9rMU1NbBVP7lJOTvUpMHV+K3YaTwgMY+Ep1nOU3YHNV3lTyPTpkNHDXQTcdlpB
ACWo0ylC0bxTuqaibC3a0HXXPxm4FXatYqewN8MLbNGTe6vMFrMSGMFFZNLJu803uv4KgZdnWouV
SXgivbOn639Mo3U6sGG6dWVnbUSulqRCAGL/gGWgUii+Xza+uQ0nqz365B/hZIKQCc+g/x4Avuxp
VJ60RzKVIP/ybapGBGUlp1J9cpHvHMuf00euhbGnlzSPjGmGzzvKGiLtUw6hIfNUBupKwWYUZJW0
9F6ybfrjFktcLVpScxH9F9RR7wBkqGsUs9c6BQgt+ioM1jl2HFXwuLm76tmazNVL3QgmmOYBJd8l
aUZS4yAtUVy5o++0AcSplKWKdfvZ/WIgPyVyWFoVU+M93mBxh1xlUNPyP/78OUTh/x7g8t5vvfNz
eMxm6jKbgEaPp4/oXNwSgdmUCGQZ2bdvOLKDBcnutX/8A1xEuR76crXOVB86WXbWYgwDzMc40FlY
YVz7gO4iIjO9gYqo4JpTzIn1GZp59wvQwnleoxyafo+bSEEbMGbqf5ysrsz7OpYzEuexR6ZUs0bG
gc8PniPfF1P/cA4TeMiIozJZRP1WfWkk7tlrqRVT4I7K7Wrl0oC43bQrKnsXiCrxsTtJ+7Ux4ReD
geuPmFvB9OyD03W1coofhekSBk/gioiEWBTdV41IA5TYrfI/vkvRUo4iELUVbR4AV5n4SPdVZYhu
o1KrezKcyOfwElVn+nuQ2Mpa82SgFA2hBGm2+Ofimefxy7FV4zu8HFvPVMStOVszwM4xmymUUr/6
ISUyvwXN+hlow3SbSM0mwO1FctW3Fnl6P21TliwDidxAnLSkcVgGlk1WCmK5w4XXUyLIg+KVMIj1
6x/iTb/JoZjA4inPPYHGem7H7toQykQZLqtw2QzHColY3UHoL+m8Q2F3KHKJbbdHxWfpbFVuzI7R
UBV2se1X9dU0yw6DORfQq1f6/wZSHe0CRxSMmslTAqhZXie25VzAuZkztNda9qjhO39DOY3CQW+D
xqJYoqsGnqbTpEXAVKQ7L6fsBE1q5+kX67VFvspkzuEgn4vji9d0lrWIfUEvncqUSBbMDMpENXwE
IpcfNEV8xKeDhKJczzzXWwP1RD261xHT/yERUYru96JWy+GynQQViChi2fomtZ8q45VeApPvFtkf
hyrP/pXFlQb0Hon4Hhr8m3R4ydS9zUK35vfAaRl2PdzGhcI+HO59dX/jWZ5ua3bwC3VmR2HsIRtG
lufNlIqrs2y9H97tTMjqSHDxcbTYoK73cLl2h8rh3exVPe7dlPueD9ke9M/tP+kbFzZxaijip/1j
JKtvu+FaxyQk5puKO7OeY6thre3fSc6J0h7oVjfFDPeK9s2wu9oZETJZvrpFlow5qdPILcRKT9Y6
6HPk5iYDATRs1DEW6luWyq9/NeSuyUX/WxPFXr/p/ixYkQ6vB2XRY9CqjbopwhWUNe5iqmhwpM52
htZ91gLcEDE/iNpYfTHWgOuxTnK+kVeXDIzJ5E/o096DWWd2NKcdlVNPEVM+ZXbyetl74cEgdudl
MJdtIX+bi9mvF9tIDpiobkpFxjGWpfxysBwiYDXU+emblZhR3uKFTKTTgCjzbfCbb4C2Hh8ACcdt
Q9oIIc2YZxqVGFVdT/yFkhRh8o+oE/AOssNFCK6On2Gy19GZxMA50GAPp1+taFVlUMmG5y4weieu
JlA88aWgBN8UzTUhYLrw8rQTnCFRkN+rVP4lqkI7l6rEVNEaaYFoQAYDoM84ku/HbUQn2FDuo0qh
UAgxAFZRijgG6zJ3IZSzdloEbv7ZN+dva8+CZigQJFk6JQhbHKglIiDHHDOCUDiy+MoebjY/T8Kj
mGNMiS8NAjDqfhTUSJ7ETB2bbJcoDmnshOWk01NmdQTsl94KKWyrH3wnxUcm/fKwYMA6ygAy+0yv
vv33uQJxOG06P/WVl3+o//n/phKygxpVNvoIqYVjBQRtA7UbPLPqXfJRoLqN58H3d8WGJzQrms/5
ByIEBaPF0+5BEqf9ug8fAVAs3elsVtA5HL/KemCxWK/D2+NJzT3bsPtLMREW/R1L9mHqZqzrn/Qs
JYiuWzZw0Q4sSIzgSTSU0B3rHCBzXf4VunI+f/wjkXSwbhM4giD1Qqg7AZ2lBuDCHVCwA/kSXRRF
LyNaNdLoA5wZPRRrtm4eQjq+1F6mPI6/fxG9eIUN5xdLaei69ZN9TSEZ+ERiMgdN7cw5YzpNh81e
2Eirsds9hxQuc6bMR6m/fqrXvCP7ETdN2eHg0TuVRFDpQ/BxYu+5rSmgsPy1qJlxvhC4UZPLO9j3
AMsiOmk7ZigsJ4yCnd4SXbEmUjCc2C7GBbYmDj83EoK+nG0URXUoAsmaxwwJfxEL/o/7X26FeSt1
s8j7qBcdSWEaZoU9luGHZ+aRgONZu+AzvkBZXALzxoIZTMSEocG5iD08DUJ3sDJFt2UJ/w8uOun+
yVH3RWpUxKgeRP7ZAIr1dFxhon32GOvhfRLz6OkpeGghb4fvRqb28gkPQQnLOqrg7UU/YmX0HH1A
Q6ZKB+5iPRMH8jS9k35A1mtyZXaIFIfzBfoXJkvAmdvkG3U18Yox83NX+IGJmdLj3hp4ymxjVmNb
bO3kueqG/nEbsegLDWyx6iDq4grBTHZ6emoRC8z2ZlTU7odLzojtW8crd+fIyqPzLlr8KAhjLe1u
XjsXLULMwZzSEydjQxGuO/kfbHLrbmGJcXtunJSzgxu9u/8cj2tsZngesc5xALqQt5Rk4/HqqJWW
wQ8NGHfKdJ6ZLIsZfw2EsWZk0JYuiubekWEPCXxpNlc6A7z5mZjGHm63q/7DpWqsTfG6rLNitjIH
8sEIKrAljQ2fbGBGclptxR2rZUShWp7sHbLqpvsAvMSm4t4qKBgt9JaLY3vISCFmHlWUI3gG0NK3
QQhvk9c3WLiP8RdlGe1qx1sFSmC7xxZzxKRsTCLC9xiktm/kRoVb1DfYWe5+LdESuYYG9l/Z/mU8
bZlU1s4QU8a+BU/RlDSuCLAFnfmg6cY/O683TPvF68abDDcjPj6vIdYBvzS+km+GZqgybk4fNs07
rcbdD9Q7ISLuMS4MvJ+H0461gcA96JSwWTvjPCYE78Uq/VSZ3l0IgmQ4r8OGtuv3FC/4ZTbcW9vz
tW+ZgqP2p91x9y3abgIuHsQmTFxhgSxdU2XXiV+7xWhCr4h84hGT4ZTjiukXALM4oh60Fyi7YR1c
/HnwdMNt0tC/xT4vjZxs7cFVhqvZJooKtgwvfYIRVZv5DM2cUW6nNQgenJVtXElmaw6fdayKy4TE
q/vnp34VFAO8GjpO3FofFprQECw5W1jNCwQPOK5CvHzPqlB6tG8U5TuMhUXhfKOlX3gzLRelbdIg
Z/1y3sG5MmwRDKpGVhXOS71UjIpGSCRR+oAzZG6FdxKu9DQElgBa0iLvFr0LgV8ORYCIcNtHS8RD
BENZf2wMmGx0BYy2ykodqfKQCEp//NQDdCZUdYmpEOkAHSZmXBrYSfzkaouJL3KjqIpMhKdsGwti
Q9X4chpQxv/ay5vVcNmUlklvvG8W9m0Y5ZSBdzqJ7xe5CZcQwTYPpxD1Z1CDkdRD1LfmMSpLy+nH
affZNffDc88mrQn3klo01IqHvNEHLYNjCvlOPJ4rPHCkYmlvesXaauo3XaffPOPW8v6UTlFoRouQ
EoHidQwuclVSlcghQvjqQv+zDW1yJiB7P2LzsmA22RgG6PCF/SbYyolk7FnhzMjoJOL9cEMyxpFW
vWRidT/iY2ImrxBMZqxbPQvvTFYSdu5d2SXbeNumSHdGsmQuWAhoKeuYCYYfXNR3qggA83VF8K67
9vWWLPBqrrllW2/kWOiXq9fsIDwD/m/UuXFcnhw6EmXrk2gUt4cgwbGAohocPYZjzIF0GTtfkHEv
Y4MevOUffsy9wbDdwfEN/uIHC/LDGlKzUjY3Kf3Vhv9DWwHKCVAkURfWaJF21A10FXUEzOfeJQSE
A4TuKedGJRRj3VlZ/EelrIAdQFp2GN4uq9KOKPZkZa0tBpnfKuzj0KOQ20pxmFhkFDyVIwZGf33T
X9DLBOxKJBCvPxx4tya6c+LoztldDZkjbJ6tQFSlI0gPBB5185XZflU256mr58q6u6pZXxCiAj25
RqTH4zt3aSpQrIuw1xZytss3GAC/hAEAqfflWM4ynwnZctjpVPihP2iOXOrcivY5OQOyXUqzzTj3
EH4jQ5WbluEz7akxByVDUa9eyeEqLpPUdk5+k9fv4biU67LfxOsa5n/zgEtTpLh1111Q5qgywCeT
BAyP3ICkOTLSTks8iqoP726wF8mGUDTTsRWEyCoaIshe5hF7LGf+vLn1g3DyM0PMTT5tWgYHaD7L
5zWjM6uaaetgsZnU/4mtLYN7izj1MeWADQt/8N+qp38csdDBG27ZQYmrH5utlkKd2GhauAYwr2RU
TdUa5u15qCtYnGJ8Z550O2fmb+wlhYt2GqqR0LhnpZJsI5NhZ6A77qUpjrBuxzk8obXociUEJnHq
uITU1cpkvfhiiN02M4nBosByxVHfvdoUIu+nN7n5OdMfBTUqlpjOSyVlrKRaI7H6o/4tI8GN1L3t
vYGUvj8ZwP+lMZDiwRVVs/2Jntq5O9Ch3P0Z+s0pm3t/JYBu6D8yVRUpHgB8fR2PJu3RtwREm9HB
TBJLD/KHxTemOVHx4esy1dm1M/R30e8gEPN9RMEAORvSDNAOJaApE5LEfNFAHUsVwhnJ7tecQgEK
lk6Cdf2KwXEUwAOKBYTEAejo9VhBQtZ+j+pejmtqk5BPsiaT7t5JRsDPev1f7ZskRBcmmmk4cEe/
lkzKPyQclc6/hka3LMwOJ2oCQUdpxBR6WkN8llqw9qV7DHXyUFD0Z6tfiWhZ0dOr5NIIoH0IdJY9
GxnYIm/bfuT8yQGDfsWP6l9XBAmJTsCfhzXRUByuIgm0c6i5fx55Uhv/SbEYRvFk7m8Vzik+y0sn
SKH4RYq0iQOw10kO/x3TxNp5OCb+9WUhliXAC+MVHCG0nOYhBHxkT9SVjVHRhVY5DHvpKqVIanJh
MeohY95hCSUdf1wwslGWypy+XBZKCMao4Zag486c+Hh7sVuL4Sf5xWAyhuqmscIpd46KMl5GbElP
amRNmut5MZbgz8mtocII6cBskYIHPMVMGYe9QP8dJcLMzolDC086pE7Jpq18g9vr4BcCNFMk9GqZ
P/NubXaCg4jwnGNG9b3f7uVuM2VxmsvyYjAbE/AdcgV9AsAx/syDnI2RWyscFr8pkrutJ5l/ejLL
OnNdoo31OAjmhFXlJjWbES9tGV6xUoR3FpU1b0rSMMuQ1Nrfveu4k10TLpFu8MP5IdXdVUExlAiX
aOOWDasrX1bBki/AU0iowfopFjJY+cxuqUEEUkTXrwDklVuIX3rmUIwYFxK6J0Vm9sESk9m2VUso
q7NOfe6yNiTytqwMJK9AQFwOhrmtjayayASNPeLu1UI5ySPKWiH4EZ58y4tlrMwbwWK2tP8PTE3Y
S5M4dL02YicHLZ1EPATm+IE7DqitIUDRgUf2NScW/TeJccg3XyUrnrj6CY+o7XT/TpvjCnzI4bMF
d87vnWMaxXCag0kJKowyH0Tf5lrY8PRD9m55Lyn+r0d3/UYmKsi1aVxBafIa+jJ/P2cuXTEAL+YN
Hzzx5JXMUGhA9m/Nhu2u1jdE2LW6G5516wgutXyn3T87vwCUF/DOrYCf6rqegVHmc+2BY1QBrDiQ
k1O2oi6MlYRqKp43hGyU/EmjdPLjXvERCUrm2Mj1oJIA4WXV8P/zu7PXIKf+KTruIGUI99nrb2EH
py+NAYrpFU6ZE9QAOAVf+X6DRzx2sXMTJLKGOR65i1GYILe5HBuXg4RiFZVbsWSKQACk7V/QmjCe
ANGG0sE+tpCI1bR+D6MgWuG2JM8BsQ/c568euz3ozfn4i0yR3QgOi5iWeAzGXSthhsuzkupPlreS
ivMX5mKGP29l/NFNO1NBX3q2zR8e3tWSFIMUi4xmstq1dyKx2LapSgnBlxVfiLLreG5Vm9cAvmOW
7ChmjTLT0Tp7BsFTy/+Xp7JjcFygHYwMbhGshDxO6t/lDylGWtuPR5hu+CkMvsJxCfa1h2H92llu
ge7+K/RfmSHeJJ0kHqdWoDAukWa1MP8pIY5esIi9bX7XTPhOVc4AlV3rPuoZ36wRj3wsiumMI6Vk
nAmtkSR8whWdrxXYgjh7Ww8uWobkQJRPFFhZBdHAn1XnWJqY5iRiMlSRSdwmG+M0mf7dqvad9xfA
X5XMPbm/QGOC6k0u9dPcr2MNHJto6QnPLzd0rcFbkuZdzerPbpqFZr/QfcIB4NU7kSsCPUjFqFuQ
WT3b0J+Yxy6BxvPBl2zc2GfoWHHKCUoYmMHCbhNQtaT9uBMZrwJyrM4+uX6oGecLgUDbtz3KXLRZ
8XaFVgWk6W4Wph0a45XgwMtpaWDZhkUMJz3PycuffG/cJg7g3nD/7M89qs0pLiQXTNLOEWrpMnVd
zTtTdl2H0GEUw34URaYzua0L/KKvAyAqj3CVn5HBGxebanSPEvn1ONzQ6yV68X4mlTLAcm0lBYZv
MGsAgvojxzKU0oHrQPpJrR8WJsJxEDWFB3bHTteBjRZ1Tyl7ghABupWa29vfL6SyAOhZ3OIkmNs1
zwOpY+tLxvI6nh6sC8kFcnPzmieDyXANy1Cdfti/LLiK5cMqVRPTTHZP/u4EMDHi8dnJE+nV9K2A
w5c+gFK4h/wJU766RirxDI5JwJ+wkt/PtwN7/TJD5eTxHufbOBf906gYmF98ZxFRqzIGkTcoUYcm
yq0szOsvpo7dAPJJfXZO1wJrCSITSm+PftRU3Qh6t9w0XNl42Lo1LSRJZ4LdLe12sNO0HfXJbNVx
ykgRVnW+4N5+VfOnfKOph1BJvpS9BXzd+Ki+BLWw6D3mP+qPGpBC7Izz5empkJ4qqj1iW7pErokj
fBXz7bCP50oTJs6NI2bnK/Q+jiy87GzEiLfApL/Wfc9KJAUPKGu9EdUgEaoqLmuZM4k6WYuulzB4
KCtma+zlgYCeWIKoC5k/uTq6zCvvDxqMdA42VTcoXK8wPMmNyCYC8gSNRfWkYPXnUabwGTZvlM4t
W24XARg+YGnKq6Je544/ZZ02RGJUFFFwDzgoVKDobbedteFbxltc4nlCyroQrhRtdNnbVbgSrH4m
9V9AqEXlyTSH7N8mM5MnujRwP4sJdCxziDwanmKnC8Se/p/dX2s11n2KFw8HNm2xzzydeprEhXSq
hi8tKu/mdzBC1OIJd28su3hL1E0OnljiJx8PgOQJSV9huiiOykS1y7CbyMQ8eZG4nLTKeAP3z8+e
PmU3wbbotWXO5+NHLPjpjIiKYMzNpt7skm01WcqX4Sutd4CkzFoFiD9ks5GNSXYnbUSayZzl74Pa
1opnaensE4h12xLqsc+2oUaHZaHmXIaNNNSIQnGjfXV2SRrsmGd8aejSfDZeJkDEjoSASIGuTeZu
TNVTDjV1diqSsg0ghc7Ma/Y3qGRIOSbat3nAaM1NRpKvn4hkHs2FpjcmNXVHaQQ1K5BvqNtAe2Rz
uFHo1XV/6Om6Q3QsaNP85EhmEOyN27TrXyX5SlF+wCorj/IrWwNJu98ibsV68LG+5K142HJZ9m0Q
D+vn+4D8AH1u8Pz7oeWPrYhmIV3ycsfF2XaKaVbr8rnD6ugkUT+re12464Fg7D9vTEUj6dIRqjBK
bwgJjU7ST1I1ShlRd9nPgUtT1aZWsltySyTxyYd9pK5QrsuKBL0ao2vhlcK9Ux9zi/KFidOLjHQN
8rh7m6Le/mbbomeMy9tgWlyZFLwv8zm4aMIjm/COHtZ+sk54BkZgucqJJ3fHTfWQM6jy8uKFLEum
FieDoM8Uv17DABHPcFTVvLmF8nLteeNbZaOTbxgj47sUtvjCpp7OVntkp/OgF2Tu7u7M2QXg7kOB
nr5AgWwWTpkqycDVRT/ABlPtBmyqsTR2ocRa/nCCsProT6cyIijOkBVQcRbs8Wdl1i0ztE61CGu/
3dmpdgq1xPiHnygHZ8j9OHlHJcEsqosB6Lb+vPK6+vUtKcmoS7lEgE8pfG4yOGJIokBmkAGy2VYp
s8cvXZfdnK5aNrK+5Qw8pfmJvqj1wFMRdqGcfWrrVXAOsXZN815hxa17IMCf9+h7kgl4WM083j2f
wIV4+UjyCKJ6kShQlzsg+TLtbNIqLF6RkzE2GLXuqkAAKaaRWdRMieNbozOKIo3byZXLEygaI92Y
z6QhBCikX530X9Yk6HeRbVT1UCEngfZWhx7MEHw3H1bvEvbh2mgzR8suC7TbQSkBRBkQm8ut1yqZ
xIEjZLSZETjl478qP7mueJtvCVjYYHsglC2nTht918/l98GqfAwhpVssWDBydxijApAe91mjVi/Q
AlwxthE6vdJ4hSRmFYotpOZEQnVhqhZm4F7PSj7IeXqvSB05PShiaSFP2iqyxHapmLo7R7CyedWW
Rs99G2bqtlZYgqrsSeyee1c/uZiDR2UHWSToRMnGgh/+gBKhZt5BKocTrn/PzdM/VDDsQvP3E7aG
0a73K+reBmct7dasMWSuWYnwnabA+bKEaeHAD4dZEmH6Zb48Q1lu5k4m0fXjJ/frJiWU6AWVwhqX
lNRqIDzcUtmLEtsIXfYElvu5UrmSM4COFyt0aYMoK/86FCta60TyMNZX8UZIfFqt9gg/GjpNnRqF
0n69uChdqyYRUZKdEKq97PA31EL2jGKTjsL4YR9VGPDcBWq6vF4RAS0FCjhzWiUW+tfTnuOc12G1
A0qpb6iJuOSz9SrorSvoow04EcYVFXXM/jU90gaOzdu42M3dxA2dl+HR9HaWI/NPKSJPB65nO0uy
H3qeeyd3C/YbQT3hdkpQ9NaThiwPELtZc1GbOWIuzn1MB0ur8DZvw+VPCgghYI/cGP2M72+wIKzd
XgCIjh99ovJZ1b3CWROgSsNjSg2WtmNnjnVhuMEo9S0F60IJJ19oxtajF5Fx3X2/lT1dikyy3eT9
2obaoJSd3n7WeLI/eIZbm5p/3kHRwsIXY0hI153mlSv5FEHoKWhTTLmfxPcHuwSkAgBVR8nq7Z2K
pnFm0DtR6Gg+nO387RECVyG05B5Sjvu7drGBk1TO6+Mfhe5s7w97Ohbex0hadHj+8ER/YhG5CTY3
i0VF/umlhJQ/fNJmJArYeOpAf1ELBwpkvHhXhF9UJ2RNTMNlqM6e0ailfdL4jeZMXLkBXRmNUYQV
fFrl1i5tXtfA/PhKWIV+zgjKIB04Vkbq9jdWiuRLqD+ftGzO0ZkcB20maEnSkuZWdAaIj0/v4dMH
blaIYudr9ZeeeYITIKFidMwYcnNaEjx8QdpbCvNxmBzBVvGB+BGCraskWwq+ga3D1cBPdHhtLgAK
JRlCGA5CyXM/KxiwH3JWnypPe9/CMndavOvzx8AXbamP23d/bx1I+6poRda7OFQCDn2p2MFm00SC
0GBCoaHiIoM1jvkwkSM7jPxqq9qOgiFn8Hc0Q0c3EiACMbjAAMXRZ3a/eoAr/SSuaTa9sQ9tfVbX
Qf19SvbrJGcVUVfJZQHP08/Ew8nImreWXc6S1UvfWQ/DJCu6E8GlmsMHas3tdqLw/fsag+tsVvcR
d/oDCXwDNi6tvBsELv/YBzxj/rPyeoidZQphw8oNiEgzyITbMXTjTs5TYMjLoGRv1zJKhX5bKvHL
x1Jw4CtCVhglqMR9/odk3LlAeFNXA21BQECScfuyQhA9EKsXDzkbv7THNOtfInnXTMavtUohr1/Q
RqrHjPUt/rI829EIKZ66U93RmflYnc+uG8T+BZuzzSSCJ7v1LInw+D70zuteCfhZCfqHjDXNBh3q
M1f31b1jP9HOgbyY/L+bkLyZEsbECyuX1eN08sZXhfUkXtYWjLnTDS/Kgz8UJvGsE8XsBNXg2eHZ
pIVWQ1hKfkmyX7IMera+mosI3vKDhrlPeTDH9DQ07MewN3SgF77lu+m2ReTOyny9TqqU/RCMV34l
biEBZayWMOjfdV5EpI6D1PratioxRGk5XioIW0vPYX+Nt3Dcz59O+oHA9QBXyo2KAZCQoPvbuCnz
5FNIncCIToCoSGZndMNX7Foy9Fv6pez9Et6nuf96Sm1h5xopSaB/AggKjvP0EneVGi2QSIjLTnOb
kFh0ZMkstHEG+khWOh5e+7DaOVLdu6x2jwQ2K3I3AMG802F7YEnxLzLTb0v93dCl2pf7tJ8K7plS
zDCr0UAqpdjrcxf5enD2tn296vYfT3kLuHclbtggMDar5LX+Oj87ULobkuqZ8R7SXsMw9q3bWjLG
I68kJzdfNilIYa3+YI4xMGU02oo3nAR5lh0DQKVVvvDYFmUMwpQAMdIHA5HtyzHSOHk8pYTgujcM
ZsoRVd18PeP+9+W9KepJt+QK8DBeNl+gOy74UIgFP5MYoLAEGxizfCCQTJmE4D4Ht99Jqej/UxRn
tn5i7twAFnH42TBefozDrlVqEpx4Kjl+ZkU2hafAfxyPmqZm0Jhix+8ryIIj5V529kqlplRu06tD
tqupqxwUhiq+pP5xNE2L74QUA4x1c7Kyzuwjv40G2yOBtHNDJzcSfzCAa/lDJu0opTFi8VuNMGU4
wghKDmMJgbu3Yxp147vsTWNNmtYUqEa7BQKZbjLHSCjNf+GTkNz9NeVAvQcxPga6vz5lFYLqWsVc
MkdVpWjYnjYw84rkv/S9sMLYWaNHP2qTJJoiS0cmAeKiPh4StcPwrhIVDGwK4EwvoUjCJ86B48O5
PrRQNSN42Dn7n1SpgvqtNwRTlNqsSs8yVQxaRmxuPXko/OeI+CKJjwUMQesQDligaeu8t/d2Wjb1
k8yUrINsEb9Dt3Ka5P/uidnCQ2q6xUc59IkFnW5abPEVNpZteHkyTaGdV1vpvZ7HPxiD3UYOb/BW
lP9TNPYYlej1MBrdRtYiq5x/744SjKAkLUbKMml2ZUhWTnH8juEaHUXBYXKQjQnIngBuqT02Bb/D
D+c9fMWTzoTsuq1MBYfJHIHh3zBjPWK9GYwRzidlnkP0+inMYeFkeu+gMp84Dl0LF3CXDoitu6vv
VQaVqcs6bcp15ZAF4oAa6r4bMYESkc0oQcxUSo+nCvZf/DnmIpX8x4LFalBEPqHD6e3Vi0bvmP/s
XMTlcI/cWq8IFqkkAQBmrN2jRuDHCFA2und+QcXTyx6gai4gqU+/2r5J594sMGRn9VqsugiIwxJM
DP3BHmhqeMXW3Ynr9wkSW0Ip+NAMmOguXInbOuuZ4XNiTA4fjJxZnNIjJ9vPk5VD7FHLc6NeitpK
GrcLArRDy5F7rNzwj+jow7IsZLJ8gpbkZHD/NptH5W1y48sMDqB+mKPapvZ2z006idqTCX80YoC2
wI/fBj1DhwYYryTl9Yr0rqBoM8I1AHKaiZJLTQ9WtRRM+pJilD8j34bPX3mRSFDob0nlRtEVe9rF
OV2roT94cGLU+NFq6lIZ7sozYL6hltLbIRLzS2QHzqrwNCalG0t+Y1kgzP/QBcPBjDe3dGoagqcx
yPaDK/wQMjkMgr19kKr05GO6k03rdTeALkMvkTjHysS0MNCcZcePouwZdJWkvcxu9Qk+ntZG+Pij
ajnyY+5M2LsuxS3Cgek8ksII0P66bExLynj5BNta5ZE+GnuF1BM96q8KeLlIapJ7ookuumQhPvsi
/rQ7alQPdvpOo4KiebgUebiIX2DGdd2TQc/RGg0zqSK+3FcflCPd3L6JJATwfHQXjwlmx7exjX3S
5+yuzAV452GXbk581fKUWKVxm1PjNKtX5eMconeoqYWQnURp+oHw+GpHJNUE/qUaUPkMbIDv6hlM
BvBjXH/7b/TBKhHZeM3ISEiSNcDpD9eSV/PkGxLCRGQkCli0WjKcHhO34wvhtzG+DM+1WJ//T7a1
v4fL+0nqOURaIbYfP/LWjxTK28xeb647W+HzXR/LwTiV6KRSEX6d4rrR3qs9oENAFUFO9M6N7xZD
YwVlmBsKAkCsRPqRh7yOaoOCVM9o6AVGaYWnjNJc90uYiSzft9RlafrMzvIhR5FTV2Z/9C8EpPw1
RW8OofJtTfaJ/REO5PH2mV0Dd0Zzw45r1PeyFieED7BBZnUb1ckCrKLDl5Sgod00L7jpWCYEqndK
wvbnPOmrDAgchia3SkxTPlQyYo/pXSc7YqDudu4+bV2CfkjwYPb+aTTOtIXw0hlUo51HNmC0zMxO
jsdTqcqGytyZGElAhWPf5DjXN8/ZgjqVsLhvRcsro0oEiYiKJ6aXg2lY0Vo+8mKcSz9IKIEhE6rY
dNP2TlqOtyF6MCG5Ouqif5oqbskHbQjV3R03gOr6MjpGS69ABwx1Y+usFbXLaSYPX5dlBSYZTYsj
RXjupdJIkGIGvzVrpWis6yQjnHGjXeP6nrhbSOG0ZEEMoN/WuJJUt9V36VUsvmHNNFkxNZCWUOGp
1HFKEA4SD6IYvTOMMHsFBDWLvCnvRkge6867JRxTwBA4IPS18GpOalff8UY1sQzklUQMvWJoxqWI
GmXk3EEcum+EHbkWjDhCXu3DRzeaPMLBDUOSmGCXVLxtERUfx3N2Iip5FyqBcPD7kMww1fe1kTVZ
oSzefESaxpMk+8Ps+eknTeHItZAxEn+igDw9KNlATO9gQxGR/IisvUkCD1uZICCQWElWuIttrufZ
hlM7vjI3BjfGKJGBxtfv2Kyszb6LcFfn7jNTX8tK2BlJ0PoP2ryClhKxDQtF6ZMbcuLZZxD9xyKr
rGsmu3UPwnAoLr3nEFYIrtCfDPR1d7VleXSeQd6rkOsr/N49ZRZm4dawA2xKPjTjPad5D5zTZ5DX
n1I2pFIlRPknZEuSnF9CyaVBHPjqyNcaKnoSIEo+RKDHer1ozwT4nSiVwIjTF37U7Rdx4r91Xq3u
H7wD/jz4g3MWPeK0sql2BeyUbZjjQHZunrf6mrSIXg2qQWwojLOnxbYvhA9c75PxtbhZCoa5NEqr
5JSChTNyohXBTGoBfRRe9AClb2wZPFi3stPwIMn0aLywGQPqxtFzdMxU9ZlesjF8ZDeR2hjlwBZx
vrnHCoQNlpjLY63rufssxxjwxwjRfCfQKo1rvqoEIzH+VsrcdMIdp+MRkMk24qnb6A0sVSJhFbvs
W0cOerXXVX9PnYOdEhxAR/YocL+EV8KOJbF8GqO4eB9z+m0uc2vvlSuYOuNC5NVq7uC+zwxn1BWV
5r1OuHTZ2IzRfDCpYuzsa5AMzJVh9OMpy20MMIIVoPeNt6TxSvvHuZflWrVENp/Ke8k6q6UWJPCv
RFASQ/ZU8x47lSPhzGjBcB9PBCTzm2yCveoELNc2I87Xi0LJ91sQwGkLJTW1RekZfF6sSfqsQjx6
UwGj4IiHCb0l2XrW4y4tOkk85CpsFgpw13v2VAX4pdHQds5zNDdNiD3LxBPmjLE3Rblc8fOPCLwK
MfSJLxc82c0IRK+aNWMdN4sHoSDg+PpMzabAmCBnT8CmevFWEDv849m5XkZGSHTC/jIGrwMeStCe
BbKKRo7FVCZsHs0RiK+k28oopJPRcJmMUvjGB3rcsYPjh7t6e9X/DbOHSf/0CDM4ZxC4nx3iMR/B
DrzgGlhHO5CGwmtUrksPW87kOskDkYXakYdL1WyDCIV7nBgYEQSvLOLp/PtIvG8KryR3UtYvVZL7
EmmlY6bsXhSdpL63XgbA/X3U5jODuVVa15MK+SuKFSmQmm18q6hZ3erE+a9u7jusASnW2YWORynN
1iLPCVPW7ovWjV+6dOba+Vsykwbcn+/J8/l6WUogg7lbm8NgPNykT9EXIO9wrE/PnSnI9SCIQhcd
yvQ0ir5F+PsDTc+0EJVeE6sSgCdqQTXCpemjja8Gx4NntHgLJHXyAtGOevD4KA6Zd1Y25mTi+bnB
r01OYD2GnLl2334bOKeZkMkBajq8UziWSofcIJbRt/IMgSTZwjl1PyLQT8ClacA0CHwzrYyYdXoS
vgaNXvt6oC7WM3gagysYsEfW0+H9LUs3rqSiI4aIJXSo1v0bY0t8zjePwwEUlVSsEkMVr4SZf4Fr
5corB7/zhQWut5q7Ulab4rzhHJHF38O5O/hqYCMZkgSIjTDdtrAOmPF2YPfvTswhhztKCvByG/DA
nB5ztgwixQZJ4MtMUML4uvJwdZ4Lo8P2nVsvtXtKkulyRKE3LyAMRRAR95JtboyYxl1xTALZox1h
BoZMXZB4X+gq27Y2DVUpzx2qmkvEgKYgc/SBZjiIROhYc9ySR4PbRIkIiMd3jBHnyJE6qk6ITthN
1kOQnpH0yGE8tB02oKlU5/i9c/3aFw1Unq9tAmh/vfmvuIcnvGGq3eKCJeCj5tOy0356//eqHZ4j
NV9eIHd/IqLKqr0i7RyVzyqezZE5HBQcESyJg0q26rBaebOnTJAOwXDzi8k/A1EKgcnmeejlb6do
xoypq+ty/NfUF4ZgoXLzT96Q5Am/PhEygsNw/1ghTd38UGKISNcDvoEoDoUmoTaa51wDdKmZXS3R
LoUrCIx4BaB+mgLTbuob78brnW2ZiuWDAnQS2z6HLOgXoz3bOjaMbp9mNSOkLIXYD9t1GldsghnS
39w+vwuhFeeozxBCF0BiHzubw5eWfnMWniwEorBk5caecc+6h8/N46oBrMWFsNJcIUllL6Pbt+kY
jyju3Ypmzq1ovMFF9pHgJ8levktXlQxR6FCzUx9XwbpV6FmzirD6ZWqce+MJb3j6N9bKFoVlnbfz
x+2QYtlJ62i72IGACfwvOAr/xoktWBaVZ9NSSFeC8OgAlSebY7SNy5z4iAbDr+yopgpN/NUHNNWT
jbhltI5DxROKMG2K6ZSWeLqYSR4ORBNqjEz5uWKP755fjVMn/4USGJqird3DfoB7G1MnB5aRyiiq
sHP4xKApYsZ37uNf8pGhuhUegIP8/zAX6citC2hzfazpB7XoYxBtUhLidR6tv74TM402naoREF2q
slE3+ZAvsnY5LPfEhx7Xzi5YJKnNkCp0apHEnPDzt13jg+h+/u4Q8yOYweRY86n1JdcLkxfdC+K5
RLdYi3oH0+drVGkHb1OsLIiMwetJ+io87hIlBYxWIoLeKVBuNS3gzAzixqeviKh5F5qNfJJxkt+s
OqSsNnBIL2i16eTOlxtEWWL3/3c2zyVZaKaCWxONw+gAltRxofnq4+AVQpdHwqZhsobsLy/mvoJe
A/409NyqsgZNRz3YHkF+kfpBGTx7JbB76HqbdE2Rds1BOEQy2NWbcfFnUVmq01yxZcYrtjeNx0xo
iH6iOnCrvuHYXdM42Mg+SRNmm+8IO5b8xdM/GsLzIpCSYYOGskKBO8bDsmp4khPS7pdLXlz839KC
d3jkBY5w4QIE3dIbP3iyImjyU40cO4cgDCXSr0KpZuUFYb3DMdG1NFrBVADnUTEz964HOhm0okzU
PqTckbrrlqdh1NQ9GIUoaBC9qzcNwl3woEsDxvMSdrvAmWPUFeL9NEHXFNdjLFbPgLuudYBXUI4f
1D4a5kOWaxO50/H2rXIWvbOvKUVQNv+iJNhsn8/m9NbcWxSyXB8ttdqREFVstCAi3cNzqhFKj5WB
TVZlK/UU5EThnqqDoGsXd+ktr2Hhce73xAaepi9LMDjbA8Cy7N8tpUl1QCYlgw7+lzShYJaN8OOc
5v+VWe/W4bMgRIBLK5ry9F6LxebJPNqgZ5x0RDDj0DnBsSO8S5xT2Bc6KOqhcFrN5SRJ0yn+EzXc
+uYNvqWtYvjAD7t7ukBauPnYRb0vfh3X00NA2sLjxD5GoJhbBnMXJErRqfSbFi/z4wMMtGZ38tvX
7EmrceUuT+abIQtF/tsqXHGFsQPMwzZXTCUMUZH44Qtqy+Vh34vmFUSLoOqeE1sm2xBcr2iZOJac
TsIrAtyxThYRV6dCmyjwc1v7oITZ1HvuMBEJeuwzH+HtXCyCKmRAVgD5NoQcM2ypfE6DVTSF35/+
o74Gw/2vMvg5qQWIOAf1gexhr+o8p/Ypr+fFUJHK6D5UwycTPn8ATPA4cbuTh4u3pZCPndsdvpaj
Q6sJgLSfPt/jGwqh/csFPtrcubn5Su2txTDxjGLIeLYMvcOsr+qdPMCW6IDa5rdeO4kwE1B7yevw
NuZOBmKtsD9i4JlkY+18Jlam+oLubAVNrlxbXNRrqcZP1Aw+qj0F1wcauv7Hsy6YQmoghSroF3Em
CxSEzUjkvs6tdMjYm5fABjaAYKwvcek77tupUW5hA1zaj9snG4G6DxCa8AxLXhaGN8YmaPk/foSq
P6/rcInWEPz/z1Y3zNUXlobNRridvwadJtPTmoqfHfOS6wX0vws1WvbSl2wdRWcm+gwxkr4LABVE
NEOnQcK/EHUrD40uDPaRT4SVKc3fMv+HYmnoCcifvlpPuzqog+f9Qjz2s/R7gz9YnoNp9xoVry4f
egC3cUyMG50L8n7/ZFPNtSZt4ko3Z68hSbk0381a48HfB82Qq3QFh8ODUQ+FaMm1B1Li4CPpEH/A
Chinxa3+8tCMB4nSxP8WzSBpMdH2iCI00q6Kj6lbuDQozCjNQKWje+5J25hFOzUMINQ8dkNWAxCL
LtvtNJ523bNfDj0Y0vdfYyJOe+3mCNz7s42kiy1RIc2VPyBMk/RnovqItOpLzLiDn/Rwtdh9QscF
zLHshEaPTNdGcxUMTNp1prTFo/IkiofBoXCHjsgtPVdKS7yJmnfzUR7sEsbTQj4pKqbVONoseqGZ
ex9MuDdlrah8FFD71z/+VtKdXssMNiIL/W4pG5aL4wtoOmjgrJihFjW4aaQExdePFy8xr9zEx4wg
x4KzPqCbuGCrYyapzWskBS3iRHHim8wCKYT0zLWPxseC9+jx6yVGjEZnndOSQwplWBoG4u7EcJVT
qDrjryM4B9jPmCIcDoEqNbmcjhRWWaZrcq4t/eUkj4vjwW8Nij/7VlC1RmxPVPi5mQu1oB0dSyYw
kp00u7qU/feJbya4RQkGi90OlLZ0bsmHZWl3zWs58NCx2FsXgGhCVYYxPmS+RYpTX82o6cqHWtlG
/BkeLX5gbwsZO/OMJsiBYyHhnMpXEkoNu3Jx3TQhFzkgC7hJxqwYD+dj82gPkwb0X1JyH3e0nY/S
wSTBe6bjTv0WMM7AHF6eQqdWOsGa+OZGBV/sudNu2Qdyal8W//MGiI/uYfILD0suy7k1tcjl08W3
iCEI685MlUsrBw7aMQcanJalT2dgwSHuCDSrP5Z7KuVPR4NQxoT0Ml3cgU1zylbPzKTWv6qDaDbY
ZgsJNzWx5gs1pMxzWmGUX3CzLrVs1U3Gc17NXHPz4b7l5v+bTusJI7a4bvDlUp35tXh+67mwS09a
f3PPKkpfvwox8YuFib3Z9n4uJlE98Q6f7AB+1OKLdZ72tMzDiax5ZrifjaRBIHdYF2pHQ7MaZnzX
GivSso7O5QXAjIeUJwhA2ilr6wJypO4OQfmAXQh583XcGv/gu7G77nFWeohZEpHauzO1TR0+Y2ak
Zhw7PJlUxX6ObsRESnGJYrQlYjM2peFM+YeK3pCQMak/9B1IB5N8lFeCxCPPDHxYcLbWdI9WOroF
5IHdqvKipErK+kSuTLHZD5rRvtTg46adPJnp4msXjrOLniq2BieS+S0I+UKTGGW13QV/MTaAwW9U
mxaYwazqK2jzPvtF29YczhMAPzF/ou6pN+Q3ehMfh+eLCV2lkzP9praZlBYjN5tpyf548g2DVThx
xYu3NbwUdyQYy4+u3u/MSFDUU9XoDfAlQAHfZmMe9g6ph+q2LUtCMtjGYvUKFhvKPW0ByRB2MSDW
s3PM8aOd9gfUks9XAFobWUMD6aTVwe9w+upmarmrr7vij1OS4L25F73laRICqbbPDMrkXge0EVrZ
dGOXFJFSQl7gaYKQ7Se3PFNBizABhmJJrZ4A4GDtmCIuBq99FF8qk+PPob5833YgLaiGaJarSQBv
vXE85K80Hl9Hy7dpWKqEfLohfGOqPuJLabl/lv4co6RQq+biJk7lzvp7McZtV4rTQoCJOVDw/sQd
hJlK0WVDyJMkc4yuhsk2BmANIjG91GeFcVcsV8V63kvBmLfoX6GFD78w+po1Q5VXu3Xy0GXcpyDr
kFF4A26bJMHq2TANGr4gB3EzoDzEYLZ99+2GII0v3CDoQp/NPAWySz2Ukj0S4DX1Ds6/RKxbdIpq
f6/ETWRFkw+tzqm0+ml8XygMubBLTIF3LfaJN6x2wbu9PEBNKtUXh4TBYfmtnNt8oX2TGxWI+jGP
1Xs870rKCHxrW10dCYKlNa/DCmblJ5S4Am0O7lQDov+tsZ6vPJFmQg58v7Shpuu6LrCV7SsqOZFh
UYrXIWpANvIeUyZ/4lQQaCDc9jisSRnZ18zFJyRaJ8P9ln9Kiu3ArIYQVdmXhGFtKAAhts0N+uGg
uzGjbczCX6BLfziuKo4LxZ/6R0dLWb1LlfcX3uQQtWTvETtKmn9R1mVHxT49WaBoJjebLpPN3cbw
IEw3wwpkcvIBhOxAI048CXnLFrICenUrQdnR2RgPbg5H2RA/8XbrX6MWEsPNBgPglQQ+X6+bAObV
1qar1hQrPwkdTPgmpH4kT+c+86NRI0x9hxilMoR+ZE4nsL+tbFkTdGaEA5wGRR5+t3MrEJ2RlzDv
zri5pxXQo/SamRu9tSiGzRpYooTATNn7ZBX4E1ZmbVluSX1VRbrwsGD5RLINlcEAMKC3JjB5lwyh
tatb3bUSMmEXmPdiEYjmX97l1FPGUsMPRzexhe5V72F2eJCmoK3VoJh6+dtlOZ1k7iNhG17TrMHs
Wh92l8fn7rOda3PilDBL1BMs+gTowfYqmGN0AQF0tM4ynupeMkyurCQeDGqnBMTVIiwtItNTXMll
TTVtYh5WDoWnEOX+dWi0q9ZAthPMsxlxjho3iKdSw2SA3InP4OeVYMQmBJcMOEJMXIRDOXd/wBY8
Ae/Cg74Mll7seP7UWLwfbmeaCTzDtvcxAAJsBy9fT+zApLxa087wa65wGr74kyWqtw6qNNCmAnCF
S7cg6DrkvJHeXndzHlgnNFTjiEsq9iwSnv6SjkrqlSOkmVZ25IkXOWPBPYwkLPD0+opkA3Awf6Ia
izzIXpi70iKLVzVxwX99ERS0PZMCP/5iL0mUUdn9E74O+50iwtLKzX5iI4WLYFgg6fYF+9Cqcgdh
eGnPUokCCt6gqO+0QjiIW7qz+sUB6h+Y18EfH9xUAttr45LiEoHjJ28O4dIF10TeLGAvDbAySM5v
96iqqqV3qaP50u6gPFgOCg5LxpIIM3l3kqzxhbVKyWwNZ8L0r37yYJSjZfkw6L9/cX/heMtQGcji
QaP5qQUqQULok+k4usFYnz5WJdq/C4m7uSvmN4oB1CvSX25pzTcUIdJ3ZefGETn/+ekdVzNR6tGo
mEm2SVCDd23a1LryGf2c/Cs8aiofCLMzexaVKB03GQPVRWqMPhZT7jQUJZntlweRYUEUKrCglKT2
LfIfbFyS2zkoD6/LSMBGG9NDFKfk/R7wTTmiI3d+/Fw0v5y7sNOeC3uPpOQ6RZTAGF2dmItGdarR
lfDyvtr91wufXhjmNoE9/v5cRxqMtCtZb7G6TR2FR2cgVI00boAWjizSpLNqb9iPbdPHu+gwMKo3
LRAZwrEBZ5+5SU/Z/a0MJo4OM8wcKG9ycr8wpKFUCwj/EToQQUKz4yI7YkIdnZRTMOBPuyFN+7fi
WEsAil6MoNC6v9BlPyDmwrIGlsL3WQfA1y8GftxMC1vuArkd48LyPBA+aEO1/pMCP5jWk6Eyv8dW
bcaPwMZQr7QJa/PSkZarGaMqAQyuVkHvKCVbjyKZhnz3rwtb/6cPZ6dG9u2Oba+x/6ZI2F4mwRuO
XH8VYpA7dvF0Cphk0Xf/QRtlL4zxdmlivZ6e+PG06UEfuVIu5YFcDFnsUoZ93nnsEhqxM2EvYSkr
0ISgz5C/n9kPMV9tmId4LZ8EAEDZJ8orVQk5wdbkXWtD4n+zQ7w7AkA8ozwgpupZrv3CCteJL/H5
5YZMkvWCtDRVLoMtOfqZZRa8rm+sqdR5la/60La3Lb52R6QYkWg/4v0nyGleHKvxewV7MpqArT8B
9tkQ6Xf49Jca4ncxRfvkT+ylCC1dNtjBaxtqEXMUNJ8URMhXw5vnoJ26wfW6KKAlr+GK+zsvUNGa
pajM0VQSpG/au5ArgjLVcDiy2s/GC5IKrzDBZAa7SztnfPFYL2zTW8D94+SClltdDz1k2vKtPE3C
B5b9/4nZQGCynr99FrRvbtDzX8cCySFhLTsB+Jzs8ZgYmzVPXdRcONH9u7H8hbfv3jvtKhz26CeB
8mRLKtTfv2f+K8hRYjNKI2dhYsTpnGBcGK/JB/tk2bbnwGNdjkAEGoGuTwRwpWzhzE4IDWZMUKJc
7Ayec3696ZiDfvRuN1oCPtsVPGMBuUwTuDDJXCg2wDeAUcJw8znKE2qPv5TWPe1UIMihsu+3vWng
EiEhz1qF3qeTbQ3PM88aOAAhfpzi3I15qr1yM2jfxw3JRAHD+bn7Ag8kJCpj4e9Krmkl3nxrii7K
5hM9A3VggynBmVav1KOd/cdlCnIIQZee1NLwgI1SZRAOofT5MYocFaWwL7yWMGkQzmKnXeZxYwGF
mUyiCLFkr1MuqCS+mv3y/MVKqtVxq/yx8RLOGoYBAxVWSB2aoUYpS8/e2ZGpBtwPhw1ighcjJDYP
mnlL+ffvwUL7pYBBoJXVbC3SY2pk9D4jdLGmHJ10QWr70ExV2wGj4lGwr7pIGm8dAg8bqBFZSlHf
XiT+aHOdFfmDCfZ6G3GYRzeo0FMMmLf6/0r2+1+buo96JHHn4IC+HdyDSaMG3Hu3AGP1Yx0kvsX8
9QCgByjzMy4JKxt73x59KJZoLp3kD+AVnOJv9Su80sIRyFV+VU6YSO640mGM6NJ9Eami9aXe3vhs
G7guL3X9gZ37krSnHGNRjRw6bAjpjlUcAuLJWu/x+vZorg2BMiV6qOF+LBWCAn/lip7wzG6n7PBr
ofEB4OlGHLlKeX1m9iMtGOwE8/9/rxNF8ADt0i8Ufc83h849AetJCB9+twyqcZY8BEmz7iBcaPEk
78ldYd8wTPX4HfSdm5eHBz0LK8ALjvksx1Q+J/2bp1VyVJHsdegWexhLmLUQM7tcha9NYVSCawDt
pC9Q8bH8z7k+Z15uxqn0Ht277HyapfgPJb3W0qKmej+XljoT+voJJnsLkpircZLM0Pfzj3JtpGWn
Nuh+Gp46p/jlHFbxq2ujefQOnaR1Gnamp/ljE+qP2Zj4qdxpqH/z5ZebY3MW4dSnpMdyHLvxowqA
PecrcmIxrGIvTrOaQI/5djZmnqak7znoinFcQkr+WUnEjxaxH/zC6mDXKWNNwSNIAS9iSenz8dVv
2xTna7tOW9jz7gvY2RkUhpT+gK7rPPOrPwR92boPkrUMawEfCuG6axL9TxwKVngmNWhXWFZabUT/
AiX9FHE60HnUBg3hgDqFnCS4o15lRZyz8/OkdlxutFpvd/SHGAmf/UBDD18vuathXGgtox56Z1H9
CUmJ1pE9YT+6IODTtsUl3sRGEAEbT85rCP6Vo+E2PSO/HGSMaVOaqUwA05xtZ6agWRWYHzTdO54P
eP4NadphmN1/9rSMkmz0HQsoLmuu2h+3i8f+sFpmm3AGheDXMC6cOXygoH6JS68ulxBzh70fOy06
j8PvXhtX5ADiNdtBemrD36EUoYKlBDEE18tPR89eiy4b7eLMPA7x2hEfk356doEnT6nnfol55ooC
vVtEw8CeD4DeJTDdwnMRmH3QwZHRolK523QM2y873cS1jNFqb55SP0OpcY9x00YuJ1v3IhEiPpw1
pMzF5EHElZPhXWTxQutkyf30744HB4pHTvSweHlem15OSbQa3lovkrIKSEwlsWihTYp1v9n6pDhc
uHUrzLbysjQDkmseFirlqnB5yDdaS6XBIoe0zgzePEgL4/KvP13ktf3Pl40EoRIv86T1R0diSlqh
NwXBWZoFPQXUI9206MWoPkvwYPkjZwUDGdSNj70zYe8dnRSDkOV0bUJa8f1y2dugRpbPocm+17L3
aIZWCr1WjZokKvekdS5UxNxCeaRTD3qLX+wI3j81+vI2jQ4gjZLlUjgDRuoJbG8E9XVl2ptqytIo
ZPjQdAsN+S+55tbKLB8stPVJg5Sy5ebfYjWLBCZ3B6hJ2DOl0xpZVack4l2G9E9GRAvAneWO5oTY
5a8qtYwmwpDmJuqLlaOJYY3rA9iUGxr4eeMYqL+Q5ZId/4yLRWiSqnzGxpeG60BNCzdLhvktFFhi
/Cg5Vmc9pp7MqaAWQVPx101OBTslumux/xqXJcgRzt6mxpaCz5JDUaC+WNhGAzv9EJrgn9VgTMr/
ly+BGHzaE3TldQogXis6VSOCPYZDTYBvgOrQ8mX+sc0PXjlFTj8Hnzlm6AQ8zwO05tD9tYc7Cd2B
NPrv1UdodkJdw1UN8omUCNiBuGSZio88C+pZLSbVo7YcPPSbSnwt4CB9WJmOxeOvmsyNBgWQgdp4
cUsh+2XhyJnC8DaEY6l2BPCAbHKsAcsMwR62DDNCj1ZshvHrZ/Pb776bw5gwyQLv5oe8Ti6YM39z
ZtWmS9EX7WVRRagrl7dc0wlUOLHvkPC8vURDphHCdETxhRs0GjO1TMfBJ59TIZ/LmuClXtKGXyk3
jPmi89WKJ0H5uwdZChf+6mygZEpWfVBpPZKfrjTEa6CltuXvUwYMC8rxzfmxjr3kxu/s4xSZOYCT
+Flf9kFqPU97z8JW6maMZ2dOEdRUElec5UPzZmMlBZ0rYhBNlD+fIN/W2RjHHPQTsyijiVRG+Fzx
+YUBQbxRPYezSE0t8ZhGyJI4BzX7pmlnh3zynUjdtI2Bl32hZZ5c4W6js5eISggBn0oFozPaWio6
u9tfJc1S5SssKuq/p+kB9/XZCI/tcTsVEbpV72BCN/PSWuUpMcmC0LQuoYLYeabTx7rpoUB6sEXP
Hee4Zj8aaAMF3PX6/DxjS/mcoP3U+wOqwvZBgWyn7gJ813w0iN9UqLVHXbP84wzSPCps3KIAISpS
TJFX6+h2ygxf7J+/8tkAe6u24FL4AWXinPt0W1WYY02VFn73ckuT1nZbDKcFbx+cPO+SHZbmUUFm
ooZ5jSTsbNAkLaWfUMoAGKYTwj9QM7iSiUSEnqQD0Lmgd0HDnTZCqKzWsQQIQQCxa91cu0rcTJs0
es/t4ZYtFtMd41JL221CZbeFSBna1xU/VQffXWtD8vx9J38bM28tlv+zkFfxQht6UPJ24BBmrDGv
oNEDXrwKSlQyW6SopokxjHP9y0lPXpoVAzE9eJOflEa4M1IVznGQLI3p/+jfUUkvqwrTpObUcTBt
zhshJQ8UgOGV7zrXcvhs+EhmI74pUY/0s3EZn5INgvcJGA4CVMwupE/7T30o3hUQ6s1uf36z+i1A
y+gg2WMxk7RxZbHGsPEV+CjwZWJNR/STKyqdN8Wem6TgEgoc6JNGqF/6LMZl25t7EoSsmNMkR5IJ
TM5b/kmP+RX9b56KGMONlYKtTBW6VaDljpI1p3eyCcv9nl1Y0Ce06plviHy4MM11xiT/Wvlbb+SS
puaO8mBppnBLDDSMLlNOYPK4Fryp1VCq5RyP/8souiU/XAFagq22IsMiWvtakCjr2MRBlRfPUKE8
+9N5aygsgH57LDFQjxneAUmQpI5jPS06rbvIu26u7SlQPSkMHP1fzrgid1GkdxFNO5WqfN8ycq6C
temIiR8kg5BJDdNgC4Y2tdZDhTPaitePofsVBJh7CGhNXKgbnkVFf/WtSrQ8YJ9eMnioBQLXAHwV
fV21qEuB/EUzdG+S+sZ/du9ueRkgwFoUvgfS0wXRQXTilu3CcwX2Y+h6khg2kMqSs5dwriXKfCSx
nyUrYdSqBH+sRqTdfDxds83aMiD/5hreY8RlVmk3Hn7LHLYy57+gRGRgwra2yKrMEt6lfT2O5h2G
vYIWK4jJOBXEbcO6kEvTHb8QvbanX9LDhmIw5CTkDoaeO1UFGyCW7q+uUpIBXTR9QR4bXKYy+0cB
avmWoDTQWSW4x+OGNO1pYkDZVtAoloo9uD2chtODQ+u7neCQBlPvfpN2/O/xbhp7m/WLotfGa2iW
LOYCkhwkaryK0lVZVBtZp42/+d0vh2IUZChqF3oOIekV1hmnuWcWml1KLSYh0IcERdv4dupZCmm5
k+3RGE3eei3v0Al2SJx2dp+qsS+1v8Mrvq9rz1oivuQQLj9fBaEDE8OPpbtwPKMaiVe9MbF7nldC
edsmm94ZCWMjyl93l/CMFQJGgwbLm9/FrIdpz58qaP/QzUVDtfAceXGUh26gkAIR23bQNEjXH307
qbJyUY5NKVSfg4yaBzpE7aE3ZCsdU6nVN5qrGD+HmQsAiY10Nwb1MPw94hb9ZLVgPyjEik9sRAnG
mT8EHBc8hbkQp8B8zFubkxViIG1T6vuIYjPndkGaSf/C41BK5GPlv7iaTB0ELmVDoWMys6V2FE3U
Bwi85fImT1qffoyVQQHsi12Fvtv+NxtVpqPUu6yX6AhdjXPja/nRIb+dLMvNjl38YuLZsaUK2Fmt
/rKmGcg0T7G8KdSYV9WDUwdHfONqOO4K88N2BlmLsW9cdZHhJW1GElKLupenmWz3l4Yuke0hQ12B
2oVFshN0ctbUhN6AIi0iKCIbl7znwubXnmppRDponpz1nSC7VvTpbO/iCfJaDIWg3Uo8IRPguQKA
6fZsAE3qu3DP0UW2GPSwywVrZg93mluY6g1mQbNzl1WlFe2KaFhJq7uJuibV89DuidcEVHJeKO5s
ppllitrdMZBc4A7FqdUdOavyvEMP8gFfDO5rY5/f+ZJPeZHjCLbsNjXgtUePFp+UgolpuJh1LIF9
Gl4GGqQT6b/wOZJCToxQ01NVsrXU7sRT9/BrdrGjNZWHzG0Gq6Pf2LePc9ocLa8ax8QAVRah6GjU
cjrGYESYACJuCsCuGXYQOj26ds6zIqo9xaEPOJmxZRphj0ss3gmSOBh+dn41EM9lh0f6fB21WdMK
srgyw8yREbNQs3DZScrLhhsa9DX0UTolbQEMjaCMud76aTb01t1A9PHWJlVGNxlE2MaiRj7YOjo9
+EdWfbUdnDhSBFRkll8QZziCSF4xBGaHfoQawYnuSulj19Vby1TSsCdvn+rxUp40z5nrzWNVYBf6
VXVGDOTpyV6+zKSe7s1W9EjHKdHx6ckwIr6jgYNV392KOQddnzNBQzJg3Mfpuylv3ZqOOBHsffrb
yLc36GCX3qz6dlkw9qx/hwaAq8f34G5ck//WtRYrEfZjwB8unCSEk771yrn43dmUFEtsZriRc0Qf
5BuzUHhKcIJkAB3o9amwoTTUYZ+qUrOeWXw77RO74eZs1pV5kGEqSB0TmskX8+0bBDzpOmldCYln
TbHtdqPYRiisu6vtScOPEtvYdSxpU1Hdt2Pq2XWujS3PVFK/0KbdKtVnAGsb4jSr03Sa2kDtD/Nm
6iZAv1fZ7k5pT7tZ1KjuroqPN1plo6Uoj6Bjde351sywNbGfGuqaPX+6n1I7uGwMyYGfflzZAdn5
OOnB/fH45DQn+qPMWSwTVscryjmr58DA53bLCFuq8fIlUTI5nlj1dtP9YJwi9vDHTm0dzC4ztLpU
0cbneVdSXefHj89Ue+6C3hrxI3f+mKcPrhZUwIDaii2garofi9HBlLRHSk8/t4fkVLV9eaaW8Ups
mT9be72zC9NXOIlg/rzfKmnhanoWBD4ubaxuaHEcPvbswIRw7KP/2TLK1zJXmRUpqkljy3GKxetO
zEA4fvjSE+pCyeg5hgOeumECs4nHeuPhOlUYCL7TqQ9bx/kcfzeNcenuBu3YE0w84F+TLWoziQ2t
SXsqv1U89jxOhcKBQaoyEA4GbT8vwjM7QoLT0G8fFJkcT0SlJCkJGzC04/Qkg1LN/a8wG94PAD9t
hn+X8olDc4egnB89uVJMh1SUtR7858+mCztFTgZ6dpm4cnEP1BQFO08UcwFBVF7JoGssv/hceRt1
dbymLh6vxM4u/PIYAm3NCAa7qsTonmRpiOFl74aDlmzXIvnyoUsMNohk6sFuvJgc3nzqi3LlCZka
qerex/cNGhQUse9FBjOE1iYBgHLZ4Pev92khVrlYkllOjr/Da2RFgReVfG2G9rIvfoj9ixHA5DNY
8lmU7yW+cna/zaTXRqZ34HBMczf0ftNhsTBXIZjhw3i1BEaHnVAJuDZpfgGAVIv6O6H6VWpB+XoX
HqhELVP6XNoCyNT8T7fpJGvsrmjw7O/35NExY1hp4fTk10WNrQJIeWYDvhVZ6jakzLXAXOM0BTcU
+yytAS0kAcr/m1gH0dHGdKPm7y6wCTL9MO1r75F5KLG8P1ZoQmA97HgzdeaMczbXRToe5y5ernj9
FDFtKepuYF3tB2MdDT5RdUnm63ruPtelGi/6Q54VgLo/lRnJJZooc/alEPR6kSGZoKqz9AIpL0lN
rQImx4GdZIgiNW4BFrchdDoBDPEmUhEB+5tRbzhRC36nqPsg4P9l2/Eax4s216q2tKeqvMD1gqOw
MZvfj1d6tLqFUU2ukIAK1NHP4GSFd/H1z7FE+Jwlgj44+PMdTuT4fi1o/2wI+hWMSLHm2VwpbdzZ
djkCHvWo87Sc8yKV/KoTTnp94+N+DOi4dLqpf84AR36Ecgz/w5x+A4MErot/v0WNja9XxYHBcd/g
fDG+gunVXroZE5TwhdbGCInbUoa6jabo7b+3RdiB9ChOxPdjEb8AoAWBsxejcvdVU7ynKvF8+M8Y
+vCoqvnZYiHxiBJShpKEbfwL2wWuv0jWke1VTx8hfTN+XTqCywO3dCnzPDYkfNLpLWTnvtWbViKc
wpfTcjun+3Kn5dlN+Glmlp0t7tpuL0GDavQDRQcbRD3wVadf7meZfn5zMcg1ksqo6pEEhfH8U1P8
qQ+3H5NeYJ4RedCaL1UiMJufKO86pHSFdHv+XbqvbfZPzsQ9B3UARbMBU32lNjwc0Gsk2EObQ9B3
jhkGIhHnpGLSahRKodlc14tEAGFm8oLr9f4NU1PEKVC6Psjpa/3PG9bHrjBvvBwYAqTxXSmGKNIM
cvpVqOBjNOR2VNQMozhnkpAt8ApKbbXjm5HJOkqplHrUPRzFhsK/NgdWjlu5oYiJQvvVL1jgukgW
7jMS0bCPHBW9GqXn1cN5gj4Q0IRDICiFKWTQ5r+9m4iS1ZW30u3tUL14KPASbCWbZnTemHo7u4pY
AzvOxNLM6128DgRQ04yONkbh7lq6NTey02Oi3AcxDb1l/LPO3WWE5yzf2XjJTn4ANe14DKRb6YBE
+aP/RnKRAsTL0FCGKOhCv4lylUH0KJnlW7+hcOhcpJDx0mxxgkA9+45PrqWv+HT093Y15spUanRJ
gGLgOwMQsL693Dfj1dDaz7HAE+vLWkArlKiC22QEUG28n4XGXkMw59gG0xHgB/m4FohH3mzaGx3F
m0cahKvDqKuWsIBT/XLbWAnq/853YfjomYiMfSRxHcle5Odz4v4+/OYROi0mqEz/7nPSIauLgC84
Evn9fmjd9PIdaVZpMytNOPztaIUVUanG+tYBnt7RcKuDXer2J9h6baF49LcRKZFPog92OpE/DxeV
dXC6JBCLACkc3qTnk4MGeMQyR14+ovrMWFbMpQ/28yLfLjpL56M49H0jh1zD9lXC7SA+pRIZdT3B
8ZsJcBIZakk5i2zNxazRi8Xv57aRvy3taonlb0RTvDXP9fBuUP0KdYn3mm+u7UqLkbU3iIUZAoTw
jcfkngWtsPaOEK+00VG2aXpAHKzv45dbax6kyLSZubULnJrfXkfe01CliFRGwsuaVoMSDoS2hbES
CNfGS64MQygbOvJ09x+IURoBGol/a5PmhHiaVbhtO0KosjespUUFTgtSKz4cCbeR7eJSfcKCR0xq
9o3qkkZV0J4rbxIuWosnnumksw6pO25J1EcoxUrgfbfXBaOHfRjDej52gBR5Gmv22JOx+9HASMOa
7FUzcw0ZTZqaOMB4Qn6tPF3JY/jbPY65rH/YchoBkrCPxVi9RzKHq2jnt21+lndMX9EOqg3erYkv
cp4keXmcX8TkwyDiKny7WuZ4LFe2qZiDLd616sRzyvoAAdZbRHNmvQjB/HoyKHHEWxnH2vsjETYA
ALiOOX2xHxOfBZc3tZci9AtQr94eOGh4GCvmjgVj5N63Fq7i8ICq7UtYu865h/pu6cqrGCgDWqMZ
FCaesPHQ1MvSS7mXFAULbRGQL9p8PdKJ6usS11LkofE+hIa9U2Z3od6fkRqhrw/phNGyCXS6PZqD
sfzzvfG7SLDj65XN5WnwEI4hGmdQRk0SuhAx2xyLSQDUrWNE2CBLqFRY45zgu5GSKRQJFrMl/j83
+6VOnV6K/Zm+oW/pW9IR0MgSKdPCx7PlLjK+KjEbG2pNys6Xx8P2Q5R0TcvBADzmnk3f1oS+rv8v
TaEG5w89sA2xMf8CGJQ5RAw4ZJt6fzQEDj4mXDk1eaf45dIpgjJPDRuPYvVZJt2nVhylNfe7Tir/
jOYu12I69eszj4DZXE8MUdLtaN6Aj0/mSStzSwgeeQB3rPpWS7BSNRJjm95/dSqQeJu5eUkSp4hr
FSl4zZPN5h5KQhWgsDUyqTx1GMPIx/qhEvlTnYNPmN9FgWEAinyZuGQB+WrLxsP4EBrIucGDULWG
WvnWbd5zz1xk574VaJqjt+A9F5PFYD9cUPSMCy7KtFP7TvskE8TLDXUb8Dnjof0jBQ/49EdjnGa0
wrXizKlLQ/j7CwKQL3GxHSbVIZqYErbvwG6eo13tBhOQhZlJiq0Ki3gEe0DACBR8a/Ll+mLON4xm
CvguHLgiYhvppkP3ZvkAukWsVFz8rl8rSCR+1TIF8e1fxz5a4skYQG/E1tTW2VFDJF/DjruZ4Xji
550TiXvVOgk2WBHem2EqkBuf3VhVIO9Bc8c5P3rcQrWrU7b6vpH+cN2oVBP0DGx9QZ4E2/jH1C/V
o2m0mMbZIb0Uk7hnG0rAaQsQjeGiBTUyvlJ9BN1HQFCdHSBO53G/Qp4A33Eww3qnQYjDuS8uTLIc
GaIrrVWse/8bE0hhLlLPCZmt6ERDHPf3aQkpWNxe1LcStpJR0TAc6kE/y05kxrdVrCswo1V+4/+V
bKHsNIQlCmVkt7s4un7E0fIoZqdO1bTDJw5sahHty0CfdlVas47ksduB1LnzuZ0WJD3zmxbmkzZl
BATG4ollgBo1cgrCnsuGsPHm9inxhLOMVosJSDt8Wj9YifW0KSDAkt5YVnoR/ISS0nzZwW0+HgBA
9k3460FWpN8CzljDRmMTD4E3eNvlvnNyMR9OOMEfYPeMoy9SKNnp3FjlLTtkeuTq2kf95TAxLbci
/rh8sUVgABQQ1iq9XGYftlvqHXhz3tkeuh8RzBOgih3gwjuHK4o9e4CrlhBiaOEs2GIky0Mk78V/
wrIX2xefiC9sB9RAL/3pc4IPPoZgjCEyX+/G4vRLbt/tZKHIO6dXhg7hsdn9PaOd37x8HwYKYdgi
V1Z9CVeagB+7wG/u9tvVg/7qvQg0yhO6jy6QxfgXfSFz6b3z8tce09lmlqo5YMjG+4hIQquV1EY5
F2O6+xEYkB9YxTVMJb1RHKPkM0DxHXGrWYmJz8OBQ88PH52KYkDfUcmPKojv+tZi0U/X19p6mfK0
uI5Dwmi/XHvNU1h+FPl4Moz3gH1tcIAVeIzetnAja/K0XGs/zrnNLsji5jVUjgJKC/9fe5odPWs9
RK6VtQt4oTciBrQkymrFhH7yO04bUNnlVzCNmKPk8jRZFAeELJH8HC6NmU2/QjBGvB4SnBYM5vg3
fMbfdZ87HiLE4HAYSGS97YjCJmsoKMgVK6/64zj1FjD6vpCjam6xBHwtYImcMmrZ7YdTcjaUmz5n
/+ydJIoFQbTZ0P8ekqgXUZKlzNaRukmud2dlrx76TisZtPNm+5ywK4rNW8gqzvMewVtb8FVnZaSy
k6u0Yi3L9GaWTQI3L6ZyjuhHLK8CYZB0Fl4LKwcIXVmkEHp+N+aiIaMkSjdSvDnmvrXi79xfoo/r
+4U1c3mi/ThwLHElLhzFuBybDZvwyFWLJzbhmWNf5hS4eDfq6dHqs5WnP+WFIq2Njzn6OfP9WghM
sMfKYZxXxYwrJQYp8utJcdRBS4mIusn4FOaVBaDr0asdavtipfcmfJR3RNJJwd7YwL5l/aERdbcp
LGT6qdJDvl458ySW7d7Yi7OEiO3iMiv59CcUk+xFGT/YDBWMbD2UvCf8xpzryOiBVrmzxjSgjsxG
str6bFBBHiHQ3Y12hokyqzywuZnqaWueUgGb8cADV4sXRHgXfFXdYDEIXxbjtoUxXnfLf0Zcuy5Z
BIMDtlLFv8w9YP/Mify24xm3tWjQ/F1UmIXGBOcF3TlZpBpBrEFa7x5v0FSwzigeF74mQ6DkOo4r
3Rvt56uSUGu2mkBhFTH1vssT0k2lVoVWKvpVzNV3xTzR8+6fpLNph5keDnXkSn9oEUzr0OGYKzwk
OoLaA6ERxgmCVqitFD7Du9mNICuBXwIEsGULCew2LGssecbs8+KbI+D40+BPIG5O9h/yea0gdY7c
H///7FRba+4uIZBEKaoCohsW+XwcmnbETh3ndI24IktQ/Dd5/mwS+B1YxzTYPhAgPbTTwFTjzifn
kgNNi9DO8VQtO6+xeA8hKTFjk50agR6VxSXCkVUNk+sGVWOIb+BWX3+R+ZLBw9XJIaSNWFpHqWJV
ytOELx9qlPhR1Fo4PZjxM1GoicKexLGCbOdEEpxd9sBI52QsGLx82FNrnY43zQtnRLrCwEhNDTwj
CecC9rLyhG0lutdQ0O3Drp2vaLhEgMKk6ct5hesJvUZ6VeRPADcO1QvAFi0eNyYZTKcNz9JjMa/b
TN+FO5vaPB1fbK5phSLe2evZI0P4KDjHaesdXZOoeNWRGbSfmDeOdsPsOqwPC3FrxA6vCiLvxqEa
zy5lWqZHmHvURM390Q7Gi3ySbLf5pVBFDcAedzEUPBZxRxrVbiRj/s4v8Z1jQ1s+k8jpnIrsECP1
5RzuOmHkshZYtSeakqhEwluekmp+HmFydQPl24Dlh/N5toItU3Yot6QLeDqsMqXVcA0CjCBEx3Bl
spAbYsKLfMyAGOsLF/yNLSZNfu3Kmlnic9oCEO/ZOSR4c8Avj4PdeAE9HbAW6NlBPrn/yO+YCRIO
2t781OpmOWsMWVO82Cq3rr+7SW+72B4wt3j527Y/Vxnppzg0YHqg5yKojZrdwpiUhztJC0zVlKoX
DhmQyBkYa6d5c5c5bCeejzIC71v+yxCj86b8O04OCue4I7olO2kD3koaaU2CGGZ6+fnLKvpsRSFM
1/Qc9uOeJQZ7ZsgwLL4YUgV+3aZxp44cYH0nZ+mOvbLnANZ6w1AgSOWGap1JmQ8dnaWCdbwm1LLe
c3Zl3UtWPiwByLWcPg/XrtiWioyIocpKz1a2RIITnz1rffmIUAs8rcoJgCIN6LH3EggaMfQwLEPM
euAZrK4UmIg5AlHSCRY66DbPsXeSsoizktSJDShcJwI/hXFPZXOM8zQS/335Tah33VzrpE15Ar1V
KUedKip2RvDaEx8l1Z/6TYoaYLMpLbQ//y/Cwu5A4PreQvRFT7gsdZRjzCiACQZ66fbqHSw8DhmO
SZkUhkLd3zY0/+qyHPQBBOH1abFv+jEMUjyUC1WLEtpD6GuuF3hTkzfzVKPu4Brv6D8zXh67BgSj
ZxXrlPkTcUdg/tD+rOAAcp4e/oYEw7GjNi/Vq5EiWkWaJBg4ln6EXLf5CJ/si9wYjiv8bQT7y1FC
+JF9EIRYIDqBryCwdCj7VS6s2m8A4Mq/aqBoRbD0ovMJ6dohlyH/iiVKc1Mc8Gr+8oiHOgc9NOzP
kNRnpRu0qyPU19Ve8X/16hE78//gTBXZAqbc8xmpG2vJ+rTO3xCWN6ikh0JR7HuIR4nnM7utV/L1
6vSjd+D/8wnnUGrdiCAHAYjAwh1nHMdoRY8Y1FuQ9ckZMkkdcqvRJDh82OLq3zsDFjTwATIQTQ9i
1FThrXlxuALSs3LJBhZHKH/EDBNgZ/e6qRJWXe9CiupZJKhDkX0o5FHaxCIGATNewdOU1ewa3JQ7
CUqT6HQxCozGNsSds59DvYLAz3KjvXU4l8buRH8fO1oUg5fflYk3TeqEBOMCb0fToUZdHg5v5kI6
nSVZjYDzy9TKMfp5dPJFZ6orzuRjCBthcfubfDzJ7tj4UfpwJ/2+haDZ4zeV7THNxHjiNBk+/Y82
7gwPBoSZ0KMSVGbVXvz1Nkbr5FaPGazFAXO6DRLRlJXnOb5jpbqiMU8IF0HKph+owH1+Z6iZapJD
07JfSoMwg8Y4xSvzpBsBvl8a5eISdBnD/p+4b+c/CHTbSQZ1ul5toMsufDrc/omCK65TKvCH2dSF
ZvA9kDlwpnNf1ZhPTAWprkw/rSQbkUW58zoDP7W19BRGeVw3f5xsL9evbxD5sVNc+FswJTpCpeQw
inhaitYVNBmQntc6RCRI6M+mbk9liJbNK43+G6wgHRolBAA/ogfdbi4tiNW5L67XF2tCGvxC4NR3
huyn9p/nhZgOuyCAUEq1CGofPMz5508M/+JgXnJHn7/hgOa7v336lC5Vo+rGLhWCwUtgBYmCmRae
/rdttd0Cf6DDPA1a7JxlG/VJ6YOlbpd+wBIomuP2bPkc2gpajMBvm+z1vqpL90JQHFfkrGBCzlkn
5uSEWi9iKDmzNz/e4dPskfgmNqeV22wTxOrkF3o9Ax1++qqTf3F4Z5KsSFRat873jJRICDcPOXhZ
8mXrg7f1rjrvDZmsc5A2TrGuLnMvbI6sTJv+SCbJuIFEa1H/9rFrzpuL7JICZo+jjM+GJ0QtSTUN
472SxepC+9YT8ulPy3vEUeW3IgRAhYvzZv8jwxzRCeLOYtrxCeljAGQv5A2ZXXNTZA7aCJqYMeJc
wDZnUrw3q6YHLqhQthtno1BDoZcwwtcnI25QrbaYaKCFE9MktBIyAEXE0yc23WbirqxOSUVyJnR8
+wRh8cjhxKPMZVwh2jlj8XAQNspw6562h/FO262wwSTzxy3nF6ePcXeu3Z4UuoK8f7NUS0fe84Jx
ll6yTgIgTo7vYwgVnTuvVmjbeMxiOOvkABdzuqOcG734Zbr2X4aKOuH619VyR0a11wS8J9qNeqIV
G/KpkFqwnotydibl7rBmEGuxdJ5Xv6cBB+aKLDmR87Qyo+tu7v7NH+v0Hdeyc5xV4c+k2Nhql7JA
Le6j46viLK7snZoM6Y5kyusPNpwetEUZJE2q8FSYKa0hy5a5vrNqEJAXR/k1veJDe1BE/RDnQv92
bKtunm+Qv4C54udMcUwC1qYJiiXlouA270zmElzUgLJO2/oi4QCMkdFAx9hBOoqQQ2FLjucI/8/P
tjbJ623KyC8IkmIbgy0YA5OKxW+JASictnERkY1Qcv4twvSjMJOjFe5oIiLoOihLk+6mFDOJz6yZ
muFK1UEQz4hkSOFErGke5jkjUsSWWp29TS1oKqvg3WiBDl9WjAT5DR8lDQF24xiQ/Y/3n0p4CTdG
UIIgKbgYxmC5efa0n9H+s9IrHGYb2DHkKA4/q7tmRGbXSTnxEoTQDFOmATtR52zFKsa6MTMmyvpF
o7PKBsy9oexU38KZ8b/jpTQpxcRYSp4eqKcFnCjnZirRcYm0CKJaZZ+mAAttXyDvCA8/9cSj7TvU
SPkAxddy4+WAh2gkdk7mKkMtQtYuo9A4vvX+56ITLEkpAOH4nBbxrV+cKIW6/nhxw6QVQnFhykBJ
FKbumjnJZw45Ku1jmsgrc4m25zdYD06L8X9mJM9NObuxqR7gHHQi7ZeSzM/C3V3NYWyQ5SchiIWV
uLp4FzHqYcSOKwRnzlK8ePArJqaeMqBVyJyTQ1Qq+xesV0pTnl4M7mY7YI47yeLmZOavFIaXInGq
xCkBKe7lNpqQwFXrpOmdN1RXoNMO5U4N0RuzsAhrTtYrgUwUDmehbvuLPPiFgV3FCIkTSXC9+S+C
owUGu7LxNcn6dTO3G24Pzd4NOcTQE5IsjKNdGWzNpJnPHxguQsyOdYiZWrpbhxUHkI1IqQBpgLoy
DykJIKcdZ/zsxAyamMGfqYK92V4IsM0LkiMXCQnxG84tIJhHRiGFpRpvVH9oHhyJ12wMuPYLKynk
RG5Rsy/clLiPsYNvutuaipNo/ROmW9sOUUHR31BHr1Dj9CRixDqQE67CcCTWaFw03vJyvPs1h/R7
9G84ldkIy1rjbw/Ymd2Uw2SuDmCf82JdkNiaTG5BjnGhIkWvcpmMntap43tbUZaICnFf3zlEEa1f
hN1IaR/7JhuM9mP2thvwER+N0Dx4W4gZihk7/sc9D09VZvqLjD7BGwrRjSV/qwmglZu4UlMraiv9
mRgdM+UHFpuHVeeluYE8VFM2oLKeNGDshq0c3GUJcMNChzQvyN9JM8mG+s7ZKRE7jxvmvDe+pSHU
gY4lFeMxBisPFmPFMyI2sm50LnV/GyffUQ6kbzTfAdU5rJPpZbyWz693gPIXSMxQUL6ppBIiuMWn
Yir2qR8XM3KZJbSWGH/Gv9+AYWOx9Hm+TMR8ndg7X0H+Ztu+zLzFbHbgbLUOU6cKZEuBKnr03/vR
vdTRcMmSlbc0WWsVZVshD6nvTXueG0S7NTKOE/fQ8oEBPyEPd/3ZM3d+J/qwK2SumCITuZ2j+4u7
dU6Uhg+tHcg2N9Ncx0xJQrPyAzEcHHtehVaDUbCUeKvDe2fXsKouqRPUyyRHeDwSmrtQ039OGJgd
SoZ7sqNJ4PBGpT9AMT9m38KtKvTre0MjxnEvKR7sKR8EM3Egh/Pe2WY8+sdrT9KJP+bCCA9cFRM1
F4bxyVeVUHNotKtJylRO6WGVZrEt8T7KWPS/34zw7zhevWB3iy2itfYHt3FKuryH8OyuEhK12mSG
Zt3y36JYDzSGe67bgfIte5TyPVoA8x81+7YpyPThNlr7Ck7jDpDC+gkRsS44AuXOMdetK9BYDKal
6ZmtJq6e4u+jSGu2wB1DUtaSoFfa3pRLX0vhHrVZd4EFNiEC3zzQ2a3osVzjjoRaF6wrTBGjqTEM
I8tJdWYKQRmAfXZsrtRDh9dyg5TuuYCDEBYh+XtEKZIY+jFXDF8l5bCwSiDjujEofuWm4eTUL1hK
utBT5286SW4LkKMUo/2NSe1geNTxeq957cLJi+l55RiaDSH+s086UcS/rGI53YuMXY5mBdm+Bs+8
e0uy3AjgtNp/hJA0CPfKv19JbukXIbJh315Rmjv4eDZNMyZIMs4hPbnCeMoEUZB8CCah8CBf0/Gp
Di51ET8Hp6qKTgjmM0ozWZd/KfYgScbsFqMHZrUWVvfeemHBXS8IKKfvRCWC1W1NjGEtfnJvZzoc
ceJyGu8xylNusKQChozSWjikWX/Uo4O43o4f0AMnxbVzZgcO5QvQooarpaRSyVGBLWp+bHTAOoPB
mrzoauyDE/Xv/om9Z30YMvGln1khaQX1MZx3U30PQh3MatwLPqBHCqDzhNsD7FeYZCt/bL90cRaC
k+c0DIushIqmCztKg1uX9AJbYSaFhhfkqm/SjKrToiLo1Kddv1FlkkdqghDpADxnd8tcEZKtVb09
YXpirD8DCsnJQ3cYGUlJzu0lfH0Oi23QjthvR1LUPLwNvQi3oX1DZXJNpzmUNQ/t+WUADu/M9JDa
iiwe596mMOXpKYR79XdhJzP8eNkE5v6SIKXjhNOcqPXNOyWK6p4W6QYxEZrzIxv2V/mgQuIymmAN
B5KH6Wb8YTvPO+nfLeNPU5nwbjIDDqjCmU5MA8Dd2/8NtGQH5E6J8Yx3A6tO3nJYhRF7E3UGTc6V
r3gx0L39h2JFFkEgsmu60ENOEWMvi6fT1fdnvrFr88Nbl+U52Sl8vh7z4T+QQt3ByQ8EWzI9WjQp
YnM1z6dCfLRbUzCDEjY1Q57qczBXfltYwIf7nMC7wDmleRxQZNFIYSdrwnFC/OoDifCURKEGp4nJ
mDH3fpOaYewEhV54A3G5tEE10iluu6GHQx6cY2E6qAb0g3Q2QOths8fBKt0jPrXKrv4mmNUM/vAe
xa7B2Ewc6+UAkPjl9UcreLhv8U7BPfv3F046mhu06UQL9egJFpfIigzUNyn7DVb4qr+/DJ6aRPbd
LPyy7efR0oOGj9nACD9VYDedr5TrxWacsiNQChQ90Sp5PPpFokkGCqBEZUBLtNLEGlwcAUxuhM+7
7n5S42TIUhJre86X95XQFTMiZGzHK3R9oUdXnQKhmTrc7Wv1Gii6+mQ9Y9jfAOvx6UDTH04AEMq2
uBF5HVy2N7kJsj8J0/qsizSTZgraVyxqp8N0WXDbBkcyN6+7vLqyuipTu9i/u98LlY+Leqm/J6SZ
nh5OJ+59U+s+xsEplRA0GPzP/20srTVQRWzNlDNJRGdgSEUydwxclsYcvC3qV7EvXIneUqP1ilyR
gchhCns7QQdt4+MCCG5ZOm/I184ci02HHLFzMxgf5u5lLKlsUGGTrtittfW/ZQoUHOgX4XgCdKUk
pqA1VAI9KjjEose9b6Y7WW0JB3lAVRW9pQoWOtggCmzHCw/Wfyg81E2E7ORjaElQ622k87myTMyA
rVuJ+Tgf3+dbGuIlaD0HHhF5jtR/fGsB9DjEryg342uoOx98LEVWAM8RO+L2XaqwH8CuO3AUAjNn
T+dczJpbxJM+IMbifqXnYBuGsSzPjwSiJVH6F093dal2insVS+HIzn9w/sHGHDxWPisNBrWpexFS
zG/gecvl/S68tHFFltHsgN9W0u5ByOyhxC0mZN+RrI4VFZaXYuWNQrSfeZJDlo5BBgdVXLdUj+tT
7i57OTACc1DEYescvTxhiyarYZDxF2q1q/BS0nSZMLYgLb+6/Nm5jdvzr0umfOv6oOZ/VWexBqM8
UA88+9rG9xU3/56/YTPvypC2vezPOWOCWb9fZi2BCqyFc5Q+SuskkKyUaeoTV45bnSUhFGfFu5YP
j2BH/jMsREM4DhrEBLmN9qU9K+aWnfi0/Eu2owhc8NbAbn7jNkuQUPx0LbCn2VgRdyHQVxKXGoux
LkWJ2vi7WTXbN9yGcjjJuYtyVv4qkH74aDGD1UDN2IQaFhI0qHDNsXIQHDDricM+rrH4uSLDinrK
XCOa4xtuh64G7cl8s91GNSzJvlEMzPkwnKYaxF0ryRZmg4AEBLBeuJYv7LhBa0yimN5G2i3RO70C
VbisyGmD1Vxoe2EoRHsVwIftMq4y+BiCrc9/yp0jsxdKwoXiEgKtBabk3g7vGUv37pCTpuHbxV6l
sfoeF4TL3ex5MTeFm2gzhgdXIa1QHrk4YOk51la2cpMahXCZRgY1HgARITIFsatqW37bnsoDPVH7
rvI/GNp98zOOcIcEigCGX8UKce6WAKe3FdRNIBkqgmUNWnjpEvMyFPWcuMXcZA3AkdtxqgMI6C+G
PsAT5J4rXSgwCwJAfh2nCz3ZxTmPiybUpzgK4Ck1XgNbrigypa9U/jHbDFQ3aofgzI5kdvNRnKKt
oGiiJ+PW25p/ia+RXhSL6nAS5XYY+QqEOJEbfBjMsslhsw/RaDkGCM6epTN8QIomGiDS06BYLvTF
nFkSK6z/C8Iw0XlYaRkVkuOyRWW9x0QoCets6N9S3FkaihU5yxG2PxzDhQS+Zl8/MEprt8Vpf5Oh
vocleWeDX6h+n7JtTSriVFo5nXxFmjR5357E2IODVS2x8+VBGjQeqlPAqir7HR2yDHoWNhK1io3G
s89gTUCYmKFF7+LuQwHz547N3zKjqvxm1PkzD1eu+X9FD1p5a2N2UFYG9OiH9eKRvHXzV2VGKxUq
DtK1rQRCaqKgp/MtJNs1qmOJO0i7lFACiSUZfhDQqpeBI5foqJuj5Da3UUgd7ynYn2BVzwPneqOV
faGE8KukljMQsqchc/t644XoJF9B9MUtUrmshOQadHUJ9cLO6h+mMuVQV5lZmB3vJT5j6VUEud9T
Zd6xaCu+ErweaQZl153VSVU/6UGqUH9soe7duyuJBrf5ler713T95dyNRqOJ8ZjN2lkGKDcpS0ye
tCWf1FEusBxlpWciGYPiqjibuJk4m2TSvPD9pgTtLechGSpvE/c6JzVvdZkNc4PVH6IvgX4wBOqb
t/ZepHnqDBWbKL30clmSILwNClqNvyIqUZAAcAd3XzYQHUs/c7D3VcDGz3Pt1NI0rViCZEsB7r55
n08Rkhdc2YKbxG8lwisFiKC2PU4DdZfULckWKx06hf7BZNH4AUMwmsoOYpe0vLwgaGSh35rrp2kc
vdiRPGE5jXBGrMgfvUfhkHRuaMCi+i2Xybxp6tUVAH+f5JduKqjtkMoTSGJgD6V1zBSTjXkc5TiM
kfujRU2QJoyYc4gzxKtFb7J/jrZQUZ7qQR/Kx1nxUIRoL4goaY+uY2kXYyITi+zICxCg8vRj8GPb
Tf5OGlb0gOAbmaCb0PR7Sd4ZlhWUIfv7YXH9Dpd2yXUHx6iM2iekS6mYKRFpo3ctStIvcoKJPpdo
Tkjsx2Ds5GZ/UqzunukALVdGtpv47BN8kA5OVMsWpBJ4Dk+GfjQL/irXQheV1B8/jWxKV4Ak4arB
VyJWqUTtkPZGXagFUsImKWMZUL15AEApUl9DfWI6dBiGdpmIzBtsbHrGPLthkkRg4zlkoeeiDIav
4nCiV6y0l/fjTDGn4Yhd104ZpQySj9kPF/6Sm2pWFnEzI6S0rTZiNgRmzN7T8fU1X9t11d8l+gHq
GlicNEtar3O1AXrCFm+IIQaVYztpc8jYphgLdnNoSArRpeC5bv5FL5NquDc/NmliTzcy6eEW7eQO
sQiNbXieiGI+7VapsaZoBjipJZS521b8Olc0D+h4uuGAkEu87WuGpDR/9Ikx+XyDeIGzHg2x9f/z
efK6Lkky/7YqlC1dv4ajF6z85j4uIzbZ7LX7broQDml4cbOL6cOUEWmG/pHg2QDgdT8GPXCUcNqZ
tXD848yfeiChCS3+Dtn6+aV42Ti87FkO+gZ/jPcGUsMQrzhLbVNG5D7JOVtdHAwAoFFivq3lEdJh
MOW0AYmPTeHe6FcZGDkvSC7tMdj/38V6puInwBhLjAJwqGT6f4wA2SOLEd6gpQ8lasFDLzkMtGSW
W63OG7bHb+YGITB5JLnbusXhbPb4bUwkG13xK45/nao/nrATiVmrSLHpGL7d9tTV+x2xEwUpz+P9
z2QN16tCDUCzde3diFbURyKKT8DOSqlnV7oNd5DRHN6L/u3Kin4MNQH5/vFTr4UpqKGTuFKddfj1
S7Z++ApitZNh170Th5fBqTFKGEYI+HEaE3NuabI6d2Z6GW15g8z1SmsFeWnDIXvgQ4Ax/VDClNm2
ZPxN3qsYs5bdlHjOM+WLqNBElTVM53EVRwkqDT1+BcwmFnvsqzQIMzSbzEDEGJCYxn4zG5Hm5eFZ
1kdkE4hpoB2TYieX4UQOIf59WcC893bEaSDk9sDXTST+QCimcyJbMDXNfrLvJly0GzmDnckCqSw6
lAfnhlx/cCwpwzJxI+oH2qladcCOev2EBCQ8d5q9meemaMwXt7ddSEOH0jt2g2irl5Sxdpw6XLg9
B+aOWb2zpzV4ZmMOHzNKTynvEtjZB3QEvrZZCJpdCjn4TnxmGJF4CfvxrCrL4K6mFyfy0lLA1QY0
mMUqTTxkHuTDbSQzSJexKJDx/AZ3/WB6dGgUKTDUpzAFwYt6AxcgXr2s6V1PEDhMCvpNy/jn46nZ
T4p6iuqAQnOmKeriEicu0AyyiOu0p16WtLsIBWLHwKJjvulTEQrz0n1iYW8J+jIQP76JDvbS1kEX
q7o3lv+1saBwnm2/fvehm7sqTZYSUVK+diMVbUd3oDTwW+VibyrgxwlmeM8mln7drXFf29H+E8hO
WYs5bujsOpmB5Hayc7wZIrmQa/lOJl+E8CGlL/4TKUgrIlq4AmD50IGvDPWaXz8M/l0/kZJU3bHV
GoLbMJ3M1qKF/au2ncYO9VCRHKZJnt/msnhPwnRuohW1ECypsIoJis9kdt/XD/7jIoUe4ah/2CvK
CwYjmxmY0HYzCpOzim48u/Tl3fmwbRNcZRApvd1XszG7tdwfPAchGwRnQtxMep7sGa9O/4wCtqLX
kccEvRqheV1YTtr69VjGqzgIKM3D7LtG3ZQvCblMLzxFdldmrv0pZlZUe2yAfkjQ3NA7fLOy5NU3
YCHCs/zmZ+m2czbG6kgLu2H0/y6cIYPI2Y3Nx7zUe3hxexikGWKvYLVevoA4P4DcDX+9ebqNEma3
ZSphnGPs1+rBE43Q9/eOO4hT0igUEXSSnq+K1rJcCauYGMjZj1dQUFOit3xr7SHGtIIN1gJolBei
Pyx8OTFJDWHMhdnpdRAwoB7RyWDMRPoPvbGRpG/a/AUNEB9uxeCvr7PlqOwq2/d1GU2KHsDLogAF
hdSMZt8Mr+ofVtYQieTwcmrKHMdgZcitcuFrMmp7RgMEkwyix2aTYPdYQPeznz7vq9uoB1Olo75X
ltTYFJBB2UnKfXeZKR7srSKuEUFedYM/5TyDSOhIVLDRLXdHEFjqQ+XsoOlmBiGiYUSNvxFyLDIi
GaUDpFb3qdWfdvD0MorfLKdVuxcLSObpBSVLhxQIa6OAzt7U+HVlZkYglizNBYMKhrocoJOM7IJL
fAqcO1cNAWnSMkAN7v6DvkIp8YfCSGvZPKXivwS7jk1SpAI3Sz9pNsa0LoqskJvuDzBrAXB5NQn1
5xpGnsn6CmWepe2IjWIsHBgjuMnFqJFVy0Puw/omH/OXRhxdaFggLCkqhuQtdKIbrEiQH6jOXWTt
3hCHMnGNdBoxsQxldnDGKYWM6zU8MSIJifJnbLcSoU6TTzcIWEjK0AmxIy6D+VWPKrCbFnhplCTM
vM+/T6H7DY2Gs0gTD5NZfBvRQvdR62X8S/Fwb+BJXCKfEFCaAdHYQzQlPk1rmRIhduJR7jAW/UsT
Mu9QkLDeoYAR0Ty1xQncKhSYKSOa1SuPjV1prZU449FD3x5iNvppu6maQ3nZSLHVm9Dt1xEzePNC
j8HavbyWW89QboZakCqK42EkvOAle5ZGfT8OGzaCRMRzUX/2u0yyqmKmKWVtROkPWWFA09viz9X2
JQxa1uzju0ccFoxWGK6ODAyt2JIPLndARqDxEiRPGcwZGQOJF1RRGQwMUMSgRYIcytxF+WSn1Jzs
rkIvhhRt1DVgk25KzjkgvSWtcRLBWzc1RgP03impXjbBAvQk5QYWf00wYd0dFYugscW+Qnjjs2AN
ohaqVwUEz717vCDT7cdRqg5GkVbDoy7V+gNDvz93PZfIh99fBxWRgrWExP4RQNKC/ITU2k5vHAUq
9WgZLazXpe4Rr8fX8gX2lf2cxn4rTyWUx++JeJMwDIRmyUALd30LD6qq2SdoJaRUBDI1rZuDC3oM
Nzm+F0IuFgTbPWiaNxDIQOpjjjYHvqFvLMUBlVwVEkDEMasre9foz6UbPI7i6Hwr9KUIfqcAnazX
wv5QyMF0WxQuMd/3cPenevcnzfsgIu8KIBtt5uQZGOL1oXy1wkEAGEb4T9IPH6Trk22iWl3mP2bp
3lKrhdU+TonA0hIFLvG9G2XdQnB99960BRRTowhyTClnoPmhLoRh8HC0MdRLf8hqkEuB0rIGjg0Q
O996/Edj2risJZczaJvhoUgfVxzL3+z+96/KJsKAqAviQdTLLpQTWPvin1MdqdGJzQu35TO1IAO3
jVr1SKNOISY7ckLEX8CCz8sTn5UUqss5eBbnz1XFpwc04yfwbtndEqS4KL3NzhVPRja2YviavbZw
fe5N5mhW1iQ+JUIWJVxHpmacWZ0A5NzoDOh+cz+fjv16R8cOq37G1IXmRiV4RXuz0z5o8hS80mQG
3OGRzn/fxNc4b8TVYobQFHkj/6cIa8Mvgkr8+lWaqBmGhEooORKNLyDHKg0v2TBOx6YohudCIHF1
JencVYhQzza+M5ZrJl84VJt6xjnFsV2Z+4paAzVEHGolhIvOHUikpXQqUrc9gCvzK0Zbh9TZ7XmM
bj2gYTARqf5y3E1KyhvY6zwQ+gxVjIilvrzieOt0VkZ9ZS4rPXsX1Z3HwHSsNQ9/+lBgQ2e7ifKC
+NxV/hk7HJhi+Tu7JcjGqyTcRcy7M4H8uezBeG+j/hQdgmv1SDdUFcpncj7HAf2JVql5RlXvPI/x
zE36/kC7zQBJcVmPMjtiwKOTD+edvwa1Alk++9KBGtiKi+FyH4ibsjPh5Kx5FS5FFkRl/VK3jBBV
C8imTVhgxH7Egm3VZ1HR3pJmeud9GITwyPbjrtPWQMX/m4elDYLWnm/Zir1KX8RWp/eJZJu0/NxJ
V6FfFaAn8sCerAKrfw41GCcVLBeQtYY88buCIfz1vTFegldJndCQQlSH4yYtdiT3PIxJxBvSz6lV
nhdLlrLcPw5XG8A7HgGGu6kTajLLJFwZblybUv5FgzfoATvX4T2avnkThMDepfx6v2ywfqI2Pl/K
LlIeiAFGO51OcSJLbslfH4hzHX7E0KTipa4MQg0z1vhYjFpEzt6qcNd3bkqnEp2lLC6Uso0Q0xu8
S4Udwjcd4AsrQ2/jazZUxRmhi3iy0z3wQ3iNddaMGq8vkaya22ihmcRhiwlJ41nSgWs8tn2qdmVF
a6wQuJI6bdiUu/CpDkOxNleoE4JuOxbiqh2g2DOjzuMPVDtcqKSwf60It7bycxZvtpLTtVLYjGdm
vn0NDyqclvO1bwlljQ/z71ZnOr9gwoZEd91W492mLDPQs6hKEKjoj2Ahyy83IOzFY970E9CmhVWq
Tp7BLEyUolqkjMh7dBurhEYhv5l2Lt02n7d3FbwaFENk2iC7CsyptxjBcrc61XZcI9vaoWbVqPGr
u6pA3M6D8eDqir7CrO+z658AmKzOY4vLzZuGcnshZJboXI4XK9Zv+Etw7/xPEF564be309u+kmWV
88xyRYiPF6Wkw1YpYWHZvUOx5T7txQHRuCp6ggbWmehNEL/8RsyOUE1puuMAShifFfm2T9YJiFmp
GC3oQ8ENJ6X12QCVAmT2ITyYbRky8qoB/XZRcaPFZnR1lcz6sJQEGI0kHixFmrFRm4zWPu52FwlR
zRnNbsf4o/ShEeEnDGAcujEk7knj9iV6X+VHZExz+1cGibsjCAnZ13wEELtQ2BDygJandG6JHcLS
NOaMYv+ed2cFc942SrMoY4zsPVBj3GcD7YahXJ3nOXXM1R8Tqw/lLt92/pka3mtKYxEhgqFhwNxj
U2Eeg0sgBV8h10E4GAgQsJXrTMMYxrLXHkCxchU6DpCQQ3WjgemLZZawLS2ZWV7qNIzOQoA+2hJw
JN1ld/Mc2ZXObtviuuKOTx0NZuQUIseiykyUmpf2viHV9y7YdJri0RFWNkcJWW8yCUpO35o7F4ec
qqAEyVXRkfWANwya/FtwOL1fybHZevbM5Yrr6zA+ouHtB8hrFxVy9uGw5u46A/TuoHRObMnqwUFn
g2npsY9shwZL2rW562KdvO06kqtYt5bVtQKjudBQavfpIuqgsoVeJ/kPUxDU3MiVh4VlnQ0wFumr
WA7g2tFVdJwzuMEPDi0ajRFwSB1eBRocCfUQcRVxB14z1jA2V11C82ItNNMYoZuzJdSZY/DlWD49
MDXg56QvJDhpBeIv0TEK0hCIupbg98i8hfysm4+jveZaPaBnROLlY9+w13NKN5vAJBJ1eTUz5/pp
hO6wAko7iRBq1FcHEyrNYtZBEO1azvA/lnZ2UHWA5QcdLpU3sUbPf8mgBYmV7vZFC1bxgqmtYgzs
69+ZPBlIFCXGey0/5NmrE3MOh2Cvkzuw4o6HoEigP9F4jchLF8Z+8s6rrG1nR0ipQXc0JL3Q5wrO
/TzJXGd9WdlgxaT2MWIEsBNtXmnM3ThLLxGntMFPAWWXnQTXSPPXDvvEhSAehM5ufdXjodx0t1Ah
UjSKfCfibl18ROAS6WAE9Ptps7FhxvPyvGOgnBsvrHmB0d1sPWL4mHbZPmrfb/fxnu8EpqvD++dS
rWBHlZkL3iEJuZUK1LQK1xZV7ITSC5t9qqUkEWPRTxkVl6HVP2ZZ1JF9ZT4oNXFktn0qwWeIxlrn
Z1BFDz029LphC/5jStPsyY86XM6VL0zhSACvHlsC9sgsH5j4lzeEGAFVOKOz1tt9aeaZ5PDpAIdJ
twARv3fUrsNuDFLq6gBN5zLRuWwO9ZvENXBIV7zQqHcVVv1ecJU748Ev1M3pKirhI7JqPAlYz2Oi
JMTJLhWtUg3c2EEdKdHESb5roxAgA5eUwt9saU992CRD7MncbAIkTHKeJ9TNNuUwyQbxOcdYJhdL
jBtzPhS6vmmFoy79G9O89jUri+y69IEvZOYevCFP00BYg1QKylVgByymVImcpJSQ6NZ7YCure7kW
rzOt+jGQ75w2u413cBZ8f6EULgbLC1hvhJ/TpVkESkUIIU+665vSHd0vbXPjfvMrDhdi+7UP9zmB
nAdpvyB7JYRGF0qfpULJcYCZQfUMB3HixF74DSX5imUMiA1cqW9S8hzEYP0X/nN0rFW0C2PYPTQI
mHX7ymHjnqGfUlW6qALOfkFlq6RALam//63dusCjxBuCu26WjMEEIjJEwSSGxaA8pI6iS91e2KL0
8Dfc7EAXKkE4YiERyOmlTIjUDdVHCGsbQjZOm4iTbArJXTyfOigUxIxSo7rgNdrHydDNP8KN++Ng
3RukdWxQISbThOIM15nsdRpF0gcI9BBdCant7x/qnAxcp9xlk/3k2+OPi74RFbnUZDZ3yQ7eKnD5
F7uEa4igHI37V/vUIPOwjuN5EcG79L8wNcqOSmyEkXXLzfV4ZiRt7avS3lDVoH3GiqaobUb4t6CT
JzZ00zFDSVH1Kn5m7XGT/Huryui6sCDWWRt73nhJt2rkAfT0/zjATohHTRNxko9beH1U+pailzsp
3Y4thVYePfp0mzRlk63gTO16B18qLzxXScXfqdUb28midgP92ItxoygDW7mQ8Z10yDOByFlDoGGp
BQE12wmNWbp3ADoGgVgIBsG4tGlriyABBhSqJwP8iCQ9cmZ4UQNsbMby7jxL+orxY+na7mUvLn/1
rWlkUaFBbvT11WNa85y/9FRGAlKwXjX2q6Idi1BaKkrBVUwvM3/rnMtx17/8yTqh9I2C+ggD3t+u
cYOlvZEwFuLXBLqSt3WZJ+Zdwh4lFWz0Bn223sYhQbqU84EqaMB551vwCRUxnjfP+8Kwz8rvlY97
CZRkeavFAwAdYTkDxsT33G3H6qbGYNyMif/zSn2u0S6QjUTArJDYC2bMxAujQxFX+y2UasaqpCHx
OIwKhc2ZXyCfMeBXmxxOsOIo7eMr1EgPPvQXWZpYqcSbbcKfI8CvxEBv0DL3YQXNhau4+/+jTlNW
Np1/EJaO3C7cVMHmHM55B6hhMOkOrXRDp7LEjMtxhnZwit8zJQDSjvZtrjwtJLKgFPb5bvuxkTVz
kcBjuRxgYyroz+TLRfddV3IYysyZNZdgsqNlqpuOboQLdINeqq1hvQwYeUGRbQpOCVelmW4C6p+x
535iKuhXXtI/5yupLLIzAORS1eevQyvvfCX8jsAXOKno7ef8L8IcAozv6pwyDOZh33LLcP1rjtjd
9yDEXbwOVvxZZ/tsYFC/5hfgGNVoJrXtsW3diaKXd4DKfChHmQrqcq4i1fonFF8fldERoCjurTgX
fUOHffOjGG239vNbAwsl5uAFFl4jtQWTLAJ++mNeNSkQe67INBMxn58Odll8+AfyjCqlWPB7qiNK
co+Wr8uu22TNvYjz4wprDkrC5iPHmk3fhKxND2ueyDp1eE5IkwWbOsqNc1tZXRoIcheISaWaG6xV
xeTcp9ZiAaJq8O5flC0iL/qoIGloZl6N7Y+ScrWk/L37t3t8nnG1sw/d19b2KOkUWnMGrwprLGUg
f3e73tYzM7ER3N4kG9tTyWmnSx6xFnOC7tgQuwMNB89IB4cBd8QsqgMpVg5py7jx5sQYUFyQLMlc
yF12V9i4IXm+3Py6GQdMC8rtFIOEgj/Ize56EOJwLaLOe+xJa7wO4z6rT4XqZbDA47/aicyvdXWn
neCvy6NFS9fvZz0OUvclADHXoF3qD//e+lunJS7y8LS8Gk1hqAVnMT66y51Y2oDVXe1BgJOm292v
ETgibkhouq0PrvBYegH7mjbigCc7irP7So5m1+qwxZlAHWrH1rJIpe4qat59mqCAqU3hHSs9Insn
GPEF5TBYDbzyVMgwhWmLb/gVccVjdM1kDN1WZxVFQIswEHeGq8c5C81O1n5g+W/bmOh7QqMFqpd0
CDypZxwNH4ilFtwRNy/MSJDp48trINltp35nhlZHMAVCVkOS/h8gxn8uhsuO5p5GMaUKn/O55Z7R
gl7MUhxMsosNPPjxB5rIHEgTqC9q3MITkemjaxt3cllLAZp8rWk+H5er78d+VqI7UjFXSpMFkppc
oF1zf3Ys70P8vhlOqYlplilqpu+ekhLHQnNjUejM4BJkAgOCjrkkWnQgC9C4eOfHTaCpPG3nPVo/
YH9+m4VfzA4TbTk9HR09s/q0w5CjzVMdpvMhjEfV0+H/1CObVdGAPKFJ7WczAJkd75DRn2VvaBm4
Uxh2DhEvc9r1qxtlV6MDbERmlNsU+ZyG7SSHdWzdR/CYNl+mc0Nl3ZvI8qyc88C5fOcT2bB8U+HK
iMcuSiWYvYfKXIUsJO2FCdhL6D2uVi0GbLgcj/T+GiS9FnoPoJwNHEUeH4FVASESiY4LpU/zNaAp
KKZo/m6q/64NU9ZntWRLqngH2D6g9BQYHuq5J1MR6eNdSaiG5YiT9rhnntC7Fyk9Ca3MDAjHFMb7
r/9jBZ7C7K5I4qMc/WdbxUoo6C/TS1YHqe7U/X3rN73+mgMM+uLpCZ1DGc8rvd2Gbk6iEavBQ9Ob
eleBAfAQS1s1hyFbd+85Ew4dZ9whWDBxfNg2nZ0t7Pasq2V5McSJhJDz6QXQ223DLtIziW7B6jtC
AQggnUm7s+fIRCivDeDallYKcWxykQLNSiT5781S8QLR5SLaIK15Gdb8vpwHF5an5knuPisT12Fc
9WHjpkY/y7NGWDF8+IEhyVv6WB0adPwBKD96wxyIwbA/FIDPp16MFL0HRmm0ZHKZ+rjxq3KqNxCO
j21GeAMXQ1gRv7DhcwN2oFBbDgCrWchvAFuKRxLnfDZv+40x5HVyAOcEeGQZk+i5kvdVeV3YXfZE
+gxqnXUxkKpS9Sx55TJ+Ip29YyTtrMAjH7o9iRJKoTvtIGQKmEProvhl6ZytL4IZgNe+Nr6UgA37
u3nN1KN8wd8zzuWsHtzelNc/YH82PN1WumE0qnRyZcDyCj8bvAJrqvirhybctvkJK3uMV/f9o1dM
h1BMfFtv82Ebn1zQl9um2bluKFrP7LlsF3yNHklzpS2hBc5PgO1oZjMJFuKsI8eZjKpar8T2u5sr
c2c1/rGS3w6wbBajw2p8ikXThTEf5awkjXsx4fVU0AHM4fsnL5J1XHh45SY8fn2KSIpOp7j7Elm/
PqsvGI1zBGFEjcC4PKpMueywecRDj5NX8hDW7CF3FMGXW1yiQNU/3aGQS+mMQo1QZk3r8/qp8qlI
U/Y05/iAR6qDz6EeUhW/oZ9nm5/MePIGtZahGAp8O1iuTE9o2enZUB1+GQQVk0swXdSdcjr/VTFT
C6p6lUsUND/cA9K0OUNBfQjMmJH48UUOWqyn32xfiDvwJn7jPptmT1MPSYXdvHGaJvGc0AypvFCF
K0FxUMA1hn8d3Fie9cyJIu6Nc/oVNvDMd+COCd+rYhp/V3zXCZGEW+aWME7SXulelkUQg6XYlr9V
LVFcdhm7LGfsEyFOnwiLFRK6SAkwh8l60GAgQ2CH+LJLYeaJsoysIWM0HhrJ1LcKxZ/+efbS/zIw
MAAp6Llwh/9BrVydwCmH52vhyn29+XhwE17qjI/i/14BQdU4/oL8T/aRcO6q0bxecw4TlFnfz1fb
a1J7HrjgncA67k4OenheRAhmRX60XJS2eJ2cOYFSXy6e+69B1aLLFP4DJoiv7wsbqy4h6952c/QX
hgmHbi1pXkKoiIzAtSvH3R1l/BZEkQmKLpllvdP+fgBubmb63yt+f0vqtwgluay7jpkYuhuAb5n0
7vsme3zQPuvVwBSLqavPzHeuHQ2dwCRmUGc+JXWFZNELl03ZvPtv4fci50vAOfmhw1k1f7t9ENT/
8OTcaz3HbuVikJLqIlevTymjLj/embFXSEk0O7My6CMj1r0fBucI4qIMi2aFCUh20VIqVsgDMrLm
nppGE6vcjrGj1A3z+2Oj9tWztm0BebBxpbkUzc46OeoiZh8ER9bebkIwcUod38V/tOOxvVWe9qbd
RKzjPLP+YmoHNYSeGGWXH4YtGtcNc7i4hUQYCYwj/Une3ZZfihIKplQV/KyJbcUB0212GCsC73zL
9XIw2fynIeIqPrSVthdDutge6gwh8F8Xh5z+Fy4JFwzkcURcQ3FnKcQFAtO3AJvOaq2VOu0nNk22
kjaCd/oTykKpOEkrHeOxBPCgmL8WSLHlsVyJziyzCI0D9k5oqlClybL1i/+pRsFhHrk2OUkVJGWb
bIi4QS6UgNaiZX05iz/tt9T3X+BDDdd8kv6k7mla+XC/mBkZPiCsjphdBTRZt5blj0mSc8oydpRo
SbONV4dcOL4FkdVAkHQoyqpUnNjseJXvRS4wPKqXjcPGdTPgaMvfgqQaoRIFpI/ckATQsgbBpmwg
9FZiQYBx5GXtvD3oJIbVZiISgfDK3PXSIUEgIkdG0uIlPKpJfoqVb18FmSL4RyBg4/k28VlkIt+F
sWZQ6mD8pUTGl+kpYXe+4m+n2P/xKz7x02x9bYpiRUqVYGLtjfGcXvV1hwQCGN1dOkx05kLX7XSt
CXF+lzgRfLWz32EMKfX0ZpHVsqBtG1nMdCzfP8/luTeNO9fJm/ILWADJ3yeE3G0aEwuQ+2YX9drd
5bcNMvdvPZfXMNTyrqTEohy0cVxgAYjAh1W9aMSkJN16Q6MnvHej2C/BMYJejHDjMFL4VLWW4rPs
5bofnHfwLPa7pNoJYQlotQJhl3PaE5S9zNRdENoES33xEXfGCZt6GEk+3sx3IqJkTVowAPmTxC7Y
cwKTol6yL2QeaPxbVUNMk2h1waPBHHMEVa6/3dJE+DGBGK6GY9xJ06g5TZH6QLqKoVut7AFuayAR
DdWHtOqgC64zHST5q42gTkaON6lwq9esxwuOAuwpKPMKirhirlI3FuOPE49zekhzN8Atvq8jD4xN
oReW/ncTFET5kcBiXfA6e0xpIe45t1oHhFGIP8r/dxKN3mxpeqH3Afo/2DcUvusmuL0UBl5XiTSd
qx5dLqk5HbRFzbLJJnxcvRtlgJ9i5JxQRfgXFYGAvcammjxNz/2Xc6jZntzOY5G2YMwina0+3gyQ
54vifIoMC8ocPtEuHQkQVZ+x6qSKX2DYLjfsx1QTLHgq6uCh3y+GByQacJLT/q3YCrfgzaQUOz0c
Olsd2S6GcoKnyKWQxEdv3bJ5soXVUPooIt8WOD65sqvTuPhH7BX6OWJeUr0lyqYvUvVaEfxYTM3c
Dxrq8TQtKfUHYV+D+Ai5QFS4cEz7v5Hlab6f3I5HV5eLYX/tv673okuNQSD4ugbgjvfZD0W/9oXi
UZH1juWPVm/6ZjW44dxqDRC4b1hXlbmNG5jE+G8uY5ZSKt++lToDodvAq/ROpJsbXwszmzVFOQFn
Rsspa1xS3H4N8CxuZXwWj7jOHR/Q3ppUHDrOwZraBfVVs3pkNQXHUjO7wVVW4aV4S0OZ+HwwW62r
9zTWmBp4iBjDr55/6vC3ydn+qq80wsCuVAmF7Kx3Jv/6TCYnTEgxTj9LVbx5chP4XE6FfwUNBIgs
b7YK8aSGGSO+48o23YNMahbGlkSn5x1XCoVVeufgpWQQrbBE1YT4G9jf8y/yO0z4KA9CmLLHacF+
jm93Hlc5QEGRauoXa0WOBys9C3UmCDZ+65SxKQ+NlyKGUL49vZQVpMz2GZUdI+++ZDdh23/OLF4c
oiAFKPM4EtLRokzUDjs29A2oQzJkyh4SBTF+YYx4zs/vmRIXyg7gAVoye/3nD/n+h9PzJl04OqRF
U/3h0FJBBfSb1zQbi3TCWFsX3tSkzxDfkPsB1+Eji2EtlzATvlhol00daDWHnVSwRpB1ibz1EAtI
qiuJtAzlFBNZ50MHLcqgoT1NKjhES5zvhj37eenGkU8oS0WZseg1iALgVs1mpCxufAVdzUu8AnEL
v/nwXw85MOqj57n2hTULll3BfE2pLRJXnJ2M/Wm/l+I1QjFfP0NcUt8gmOj3dFn7q1HwIJ4rpy7C
Pfax4bNOnVRpFIBgHq3yCYs04iQs+9JfO7qQ3opx22RocOHYv3UYZQeyHPLlzdA5pCH9oKt3+B3+
0bZl3ZqfOxno2N+L2QHpIF7P7+F+rBNWSicpvgPWXt4PN4pT6TxBiked35VjG6LajU2o+ZNQJYUW
kuvY0konI/l3lFKUSfiPYj8X7+cRWv0TXsBh/kIIjWVatTVTMYHWa9zMWf2QoiGehEFn8WVdvk3k
NBQ0hZiBaSucV1zJTykV8G9UkgvSYLnexk6lBmrNg5bxJsM3Ha40XUaMIDcgfj9HByyBm2B5H353
PWmOvZbQrPcuN/ubBNrTNWLGgJuV1MoNfo7gMqN8tqpA4pk0q0et4b9VC0TH6Q0+iZdpIblTVn99
hcs6Zby5gQubPdBSAISueHK+S7b6mg0Q8h2vVZYK8UtG3UIVntzVL0tyZ3i0gJVlZR1RhZxy57XG
feTnLUQMZjfs2KkTbmPkIDEawTUCwYshjeo7vOpGMc7ZEeTwu3bNnhY0FUE8GHPduPbUt51MA10u
B7H+PthPMJtbJhsRQEypsxJqmttfRLGvZCb40NL6fAzBvfV/wRdGYGMTAGkk53fZmZlCgsrAemSu
JfeYTMFZwQ63VI7oqkpzOW6+owt66dgyOC4K80lwNT040isEolT7+7ziiqmtkWjMvRCHx3wNqGbE
okGI2Q0R3sjj0kn/6pTc4oaPNyPIirJw7jwrWGMFkgtLewz1qJKKbYgv0KTMtgoskTrpfChZVciR
95Fddl2eAQn7reDibd7DhyJExjzuiZw9eSTX323obPlNvOxAxFBvJVAu+lJmX1DMOa9Rk96Z6wCr
6u3G2SBB6WxW/AUsXIMardwOcq+2QsaM6s+giEaMEQUyIgbqC7i0RiKH3hIXrGQeVrQgmdQYkyrg
VovvamLX7MmF/TJ7AeS/tMBzbL+GA81U2tQD7GbvZw1AoTwEeLTtlArkgo/s3oVyvelZfApseX84
txOCz9vAwh/ac84iNjF8DjkX5x9rPSlUcES6BZgHUQQZRgyQ18bIoPE8ND+Hdpp6kgDxiwvYWf9U
gw/IU3dtF1HkXqHps5YsRRRJ2ucpHLC/EqaIJ91VP+ypnsklOcf0CrVMOoRvZg+JZYVdaPWqRpv4
c3BOgHKzQY1GdzPY4M2N8NhtX+RWlkMYzwjte7ln/0adoBKWKgsnksDK8RXztPqBfaiaZCjD6fj6
3g4i3DsBuPekrIgxR6dTwCnzxsGcW7gVhaHz9KCvHOB+TRzTL03X0PtOc9d0pgHBiZKXRA5xna8r
5HndPr7TSAJj/bM2p5l1nl8aZCRdikQKSnpcB0ZJUEaxcpHlv0+4PescSw3z3FZkDfuazw9gGX0e
YPulVsAtor/ojazIC1Yb9Lh6RxtC1v8B1hkfyC48lPzmBuV0Aw8sHGcNzc7FjaEejuMQhlj0efnp
iWoBgC4OsNB1ocmSZFgywzEosUuoUWAenNTh1Bs4XXgwNoPOhkB1dht04Cr9A+Y+voFOPG+vlTHe
z8tt23RBE088oVN4Zv8L7P4NRf/bmNl+u+vOzd4L+Yf+FiWjMVvITXDGglZGcow1tAFnRyNnGU92
3gFJC/TSwLnX1Jd35tszrFwdQ76hgON1QFZPmIguibfDi3DlDkCqFnNT3k7D2EV8GsZS2di7odQn
jldXXJYcpjRb9vFDb3wWiGVcU+5Tl843+9WfcAJx6zy/LpR95n0ySGQZeeuRaJBUtvmvQQWBQAR7
IBXJaDLb1JskkBwzMB+XL2dk8UshwfqChWlYqFYdgqBYKlCSYUNPff1ns69+v+qQxeE/+9jDfYnK
FIgyyjFQQnQZ8xDFyv3duJf2n0cNxNgygpJJe/TxF0CyfI6XORerczXVv5ECDCzPM/hCeFZJjt7a
Yarq/msVz/FuMfnwmSuzsFUXi6kR7umI6A0y1yc7mtjhzq2QQou2OD/BcKcCjBUqZtwiuNYg1nUY
NyAARlFsFFTRI5N5azvUuP3ydbRki8yedTDuFz1ccrMcBgiy/av/B4w4IiYQAnbGTjAWKYxOU8Ai
riI+EIfAN3uCs9qlwCtjTwov1ndwFZFY1HvECW8AS9NOkvCnsPmjoAygpLphBUR0YfI9ONM8moR6
IjiG1XAbmuBFh22VDpFcuclFOKR0qhOLpxUc9Yjw9cfXPHTvQ/fmFUlV4S8OCeTm5U54b1MWtQKt
9P/4pxilfAv3WK1rnFZiroMDQxK3Fi51e3Y6FAbTyTzvvTVdL94SudKm+jC0UtPYxNTnUBWhADHg
Kl8Wyzl7+FHmbS+Z5/UOsfKgz7Go/3BtXHqwR9hB5YgNTEruDpAKXP9IYOXqS9aAnelJ3DtTrARQ
RswbshoUasgiONgkVixMqGFWKTS4TtbfSZAmbhetA3GaI0+/ztSj6tUF1HQPrSQkVkWXmbDcslTw
3eFnZGQBrej32zxD1detK1hJ8kBfpNRR77eJ/iDc7sW1Cs4b5zYFFrC8Yhm0wEPzIIYVAg9pSSc3
gDQREOmzGtqSE8ej5HXUVO2Ehpnvy4FkMHGIknBaT7ILZOI/yxOIOxf1U+uaMwPMGIcy9G/4LG+5
74N2cXSBgV+3dvRNeQla2wquozXDDfI14FSDOPUPBwL0Mh4tHyLuIpRJHEumYYN5QQzT9y7IXgUC
Bpeu8TSJWoweG8+UfnS1Oi0H4wF6iSnwYV0LnIYrPS3hFOnt89YuPukW9Y6MXMZC2YAy5MooU0dX
YIxS1hE0JdtO9QwSOZjJfM31crnsmbKKARmOvZLW4xOUbCgeDRJB+k3eXRnogkbgrc6NQ159RMTs
Vobj3y1smrehZWd1SFiqNeIpJQYL672i2PMMPMlZIdfaGIE5USRUKWAscnhH1ZKeuhXdqPQvmKuH
R/rWx1iTaP+3Tr+bdsx31i+suDJF4t8y68szvk44dOWGrOl+LgVzSWXwXZDnComH5XsuN3llu4QX
JieoZAtqEnQ6rNG1Z0wcYThberP9oyW9m/Yj6fJhUdYTbu8IVqNB9XzfvOo4UNQb/tA0QEMj8LM9
pFky3YC+MEWjeME2EbvwiK4xdWRyF/yYyhyUgCG4ykCEG9wk3Ow90NUUJ1+0F1H4KOBgtuFNJtpZ
gMW598MmTRPysjdnetb6r2rptRtNm6jnKVoL7yWb489+nSOzWFg3g/TQvXekAg1mpnXZtHY+QloO
r1MGpQv9ZH3Szet5F7d750/lDf1z8oN1+QLw7v23dWZ4OLqitftvVXH0/7O3AA/zTUeNpbmUz8o2
l6p1h7AgCyEoj1NJuEadB3yVW4ag6SLGYfZUvUwjx6e7rBw2nh9uYcQTKQ0YTi6cipOZS7wYSfXZ
Pj239CTKyICBToZ125/5yWLFOsUVnFTTo6Wi5MF0JbQbc21ImKf7QL1sE/ClEiMW1GnC1/Azaxn+
izoHjKC0AbHXarzmQ6dnY2fp3MphKqZAxdcNMz6wj8oPKvC/dHwO+dvkA7l6d0L6kSKZsDBsMRNM
xuQKfyoKjKkEh7KTVdwecUrIZbU6AOsjeuDG5nBevp147sUc7T6Nz9FEndSlXSWdQhj3dGk7EPMC
q9cToS8A4oRG0RZM4tBv6QpvCPbj1ycU0qiQ4uAZDM5RkUicV3B27G0PBk1d6xCa5KOdWeeP7Jjr
kQp/8DbW2KioUH+/UFKOw1WMRHOAKW4GCvb6ekw1XjtmlQehol6GOw+NY7fke5gt9W7DCVDI8Pto
IObryR/qpsAeF4Cz97fYhhsAajQUgjzewvksemUZ3jkiRx7t1GdHNwVCA3TKLE9mXwPNahmj2dfF
QEv+gvHfkMIQlh+zdBCiJM4DJMQ7DBX6BSIh7j/cn3qM4/x/dEJlPIFFqvzrXqo0+xo4ICOKDkvd
cfchDkFhmiJmBXPre+JAJJJSWtZjrEVkzqugyQSjcN+sgHdCD4hxwtMzJwi3NUfajrJYqnA7rLbq
ZX3RRDcr5wZp0xCS6Nre+se3/m31/Oz7dtLM/Kf7tDkbJLwvHVPbWU+YYsHaXH7CZBaHTNK/4ll8
MRE/fxK/DW6GrKbTLRl5SGqatQeWB2k7MxAQ4FwSsZy1sIIXAxhJbtZrTFwe3aEC65GATMbFGSRb
0ZuCW2rAj3v3uCYT7SX3ru+KXtEZSMQ1Z/VsPYVPtvFJRYo0uWVnQ6dD3yybY5v6U7uSEKChmGB4
tAC2i+h/b4zB2/+21BOiTWJmPLLRw0Np1vYY0M1S+HuzyKOzISajxb8YXrETtSAjlkfL15Nq+EvH
XgtxodXk7S0NUyLl4uXHvblv6k/R2mGk3BKAw60evKmvgae7489XrmXaTe6m05zjZxR3kjxFwRXr
TWkjuPlfVMWF2YR1hHJVUto3/CWEk61X7mZ8Saq+RJei02xzUlrCFaEF3RarBVH78Bh5kHSLaUr4
M+kZHomX+TR4THJgQ/XlYqyFUtz2niIRkc1uaLxki1/aA70OAPPKYw5tYFFQmuRzcaleh+mpd6Vs
KQzz3Aqabfv8vTnWELst+6977ijXzNyW3OnJ6dQ6ycgTqxAE6bnPe3FFq6hbQAi3hOqASnoKch9X
o9Q/dMZO6SoaCar1jwr9WP2sogZlH4uijjvcZgYs6TaH05cGFMOVjEbtXukXhTadbUMHBQibcaJC
tUKlVwpLyx9fVVglbsEpBt941AHFwiS92T8fBZYSMKa3gXRQfeE/Xa6gguy33RzJ78r4kOTWjBsa
6wlir685mbnfKrs6no63gXAijrxoCysaxdcBq7Cm+UGpj7GESocIhfVYQyRnZEH+EuiXIgfvD8dl
mC7IFmpQYvn6aHgfE/S0Jq/yq7IAw1IHbnYVO0zZiY2SlZZv895y9laST75xzSeqmX4/LGby2CIH
usi3Gk3a512EnorPDaZyJFw8JD20tZVgp2ghCS5h6CH0g3idSvL3BsYWScL8n+R89o4fXWjkv6CP
UYFrx61e5DzF6CY9UOX6X65GpWkNqAZeU3NGDgUFNVEMR5NuSbhd7ej9VXOpywPKVFjAPBtCMxLj
1o3dHGAiHtzss5kSc+8MDZHeLFMnEMkkNK6hlKIBDqk9mDK4tLqP2KF47wHIR0QyJhdb2a84Zfnj
oZK+ygup/b6fZI0YyyVzrD6BDvJyiPy4hK/1CDul8md0KCQS5Enn7IQtfe2e6TfKs4XAgNW+KLA3
JzhODZYVy1P+uncDgoOb4eIYNE0SxTSZdSg++gWDIym/ruO1GX+wlB2VVmg6DvdVjrpzmEYiY1is
JXPbBbsHnnEcNfdvhwcMLw6fJjHyiKyGoRIDImNNPgLYe18P+PWc+GmFnvqu3sW2k/VqhpGnPlDu
08M6rWRT8zmunT+ma6fIM/D+8cY5Wca5/8PqVlgwlbS2q4nmOGmzv2DEM7sifOGqA1cWgM0wLcbE
3cVEm8SHNhrVy9slwzvhbHIZSkZBrmWCjx+1YE3bxrRMz0U48rth3NJ46RhjSVeJH6fa9V1IRcOZ
Wf6MouJ8E4l0RsCv9Yuvg8F7NDrNzHfzbnJ6jhHlA11ZGFpjGniy/h24PHRNChWMwIwgX5vcqhlQ
DN9fFGuTYJ+y67wzTvo3eOJPhq0Pxt6IKRn/26FhlqJoCaTvoFXwsdh/cNjKCGwUhhB1r3+lDKNM
BNGbpoysGPzBGwTYsJuFSVw9d3K0RWgKKixnDFB+dfIJuCfbFacDMcY/S3H7RIWuflPIcg7fIvSZ
u+rYCjtKNkw38l91FvAGqOQO4Zd0x8QM7Lka/mDkNmkcD37mOywlThYUQdBHdFMxJG1rH2b7TtHi
3qPLL5YABFb1yhfx/PFdsHBIolKfRN8ygRrbTr+SuzNVu6UpMT70SEevsixlMwZRbjhbQ8r/zyKr
elwVqlpRbQeoSvpFOdD4Usj4ltwoZ2dUPkPohPB7tc+Qn7iXDlTEH57f8PXUIe7LhYABThqYc30o
MZIDoHDwigM8tjQTPDf9b/CDFxgTKIDe5vfwpRjyoozfgjSnAn6Ds34zB3ABMfGgM0d+1fLByo2R
efD4HNwiQE0zjpxjTjHujZ4JuTtZsIJEG/HgeoY91/yOyXsnhbJrsp+nUQZKDefJxfDYjWB6PqVA
ts9+WabbfAz/+JBGm7/C4/clY3YaBleTZBG9nbrg2msT2Ltj07c+fLNeufca6XIRwpgKdht6Wj3A
gkxlH47EO/CkH3m+gdbYbvqGohJnviTXJlqOdvYlLMslrfaR01ohySMAzkGx3PfPpSAEBx4DU02x
FIALJayJfATV106sfDzsI1r4utKtsyz+o5W2QHeRV5Wm7tjzWbAm9it602g5Vt49MeQ8xjEVxBX6
9gRI5bMYti/l1NtlA63LccNX83E61P1+S9qGGuNk5xfp6LDYSschYxndwbtsTvvZLM74Gs8L+shL
vYuvQs00CoptX87G4MiMIFJtWJ0wosRGR4rE1g4oNQFUNDW26g7A/ITloELVOcXpPjVNnL27cHnT
+0pffZem7y3izLzcK0jWJGu6xB8LfADlS0Uxx7FtpeztP4DpneAIRrwtrezyvuQ2S29aPD1PsoMj
JUX8gSiYyCT+bel1+4P8aR5fJUS5ZwdeN9IbpkYzzzO23X2dusA23kzW2Dzou80duhdtnWDXBG7m
/c0QUGhzuubrdcbahAAd+4HMBvzjpUtAYR7qNjZP1FE1BYoEBAKbn5EDaiQScJuYOIVp7b67yT2M
cUtPiUEksBJxpWe0NM2nTFBGdV00Y43NIPkBt9NOYrO96Tqvz3QV9B74erHBHipz36Ii1Rnv9n7l
yg769wCG+ioYoZvM1dpKDTgrL9Vk89pMLEd7itFC021FLq6P4AuCVvV3rHvCBU4Ar2YVPK8Q4MGa
6Ap1gGzaqpNMn68n6HAKLpMhGK7Py+XTV9Gpa9L+oMU1eDdLvRzl5uNPsF3HbYDG95okRT5xr1Vx
NLw36mGcc5vFvX/qSyEnxWLKLEdpfvyt7RkMSPPu4ulUERqFBcUlW8syopW5p59bdoo1Qp5zfESW
BT+vbM6O6XaMVYU5x3Mec1hqIDaE24dA7TMH7vB5lbPWvK81Jq5SVk0sI80og94pUOPdsvfwqOF6
UDbE+Pb19rFjTbcfsZa0uIOg5Rr/ZIeJwBD7smzHFERvHG0QLhtHYwzamuKLyusxll0ZOzsZ55SY
tCbVSLwMtCGSNbCHBr/tSuAObQcZDKG6CCaN8749xwL01V0A88bnVZRtZOhtZKjzYDN3owycqhsy
myLQBPo0sniepmqKgxz/HSYywETKinF0+iLBy2U8JJ+nFva6polnjhTGlqExO/GFzMR5TsrObJ8j
s13QTvhKG51mYUoESraySITQglzpyxYeW8z3dv+xN07l0WoW43w3fDK6wdiXWzxIYY4XIM+HvaI8
D19WfQc3GVTbhK+usruAuX2pmboixTywmeR5VoxA2wOqvIZsp0DRr4JlvrbCrTjhZvHkSgig6gvC
xe3Skea/Ofl4aU8kUCgFcL88+mszMFbQrY2uF0lzuwLo3rT5jRef9b9iJO0ZAzqr3MqsrVSP7jNx
vf1mUTtKpzbWYruCJSlkS756D+kLxNBFNKCxo+qXgrg0B5ImsK3WKA9H7Kl6PU6aP0hqMSYbYwMa
OLGaVPHm9vLz2vIqwPg9BlcYDQbcJ+Jo/Qf2O99RMUB6PGsocNOgrx/TsiLuQEyW1hQBiB/KG1Yk
F5OJhB2DLL8yVjMY+bLrBdnlrUJW4uyZnIWVDQHBQ0IaLxJEL4d28ZjBWTtsoXOvEJqu+7jPUEtf
U+gaGjGJ+4SQJ9Rs0h0+u38pp5de2qWCi17ZooK8j47hLbB3SvwJVBLZveQm092NZsmRwzRCmwLG
sZ5nAm1PIlSvX4EeOBElg3sOJPLKSgbacLDim5iKCJzr/XKVOUrPfKWbSFymxmlKCKMZKgfm5Jha
v7z/VUL6hWk/1S09rizcsZDPWzBs4RxYyaopbQEjnytPD5Ubl3Ta6KRsWN5GOgIb9cHFLL/9w2Os
5Ku2kCesUEY+RvF9bQX1BIMRJ94iMgYsTpKQRrMANdnAPlpYsn7zdQSP1U79/wXI9uOIgE1id5P1
EwAz1uTyo8py8C2XES0QCSOnpRAaxbDEyG7jFv8ST0SKPPBz6uqJjQ9ehFSO69D2dXMp81oY7gBB
W1TlY8CdJYXPxnO1wVHu29rzXDyoDmwzIAKBP9YC21TeJU5i6M8IJdEb1vKbF1BjxOz0RVArdklg
hgzmKpvT+avc+YNpl+youY1kCYKKsQAUG/4+voQ4mmWuzJU/t4O2L3vh14lKfwsNqYf2lHFVBE/t
ieMRXbcTQxsm1HZAsiCv9rUrCzYAfE8DB0W9ip4iPfhsch/ey+mqQdMTDuLni5/yc1H3tl6M2wCA
prXYqWGptlJ+fb46JYjQP6yaKAMLbPSlSo6/aFcvpXaW5kVbyxEO2OxGhxk+en0/ooPfLrE4XujG
IWvXlK4vnbjHbVvIp3FCzEL8n6PjAVu0dHPleGfaB1kYF9UWrRhJ4mbjAlIqgYYocgVHHjLbq6Fh
e3AkyFsfwMaCXa3w4KuFjAbiorU3QsHxwnQmiNzA5f/8CwbYHVE6rO4v3h5yCDuXmEVkUyGsH3tP
UaZxdyOK572JZgmpccYyADN41d451soXOYU/iOJCeFi7mTvxEOC2KmPRIIrJnhYcU7txkGkLuxTL
jIMMOlESA1vk9ZdMpyd4LcQh76gCF9g3rXa3UAe2+/6eEICzthJGsfHb2m9p//1iqeXrm814F5Mz
2RH+v5vfbRd8VVNPWd8dQuAhHyH+8HdLfTqI4u4A0gS7flnyVNw2G5hqHSHVtzMWQccbTkF8ZDz4
xXSqYc7sVrmUtbICep9iAO5TqTtIjjQXQXLso6wvY91hzUwAxTQysFnAH3MzVFHY4wnrxjnx1cHX
gfn5ZwKMrV1jmUIHcOpP5j/Ua2DpdWt80X09gf2KNT/2Y6W8fI/P1nxv1lJoPTDy2ao/hRC3WGq1
PWnXRIw5ubPJnFdfbEmp1cKcMZlxHKdl4c+axN13RwdmVIXXdIPVLIZMKYng0F81IVKqMqjtN0z1
r2pdPeNDahTUgtfOc0005Rx5ftscjgPlNJzhEU3DJZet5HGbj++wmJKW8SpA+aZIm5iZ374OArSm
kvySLPRb7UqhMQRh2Kl/fr4NjVkHgxW8R4PVGPHJohmfbDtXKLdTjzxatElm6HLJmJrQSQehO+Pi
XtPhskCqPolNSpbSbcz85UBS7mQUHBet/Vx1KqekpLhW4UPfee8S5bkMXEO7HRzvoyvh6ZmdEYFq
I6UEDEiTwKL+HZqRN8Fj8cPzhE6TdE5TKIk2PBiayx7TCzYOse1hOjGmo0nul5aG7DYfZ+XuQXok
GwQje/G6rd9aRoTJjeQ93/HWPP+Vc7UtktRSBJaLPq/2HKi+UPYZ/j4k2gb18u2XYlV3ababHcDB
YUMWBBdCSPUDHLCT8+Aksx9QLbUMS4TPF9kQt9u0MI45R46K3XAVYO6KDEAMqkbPH72PQ3bl6ILn
+Rc5/s8xhGrmZaZAAm37BS4dpa9euBKtS0F9RmGCC7mRtPsrsJJruyMJ/EfSk3S4DynGlePo08Ar
e7zN2IllJnX4QGQZeFw05C5z5QdEvRisMYslekYqRodbLiJ+Zjk74O6j9OpWjYLwWbgq1mEB+C9B
xHUv0Vt9CkgPaa5g5T/aBCD1AIvG0gevB15YuoDB4SDofDzJ1+NZQULelRpFy9AX8ri8ki/zuN+3
1E6H59ZPpZ/y31799UWxoqzhNQyTWbZPGBCMrUPbWx3P56Qnbx4l12nuLJtBitGhYQyTB01qr80/
FEpLZGcIxvSzTw+35B9PQcuHc8vavIiufZCFc1uYakKjwSCWPh2ewpY2eOkO17+gJ/oQHZKUQw3R
rajKB50db5H8Dqi/iQgZ86NXmrmUzV/ZWhiwTS1FAPgZ9hnDKoS2xDmQGVbkgx6rktriWBByLEAA
G7ATyD+Adv4arMr0PMM5gU20qU7I0yzVSGV2jJ2tDvujsswR52vCz6MYPha5UXXcsVNfyyN8YwNt
ABOCwpiCQkFz+sbP67BQe3cmWMgRngt91Roppzra1XnOG4lriHJcjnZ11QK4boZ5tAvh5s0EkQi9
RL0kmMs7Uc18oYjHGqiZ4hKhUdBKmbM+z9iVOWwCp8ewTFCxDPTfBL+bemqLnAf50c6qTDqPylOO
KB6an5NjBpinKCAMSEDZaS99DmXYPOHcrtiGYo8DjHUBEF4Ack0rb2WyMManqgMK/S7PoL0VjUON
dv0im7Tw9MFIaGnmUifamVPVbMCqXAH9NTJuGizr3fl4GATTNbgPdTWMfesM6IsNV9Uf84mdmNqG
8xVfNxg+lDs8GYwMwA/WS07ikzEOfQq/r8jxYtuH8jfSFyK/mEcuXKujgCiV2XGxN4q8NlHK2M0e
/mX8VaesAg2MyuaOwwKwq5zyog2XZoroio+N2h6l+Qj54NKonnzGw4Kn9WyWyCa7whK2uSH+hjLE
Y8XbCkpnonDWYV2uXj8regOPNDznwzxNkFYMx5PzrjiNeZwIrQPdfMZDPZkcwih6PJ4wiv5AsUwg
BtLasLuUWoVU0+877OoUk2kogw3A8Vxj2bEXInOzBttLRr+Km7zabS3p+DQK52W4RBMT0njJZbsv
QfiPE1G3DDaluINgaMcIOiMOIMHONEOt8Ev3eaPRSXBGf6gJc6Zw3vh3Zpz4VWOcrWasEq3VJUZm
/VXgaIDA5INcHhvit/DFCoB0X9mW6rsOeCWuzjQ1vFHxvz0MgNnGk6nJPqmWEKTpaZr5NMNdREwu
iHec2JcOmWullZbUUZU9aAH9j/sdbPTyNEBGv3YV/V1o18nOUDWh0F2iQONZhBSnPieydR5yItoU
u6N2YeAamxn+ksfZww0po2qkGwdbvfdAWxDE2CrGufMKNqV73beXETvnn8ezVRJdkm/cgIvxTK38
XmpEz4uJ1C/ROr9zJFtA9JOLgxnNOCbv7budo4Sk1N0bPPQ9YqUo0/rrinv1cMQdXPSLXJbXVhr2
+dlsMnaQ30fAZ6hV9tpEytLu/6RcIloOwRHs0YCc7YkoSPDSuzBT0xv0AwdT1j0UFM12ugWYBrMT
ADIgqk3x9dDElCR4VQ5ndUvfjfecHJm4RrDi66nxo0vfQ4QMF5W7Bmjm/5zKJsFfVEVMnIVnQcQu
UOvVIAV/UDsp7S0h+dVW5bw0HR77+MqvGT4K0bIYzLUbrWbFxKPphgDbXDxwGU8m/EE8kkFNOdnw
YO51wsnEv1+sbnyM6tnsZ/uhrvyQLq+r7qoeT5ZihkIGbRwIcnXEB43Fk68z7Cl87xsTVzfRGSXG
1IcHP8MeNLYaDGXkWjGmaXG1N7woDOVR+q504rDuWJfh9CzmECaz7bjL9malYV9QRiGKTFgO08UP
MaBf/SbcDD3X1rToekUxgKx1lYxE8R5ARX8VmchaQ7Lr4S6RpwNq/R4YUqljNzJEQYKnWFzQpXBb
WN1KAKz+rSfMOE9SqRWWX5LNyfdvyTPD/MYNnhVDYfXj02jjxHItUJJfd/69MT03vuN6EmSzo45P
g0Xy/N20Sc+9n6m0Cb6thnaqjNkoT9lY8G6uTLYiXsbFurZsFE6p6PiYEAXyWRFPsUYZtAA5DHYd
P89TJnqsJjFoQkl2nSNxpe8tBpmpuCrJwkobcRFefX5F1/DQs9o9N22QjHfKIbYsJnUTPTE4e6aH
ST//mApGLtkwjMJHvWJKUHuT2ZFMt6vcjzGBZ2qBhWqzEzXKtgmATa4WPxLLHhqM22p7qjsR+A1b
6X9klx1Gfn64y0fzA9j+fimWKgUAushUqPGuH5Yjc4oaJDuqHuRrKQAuEQCylunDtGPxdBeycEvh
gBDF3wnPeghoROf0cPHjzevNfsLax0zsVwviAzy5yrRes4kvIIdbt10asrdCoKfzIZVEaqqdu114
kMDZte8p8+X2VkRQLHnBfKD272H0kEwxPtbIg9s+sXNEKRN0Jkxb56PdIQvN86g9Ol7XU0pOAxWm
uY02Tg487Ap06otvsyrxNElxZNmkCNcMqXJfYoj/H2wunXLF6XaOpf53aLAHAq2HvZUo6KMfRB05
1ATbgH9eFWxmyceByzpt1oxBBrbeJy9iNbu7NGPUi4mbTaK8FausS6XIz95waio6zb7313b7SU8s
OXTDaijFnaJPBBsINHb9B2jpSjV5/yVLsKNEiPjb/8vaPCqnkN8FMP1bUJ/srY7X0EiJsMVm+CdO
GCckDZD5v5ZA/BdnSdGbHNDegkEJW6jWBNQWsatlKwCiW2X4/0jjlGyoNDuDPnTDH2Ant0MqePSS
tMvTeA5qD31HJXiN70pjGvAtaozxYS8K9BMNtjbZ8eKW/4Gum/Z1VDB1RBIgquN4iRMdSRxaqHiI
QrI6IhEznUzc2R0WcJnYd8GoyvEa7yZuW4ZoJyl18SmbmDWtqS6f45HWk4SuM0pUw3ma6UN+eyZt
SW6NlI9Lyyd4ASyFSzYK8Mq7BZX8esC0HJ7Uyug4cZ+TsT8sYSAGz3AtXlccPvHX/VkqsTY/338O
VqZWXOBY61jgR2D8kUPvlifbYtpXFEfnn4fZpzA1By4+uS38sJLq5S4Tv5I6eaRpS9P903y4dgi6
FUQKuq+8dip7k23K1mY7iq4bzL2TWvJgwWtTZRyaP3le1CCiYlKlBPrlBANLkiGleaJjw0czi2+I
nNAVN/5LwQYLCyXrCYQxRfyhMWGq5HSTdB02IB0XOFtoKobaPyb5+Rz2QdvmJse1E/Rr5eXIDZet
Tty/huDE2YqoEJuMM/CA6BKnadvW0I7w5AGqvDPLn95z7DYT/+lmEhnRxAy6KG4bpleqhOnyxjFV
yuZlHMYIStPIuhyyZAhRU+VtWQIcN5J33XCF6B95+t4UntblEIhB/mCl7jZrV3Hq6nJC723KILb1
wvHJ7MYSH9dLbuIg50zRObwZ1OHfMm8mo78aPX/QkjPBCAVZnvP1/Lp5bgfCCxvxKVDVaixh1OmI
EVi8MkDsxQEfWiQNRAsJWEV7OSumBT86GhgC8rmZR5H1gOcTSYqBsMM3a5F8n1Qql6BoOeOMWl3C
rz22xAUad4l3+/jDCKny5fJwgN2X4aZo8QL7ywPtnEYgxAW5Qqm/rSnUVcdZGP8o3Fvxqe5KVNHt
6kedoUCVgjp5vmSVDVb9LeM5Da1q+aaZn1mfgtYmen/8VofXUtTquVJHI85G76w499I5qaLxwQ+Q
vWnk0dEzHPw/E6YcbS7N8cBkelDsmP0yWGUYM5gF8KIXO669RIBSgP7A3oxLuuTKyS8nHZo3O4XU
gkdTSf76ZjB4XBAuFrjWclZ416huaBQp6flneKYnB5R6oqXE76fP4l9diCq1cSOVlMnRrKD2u/UI
vl7rq2+Pkb1EKvc2GW2tchEWGGllf/UCOIA2XjnPg6KVwh71rMOdAUl0AhQ85IBjf/ETaSVbx53y
K48iIJY6TlqiQz3y/ED/mkgef6Jo/2ABVwmFE0iweJhH5kGbWnaCTLwmI9Ng0VXjA8/ON3ye4Xv/
hxQQiMuS+qOBTG0oHIR0j4eRjQGZxYuFRM/KGs6oaI9mnIxlHCz6U+2fvFhldszCwdoj2eswGro2
xHF4v2s2jWFJvFHj2tKnrp7pCNZMRlq1uCXXL2UmWlCpgH5AN/EkgprQ2aqiJLUsE1VEDFVeLlT9
eXjWfa3htGkZGFJku32hV+BJbxXHlM37vhfFVwL6NR0JGpC4HWPdEd8z8aA9h4jF3dMhP2ThZIMi
rBoFd8kgIO/p+1Fd6SZGiXF0vS7+nRwN/cN28euSh7/tO02QbUf9lh5j0CsEHwQDkFCUAeRcvxR2
XdsPPGnY62HhnfDVza4rX37dTiVOH5EDtucEBVJMsH0aGhUuIbBlAuNLNUYaDDzMh25jJzfYxbfs
wlW3aOiEyD78avUzgr1uJpu1pdjHtscZg4v3vOkxFL4my65DvneOM6NveS3u82chakKegu4jMMvr
kLQ3pWv8P0iPFHpcCYIFmiVzFWpsZKU3QncJ4SslKI9z1H6MmBVXzA6tm8QFFPP/jFmVqPfsaLGI
JzTiSUSM6tICdTU3IqBTML4lmJrOfItTPUajzFBcfGaVqtkQl5MWQsC4LbtAFoDjpO7PKNUA/Fnm
+gMqvuKst9T/R4RiOn9h7R5+yqsqNESkRYsTvnyb3nym/HUk1K4UEvBBJdY6t7ulgDasIcaMEFIg
S+Zxo/GGUyfk4u0GgCKWzIj/mTMncvkFSZ0L8AFmLUM3x2VVj8b6K/J9BSIa95OikMQjMPw1OIu+
kl7/we7SRl+9k/B2KMGTM/wepdHjoqMUDUHsI6wQeQ0zNZlJ2uFDPvrQdKDCfCeEh36UBJ0UaasZ
X5I9Z+s14ZZJV/IR+hLDg+lr1LbjhmAzuCWCKFwmOt4rccXlACJPGv0y953ihxEJMvRdaF24mupw
wGpQg1tJFojydQCk1XsVcKl/eSkGDeZxwlpkM0x8OF/j2EICiYdzeNq2WIZg9fWNRxCgzxvjQFH4
XApLutgksVtUElyBvFaszaFhwOmVnzP7bNco4ecRBIZZ6utmPRONLHzK5gvJaPbKodzYrqtQ3IIe
iyZVAcJI3/s2MDKVe3gZLHPE2NEJl0CRVFMTMHzsRf088arAgCjpOQ49iEVUlykoKDc4z8vYsvtG
66LwJ6iRorFEekuzZXZ5c4Hi5eaP5WRYZ1gUP4WUB1aoH14IhB9AQIN8JmPYAA2b95nKr/Z3mAkv
89P4fcORoyrvYtW6l7DG6WiUSF3yHKWwJcN9XhQCWHhYRaKmRIARn/aDvjdN8Rkpy8IxLArAZ22G
tsnw+83uL5K0XMNLHddtbYgPTBUz0bJx1JldYgASiiR1MBQFDbeku5KQYJyHo2p3xvMR9ZCYEO3V
m2VDHe4OuuI70A3zEZQQYjalq0EvKx4ahdNNYcnRrJtLFNQwcR9T1OcZAewlVyUFbxpTYEjgi1a+
gkIQTQx9tBYHg+6+KGK2iQVTI6RKC6lFVinSgFGiy3yhjNG5n3eCVSQk5BE3ar/1QjtfKUxvnyGF
wxO8jEIBFEx+AifOVlnC1vPvUN0T3ZvgZXKPxra1RVOY6lqVb9RIiMD+cM+sQc3lo4M9A3EnophF
uVUEWHm8Sm3g5Q1W0QE/9qkgIxGBoMWQXI+0i/kkYbNN7yBI//ntcPQ5IL+q35gNBi35sLkULf5E
s710sDx1d+I/Im8npjiuCqYU7e1m8UHLrr45AUzFjA3psGSCW3e5VyvGDZ7Nd5iByCKSV8Z0j36L
b5lBKar0+cwAymo4QOXcEGo9jml9Q5bphmGclGVSymk0Jic5K6pGVc3caURPRcCL/0bwkAEBPhy5
HUK7jAyOlU1V1UXkaYtT6bXYkk+ysfwy1lVuDVllkevrMfOfhQ7QqxrZzdbvYh2tUIrxlp432AHq
JbMUZxYZH5jbggbZ2ixPbg/hcMBzm9PQt+se4S6u1WxEyR8Rm6XNMKhd1rKgdALD1w2QExWaXVJd
l2GuM3/YcH5oslvDlQJNDmG9dA+6rnqA60YzvzDP3+3IrlBtCOdNVxrhxzNbDvE5j/g45dKdPJpS
LAnqLvLW8bfUiJ+ZRBqk2hOD9jQWEsYQjmXRoWt1iAMDli6CbezxY2fWOvByod5PAloQ9zOpq7dt
m86G6/LBZiPSZ231omXK3Ewc6eJyTDSLrBdxwHky8H9pLgOLHmb7hZF4KrmBQezLead0bQ05dOyB
MSJ3EOOObYooeosWYvJ3A3+rOi4IA1L+mhEZxYNECBgRtk03093iNrc1SYcCfQyWqax+VDHNbuzu
7nmNUtaZLdqfVbrgzgIIU6uXTPU7cZ1xNaOHYs/4Uek4PXNfN7JvQv1md6LPkplhEu8JbY1viWlA
V8KQptCTRVageubIyjdOdsrPoIpvb3gqULbvLi0ukJlhfKsDXwswy2uzDba2UCQTmGhiwJEV1KR2
iAZ993LW8iRrDXocVbmpj8etNke2n8D5hdh/AQ3Bn6gIXeTWPXl+ZIU5zEg6g9B5W+HhVvUAXak1
yFOdo7U/2v2DLIC+KWUZFhgekd/oyafGjQTLDgnMCVA6CAtwFwsTkXV2btuD/rSWd2JpVNClqz2U
+Dyu8vpTdzAAftYFTtuwUwhgM/ZWOC14hvs41acZzQeAtG9CizcSOz0lyOihwTNd4vkBR3z6DEN8
Z6Z4zdOhy4YFzfGNWxcmZWLrExBDALsFw35+AXh6K4YyRkXHcYtZmx+XeExtqdqPXWZ5qZmJhZpe
uOK4c+aIXPDFQaezxLoqNycATDSUx+VpGt3flKMb9JDq8ALl9ONURMlx2+qcMDmB/2V97Jammk4X
ZTEARmIaRXKP1YxZEsoS9BGdERTb9DO/+kiiwPsfbaLpo/GyEEFwPWK0HZVQOh5YGO/k8+rxnGyv
OPQnhTufwSJ1cpk2DArv5PQ3pIsM/sVcHH8/WBG7UOaD1LR2f1MhACZH8baITgiH3urf+gbf4uNU
KCxwkFxna3LCWB5gZQOLUhFuzA8CuR+NwoxfgkrwsGJ0tu7lvMlDgYeUOt0P4M36lFUnZ3cR3o0l
S43sh7vl7cOCwlcq7XSo0O6qvVzt1689iWqZAbKzfOFkUAQxJdSotRn7iJT4v6tik2Ws5JdyNCJM
QTgOYbnFceXeQyUu81MSjQih82LXWZnonYzg54nF5OyrgeIA6OmAVsTcJu4CKLVntcbomj/9IA2V
MV6JBMNBc1Or7b0AiHuWtRbUA3hFK8xICX2JMPROZGFG5ZXPLmztU6rRBv8jfj/V9uLFGF9iBCOm
ghDz5WjZ5HKU1IgsFrqYQTtRunjomG+Xdi1dNr0nmlQwbGwAt2B74KVh+muO+YXFnybqrP32WRUi
1GP7vj0ZDxyUfS4BCfPJVe8XtXUz0W9o7c2tqSkCJtK0Ry1ilJzxYNKA4u8u1F0wimjkyY9RbhEx
hWh0vJllVRofDtIRIum1J+VyQlzihXN9eKD2VIZ03ZUUQEyjf6aXQ+xJYivkWqKK/dObuEPxrvyY
d+AhDVkocnBw6zZuG/jwdyKzWaa0QDqY9qnP4Nw4cmNxPr5b4HoJDy9e54mCBR/vyN/E2+LO13Pl
PpbOqPgEoiwc+vcPy76bOve/0Xq0TkPb2iQJMkdRudBjtK37+BlZx51qnJTOPCpRdQyrEoXtvhGT
36ys5GkIWDJ7H0s3ae0PgYxX1xirhMU35itaa7wv2CjuLawMnC0Kf4+gZGjsul/UmCmG5SDwHogK
YUMMqnZQpdwFZplhXV8D8/41gh4o98g7M1e/uyIifXUHB2VcGnVTzxcp6ePvxgPV4UBEnqA5q4BL
pDI11/GlMCdre3ddo5Qs5y4CDJIMO3VL+2AWhAJq/+MtdQ7GInVHPa6viqU5+tuZ/x4MacbGiVai
Bq/ngHv3W9dwXidduEVHNr1uS6jhmD2qzyi3SkGtSfvR9cLFGFrGZRRcXh7+8Fd3p75Bf9tJ0hS+
JGRPzZZL23BCN3pCJICZ6PGUoBbGYRfQwKQHOunU+q+bgleDIKA4Y7ZEg22qFu763IdXkCwmfzPF
3K2a1rt+vweZFS1aXKuAzoYitGk+0X2syoHNre/qkt/vwPTkReuKSjMClCk/a3cEWytNvpBO8xWI
J52dSJ+3iKBwia8DeHT98bBlEqSYtYeNFp31lK2URi1Smn5Jj491aSWZLI8lHOMUyjO8NOT33yyA
ANgiJyTGJzr9mbGDkKRmGUh/B2/GWVAkqItRrPPS/ihd7U7q5ssgeDWScCoY3SoANuN8ArkcYvlv
AYcDSyRYj+Qnkc7R//aNo+vGo1xU0+og1JXiG2xkvgKe2LwusrcrMalH3ZTMhJnRXQvtXICMQf8l
bLMwyxSUO0s24juy/WYZva2LhNlrNj1dU1xD+db23ea3aUKXqafu3RqyEPgWfeT5CJwXarLEpgIr
VQW5vmd8se7OrlzqWIp9hQ2Mq1HUJFqlAdEDcLHW3s8GXdBYap19ujZ3jzGDstDfiVXgifcdBulG
P4pPe5LxrXLAMCtfBJJ3mAFtGMK4IydMcDpLIIm/gi8ShMs5mK/EsonxzMn9EROueaHTyXlcFTAo
jv+esAeoWWCmL3nR2oovgGBROxFTBxv+RfPl7s0hY+ibrmOlQnA3t/CG16G2RDSeFtTL85b2+5cE
32OkAiA0QSWt4IwQbClbviM0WbMTMp2MsVz9U4aAdsnlegwLTozJ4nUZjpZPxerceCjn/sECAsNd
g6z6i37u4/Oig8M7qryh6Aod+uHO3vsTnnFSsipcegy76xHlsvcnBD7fp1sgRRTY0NfeSbuq6JtR
/9eEWIOgqna5esHDWiicJoN4vsoAl7dQ8l5VL3/qyZH+gVvDPsMCzg0zsEwTNWb4PAhO0bleh8IQ
ga1GL3oRdfAgiAaFoMWvodDQ8kQDNUKj+iP+mFClLFjXANvRVHg5bCHcdQgQ5gfBFHYvSDfJPHsB
h5+0KqYYUIUJC2RtqzoSfUZ5+VSEs8/m7x3bJA91e3Yfu91EOpwxHPiFzLat6VRNEkBF6s35ucKM
+Yu2a1dVHx9xX4Qkd0KO49haGy26/MpfYRKepUNeLOsIgWSahXIRFJR9pvP7o94HhZtWJG0z+x6L
LhAwybLze9+fQduisFD7vWKxuta/oIcfwkY+SrvuNm9b2OXqljvnLYlKQnMooBHc/fgMI7OD+vb9
xKTpceSpLq87ciCw+r6L4JwY7JrtQtLK5v1AyfyDTtPRHVsNIGcOb9Smpde6Mke3pDZfde3vINrh
B09MsACG1XR2oAYK28VKb5jcg5ycGFu38w7qYrbNzPBYJRGaI3X57yWM7GKtY5apW4x/bI7NNCpk
gKsknbdRtMTZkj6OsyoFLX5uNJPaF+ayc1/n2mc/4cYNYpUbD8h5qsWRcois5GY+zwDaS96eAbbm
0m5hLZ1EbTrvyw+12HNghYGW0YWtUWd15VyhUpWe5rP3JovDs/6+oIWz1PSKJFrr8JeR8s+Sbx6F
IyYSVr8Z6zdF2VQuNJRjspKqqcaYMC/ZUtZPCOGt/SK5NDyHfMgUg0fppJm5hMKB+8P23egsXS9K
1MYEkrER9SE7QIp2nxEbRZLn1zos7sb5jQXoo1GwFZu6etldxhMMKIEXF7iAeKG6jIor5lHdOTfT
2jpwlCehKDkImJftdQGpGIGQFdgeIOTvRCVckxjE6/GhUlvnKv7v/P5tRtwP/5ShJXqi/6FcpK67
n5nkAg/bhyJNLxFki13wJhdtdqemOB7nweWHKszsgQ2BlypFI7HRAJuzlm77tiiNkaBayBQj5pKf
EZVcRKNiV7JPZeirnyGpwWg1Zqe21x1dFazojJZRzBHfLJ9GDPZoMLjWlrJoVO7WkTApZlPlcDVb
8FMhEZF04Vm9hf4CdedZb6eUNm0kW8xvo/16Ih9xaxxVnfT4zCOlsXnsRrswnmHBIRXuuROxstG8
z7Vxq3vtTYiVeUvOG58L6qXid/YpECxaUHAXhTePX4K3IFS1/Iz6/ySXEJToNBnh1M5zuKltV4PW
s8nOJz004eIPxn1VDWnDSuOPymi40fLGaQfMkHRFAUe/2IWd4Uf46p2hErF1Mo6FJcEw/KCF1MzE
9/wLiZfJW9h2VqKLHHou8b1oM5SEBm0g1B9hGjMcWBCJ14RM7fgwGjMQ5wXIXNoQlQxn03Y6kB3G
dJZ8CNUTf6YsFL3Na8cUIvhEvR5Sro28hsEo1AO1ffuViYJSDp5Iq4X0P67Vau16vuE4ZGubHCaK
LAP7jmKBJ2mixDbGa3P1sxaR5oMUgTdP9GzwmdRlbDdywybPAUUD0QQnkDN4y4pBp7boU+MXdF+u
rfcubfzZXNK6Uxn26889BB+ZM4I+4XkWDZBHaYyQ06aOrUnEugydFemV+ISQ2YggV96AnIFkvZta
ZbH4rMy6BGsXht1oajRjGWqNHFakQ0ZgSXnug2TNVJSnQ1LyuzQi6/q6IIu45RFwPRWubM/YKIE6
vMxm60FB48XmYP1C++7p8K3RWv99JJiCsqpiyE9p0YHx6AXWElfLwF5GwqaoNbwiS071h5IoD1vv
uIT0GD9uy7d8y+JBlltQ+9fWaltyC768aMroWjSsySlB1S2FOL27cRDNGyfuD8C8Np9wwyDt/4C1
BXzziFem0mwP6OT7WicRGQ5LtINA7Wal1HX5XuNpiimFEXCHVi9gH7WkJznTdOMHs3Vcw0+67sND
RWIC8/K6balt9KwaEtm9U5nZ50hXFfyP1azDVYAjUknhvsktsUlMcMBopIsnJKnelAR4HCWZIXWW
o7lJa7rUK3pST5BSaRQadYhoPj0+SSPobvW4QmIgv9UGNxh/DTbuCHu+Em6NIqVYhDDE3F4o8XBn
tVnl8kF+DbaphhTQz6uSe5FwEORMnerDNMnmh3T29EvjOjCWk/Q0/GxxBFVxpXrTMrkxspNkkap2
EParIzOuI3Zpv7V2VE912dVuzT3uQnqSkPFyIBPucs0Ex4PLUCMmWA9Pd5lAP0x9OoEYTYzrdFU7
gpv/aJR6KzXnxWkrGcWoDlRQLYwITBqK23z7CIwpBr+qqY2NXIw+yDBS3vz28id1TkBE7i1595y0
a9HldukgwjZaqCVKwkvN1f+ZB4idNAkrbFOMu29ywYNZ0dyH+KIrPXmKDd0IPGUyPr1dZQawJGiy
MDYzw3Qy/MOnkubjjfSAtGIVyZI70LFC3nz+T2jq7SA4qU/Ah7EnCFAi1ipNCSRCMNdxd+ZvL8bw
+iinmbxaO++jyfqR/nJYJllOpUm1VXmtiQrouBTq4Urj+ik/Np62mHIveQf671P/Jz9Efdgx1ar0
iweY2gC9iCLqNy/yPk3PTmNSm4fev+Qr8jweU57Os3MUyK20KQEbM/C42LjGAYC+Tmkz7kETrLyh
6FCANnfN3YIgveLzK3h2uSwFrtC9Phhfp222upLiCo6InCSqXs7bAuCf8vLl2KaNdxYc/n5CcQ/j
Idl6TDjx5zWP4zsqKkzMymwYsbOOfmF/CfF4Psk1iqSrTL3ZIgTIqlvAHfyHoyfHDs5J84uS+Yy6
BLyAS/EUhvMFem9rwSAfccm3+Jass1lwBQepXDNRSZ0Y1esmIXd5OCo98796bpjQF84FLSeqlCFM
UtO75jsuiSy4qQwn50dK+YaDVxaeXlEb5rZGIRfQrQ+iQuxxUO/h+abb7nJ7806dMdsxtSZDirAB
NnRkuoR+pOW8yPD7X2FPz2DkZV52Y0I5TkhLVk9E/k0VTraJgwwor6L5mJB16eqXxDEKtWAFuq0A
GRpchHmB7Uui7YzCpfmuG0gsS07Evju63quRHGoAeLa69Lr/NRloQ41VQWaE4KsnEJXGiLc1ydzp
n4Hmw7M7gaci2IMAap7KF2Gbf4U7M63roznpQAKlxyOqaBTC5JxEGatcyyJkX4Vopk2y/NoW+V+p
RfHzNPa+iDB2KNDBVcd3U2LVuQYmEEB5lN1G9SDHoSZDbczEz+FyUyIjyJpFLfBBncCVySrI33ml
2P4bSHQOp39AboKpBwLop4BqA1IHsYxFQH58twKxhu9l2jam4nGw1IQGwRudUMHUxL1vRgaP4ysc
fTXbQxqO4M+rUbTULVuBleqUVlA2z0LRfWcg0f0eKLnlAZ2daxM2oQZXH0ARyfPN1oypI06BbIwo
Lh+zgyHHn5LDhSu4H/e6MM+63nwiRVYGpoDN5MFuR7I12wEIR0mP4fzzP8Z5WApU3Os1SdqsHpKs
LtpZmRqBWxQP2riFnTSnlZqTVPOHCI76F6WdaCIiFaKWbtXAiCXd/2GrCdrsmXgjc6WhZHHP/Who
WxkygXZcW1/e3jpAI03nykDDjgw5/S1lvQO0yiD1RYwYhzgg3iWQowOTvzZlOVvDm5j09QV1953y
1GazCrAI0bZE55ftGELg1iG40BTitl7uI/Gu7vU0Cw0hEwp9OLcXau9qEdH/7Jb659bBk/ajwcL+
RXxYIv/PUgCQ0/cIBKxq8ePR+582McpZubS7R65soWBEmZeCMfc37uWf0J5r00mtP5eLAzhpIgKz
LgUYxcr6Fi3unrOpYHUD5Drf8oascatL/F+AH5ukPtWKNmK/D8MVo+u6UyNjTmHY0jZZkRGMYfp1
svIdEMTh63wgRXRRUrYt8ejR42+fip76fiFoGwUJx3LBinb1KsDBYL/z1J/coQBRzeLcjfdIyrFo
uflfgmo35P7FGhyRWbsp5NnvsSJddEu0UAix31bVbVeiFYYQQp5UjHJw2IeTGBb/D6mSYzSJUrzV
LAHakcnJ8kAxX8iFUdZdE/xyFis3K8csH8iRoGD/haTU5ocTKxtO9DdKbMr2fcLTH7MYIPinjsyb
V0oIgQEsXhR+KRX6dNv1L4OH38g/ygooUKGtBq0hxumCfK33OK/H2v/aCQyrBhEK/4alWphTt2yZ
EiV2CgIdmMJxEPJ0lS9nMMtIuLLyKOc2zmfj4jKotw4mBOC6NphKlkIq7X/jRZotX89Z5QyfgeZ2
HwE4/W0XnkOX9ATK3cebxpeQPFVjWzvEOFo5KLUfR9XTzsFcjD7sznDovEeHZAWxTRH8Uh2lGsAv
2oy+UGVoNMN/wYC8DM1zmsLcuuvRApoSXxSjNbEcjPjGCdmSjmMgQ9yPaCFFOhTl+NXwJ3068r5A
iuWEgs5YCAG81zy5K7yfnWroQSj6amKqmceUK3qKjPAyF0foPaaAPjnryo0XIIqR5N3EXbDUqhvv
pOatcKx71RiVHCCizv5djJ/lDHZUGRkS0M6oyELGLN6V+HaGmvQs3GupM4TjnC6X2+7PQf6qW9Vp
4spu7tqZaQwfX6auQ4IqmM5KzLjjANLzPRbCBOe88RSsUF/5If+pk2oEZxRwXynD/5pCis9/rYJy
8+oiq8Ck59+b9ZovkIbKpeVAapnlnMKtYkGEBsoey/pvHAUfMXH5QeSCGzMWFoe8O0DA2YrNJcvn
C78Jc1+wHz2LdD8rFhKeQv/ZAUbPNRzOEwUusSCYYcBVnEdxgyGFn+1qAGMFmKz8iSh0Ff+t3zjo
wx6OwgIA1HyP19+SMdS+9xspZyGgRpWdirjiQumCFO9nPJe/C2i2d5UrehHPnn5uo5qFHJW/t9jc
F5/OezQxI/XuJaY54PUAqDbh8r0fznx5DBg4ACHx0/UEAg7DU1/961gB3V5k1RfqSpqHt7VO9xDj
ubYrKMsbzz7lf0oewsvnYkfG8AN9G55ZEGQz3/Es/Z5vYUT2MxfqjBo1IJZw3coZe/93pXRYWBZ+
KaM54bKJWM+mcnRv/rtVIVKOj69ANf93esPc02RvR1DWmo7lLdBoNZz9vLcAycemb1Y/B3Kwr+dc
YLcZoLjJaBD1XolG8R5I6wrAZ7BbNqvsoqgoD8HPBCl9oqkpNPid/k0ITpZvbOaGZKqfPYpBVgcZ
PP7QYIUvtIHbycw21kd+AZ4XgxUOVvGK7Ji00N5YNEnIIG5/Br7KvVABHJxWdM7/651Zv4j6Mzz7
LOz44sdj6Er7iod6MWsElpdIqPz+giCYJQcWTdNA+6kiO6wXIH8IJNlMychJv1ntukcxAxdGhZuC
nQgpBn/ppipaJg5+Quu18aWNDPRvNxafWF6gEZSNFtLxjDq+i7Y/EDlpcv5+z5QiHtb/cV3M2T4G
DDwi2gZivkCF8xWncbJzJKby8R5TaYmhEKnKAEXZ3oOCJc288P/YqLNxppEIR14XPnBLI3A7P8Xl
o65lLo85vm13cfQfD8FckBSQrZRKqv6Tbo+0pv7Giqxwf/b1EObZS+XrRjH4EEMPWM1lKTAhwF+/
KprHqLW6D16B/nSiXzYjsgN0lL9+eEWMUWeGSfN1T0kEX2prSx2E+OK0bNy+NSAIN3zM3ct3+FpG
n9f1xoZGbhxEPGHjCOw91fX0Nad3RXuvo/Xm+tX1Ig3zHuim67efBnH8Lkwfi7/ixJtTUPLObYF9
ZIhMFZ+3YJ4YZUeHi7DH7gLFUCXS+pFra7lzDFFtpR2MztxCaD/eQmz52oPDN85dAnJZEDrXmTu6
CsyI60ksikZOacCXnOR2g7WWkL89copdOxQPgk4ag8R/jQvBv1v+Ny4afisfWWx5nKZpT+xGInX1
dKzIYvdAgDYuX7v/djCQ5UEO0EuwEmyy0I2NrgxGHTEwel9dDhhzvmnVHCKeSiLPYPFYNeA+3lAo
TGLe8eZOr5Qgz/26VoAq9G8W6c4bK9vorKNnjaldtnCo0HLhnTuPJ2NELUdvUzFqzKEdd2W386XL
+47Cvceh1F0GOyEgJ3MJKJQHRkTzUzg6927u7lXOniDe2rDx2Kn71Ufos1hiEciTUdxYoWB0b6yl
LVHQza9WMh8+aYer7HnFmDrHkk9giEyR9EX8nRd8UDVSxBxTrQwwaG/ZCz9XZAGZSOY3uxGcapTx
CUWFZcEneBAQszIf+Lh9jn4RdEQEtu8tEME9sX32w2jWuzrwfD8As148AagkwglwiKIVtlsooNJ6
v+/T8ec7alyPyTl0KVzU8jVOAmkKyoT+Kb5ztWTbJuvehW6h0xsyzNfSUNcxFBYUFxQNdAlsVqtD
Geu0TDiI4+iwNIauxGyNdeu6lziMIq4ZnoX6pzRN2bgJBkPqatxE8PzEqgd2yGa/1EucisG4QPjE
JF3pn08y5aR54+3+gVgZNCl6hnE4FPYwkWpAt3980B3TCmJ8MRDAgvlDiebXHT3ESrHLT4EoVEIr
avEA0sq5Dy+u73a0r+WGw+o6GTdcDlqR/pKJh+MVyjvwmI8ieaDkf8FnEjlmHY3K7N7Lg+syqH0i
25HrIuLGL8NBwrz7Uf1wxn2IiTPKJqh18ppcO7nZUVmYVyO+hYMtFSRYvVmCrt2nl7BxOXe3o5nb
vt46XGCYa0usJeKp33tJnHEr0LA8xTpB0Mp58TokgKY6AEdu17q1iUj8d5y7nQmCR7MIyVy3VXx9
vyOOYlsc/6byEsFzf1llrGg2+LzRqnVP0Qm046cO5KtDdO/i8OHHAAgaL427Omw+PRPq21UEW/K0
u0gE6t5SIcf+nd/5AmWzUbrD96ihVMD6sL+28fUowTx5TW6/k8PT4mlJKZ+8YpUMGzyNK4KtuHcw
Yc8o/o4gNHV2FOdnmOHf/hRiuIXMDTAtwnf+QUrsF41oLZvI90/7oq65ZNGQcObDTZv5ekH8ls73
KasVHkoMLDubCXup1JN/Jh9evve885xBXd56CeDjgj78CjJ5du2icjoehrlBcw8vf/38Kml9Lc7I
QiYt+kVB20DydF2XLr4lHn8VPlsiyZfVghdZdhcgqM8gwY2SGY9wtuqMbRcXalaXpjI9/XIohxC3
L+hOSpe2bGG2d2jCOj+limLura+0xKraZJXkmzWXVob4TpYyadGtkR4a1+fmgW1L3OA/ZgKQnKki
V3cs+Ytq1u/BDw8AlM8+iZ30ukxWkoXERztj1pfTSEZG0YWAJbJ1g2FlOBuavbUyyhVUvJmfb1F5
rNG2rR2JJUx057bhGLFNbjOcjBvQVcRPIjtD9N3BLoH8oRoCYdsMkTetNtu7gqmsS5yUbyWVIyKB
Ui1ri4utYhtQ9H5OVArct/3tU7YTMXYPv47N1+wLVFjEtQbKS/MkCv+5OWbK1Wov7U40hUrWHKee
EkUAQm7RsUI2O/sdLGoJacy11X7Mdvj4SSkl1MTJRyCsnqqQR+DF3Oktu7CoUrezeswDAJMCiYsP
PJ9+5zsaCPOokZVduvwMoWfYc063M1iIyA1E9CI05jd3wVY47T+QrowPadWs1Lql3qZ77mlU/mvD
ZqklN0wSxu8uonIIXjiquVfGehoJUU6WsAXkhfxyDuwDy0iMluvzZBnk1nbWrSlQB4i9AcYx5E07
Nvz+5Rpr9l+1LqWiL+Y9wzxAATm/VNc6UHBL6HkMYVyZSgNtDAk5G8+ODQarxAGW6HQB85ASkyGX
XWhXWvkw+t9tqixoAKOkaqMqSTQJb0o6AGsEetSjPuV/MsL35asQccFhnEr06f/8Yp2XRd0OZDvw
qAXWTxNxo2Uk8dEBr9BCuM8rx8jANWkHmj2bfaGjw/W/KULFV7NRK+0MejvEkTF7srXEAW0XHx4E
kWg9sxGxzRh9C75WgteidzlQpSj8odMPbLdl2jpTtRq6+k+Fa9+lkCfG6zwhjpgEEL1Cl/qOUfqB
n2iJeCBL8Dogdf1Ebhs76tCi9FHKnOQf2PGTztF+RIBxaAYLYFFXZ8d3nCHQo5G/6VEhU4wYgRvm
jAdS4y+4Xu0xv1NQ6xGLdaOjO5/+WUSNUluvQU7jdiCSaDuSn+ZcUXBa5jK8euBGw68SBKeCe5bt
No29EGHJEFmqM5FArpBYz5St8umYhWnddVOVHSwA4YxxzapbK8paLC7aiMGIEKJpO8YIMV5RMtqA
54/Kebwc4lpH4qtbFzE1TkjmnxahMkuKCEozVRq45Ucpvep10200Dcb1Ocwn2gXmsAhI/6eJk5kd
vfdYAfotRI5dRnwYA0sf+DXKXYZ70qmF18uyyeOtTfky46IJBGlgkSyi19Gj7+Cc3kffuXj8Bkkb
F8WEOBxMPfbW9uJmd4CSv8HV+gT3ZKPTFClpe3h9Y6flgBzCi8FHwRmDn3vHVZj9OS8KP51XAItL
/rrPM2Hv+JUzqNPZf6XzGojhTKxwm6DLKFhofjlsV/eY0Qyx54Hrm526Lap+3Evb0bIz6fX/geur
oxFANY+0Q2OyTq2E9evYTkAyL64UQnwqozjqluczGRmUfJnq9Oq35B9zxnfFUjPJghPiWIW89xRF
XXnrqOpgHhjhk6Z52MOD4AFowf0w8dIGUatQzMVAdPhWOS4E6DTDgq2ePb/5F/F/Ga3PrdmsgAKg
oD+NLhqFhL2MYKrMxhHu/cYzuPTGVYkEqRKjK7eujEcvyfPsug4+3z8LqzJ01HqbzsDV2fqRzWyU
CyrkAw0+R2HD+n4E/aE3DBfl7UGL7n0+DZuXbcMR4DelQXC+D0NVwIVcGay8g5GGM71X79pBfg+o
v5qg0hFLqpG58lhny9mJXx2/hRiREKI2JK9GQmdzQJmDT+Ku0ZTJff0AV5FpELrnySFAqjPHvyL0
AxD5H1rhVn/xnfp0hx4e1tXSpP+wTvgfAgbYcr7neuQBbc/o2yDFEwWpQpoqf9e0OkVMpGFHIPvX
bH/MNCqcL7t3UjsOvUHFum1cm7LE4HFUP6veKbnhggw27oU04QvhWhddf/qhxlhO0wTbglnLaC7M
9GI6A9pbkvnnBwBqxEh2vEzalo1QCDtRXGDJs9HN0qoiuzqJct5ZJpfNHXJpsXiv4s5+rmPM2UDU
pRU+U8n5dnCWf9TwvRCtC/2UUgGhhqQ+/TzIOiGxcTQf1THHjS3Tu+6MDfogD7/fPNqgEdpv8ITR
2SQ1Wo5pRramVykvpJcWE6fnaHoR2ZEdQSNQMpC7T5ONe+e7F061b/qVHarto0rvp8h8R4F5+ET9
pLmBzHlx4sMeCy8QTEIlx7c2i3YWR7F5AQpoe9j0FFz7ObbuwIEVHegzhrtuZHpMqndMy6dYKb6h
8dPdRDirWXtcpnSB3Qc/Naqu+zpLF8WtxYMx8IOEiDRCVBnueAFxt11uYSD5wAjZrYc57TbZkA4k
1wgThpri8rgLvQSOXbGzoU6PvtEBxuFw7XlYotDssrPS0UYIdk4jBB34Dcnfoz02VNa4j+vd+lfv
9zaWUy0rj8YHfFn/jhx1d9eu/PxOpeqn+13rC2oYVSPnvhr2n7VcslNUFzpqTKfhPVTKLiKG0+xT
dSpIX2OYe/Sy7c0e9VsMN66YrN07x36V9k4QFFI1RBqzyayAAfyN+Pdu4o8AWqo6PW804JFS8teE
9srBrMm4YpX4Go65zGAVHvwAgwLBVjwRAPG4pkRA8300ygUn+YPjr1d1p/yNr+FKqM2rGAELehNu
nBROx2n8OmBWTKA+TWB8Z+2/YJpn/OcbHNtxG6raGjTz2oCXtK4bJR9kmhsB7Fdju7+6mWAT/Ia1
3bY897EzzffpG909UjEUZWETUPA/8dbn34BYDQMgp31wC5NhMyNGUXlDG0leeVj+WdkHrs3mHKgL
KHNasBDW9/m5Hl6kPYvPpzUcn9QBhUrV3adQySLzVRvWv6Fi5LFbkWglhNd0fzbh9M+UoHPxhuer
eXoGTFPqRPSl7iJ0FkwCfqcJObHVOriMv8mDXz8TE+dy9AHQS00HxDiMDqPYHNSoDPNRUH1mHUZg
TseF/fESb/bdsiUua/oB19goGPSKM3StkZOuRAQ3r9tQRMyPGOPpxZ72WGjvfSzrAIU4JM2HpIxP
lZte7OPVG3s3s2cNhmyXsaKeM9ps25pDCdUB1s5G29Bdejktufr0odKxh5/YtcjcWnd0DtU5oHKN
KjDin/1HAHaO7/ZG04kP2nBKPfuqljsta9ypZpqWfPdV7iElAnV9ToYjwOEss6QNWcI+URpUFMxw
D2t8ZLGKBhkRJX4NUf6d6QOGnqne45UWUwbRT8xlXc/FcyRJIie0HBBW84riCNhhzkGtSKbAZuqJ
weEIcO+WxtqIkEcJoeWmVQbbGukbwrRhMYdzfFvTvsuFGvhXGCwjRxtIoP0Pd6/ShcFzadOqd33m
p2jnEHIa+UqLp1kC/yVet+hVR/CODli8WqU1hRGl137JF35eopGCUvpo+pZPEl4w8y/xTo8MX3ew
5RAiZcdmIY3NDWLuADeYw3Lyw75YEIs3/DdnCWC15/Ylk/s6gmJnf7NtmvxKRF7Yhq7XxR7+a/Ne
KgM0RiGaQjvpVpJk8eRkLAkHlCskmDa4MMTegUo+0n385U3BkXPcmzrjAW3ap+fVwT6tooxEvI9V
W/GZ+UigTENWh+SdCpJfTfXcrB79Dl/o2ZvI7eDNvmQNB50KFionFwHwyLjFbJK2PffGDPWCYyER
wDnbC1Hnx9+6ynpY7uQgh9ZXw/gzStlBnPp3TxBs1o6NoCvwx8uop0Z++tt3osdKtjdKKMrHk5YS
9QOaK28Zd5iIDeozooaiMKjqfy0tfj6mxSKFLg972qzr2tKSi0gUhr6JctMoWD3NzJUl/hE8+a1V
2J11cLIGZhELmvlO8Cfe8fTOG5oDDv+9tx1qoO10LRYLxiCg2BpCTvwH5PHiPbncZQLlW7eruz4I
Kt7OzW61jKRLhwcOki5LfZdZ8HCBTRyMsGkGMOnME4DuH/7mPxkQYj+BgtDahhSiUunUKM9jRKYK
to1eUqrwXVivEQRetz9XsI0akNhCondZiBl1MzNWmvZeXFqPb2suHH2udRyI6hHEyDo7pLJfRb3/
t9Ml6LFyx6cj9+kmNzTkUyXb8UT9Ez4AqhmML4dKd0/ciUJbvv8aFbKL97uUxrH5JWBKZRN359S6
dmpKXBLIvyZ9o19t+ZVjOLk2r8p7zFk956AmcEVyERzilH8SXGMsv6dMyL1GAwqr51WMo1pBqi5i
EbdkQcfDXCOG/mnLSuaYboWCb3XuXNfBaCcdBb0eMAtGoUNM2bCeef2GJe34pozyNMTBE9VYfq5L
mNe11tl0Q244buBAAYe2+DW3Q6DVZkQ4AKbJrnUt2JQCMuZcn3LIhGBFpcxQ+eV3SGaHdKmFeg8b
AmTh0FCebxNUk/7SMVIYduansQNBzlzIhjsZSvGST11hgfhvAulzt6aGPTqasu4FbeBKRrpQidK6
V+Syfzax7eUY80T0sIKjk0ACw+R3yTIJZe95aY/PjYCTxKcdL94yVmyQTlebUDcdccZTGTzVCvH4
Aq1guqfROlBPGAiCKNSn4h24PKze6VXLj/AzZ72VnwnhfW7S9otpq0okCl1qZs7SHKSSzqckpTbZ
ysA5ufjZJr4RD2be+rJ9aOeXx2XN9LaX+sa6oJtDtt/n8RUkhkZDEF93bm0cKh7fyWLk5MDFa0bT
Z7VggT6zrHbS5Cd+T1B/iiGcHm/BzQTbBn8//dLWxCRgoyuMPF/n0hlt/Qb5qTUTo4hkCZO4ZSv7
jf3y2k1tZVOZ31kTDknHPS8nhiGJzZnqMtdKTnyAhbSFg4ht0hySUifiuY7KWshmSiCAZbGDj/7r
A7+Ts5hrNthn+JYzMIs25aqvlvg6q5cwhC6JBSWomX65Ui8g7z6aEzcvNPfMRr0ktW2JcpcUu42U
Q9xA2eVJTGFD/ZvC7ppFsRxv8TBCt5tKpcajXV7DEdIPHhDOaZ2l2PPh11VspiIqCtavRAHln/d6
FFGRgYW2jVfkgq2akJNyjs5VBnil3+aqTfSJW2DiuZ1YToElFnUr32zMi3SqYUM9pFc2/lB1RN+z
Zvgidq5Tq9O7tphOo/VxcBQX3lCJJW/R7VznydtBsAEYbiKnrCw4Glf/7TVugXxnvHRL7u2Go2kS
IpMupaEQ9U3y+2iojFSutaFxX0kvUcjQdwx8nRITsuFX5pTLXpZ/tvqkAc1CDc4Aoa+I1YfW87L5
5fb6/EdqM6bX+1cS9MGfQ53qLDcG5s1d5MB0xw2Iu42nilykwL2Y8qrKqFdokj6P+RBTipXVMfE1
Rn+D+2DnlI+EgkVnbv4imfFGnG0b7LQEMNxg4TmX/NBdbgsBRMUUgyC/U0N7OExv1kpHGXmyj1Nk
4fs6gxVoagjeIZx8kSsxNKcxXTNh0N+5u7dGY6es4ogay5NwuuTlR8cN86K4QfW6Av4Lb+wblIGT
WQEFZvO3toONPbeVuRfqlnRfK5ZJamo/uthQwahrBsFBLNVxitBEKRD8CyZmVrZMtwLW88a+Kz02
HOVmbtM2xUlqLLcei5lzciDCnKZjJs3q/q4tRZruBctTrOgEUg7JE0DefuuaEXgiQlpCb9v0e4Iw
wcZkINWF6xgN2Mk+OMtiNvA8Q3coYaRg1nmMlAL9QQZtt3Xh4udI8D/zh6OCEBmZjtI/+1k1YK7r
GUAu7gV0y6QS+UTeNs8rU4C0d1QV7/o5TUhBTiA37mOc2Sv+GKG8yG+9ar/R6z6qlc2ofxrRdZw8
UsNiBUkqyfp9nMPIH4kSDlwW6wp/8Pc8yIVM+Q2xTShd+0P1Ih8MGXcJhAU6WPAmD5WLM7I6LZMc
EfUf2U55I/x184PELzLejKUvLy2Ep8HRt3pKZVUN3wFtDskOmt5C+zbowo1uSeik00z+pB+HJ6Jv
aurmIoSX/YtJrbeRCTZhRkdo+CAz67NHtXjLeLJ0EVeUc+VVCpn+5U3DvxFHR5kb1dn6CHmNQuX5
0dZXPYX/f5jGrpJWppIn4bp0Y2La1SpQvnW1E3o5znTXleY2vfPmEOJ0IDP/ndVZvxFMpLEtmDs5
6gUHM1eXsc5Qj9y9p4Inm3Z9F6tpAtUxSsqvtDmiprvakU7jAeFGr0Vq1GmTbiNsvUQyzbwySXd1
pAB8DdYvy29J0Vkr0MFEbgaCt4XQqOI0ive5nECMCHp7aTKmBTJybczorZAD8mieaVDLdpsuGBkr
LOSvEkrLokWhGhN8tHb4pOqNO3VTgP7uWeBhXbtksUmK0fL13o/VhAHY0RjIIRwqzuZsgcWOafeT
OtwLPNHFxd6sqoAFK11449SPjPwfMrH3/Mn4h8RCig+mpFIBZJuTo9QqGJsmjquZU9qanqrX0zGI
lTnKpMJGNyQsRuNMpNk2NNSfSja3LbIUq6JM5rxVWo/2GWR2UNikn9zXziFODJELRReg5+ROfQTz
BhmzNVwn5Jr2BfRMuDaexa00AZRNUnfhopdNHpwcA2Cw6f3DOh7uU9xyzykKPLQlt6r1KE3TeMzv
ObX4P2ko2GMEOM8/Tybynh8I71WxK0VGzHxhQJMIT6xVQpmnqH70R6cIY0tERtsJ74QDGph9yXfX
92d7R5HzQO3kcJnwZjwxmWPpZy/8kv/HrysndCnF++VKQxgoDpwocssmwUvSikGaW/pKQzAULgxm
GCc64hSzSbFQ+ymbGPj8rGEjUgLhYGxKuj2ffbA3asbIAjd7P2DwrBoHgqBW6kBjZmKPMn9SDH1b
hyTUVs7Z+Eg5QgP6XldTbpK3GyyEjAD29GNKR9/p6XIg1zoBNSB7jhBvXH3VyvVNRq/JdN/TKG4L
i6M9GOOZDytqzGtf/BGjegD1S18kKpa3AEOCzwCchYBURI2bdJ8UabCcLfHXclYg2f92DoDHW35+
i3Oxa/Z0yFVW01MsJnaUzEmetTrhUawH5gNoD3VHtUULXAsXMQySnVrOfOPYAJ/WkTbQAa1K/qj6
Kl72gmYalQmyzxT+37/bv0eSZIQlyU0xIiRn9OGZgZVHA1WGzHIWtPG5hdTaO+8A3ObUfQ8YlEio
6DNzkiDxFt8GayYxgFakl1ZC8JVvnVAmMOFTZXT5E8mm9TkbVwKA/6epKSa3IyjEhIaM55XZ9rdn
FzOGZw7jwE4Iz8AY7PUk4neM7/z/Gaakc0DNLjXFwfef5uF6qelRj+TXBWsSsK7+vkdFFxNWnY7h
8fgw4gbSfZkFfnjVq9433150wxyM9aNPzZxP9YvMDbij7IRp1j3XkssGDCk3MQ2tnW9xHgfcgn8u
81ZLu5RtDsX69MpQwa5hETQq3zSQej00KMFnZTjj9F/xw+0HCOP1w1E2qe7FL63z/prhxwFRkNFu
nYvIoTsZaqkrOnqcA+G4dUh62G1evEMynxZFUZNr9ew5Wx0+HhCWFW/F1NSmCJEdP9VTh9la3ilv
s8miilfTTFryu9ZsaGJoUoSYI3hCjaTPl3y2rAArORcWBfCZAgfgnQd4QZODuSWY+Ft/4q5uryXK
LDGWdKn7/nt18TaPacFhMsN2VGvSCjOXa2JCYjK+YBfQpuwXwRvDRMVRg8eitvyLWqulOOgzxwv0
tcbm5uFJ5VPU1SOVfjX4x8lzHw7xGvM/rIOJqNDSfnaAeAL1CU/1OwGYIX4kSr5TW07wKIZ8szVK
0GsWz5LGnvsDdJwys84zlwdbK7MfmUVtWghVuv7P4fFXCqooN0baL2Y1NUyg5KgkmiafC+FeqAuh
DURsXx1aFs7f/n/C6GAx48cMH1YhVoj/jeCgvwzh4DDajmzlq/W5EjhYkgDX4GYR7pvfELuhg3BX
mzgeQ9vc5BMtDvXsT9xkh/EfM4AOGKQr78JS0/5l2zN8Do7d4a35upqhItjInF6IWDG48wKVdSRj
YTeiOgAmtQzjORsrzkA8Z4nXB9vkJjI02HYpsEhaKWdL0+KBzakhkyH7t/fGXrD4rZyyT4P2M+39
+wXH9P1ik2/u0FQotPHh0Ox7GSGk3atbF2yg3Agt9V0daTeIorRRTq+Up5Px+2noFrAfkYd/O949
mPyI2ygIruNtxdXfh37QxMhUeYeI/2heaaHL17/BhcVtgRl0TuKk0CJhleVh0RkjtrQCy9t8DoNs
aL8MsXQndR0kPjwq12/tXuuDwkdvvi6v/hAoEPyrBDh9lOJCvZ/S9umX1QmVA2fz5q0D0ZvWd5pS
422if2GUvpCSOfwTPHZ7zEz3NxrvuQfXzGUP/V48xdWJnnFPAvhBbfI5XDFLSvtupRF6H1b1bRpr
l7mWA3FbFPBAPw9wIeXlJN9AOj4+RNZ/uFTKsRhU/WOoslmKrivhoqUO+39ngfDUWx4R+QPd/aDu
auPjPi0hLbvL3NH8B8cKSi/rYoNOad6N5fovZPVcvAoJtFr/8AtiSYXkLjZI446GhnUyIYl4S57D
28OuH9x1MPCSTDpwfdGqouXdxPpgTqpi2WReFCWv4XP+88XjnuL0B1llhhq9Z+RdwLsrzAIXEGfu
tgxW42f5FnXB4A6KVQ/lF88Zs5PYT94Rnrabd73mJJ1SILYi7b9pB+JWuyb4KhRiqIPo1Y5F6/L6
5/yPhd9FL1xjvCK3oO+MP2is7MISLqoXHcVB3gtP76lnNoAV5n4v8ndhOH0I5FxhBenZfeCBFb55
biypvP/Vpq9jxbSP+PG+dwImmeUcv6ot5vsN5nd4onKql/IBLpzLIMTTBSQ9eejD+kV+jaQzN2VO
Dv2zrquZ+3tX79rKcieAN8IKVVVox6Dj4J92jtfuMVh939LoMY8PXTV/ViT/mZaKE+Fn/uTaU1FV
NmT02td8hEghecNPkD30Y8BIE/jOO9vPcSodrDYdwy0KviD5I5PQlzeC5cu1bv7anud89SSL/le4
7dsOCWFuLJs+vILc7bqh6xYszTCiIVwQjxutI5ZtnkskFUwtMMijYiOmikhs4lM7R9tZhWMavd8T
/fdmnZ2TTkfDPdpW/OK+80HiTWBnWNz3FSPXZ8AR8cqPfBIMud70TyljtrqTLYhgTiJTD9emX7w5
9+ZmWZdqjir/DP4TGT9TbJdUJ3TGJHLy0oYNKLUAgAX8+3MNKuN/zsMABm6Mk8bcGSt8YAePTwbB
w90lOIf7h+bbKqjR63YCr0euu4EiuqEHEIGOR4DuomYGNGxOn89ydjp2FuS1ZHXm6UBrfDGxVqlT
P/uojyQUnt9lcHDIMxaaAC66B9fZuFWWw8JAa+36vbhYOajqKAJUwoHxvRLwhqucBphcbzvLhysX
c9e/2qm0Npie/IPr9X8zHPMWIaOa8K1lg+ElkfYy4tgcoD7xZOCBWBhZyz2acmif/1OznoCQeuzb
c5nArchIfx57pgYHQHtb25LJA7CrjwnirT9pLFNJpjLhMoUOJupc1JDr97VAI3HSAc7WwW45Jsii
R96vY4JrwPc3xv/L7GQFpfHTlue8/7J3A8dvWQi+MBfIsLM3xfCtz62H2sas/8t6CkNYz5b0XQXC
o1NHPncXh3CvfxzXCGCf+L89mKCryNGVWabH+JBWPpEoVKOdrEKfc5/1RHpKNNwaNJVSkl4edDiq
ZzjWZTwgkafqN/TYn7q02H0uBS668CQqJGcx47XodVrdxHFMZN91E+G3/sBKx5mIqA7Tf581Ruw4
6Ao5I+LhHW7PYftxKCAvuT3A0CssQqxQEzlLxNs00dDMvX34AYZIbSQMtEcxATRJfPILxCTjYfSG
ElZWiqvgmCeTr+X6kGg8A53BkRQAukqhGPjy56vE1Sk6edHvf3VrnJ9BlIDptvX3cEi3jS9I+6Mu
J8jMiEZ1UnYqU7Xg/p0ZNLMNSbFbe9KDD1NkyAMiY8IECAHs9t5lz+tEPtgg151gQex7FvkkJ0QN
6aODtuxJWAt+CAq5UL+pUhg5WenRJHTfvRhe05/UdO0HzuErn9BfI9w+OEQ7MW3Gx7zjoJdoOp4+
O1Zl9w4jkx9gIitbbcy8SA5C35k/YI9KymReRk2gJWfkpOiK+H8LH5ei9HRVEeQEcndJu8WKzj9J
TA/WZJkW0qFpY03a8VIj90Ypts1CStEID/id5iYWUg9OwHGDTjDwSBzOkUilmKfbPfs1iBZKwwh9
qgYF8N+s02L+NtgUcDQVbNHQeGt1OGf+voQzvf7RSfPvTFmbvyoq2y28CVAR6iyfYwDOTXiTyv67
7CoT2Q9Ea5Nvz5NlKIXAbTWBrTVyc5iRHB7Vw2J/ML92LFKlSoWiuvfk6S1eMgNkzIKVEsohBshz
TpGVOyIOsCiI5ELwcEyyqDY9DN8ft6kXPAgdOpydULEuSVpQXk0U/bcyaVlfRDAP1TrtPQBVNfe5
63AivijJjj8anwvTJhvV3O70C2nbL9Yctgd2fBWAyiSAHxtIVLIxLw5Ul+pEbeKgmqMjjwTZe37v
XhgqbVrCwUeUZkaoCf8/ATj8XzFOqcJCKxy0Q0ckjfZHg9Jmpr7O5SWIcRa1qQO2Zg+5rYKUmE1K
NPStRsiU3Mxu9A89TEW+KS4wVpcUbE92HYqNtR+o/o10p4thMFeZalq/Ku4cyi6/VtSqwYndQBE/
GKbNw0SVAoyaioT3z3xqyi2pYOoUoxcq7CWPWIMQoV4CVSNzYPsR+m6wzci3915PfPzimJrv8YOA
M2jO09ofTFK/Y0e0G6/YB981+l3KUzJN7iVS3k1PDAETicjpzbIzQp+OS8blmMumg/fMtzFbb3e0
33X7rCZibkkCCJXc/OYO5Wi8mG+q3KQP2E+an1G0yN4/i/KzQJhwZibH+r3/A04nkqyJUF4aafBE
kZEP/Ag332zPYRJUSZS3c5nt+mXQY0rzHd+VUAv0v+wG5mupuLuEiH5UyT5eM88Md+hFgw7caD74
SSWaJVAaQhjaznDRY51D5nTKknjyx2zXjAx57jRQpVZCtlo0nQK6ZD6xtIc6UTfxpmEFGB3a6/Pi
PFI1ZOvT1vRigTCH3oWoIEHW1zSsCSV/CXzjVKoGoCC/TNkAtuMgrpEGPcj47WK6E2FNkwOj4QeK
3nrQUvK6bXZQKGhlQcdEEkB2E6r7OQ9zznAJv9DGNg+cq31barehB1WsWhWIQPYBMGxQf3V8iBic
vpSerSdx+xQhVwGVLhKDfpnegqvH0gvr2SNinCs40fCR70p4SIZnBAmgEcFTovE0E/cD4d8pZovr
+0YLXfP/uDgviV41qtieOMOoWYHbZx3jsaV2Rn635S1inC2mwygAMU7/7x/mhv+shrzhJparPqcC
3SoNSNKFYIcsZOmFFt11fvQ5uzYw/XQ+BbCFQXAyP3TIyyRxA3k46oxDcB7zZN5DkuyHq95n9eeP
OKxqKmF2WItfrSCuBKVrTAB9iEGtfm54gB/4cv0QpxnyqOy4XI67Twr4jdEISgoU3EMnao4NCd4F
GMWlvQFRikGZk0e0IgvOGqshNKwbD2K1nJ5XLQ9/y+b4xX8dra/eFARK6RIQ02ZjlhLsWfoeQjYW
fAutde/s+CfuEFGgP3AMuKpyfr2YEYLGO8kEuC/v37UA1XD/qv0fH4tXza1CTHuMX8VROp5iHRkM
oXXPKZ9+LEIoDkENaNZIb8Oj3allx8mNtTgX/Xe5VjRxOLBrj7Wx27rLBzug2oMK6uCIHxMKzM7a
HBkmA6VtMA30l29ws/cfa6gY5633Q7jZG0SwN+4qryd5E4nDW0dA+SUEiVms4uOPRhuuc6TXrXud
G1rK+PdcbDIGowCtatMY7MD6I0DVM0Iq0lmu38Ot3WZVWcSrx4lNJMb/OFBDb5Q7eGS+7kBTVi/S
FMhgHTug1qxxXHMaqYCOQ6Eo4htnrRWGCtgYKO32HuqL0HNwWiJnXMaGMOG51j6dNmp91e7SqxwE
ijpXfaQ6OaBd1kkVRNRjrR4iUBrlggkvlYF8GOBxAjzkP3IAzZ3uYpJTSMxAfYEGGSmJPwmhBH1d
duw/OSvUGJmoPM82kfsqXVa2pqwJb+gaQ33XcwLHKN84cEfL/J3yUyFpVSorz7Qsniqvsa+YHtbp
4C0L2wQcbWJu7GNuuci8WW5w+w7+ffbT6KoYJehWkUDkL22k4/21jGf/kBRre8C8UPOv46APozFs
OKCZBZKNg9xO39cOrbE1s24F/A9Zs363MViXiLMc5x+ikDZ9t3zNiL+tt/cTv85jXNSNHULN6YAb
eMqWGGKL30KZlAelwdJcBvYLntMT5Q+A82TuT0HHBJ7BN6+1OaxNJ1V0Ncx8rbxuUlK388ZbObp6
FQRKnOrtw6WKx9mo6I8i4145g/lK+X1SfuqruhLXOhW6YjbxPYz6M2jTmJeEwK2VFoQYEAP1VG4X
HidVBePx8+56aMcdPrvIsA3dYnS8WBXJdin7goXWpAqH/vUYwF5dQigNJic6W5063DuhMmnrbid5
hs3DxgIgWftq2F2fPHcd08Us/b7tzjH4E4vAaL8U3S7FENgR9TP/fIPvuoBOd4z2bIt4b9gH7Z3Q
otxeG4Y5Gpvub+eBJao+Xg6+dfKKdDrcBUIC124eQmui+k4Q83O44n5hOtCkVyNGQ8+wHHrbPVG1
3i2E6tM5aRbW6cbubc8xJ8S5wFO9UKjhyf6esLDMEtg4cvTbBeuOx42gdbz1Xpv9r95t+6ImL0YZ
d3aS6Ps1HQzfk7hZmLm4DPiceBOJCFkqBfLav4mk+0SEMvDtPAIEl5Y1O+guI5QqarCq0bS4uRLV
F6kSqZeGnZ1WZJCQMB4thTDCL6yoTasCbhbijfMozgLzYSgNzZQW1NZuVRkKNdZMrlwbYey6M74V
KgBXsvkm4Bub+QZEPO2x39+mpewjofzd+tPNrfVThSndGuPDLsXBJuDKJSiQi5YIU/AtZJDNtrCR
v99uPKB60OIL2U+qvP5hElB1LibDsfh6a6eJ5TLESJgmC3RXHIsyewFMvt9WzHgDP4bkL94Y/Jue
q8akZt0VfnJD0dqT4TgRIaZZ+luBqWD2uFzyxaz8QoYqniDXwDFO4xPlnSAnC03VlgNF9es5GC2V
I/DtLNFORGa5unrODAicUzXPyJEnkilLFP/vkpHDF+redkcYw6puc0bA3rGMJZaGSZFVad/KasHD
CahosV2EEnOodUAgKQC0n7Oqe9evBpoxsPwkJE/7Y9SWZbqYM5bHRNog4BSjJpYds56pWgnzj7+u
M62Jy/2CVOhWbIeoIp8e/Pave0RdCaKcm4z0/LWnvpDJIha6frq9LkK5LhuNUpRAxe12lZ3fNB7j
8l1yQulQP0z40b3tnKktGBwm1Z1Vk94n/qZPEm96M0BsXpBts+mAlLoNb8TPo3lRYZZyknS1jHoE
Epus41hnm/94gg2/ITXbR7K/klU6Mlx0pGYYfy35B4gtyyjADV/bLgiQ3vQEpop04CeoGoyTKKhr
VvQ8TwRiWfdr9xZ4Lz8gXZwbdT0dUNoBSptayuzueqgcwwGkz3uK7g4xE4pgUTpnHlH3yA80kfuc
YVEiDlmQxVSp07Sj7SdUpMrYi4JB1Ms8zAgUS2ICnYfOCGv5tVQkOiqj97nsAq9DcU1H4Js/3EXE
fdLKERiTQkZy9O+b4yRTCMeJ2Ba8vdiNdGwCNExKUkRzc3psB5npaARGGglrIEu5oM5222bRAFeY
oHcoiFGTghhfUJ237basXQYRAogXQD3QTaauTh4zyy7UUInJt6PLuYnixVj4D16StrMCWRpuURmm
4+VWW+4ngSA6g/Bs0FqlrvEuirDoHp1XqkiSlJkMOLEEu+PbetOmzxedgq5YqyOcu9J1Go4N74Ny
RefmofL4h6jXyrx4E1t/Ioxf89jzNyxtFOFS7hkvP1MAry6gd+ylqOv98C2nLLp8PLjWMIdTmxuE
4BCRjNgArctapmnlot2ou7MiQPdqgQwGVgAMD5JuAy/KINR77WCqyol251tEjKj8bEfIr6YJKO+1
Scy3aQmWXRTi1kwMsHzi2m/v8M7kgTkOOCxfi2g5DaQ3zDNYEVQCzhOT9tAZHG2ptEzcBXOuJ7Db
7zJcLt3YhsRV2592io9ytjNHdy942ENgKeePaLsCseIIJSca8WZwLH7uHYEqBoE3YqiJi0otte6M
js5ZfIm/c+1ieRctwMXRJbtlbR3occH0i3nty00OY6LbdLwW87XIacpVYHdSQtyN7n7YaQZQvxA1
dmgSgCSbw4nnp7odbjkyYDh0Mrce49OBp9eladIfmsYs/yT0apHOl0SNQ0csbPXIOc2R87IGAEnh
bJjYjzuBujsIees/bpQj86phBSkD4ajDBBAa1tjpQzePqURouk4gEg9sNsJyWw+t5fC3GeUYZwBz
xSebOlLVv7YoE2qfMcY75ex/1JcQJ4bZASzNdnRZvQ1o7xRMvhiW7CVEyuKumycHtKeZV3O/41Wm
ymtEnDmM0qKc8yIkQvklsTdkVB5jKWcCjUW8OZyMusOUehiCnRvaO5rVwdfh8a64KgwWw+8I5T3H
QhvYBymwvBTNlYvBLP9mmJfHgRqPMxoPf5i4uNEIyI8MCMSTJUsRV7XF7b7XWHbnBkZs+ZSBwK+8
SHQSzq2pKja/Nt4ohWNmpVoVBWK8M3dpBvz0jsaVObIohXmrSLICE2tLQ+cuN3PmKScYWHyJbRNQ
Tv//VuYw1uONLU6VLBj4XI05RF9yCRON+MZ3Q+x8xo6AYFMxyvaJqjSSjMOF33M6l0zcAHoCD79Q
eo3Iw3JRej6+Tz65GkzKUifmkOH56QhV4GqvuTHV7SLaMGJE/rHmgHrQswtBsDSpajDsiTHd7UwU
QOS174kfTMTaO+wdTJG/mSQ0nkEsrAi6fXt1OmjN5AWcjFZedlFtxCeZDVk2dHKf9cwn9JgXBYhA
tw215kvF4VpTB2wJylbLdKuXYuvYMC6hJjUxMaGj83URZgZ7DlhS5OoiJrRcfCE+7/gnwtMpcJlO
VxO9biWZMrYlNjIyDuKF+4Sr9fyIx4rwaD71H0AtbwT7VR0Cv9fJJjQN4XL1kAf/P7yddNRkP+ra
2MegISKk6IsuKW9kIdr9ao7EBXb5tI3d2KULTJgihFk4NF/av1U9sXFLeif02xOtlSNGglV8Ph7m
coGj+/nWVL43sZL3jnSLYoCul0Ti8D91bZY/E71z9AdC270wpVNDf0alzBE/R7cAwRdIwka5X7SI
0kGYGiV0SiUq/gOke4K5ekmH+FGR3cLFPWAxeiMstSWUDEV/w0GZkNohaR+y3FMPnvkl54khB0bL
Oy8QWzC237NgdnyoLIZkTp1VQXU1ys0fMB3ZAkNPe2wkQ8ClZ6XVck/FpNUFnYWIbcFeAWlCHgXS
NOV86T6P9LYDDBbGnYikS/IU0wUzT9wFMA1fh96pYOJTTAgw6DSy9AX6VzerQmApJYW11RihCTVU
oSL/Jh5dTFIkubFoVYdRUPqvYLai39H3Hzp5xA3c4DORvN/9XhKOoUEwksZkqI9YLm9NXKfEtHkI
EsLja5a+VRDLyrzi74Y5t52z9BSazeGH4hz4wWh6g7lgmSJFKPXOBhKamCiKHsjeGE3PYJjRJMqa
6MMPzssJ3wzlBg+zfc/QI9XGxtoBrG1oBcSKz2jURvWZ/uM34E2kz0DTVusDIx2tt54eE3A5dUQU
v6Kj89BJQPcmzZGrZoXeTbi02jBTdvmyl5lpoxuIK9espTRy/CRFWItri4z4jx0hVSKCgg5v0bkY
fW9cLB6GLl3PFocIZipwyybVrctnLlZv3cfCUt+JcXcJset0ot87OUtlF1rBgt538YDzNLSay9ps
gbIRH7xvQaj2HnMCoTSCMH3QdoOeYvvifja7UvGYz1k5TtGl1f+eWOJ9aDx3z+6qwC7nKJtHZjDA
dB8JiDo0F4C4yQum7oT91Yy74BRAriKvKCCYtCuRvTpwJ4Y718tUgcq+SNDOeLiN5pm9O4qe8B7+
77DCedduaE6jyQlDhBByKdd3pdcks/9UY6XbwCcyUk1KYKX+lxlv9bDd/naOOZupiqY0VsRC3OUq
e5OTRHVuQB61Lw6zjNJuuKZ/rlXLmiIleU8bs6wmjxRZ0kVywmfAioztUjbnoUQZjoNI+QwLNxmj
uSCkGqM0dtvvv0mUjHqt86vK4VnMiGoydtSFGSa+UotpQj4mh8hiyuRYOfr+oeeMpkQ9TzXXQgaq
LR8raTULVZoOM5ccpS9YLCTK847y1Eeg8LMzT8IPM+cZ0ldJCAHbOd+IWPfY97AObUzym0eQ3oQP
a0FGAhyHwH3eJ1//KKA7/ct4ZKC9IsKhZCIznNx8NHrONrs0+W5YdUQSr/tA1S3JDAA6XswX/ZTl
5SkOxyRHJ7k1uygs9AjaG6cYgGM0+cN3zUuAa+vciaaUdl1YYzPkBR2M93l/Zy8jDZR6EIwYypiR
DvUKx+vH8k4oR4zTO7nnEWlU8CGGrtz0vT61rcPy5F/t3mXSFsNgdro5XfE8DE4xF9hyFufWv+4u
+cYfwQJWrjYiXkk1XXIcCGP1WF4q+Ak15WvgXskSbOqy9yCxD3kdHYO542psu8Il2xgn5fLdsX3h
a05eVy0g4VGxqxEW/2a058clhGTUMvACARrdf4YAtMSsZS3QMzHuoe5GkNE9Cz1FGYO558wwhNv8
TvWhmJMJbJUSZgPjcd0CwmqD3DdhnOV7qN4KZeWj6VTkq9ePvfxA/7f1vdBCaEm+sbmDq9+yPwiI
u81Zq+3yWfBfV9AXkules2Gac528nYtR2qJkQ6xOTc9FE9hKlZYUy1EKX+KWz16piHtEChOECilN
ypoTeHzv/cSayJNUbVtzflXO/0/WHVonHzvWyWXYn1vd+qxqirueHLHPphEVJjRKc/yNyYz3jL9f
Nj2G+sE4tgpJDibokzruvX2sipXUAv5o1P8Kd0SL9MiASlaspK7k4mZJIYCKMhNfFlIlvxbhunDN
RQLFIDSsODGJZ9oXHAEyVZM7uQ3zK5VmEShmuinzVrB/VaKUwX2AMcOyKq12K+EbEuUuGG/Sy0cY
+vGGF5rBBHrL1hZY8l2kfqM9tsLY41mfqA8Us6lkKQ/fZID+1jqQ4B2ccPZyINWVB6eN9vs62YGo
7ts0LTjG9iCZOeyrTzHyYmXJHBBCjWWKdeUfWr2+ucNFQcuuODqs3zecb/eI2LGAGY7o/JJGAjrm
xGv3yki86Z4uZSikU/onD7piLcRp1ZLe/088AW1P8a1wEEo7CztMdNtQIc+CixYUe37HdfTS6cuY
g7YSE9tWSw7F2n8aHdTUTdjcmj9JHD2GViVVYav5OCxBLVX9+HsGIG4Zwt+rEmNkunHEHev9zxIY
9bicPeRzDAHUj+8Jefy613TRMRBdTwzoGGO9jT32wSeSkFgmM3gxm1SUbvsOE55l3PPQA/OwvcoH
ttSWTrZbwB9hKZYGzPoWhOGj0zulUK0uPhGn4s9d0/oMiP3gZSOWXjb3ok6fyXSXKygzHF/EwM8h
7tlX54ja39ciOm0FitCqowpCj7iw5AVWXAT0HLbF0EcA+hD7KkYnRe2kfxDXD9LetJK28OUGkXWa
aZ1ELTJNM+gYBdUMFouEEbOKPEBnYkKqNlWrCrTh4E8Qz4luQ0wiNTTpa9qvd9a/q/qsZ3y6sdux
385mt3CM0R3KolR0yvCz9jbq5prkZ5sxn0Mu4pSiS0uPfym+Lud2Gqc5oEyb9X7gCFT92b2v0LlC
j5Ome0eDHmYZL/s9jt4r2uS3GuZSk+2CmOX5xQn0Osrkx6rGPjaBB4Dzkvbh4HQ+dPhWIpTpSUUp
JmLzbpUv+2uBV3hM23vsTyx+Fw8oEPhVgjH2WRnZm7xLW2B/mEEh05LZclhJkkbKkf6vIYMO9qUC
d8PZiK90mwMlSF2b/hTSNhjHWmJHQkec2mv6tpP0iqiVpb1Q8LGpP9ZYZrUb51xPg8MXJA3PqUCu
/0uzUi7s9Nd6GJFPLWlv1ljwJykbgtkbVAm73BPoYcayLLCwiCMD/JZ6PfvBMrACxsse3+9jS8Do
454lMIYSFnpmRVO8emr6nuU9W6j5Ex2+dBDOHvOnkxIefg2CPZ9ULMzGOF5A/jYAOcJzcA2SAugI
Mqsz3eSyep/0uuIneFi3tHxiVZm82/o1u+b4bGsbfAe8b8mTYue/PRayLJBwIsVC1NG9gNWv/Nj8
TKmtT0FqSIuzQQf2OTsmd+/kNn6UKuji0k+pi3EQB886qCWnxcxY7O8CcmQopTQoiHLQ0avXp8jC
6a7zkgQlbqQelxcVM+8mRuNE6bexFUAfy5mPD4OzUkQuo6yKtBMMz9SuRZ0aZlB0IkzipH3N1hiH
VbLmPD3RnxFE2z5ZZuHj0Oh+jCgYtkl2C4mLAUCzXzQL02Cxbe+EerTIzYWsboy3MoxVrWE7tBL6
LSsGYwkDKLlpmKQylFpyXN9oOUuoj7XlfIvDfA1EEkGo34mpR7vQwYr1nId370Hle2wM1w3fvAQP
dP3RteW9piTDnrZTlzz8BUeBuRK1GVHDp81bxYsg4Hxe8G8sWGSVeKl7SAgpGVvhhlnzF2Bo6w3F
HI3AmfdUuCN3FyQMz6LUJzsbgJuFEZU1xNMyBMaZQbWxyzTPQeBauXUHSgh8vh7JWx6C4gUt8QXR
0V18RRessj6afvgeaQ2jPrA76soypo3rpF0tMr7kvufr8vK5Wkxy/1CaydFlppFIhCCCvhH9sawl
CLxfgk3Arsu9jil9g2xydW4H74Z8sN6MHERbqc+xc1fq3/63BonY+grf9Wf1Za7Wfo7v7xMcGcSp
7unC2F99aZw4MfJ4nUCRWWgktFU4jQWQeh8ZE51nvAa+Q0hSem382K0RCsUT9LZ6h8aEHPpmbHEF
qSu2iYElBmJ9LyMpjSpmIzMK64BTLQ3KI6cSWDFja9wFv0iU5iHp+leSk+WuusASNrCx5gnL/4tB
MJZYNtEj8I1PNt/oBdtVq9RRhQrOOF8OsW1Vn4N+EXEiOhUBvzALRjlxVhsziDK2oJOmkH+TOJ21
CgNxmIAl4vViPTdY3hWuWOKHtWQDFqOo5yPTqkI8VGH/P7y1I8OdcnCtPORRw8ot5ivpqWId7rLN
M/j541Pi2MlGQDLmZDFXYEiHOsEaHEAoKrrSOQSMWlA/ewmgPPOGpLhltIlfeiQVODxokjUasbj9
YQA+EXuXVFT8axoCM+jOLlWQ+UYjC92n8PM0bN7P9w8QXfQ1RQ3Y1RRKv1K8oX4nA0uSzktr7zjl
eq7XajmivbdJkor97XntsZM5jep7Yo41E+jGtRLgYLCJV82GrrqXrxYd8ZOjdtUsnQS1snJYUmuc
DfskZa9eac20ixl9ArqpIxHotZ7sNNwOqfyyr/YyvsQ7RNuFNBxTecGKN4Sg4fhScBgSCgHR5f64
/xfm+Z9X9t4TRH0OcLFXy0W/vFAKZoUocSHsRCWdFYB3UF4e4KKiQjimMAhDEwVIJSqZrD5KWSgg
R7aP8pk3/Rx5pg+oELRCMoIddEQ5XnakkTy0ASuCY9GYJgqnkJYB9/fCa2vWS6E3IhQsFdEHr1u2
gSrvcc0xZEaW2i3vNxJREEjnZcJI++SjrY5iYjcm+P6BT6whJ5IMUNMqcYXez3eyK3kLkbhMrKiK
E8zWsamDXPYlNup+4wke9oDIhd7YjN2gTm82w9zJap50HzMeOOeO8u0m6QrgOUREl9Cz2AI5dv7o
/7kRH2vZgn1UvZgWSuH7RLh74PzkzJLrUScQtoiov1hHvpanZ0J+hD8hiyuzEx2kxVVpJGCZ5EQt
0koZkQ3tC73gacypq+atEbl4LuljdRtSoIOaIK5KDtQ24rfmeORvHdYaKszyJdgoCNIKvcBVzfxT
h1ZCjMpA9wnztJxJZM2xVS9e7vH4H95nOMgWEGNbL4MVDLlJOfHekbay86OT4sBr5CHVrBFiw6pj
NQ5/qw4KERuHR8gAKD9ZDfL9ujSkRCjRjag9AWCYD0ocyus4aXBrQksUSkOPzzwsCLS9KN2UKRCu
KisL674oXxbrjCXbtlv5u2JkMJgvTVzbhbS8IYwp/dQS5CMu57o+fwHH5TirfQ3rKlHBh5KEucng
yy4mEANWkbENgPq2hffYbZ2XVBUIqXrdnwRki99Vo3c0hVmJ3RDBmXkGc9MQpH5R9quJqP9wV5xa
5TvyfNAThCRQpX/FlBg7ThPh9uKP7oy1pnJyS1z7ownDKibs2Xb+qjoxgKOnHif7JYUz5FQG3UMh
2LcFET0w7SDUpqLvKBk3I5CA8I5vKF3aMKRABWkwcWeuWa5Zm1BvVl8JxhpsSCTGk9lQo1o3S217
CeSXX/c0sto2XPsWcdnsEuOcx+POtUZqVT2aE4zhZ7r9RvVM3aIp7hxrvafwi1+sYXSZ2mLNfoaC
C4yutepOtcwP/YZmUo+KlutgezbQO7N2yJMOr4wOvKBhKeR1seolwu6NqWvYaBihruW7Mpag4zgi
NHZbiqDETql2UQj9gxb9HDCJcuIADi69/XLsjNsVahFZQNXhGpS0izesBKpnEviHa9fc6JJZdI2a
NYMTOWALDeJoXSkkkWPFEvg9m5mtOwuycUaf92b8nIQIS+LMCmIn8goI1o3Ny+XtUhccMPgKq7Pi
7ZHBnWcLgeVAUs0SDbtJbhFN2rdJMSAFpMdbyjkZf8XHhJnPkLSIXtQsqW7ufG3dR0v6ozy4DVnX
QISgOay2CW5rEp7SIs8HEMpE7O1D9j0DOfkqCiV6/LOJiAHWUoz9Iy6/WvtjgHkLoQ+qqhPd06uU
H4IlO+psT7lcmfD3nu+bWZTP7z+47ai84bV/WPdfCyRGdAC+XlXTDEd/FMe9VRVf2Y648E0T+/RE
NUgFHCWhwnTlSXDt0S7h4rJRVl/bhyHc68bG0geX53O4Lhdf4Slrs0RdiOlsMJyn8Sv0lDXYbNWu
+aQQjNi9kA9wzePXTNhmHPERyeSN6fDywEIgOWCSBI96FIb64TBjyCDux8CxhsmkgclpjchVhpyr
1kzHa/Q2VzwljEs4PAII3K3HcgIsEiK1MTT+cVIVgdH1y1erS6u9Zeoj29FuILEO5WOS0K8L0kLJ
Ar91PFv6fjw+cHB2wnPxHg/f3mQm1Qhn1nhj+L4Fmyp6r0BXHX9N+UjdoNwo4Fj2FJuZli6FDbyP
8kFnr1FMYMLdljwqiLLpDmLOf8tn1xFd67w74pDcJWKW624lzM77TqrV1+jcH8g1Eg6kHRJlIp6J
YxfY485f536MDIUUrS3Q7z8RwOm6Zqdr8xehkx8hbJu7SNNr0IR4KokAkQppdpSLpdpwXew0gTtQ
OQBxPAU7fOhQe1OT575i4ZbW/ouKSMkCCaDvg+05OvTIMdF5Iy9ysjPf/emiIPKZkugmgzVOUN3t
Jkl759ZjDO+cqXoFFcWYR+T22hDyT5sNmCNilF9FRZxqk2UEt0H1xka1hD3BUD1W0cdC7MlYM4HW
OH37CmFqKT4mZlfj2MqSHmAdjvaUz6UEs0SBtVvwKFvN8wQedAJeRj8mUQBSifm8NPlMrR6bkdd9
ImEs4VIAftkDUkekvzwsojIH9oLotelbzXIpe8k7NyoWl0h4f80KAMvrWzpryY4wc1ZUr4rNSWBv
7mlwVMPysm7m9kmPq0u182IdTWiJHk3lt1MfxUHg8oTkl2/2WWtlHS2LSVGga15CcOhafc5KaEGC
HKT4rxlDIlMvVEE3fwoWXO/EvS+JKXIMlZzzyPLjRwEEXBkW/u9/9Jofh/jwYZ7i/2MF5me6fFGW
3bI1kDlvO6Lhm8HThBaoXg3KcIIARuEY2H1ZU2JR2WeoEk1lMfVCS7p1bXeHtTolZpNj5kNv9TQg
xZzwRSjf8messtOMlZ8AxYITC9etA4TUIE4/SaPyVln60QJvXcpjW3qrWoac5rVpHfDXtTXnmDS8
zVG2LK/OoO5CEyyVT/wH1d8Qd0k0I70X2jCXHLYBmiHEytk9N/neq/M5f7c6JlsSdyqUSYBIkc1M
+xbWqLMefjgiOJBoLfH6aZZ4i7WIRV2A6Cf3xlu5AGUP/n1XfaH1+0egGpSxG1tCE+kdhjCwzboK
qgzWQkJJHjVQwgjjcJ0R7kyM97HKSmgdj12zCPxzDEBWWVZyJ0Gc4iyQcUFhhcQbCjTjmrEvLNsp
zkIxlqhyX+s+bfq1U5+5oK8zI5jP2WfSnk60wjMYlCxhVg3dtCBVX0SUqV7TGmwSbocdTWK5AWp8
GjkVzG+dE1+KHRQHIVbvarWYIRlC+HCjaKMmZ+2eYebtsozt1gxC558PU05J+rkQPeA6Oef72CTM
f7NC8jzJLelfJB0R5GUz6c4d1MnXw9qHD2Z4hrFB/HCEjzBEXsJ+0a/u2HVQnD8tH/eGRbHa0RsU
aLZ3bTmv5Ite2++eJue7n4bsgPzJYkJpiVGvsg6v4bBQ4V7QJqmc0pTr2WyfdOXwmtsO0oN5ODpp
MGJz0pUygXoMy258NogG6v4hH1QYrRYy54jseu/j5cW3IuoFfkZjxgDe1Z8n4n67EcvbLNJP6u6N
G4RWih8fZT/3dpJ9srst8WKMh/AwZDBAjZPr+1Uv8X1WwDseBrRDzl5GEyEaZlBhqiWafxKuQu8g
uQIk4+denXBN3wmuJnsCQLPrlfA+K7iewM0UlnEKxaLmiikZwuXbzUGy7Rygy9HBOQty5qENdMBI
BhOhbl/65PGqRkfmcxT6+ZQ+IRO0ywKA357rMuoUMNPk5q8IIelhjBONM4yCbH/3apGeiTDFMg40
y6K9ErbOiuDlbosnpyp5sDEFHabyAoHHCfJkIdaME9DZd+6QHKFT2kluWLeLVXfNsdIV7kq8pMIh
fyrAZlYLMUZfzhxkxJUKOaOkoOhchl3pFqWSjFIOZuLFmzcgAVaI3QcVixkXzQEiEIp1QfNca0NH
QPMvlX9qP/CKE1QYBGHU2BG7jQcPvto7hZMW47WAE+KS4oIDBsz/SGgBNTcJvmBQp4qIuMSv+PYN
kNtNNU14e6gwC5uiwQlF1mZmsb5hzG1V1X4mCROanQvVoF3tIk5qctiB1JXJHyWna2F0kULqVAL8
bRBEAm5aBUOaSr/018jDn5BrNiM+Epp41rvs0g8Ztole8S0NZF+N0R1TZEbRregVlBZLlm8KGUmZ
dwuXOYF6U/NN7HTTValX5EcOQQwXHDz0RVXlcrHszEvyDbi7UcKKtlmF8ygqEs63ncHI/TGaj6Js
/SmpF8aX98UUzG7t9hJGhWahIZNigAFU1rxOI82YXkSaOVFts4+zikR17dFszP+7cXkeEOwnN4Cb
G7RlwhJzfqMK4NSa4WOLF3Zy0i0iwyN2dhrQrgM2RcDnqypicWwUds1jU3KhZ+HsOen0qzJVkxhu
VMkLmt52D9Vti0LXltCgJxTbTUAriPYIFIswmekB+1tKaEpnnzULIfa0EilZuZ1Hjy7dF+Toz4XU
urMhJDNEv9TeXChgsd7cVhu+Zpgb4IyOT+wjtn+NCrk/KxogYJu0tXAGcEZXLxMPNfFRkFrhpXbA
hZHwfH0vTIth1i1ai/iYCEdAaRfQGObpcp2xO5e0I1/MVucCmQNGm6sHC5Q/pjNphPbELbeHLbcm
K5jI9SMf0RyWMUQ/T5Tg0n2XQmc/79xqmdsojjwyr5hUVu81VAcV7k7xn7bRNlYEvvsyTXpY0pID
6SGEshUNIYjC0hkZS9Tfeq7izFaGvrnymh58SaGYJuNj8cpbO/7Ekg0oVA6FJPLlskeltad7xtbr
761Upw8oOQ8Wc9sFz4aSWnIl3KwvbqEjGCCF1sDh6DO7GDLYdh/7oKpk/kSW/5y1qKYdln7A0r3w
FwfO9WrmEZO0G5Or1RnQ33r68YYUB9Iz9IGI1fMUum2zi1ATkvRMznGuRVICEOvAOSb/GXNAmFIq
ZcYhDwas3Q3KsTzX+1wJflFC1Yol9p6nnM17GdYaT4JqlG9cgBG3JxeEffeBXkyAKHpp1dOjbE+/
O8Vtd+U6Zl24t5SzhLNQMwoXb/dLrJ+/dIX4EyvRtsEinqg2bUT/HTmqoc/v9ivyt11MFVf5mfKc
wI+BObw3I2FuR3Kt8M/bvHhD3hToHhbpSOy4immQEAY3SIzzyq6Ydk3kkg2zpbVByjJaFz8gfyE9
jb4Ltt26VoE0M/ZVf2EDRiMkCom5XqznB1kF/VjOrr8pEQvpXQxEIZyRf+R/Ef6bsd59HLX7Dgod
DrPOKoUvemSEEgj/cm4aJFG7mYu2GHgns3xJaxnR9cw8XEZqu1t1QTpHE4hOSy78QfZcusWdAWgv
uMbZmF2gZNhBfkVn8LA1aQyOGYe4M9k3VEkoUfWcsTgciAwGD1HrtTpwdTPk7kizkiRKlK/8km1Z
Ih9FqmpSGWK+C4ngX/8y3O3PTfe5GKNpfCaak3PZXyL9tiCWZi4z35kcizcAYSX0NLOd3Pj3YnuC
QWJOkwwGxHXjZWFAJGVO6bUYSwiBeE1sWk0rJssm+N+G5HTv9pI8rX5PIaYU4fnX85YYQ1qq24gU
N54fZVyFzCvtCIJxWxK+/6LBa91vLPUFUmGXk7lVtU7b3/mxyXrvWUUsHSLT+OuyV7YJa7uAMrbE
Gw615q961uE41Caa3cV8LsSYQML7zlrKq4uInLjzpvMY581RpZg9uiYkTuPhv4fZ9YwCBKFhFbev
8YVhPpJC6hIL8z5BPXbtDgKD6RQiLiIo8fZ82jLZ7T+lfsilFxNRp54AioP0oC9dAvlxBaVg71jw
pJMj5v11ZedSyTy16UvqsSTASlJYLMFko+MB2WO5nc4P67/qkwYcK48tdx50salM9PT45TsN+QEQ
3KykVg8WuiVZEjLVVSqSUQzts3cH6i4VE3Yty3JZAjia/ozI6SqdN0DfrYfEWxs5v21QI44iPjKs
tUSn43VuvmTX46TBND1XaRXBE1hXYSxcIOUHo8mZLAdSsyetLCcjgAqBIzRgadsS2XexCmPQYg6w
zF9dU6teYYcUn3/Nu9aLPm0Dra7aF74xcH9xu5ysIGFBKWVshlWGZTREzDLfmzD+Lt9oV+o93I0G
wSwH6NEB+AqeJL4Jg650xgwqedQyWw3jQMjKP5/0HuE2lTswqGLHCLAoYAsxel0KY44Kf6KpIrgo
XCuD/jnI2tzQxar4D4Hx7TmFLsluYGlrvbtuEaQsj+M8aanVzQl1hsKOpcrpAbGM8u5W0N0PGZ3u
Fe/Ie7BC+zU7f1KiIx24HXMEMjCTyWK5RfX1BjTTv9qeAHHEknbngZJejPe9alpX5TVZUOzM0t9B
4IbhXUk0NVv8uVufaB0tJXlRmqBoNiWj0jtd2rxADgkmD/3V0jd8Ezc2+D8yMr3NnQB/DYMDy9gs
3Fs8dmahCaC8kG3ysTUNliDLjAbUjwCKx1V2sPTQRJgD0nnBUUsg/V9309Aizpmvu4Hza/e12Yyo
vke8yhUuNhURnY4me1mLs4TcOhC9LuMLshaFXLDJl15YUiGJYNxWF6/mkyk28gQ+Aa0JV9B9A2W9
9x2wLb4d4BAu2HWjEONuQ94TxXaB4Ya/R69M+4gd5ZbA1rYj++P3cAIdYGSTA+8EJVT3Q1asjYxE
6XBcXcdaGkrtpF6fbYSLVvOVjPmqG0UmZodYmPbs+5tnzp8B1Pz/VqPS9jpgWAArDzigM29LXEAT
HxIwumFV/8foJQ8HTY3nR+HICBZmLtkeZ773tC5rKxdfTCGZktgk2tg01p/wyjsdDjqzTGtrAY+g
eK+TOPgIDVPjgl3tLzDCYzz5C7dKANNhA+em+NhR0caD7KZItO/oZ0JY2CVInEUlJZNFS9ExMGJN
2oLXwsvIsy82k2KctmSu8LfvS5mue8Pl7ifajX6OHCIAAV3KGLMNZYOnvZa2yipdp4neKjM+7iW6
uHVmeXJ50cS/LEcO+33neYFCIKgLkV1V8SYFqmsegeWDDn/HwqKBfFS0hUKz7FDy+ZfVN3NZ2sPr
H9jezsguh5ewMKHDULV76tyaw3MEkXc21fZJr9oxC1xYWKVawc44TN3eE90ZduqignyfZIPwpSUo
IPQPOcXuKzxCxkheepWQb37r76S3fJh2kJjikOMMw/+DTSbMW6cfwH6qQFqa0GVsz+Ub3ZzmhbAw
EoE7ZKw/jmZE3hy1bgOErvpeVRux3oGZRPJaN2KaFx2jbiHFw7VqwWCmyjwsxc0G/Bj9Dw8u04d5
QpMIKcusKBl0BcTDE/lgwGQZYDUuQ9gU6wfBW1tQ4rFArn7eDXCbB1e40nH4ENFq46FUFKj0VAUW
shdXBAJPVa/6EVWeKwWEImSzio2vv2nZxXZ0GJAcBj5wlP825udZTzeTKbRKx3rU53XcYGVm5o71
UG1V3lO0boUX9ECvFOqjiWCyXNXNxpf0viITVf6Kqf2X4cEj+Sooy27k5OVwL/1+lmvxlrgIeM7r
7JLNQH/KKNlo+OowGf2SUyH2y9LlLgw/k5c3SViVpsevuySr6DgdOcnNRIk2ihlfcV96L+ds0dOy
05rRE0UVKqwj+BobAJ4j1bX5BGQg2S1WLWGiLAOKgJxpQhDzdeTMs5FEov3o6yGafRh4G9Q6ffQb
QRh9W8RuI44jYi6xTKhHb8Md12J/omBIL60n8ajmdXZiHsJWr642IHTo7z2mSdOcFfo2xl7Tvb1p
vY77o1U+Xg0y+azveuO5oOfZLGEbMQDzIhqQXiw9lpBfFPQX2GiNxMKFeUvsUnmlx3U535Q6TTOt
escw0JGkVPCFd6MB5yp2+1/Vvz3wgTyQz/Sz3xfJ14zrvXqWp+U4MvUIlG3PdkmaaslbPV2OpaI3
QMpogFaIl3i3o1g9PKler4kTmoxjPwjJA902fexuSc5MSvKlZGRmHsr9AHAmjMJUJKkt2T/AUkpo
l4cy8nbk0Vz2gKeXvCqT5j/GTe6dpLeonRCDIeY1j9ThkzQExT7T5Zz2/iX0nDkXADN8NnPZnraE
TLHlXiZQIBVv3u4BCe19hluNFvzGQmbUEvnY/I9mpBGKwvgXM5aL+p6C41S1IjQgmfH+DOJsUxg/
zzjZ34LJLlVBihALW/a4UWli0ScPJRPduCaOdlyuCm6iKPAcd+vY1v6CaSgXahs59+i9RmOrVSAS
I7RFwuznRiqOruQtQGLZasw8/DAW/7ze2DmIOZ6SDzsW2gtRmXAMigI4hYOouy28Su+J7wyBMtXm
NA/gLka4Liiw73S+5oFo+tZt1xdByKIUbmXXgs7TP42ZO2jBXOZDvQhliCoUoAmf6Ol87UKTMxY8
oxVQPn/OngN3bS/+US1McdcPEaZhhot6nHQTYqdXqyN7edAv4DcgquD22lUxnX8rGvfPDG3BKVMJ
SIh/dBB2QWuwLOoU/x6LY9m8s+dpx4e7F0R0USzDf1XSU1q6vtKmUj/ibRgMIqDS8Lfky6xV/r4a
LvJw8TuFMIkxfV3JvINikar0wSXejBdHsKH63peirhTmUqDuEGct/En6tcUwYyAJJ/Dvsoy/nI4H
W1ehdkwdwM2GHeZDszSJzwVFTFMFwuzBPiYlebkVMS3kOqeZBS0QuxUjUdGfK+OHDzmjGB27uO4W
sbHR3To9QtXfQ9D9BHcoH+od48reg8rUS+0PHLE4d57uI2VlykokNCCLxhpJTfuWnCjlBB7XXXM1
TXjPjsvx11rnwNQSUN4mJDvUmXZorVZWJdtyMydnEn7kllNQdPw0eyyMx1Nl56Q/pvkaV96XFoG2
0tgjsWeFhzjvRj8zG6IAO/sC808Yd2/bVtVXYbv9ebT+VJboYVjEquAR5/O9nBIX6wz5D/9IEQkF
hmQtKPGyTUu0qqiiEV2KLFrb+FYbPZtehsnzW2nnnmq2rnnkW/d3/N1gm/xyguGRXQaIQchvy1i2
egkni8Wy0gPA88Lw9O3YXRY8xemRY/VrF925P+9QvZsiZm5qL1/idVHCySaDiqBBgjdUrNDkIG2w
AhE2tmmNeBHh5KviWZNQI/3cPJzV9Ompu00oKqDI3yX29jn7zdHyrIYX+bGHs81Iz6r6UPO4o8GL
tU6hePcjApEM/MaSp80tbU//6GnKtXdcR0xayoCmLw4PeZPZjHZ2uNzclcYLmgYK9zllgaSSx0w5
8GTyTR29dwlNTgTJa+3ltSKqOHeDXGJy2HgwGS+KPW4DKFRs8QpuUukwooYkyTZTSncRJgFU8ZuF
RvxJyvS0g7ca/qpnJE+qyL7U6AUvAxV3uG09c5w1OC/8g3TP3ztZ778gg8C2DVxW3qbLaQlYRLhK
BRAXyLrSikT8Zi6OqfbmxODsLzbC1i5Si98Z2ncVYCb1HktbfSqfNdy4BBCIg6FF9ygd7hbY0KAQ
yvIpZs+wgzAg4Ca/LZ0iSUhfOfa3VKIx+DmgjKGKgZ46vBsRg6X9mRTeauTLs3zsmbblOV9iw8n4
a13ZzyADu+sJ93xVZEJ9a+j7Yn4hEIc3AHCh48HxOsP5Efd+6o/eQVZPyrAnL3sgrAZO0ewpq5As
niJlQjtKOn/S1BhfUgAHQEdwqtd1lkqLMLJJXD0E81rLnHzzZLQiIuprbHmAYtnqUNCi9rCq/YZ3
0EzJqLwJsgkx5PzBFr4CaVIbL/2b/GUGVV4vn0beGJ6lTj2AB9r6ioT8wSbAir4JUqHn0etVaTrA
ch70KM1EJXS0ocdTJQOj7xs9rG6AftL/Fu/Q61qr2qHfOVcmgBHEGQzufG/clVCrKhhnULnO0T+y
YX9QwDWSptsKlsZnbK5cOuWM/O1QGe+cru4SaMChfmjDKOXlc42FmV6+YC4wjV8xu6gfDQwSW5oQ
bEpZK+U6gJmPshr4/xCOuoPEAWjTF4mzjPM/Q3NWC1KAGyY0jTAxSqfBpIdUxlmzIpS2f7gBQpcp
8B2qjy/iqb0mBQzizH9aXege3FT+Mtg5s9a6/y4R7Cj6jDju35g5M0rvJziuKvTAyDJuT1KGN7FC
hP246++7BQWpJnGyqILzbdy3v1myuqK7iPTOU+IpoY/z2IcGTOx+Nm6/4WK+0BnvhG/+xn7Rrkwa
/W+BAJmh6SNXJfJQlGGJpMJR1/1aW+il3E4CIg1Ml+ijfCssXHEElYNVkiEi1g37S7WdgoOKVDwh
b4RbCklhbuqa6nI2FvCsDCtsi5M/uBI/mry0h4+mnCBfgBo/OxeS6G+o+g+PB6kwLZ8To4QFpCYd
50gxKn0nvBANZFP8qTko8RRcQNBC13gXyWfyKaw+ozCZQN+x8FhGGRHGt346TCL7zmkBgbbWKVgF
RSH+gD6Y85xKEIe+B5qRCOpOptfdROp2WRWw7oYi+PWTf26FZRt+fRZNlfJQlsJPx8fqOacNhNen
Lf+tBUZweZZZpkdo+CgrFu2lV8Rnq/aLHDKGjRIfkOMBF3vs3eGMYV5VdLTrvVdSKT5PpyUu2RUJ
xm9eyOsnv9PTTs6gb5lIH4tcbAxQbYIHjBTcIWhk32J9vCQpzhroEQ9jHlWJQPnbrHd893KadiB5
t1SMET82/q+Lkle0dqkm6KfqnXXiuxxusVo/NktkODPRMSlQS816bkHgSWCRYWnqdhTsAlg1eR1L
WC5xJ1S6RwjoG6I8c/ClaoaLZ13GCsDRLj6aa/JGwSiJOA3DBxzyjTGZdKM3VCjw/DTLgtmC7kDG
vmMq9/iPpkuIDQIT8b0IdY5rH0QbRNW/QMSG2JuRgujCqFhL1hPnjl/aGOo3df4DT4ydm5rNW7C6
DsVasXhZKtdOfy1Hb6W7z+11ziHaux4wlgCOdL2Rl9BpZ0GfZQ1zxoI97bFsvtiE6nJG9xZzATDu
nbfa/1yUQjABNgth6UhdIdMQ9PY7AFEHA9bnz1jTY+Jvtq32p+BBe7SL+/g4rEdJGxd4mE9feR7V
QMsdGOpD0tFGr2k4GOqTWkAHQYfd5F6P4vjiUoAILnVtt6xjak+A5Fgtcx3fMtcptxLfzSaTTbQU
EuHBF559psu36iKZt9UmJPyMAzcAJpu/wx1na5VbufIWW3MY/fikggV3O4i2NMLJ3ZvnBtwFhXdk
wlhKvX+dViqbDYMC0ejMtkAsjUaFFc6wPaB5YUzVUCep1UfL+ECd7VXDSuHtplH/ZH1U+ldsc7r0
4V2F3VQcvJ67mZF5lrBKYTSGEyZdspe/3FkPz2W8CP9vKVzXHtsvY72/1XDtwnVd+yPgnW7jA/by
PZzrplL4LlSkExVMnQVV5PL58OPaJN+dWRjDkg8bs8VJo4bb0sU/II6ycSQUlb3T3P3ZSmoZr+z1
uKJvTAM7SSPoYv/lKCjGEC4BeHtBixIyZNFzX1Evky4zFDBySowWHPekfHGRsm2FV17lUnjuODX2
ts1GBXqkOpH/uBzMRpOzSRlLhVx2J4gGKdQjeNaC7gGJVpa+GpnEUcixPuwzbdG0v/Sc8kbPH8uD
UqYAjx6o06MSqXxhS/KBKix+N7hxHB2RDqGFVBA2DYql6pOwIGKtvqzz/3MZcOhZU/0ljZrBE5uw
PJ6IHGnxJWMQJr2KJqmKg+bOdeJlkeloNT3iyOTXe0x8NPKUk5AsH12UVIvIHwvSxFr4Lt6PwcMI
Weiw3XwNL3Tq5Zj8x7GzdhLOjKh33fJEH7ilmWVOO+rH3dGxdUxsSmbU/cZlsZKX7Wx+0HUUWfmg
EKy7Nshu0fklH4QheycEn0T6/XYNoEyjcNTTrwvv45aZjnNHZTwdHJwyvOszq4508h1j+VyhOlXD
lXW2kwNhEz9wsJk9k+8G5upkvKA4TPbjBc3HBRYfHrXVQWarCnfHmCmczGxC3jjin/qKsELM6BW5
OUGo8mlcQrzVLuCcIlINtrBKELx7O/dS0Wt8GKCl3FgyMIq0kiHE4UEQZtctVRIr4ABUZptrfGXy
YsmKMnoTQVnk+SFumnxf/qdClYpBlMH1WpNWh/6VwvsAV8dG4urbQPfzUE8XUOCi9sFMH67XeLRQ
/r5c9GPA2j7xT31Qxr+HyF6/sb4dzyaDm63lN4SNHEEf2It0LvBT3/2oNQapbk86oziTEJcPaGUi
yjBN/DwTCiqxoFr0/vzYTY1HNqLDY/5F1xQ5R907JSKvfl5C6Qz8Jeoq2J03RlAqzepIY/SVk//t
YheHMEG/WTSL+XEgqJz1wzG2WKYh7Gti08sTAq9xT3aFsWC3CAQTVZyLcnvIHHXJQEm2ElnuvaNr
tMT/2fXjqWT2iARCrondSbxmksHeJJW/diADKKSLCN8BmgWeEKHZzxO3sRFfIepG/9HfT2YyeH6e
Y0JQsM6UJWPp5Yvo/caY4XpDQDIYp/sMydUJzgYdYa7dcAxso5UmKtRvav3QLVvj6ftB+mW1M8SX
HbvAuXjyvSgJNiNKluHfedLHoxC4oHWbPWmPnBmIWwn/5tbWxCqM+aFcdlwRG0sHfFoc337z3OUv
QDjaoA5ttZEdfblkKywHEmVObMMm01Mv9Au+bpLb4TwBd/mz6ZdpFf5cCdUZbkVgWL3dVG0xwS5Z
SJe6p1g3p/fEydrvsWpwO4+y91SM7dPWoZy++6JZcjGoe44OtSSktavOUrpbKOIJmi3mord9vWVH
cBY9eQFKrlyfCOwpNH2DdKRn38eolQiuJDhoV6CGjNxQGVyK9uZuaQWdtpiMaTcxBTK8uVuhnPJM
7kCIWNqqB6h2lkhBnMwLa2qK2yNM+WB0/4stbsIo0Ma+c72KA7ThlFlPi2wC2LzTqkwjjyjtelKO
87N2fnbVaP20VWIrg/rgzHzcl7yigHiEkD+feP6X5WV0w/wTq5K+LfakIg4RnsHWy0kCzQ68p/w1
DjpZvw60+0lGJfC2WZmfNJhwWDEotMBedJOxFWzl9Fv5aexzFd+uOlh21RGq17ryX7AQOjdE5RVh
FwGuQ1Gd38lCEkPVONcBc9TIRSNn+J+iSKysfFBMAq50N0wYRfbfxBM8HDT33Cy9DcJvmeuyFSkq
6e5YxMz4V0vIjRUj+P3yswgof1hTj8d2rjCCjanB1dHGwm+a1U0kkKMAKD0zC/DfF1lf0LWlfIdA
ZDsA9iYJciYVuNireGSnd7iLkgVn2TZulKMOBLR9ARwJTJMCGiKGsdF3rYI47wjXGYNuzq5+Mz46
xNYLdPcJx7L12GDzBqOiEsxk3YVRTG42+bq2T10fUxCd0RxKXNgHFD4ommHOoAC5Yq3gLjoD8tGQ
KIf8FwGs7vWbpDpKq5UZFV3zs4OwxEdzq8iduCETD14XSVjAvDrJH5xWYy66vz9uNqTFiZ+EWiyj
GpkIVVWF6uukzg/+E6sZbYHGcz4ihL4Admk7CGbY3rvSBFvqzCCR5DkDnCVhkEJR/LqO35W0ZEpc
7Fi9fp5DZAZNM1PVAOhsKceJ0A5sjon6BjGAPUWpolRwptZaYCnIZ2nFroQxkW/Dd/aVbYtgnhCH
KR9D3GkWj4lO/0k/GgrUu6uWf/z0jnBV80mFUHYydPrK7rkNicekv4mjV8JkECy3VJjx9c3rkZKU
1G0Zd7PqPTepSjpzZIKhaiHsSzxsqH/GnZ5C4sSVEsd9+nnfm678Xzh/LCxQU1nosY2rnQpf24g4
+5xdBqv2qE5sVwdZjsI3rSQoQk35MnxaO8uQ/0tSDQQ71zBcZ8w8x+JA9XUFOhI4iOpHq7tHw2v+
eqxYJgL3LEHzdOQmZCmS6YPyFHDqw9ZAuvItOpetcwcyBoYNucIpr7olp0/oAMm8CQn0X/fVECOp
o7juVZ9cFUqGnacTjATQcaQHH3oDgfoZTZxoceRy5sWsdX6nAMKbjIunrZdoJ4lRy4eih7c6oTds
yGeQ1y8sR+IW3O9oA56JVDVuYvP73G4AS/QPVDubcaqSMR+m4G9sOVJELO1aGtTWA6EP1K4IrEhu
zuoV5Q2fLeU0O/rcDvdNkvWozWC/EDpaBVFdBfvpwBvQd9yIB5JSRAjAfuDlPOpr49NnbmyJifSr
3oglUBnAXCkc2o+8Km9xC23+9JGvzm1QoOM+lbG0UkO7mQrs9R50oc5w4nClBAmLtXB0lohgsdc4
QrGkCT/B374nLeGmiksSarSgAjNRERi7JhIzCS14caELn4fAoyWFJFdmhEPCqs3o3F9218LnADTv
bMTJjg0qIsKqdUd0ifV8cVyvMH9fldgqxji/KZEN12rmqA7GucOlCyvxKon/RXHxC61tOVZn+GMh
fq3sQYnzQHjn264XGPbKG725eNJu1tHqr5FPDflIoNwEDIIlLvHw9LbAVFRg00fTpHdHSLXi1ggu
b24nXlVQV+uWgOeJOXJv+2bzPPai75F9Hk0eQzt3qaEmg4q0t2wxvt+yCOK99FmtHPLuXuHYssUX
rzR5N2CIOrB50350cWbNq2lEVKOh5s1pTX2o3QcSLCQ5ZUtv02NWIw4vBkOepVrPFF9/aIDKSWLR
jRkw5AipHnqgfWVrqxnYb2ODPVNLxHd8OWVvyLVPcgb5qclRPWm64VDKM5t9RLLgQyMrs/hhKVPB
Sl6zvaXynqBRWsGrR93qGjr51WVY47A4yaJIm0Qb8ciy67s5b2j0LgDzNBw+Taiu7LOIpmO5+cBR
XH9gD2+eGBEmkcXlE6tdfbiIVwlzDzagwoNjOCj5X/dq8AttnVALwBdLbpRmPFvBLAlw+L6qnape
tpKDqfHf986l58lJ8wVDjLaAukuTUjW5Ue/LJPci7vDFeL46rB6mnH13a+tX3bO66ch6dDnVinps
cFOUh9XRwGCrNmTdaZ+j0X7Q4ZodsTnKiGINoYVjP5fB+FinW28pO0xbEQckCG4+Z+t5wNlUfFHa
T248cH1GXvH7BU5RWu8+en28Q3v8L0jZzHBpFyQlgULCodEMoWoCtIEAwdSvxdwUAdwJRqG1n4Yb
wvnsUrgqpqnx0mU+laPfviDuyAf+7AFR3QzE5B8DDacKgQYycEWPHEOqp1n81OszzpjjyMTyyhMs
NNnYbuksu5pR/F23/pWq7rnujLNHXQm+45qsaRo9IWKDAcyNmptGyr7Ff3OrfLCpRJYEdqWAHQ9W
ZBlNTnOrSt0WE/16tbTE4n9qMTOfMazzwwJZIYgNlgaffFh/cg4i4cbXB6N9Ft/8wjQKFCTduPUF
QtHmEedVxmgVSYs5nP1jGhSjZ0zQcfBRbhtyqCGULkSBiwxJV5Bp/pRcecgZZHZ03fSkR7B7mSLJ
K0GF90854tuZ5UJTmYYf/ebjnh7IogyRNMukje3JqZ+ez9JDMpc9y01B+xivKVdrmgWFSqVYtJW8
6DBPaa08A8/k50AQjl6dz6Bj+CdVEXo+Th2ztQ8SE3P9v/laalnQzJW6Vny3+D3+b7fLe9P9aNrZ
SCbS8kaSx0MNKJ15HnL5hqy7KJIop4/Mj/tTa37H0fjsDpU2yjsfJxzBWd5/u7oKR3aVsZlck7Ww
4+y2kOa/GXaxrwiptdW5+1q0CIzdTG3yud9XH6ZgD7Hy3czfpyIwe23VNpvM0y50gBAmBwd4mkOX
gMkbeD6Vs7lLq87x5lfwgfKo+/29Af0tyvnQgA8DnR/smAR/0HWgCWq/zF3Cf/FGq+u0nnEmKHHI
H6YvVuQMWaUO7cJNFEWc+E+da2zCk1d6amNIRAR0l41tISCiMTnuH2H9w5k5odgrCNrlt9VNK2b8
okwgPBZic2T8PIjNYlx9nCLqtyPIMVi3BgNXMwiuRAJc1avon3v6zH6GrUe3ENRgQAgzv6xxNWo2
Qw/kVLJsjnyccQIgQgqpArAJEhrsTOSyIyTCGB+SL8os5LWEM9EmSa9nSQHQKDT0O8SnGPjNLA4u
koX6VKNL4gjVAq29QjUD7Q5h/vQby05lGahGZZEGPuqU1Rq2c5iKKzcyH7jhw5iJ1hvVi0dUvC4r
hjxrlk7Dz6SZTBJ5Mk9ODp8rsxCLARB3TLSk5ESaPZpH/wpxNhCyJYyNwu6Lzy/j19iCg27GYmuO
1HevQpWZFKjwfXX9pXbIsMBFzFGg2GuLjW5b1cro8n3RVbBkMTf875fpy8HQWkBjl+sNP0Lafo3f
oKH60X4dfB/g99rOXIrzmybrA3cgTdp6rNQcC2yWA7US0pxMTypSuKgZjD/JOFn97O47ZOBMnc5C
ovSnBazVMW6HtCPY2I9yp3LHvy+rwZDFetCp9aCt1Ys8ramsJGjXTHTy6FtX6NFOS0xIeuHUqvQu
0xkL6Ovam5w0XwIUa6DdcUJdxb/tLkWKQO6G5mRnDi8LnEsBg6TL904RQ8co2Znxo6pi8T+zMTjM
mlhpRWEseLmL0SpGcMn2FhX3WnJUS8CpN3VLq/hqz2/mzeOekviz1lAA75mlCFNacUln22SzfCqE
iTr6plxwCpW49SzOPKUJDJL1YuvxkDzqoBB+GIAvgjAVGKRCt/dhCeeEh+izZIKTnI4fdyz+4OmI
oeJzcSNeSBiV5v4xNKCW76E4kxPo1zyG8UTvxDKXaK9jm/EZn0D0bbRPhaaIp/1SF4rPgm/XnYoG
42Gm/mPW0z1B4Un1EH00WQO8CPFmctS8mcnGumQbrNGL9p2DZQWPMBbs6vRiL/YQkuGABqSCxyqo
tYhEhoRadSiiuWaIyn72PcU9F4/h9MI5qxu9zmNU3E1gB9n90XoyUrXrC4xYnD2jiRdkF6wLqxqs
6jIxP7KPUhcTKp1gDG53sk7IUnTuM98O/BoHv6QWFeXlDM0xAIeIfXALUizu5ywdUZdAYxv4CauD
aVEjgXy4oDUnaxOIBP2fNmmokJsSJs6S0OBnLrKrNTpujKs70tl0HH/X0dLYpyRzCklyZjOj/lA7
YrDrXgDbi9cLzZMFAOkD3oNVBFvblcL14S22z8m9239Ck6WA85TWT9K/hOT8w19PQr+Ekj8UMILm
yIP3KDJseeD2VivJoSF5UtgGT5ZwhkjBnI70UrLzm0Txsz2W0SbhGOzricdTiXwpg0Dk5cgl/VZT
vRGVacpuguF1l/s8s4lbnvvCMuFSvLU/X1nStxoTr7BsRl0o7SCJLBCx2HkW3sBj11aDxEYrVcqR
hBss5DlaVy7X/qFKONjW/q7fzDu3OpqsvudU7Pat5TQofkpxIj8391XYe7nrdNHLquSpc2smfJcU
IlDEv8Xb138uWYt56/RyE4qfLo5usrHRRjdQkLoL0U2UJmndH8DVH/3EwRoRww0KubMSmRsj5d6/
dqmIansfk8SE/TbjES1ZpK5nKEfo4jSIw6xCWfMEmfcHRF660Nu7V5ZHNeONpvy8VTd1e1hd5Utc
kuMEm4dWqAfgTMcE5TUzUF+5UoaFM4fu5jurueCtWL+OJm6MagCSpWHABoDqv+z76LTQpaYoNCjJ
QEkcTqk9uO5YXwWHE/KicaWozOhkGdEZI9+BZoXr05KodmzEdJ4r6vupywSnADC+tAaRiqLjv8uH
yxr8tYlsaI9okWaIezARn8HkRkG4Pqn9Kf1PkW7RL3NHFY5vKzk6L1Pa7kiFd2EPXmg2DlrZ+ivZ
auJSvWk6iZkzTtWmsPI4jHWXEgLyvIc6eXPm8YRaXSYTAvHHas3+uI145WPg5KORKWbjiLes1SBn
39KN0Ey9jbOUty+jRTxK45Nvs2cHpzTnMFRz32ZkNn1Hv7cfnbtS97IzyrnYipFGMqOJJD5i2eRZ
XxzO5c/6yZ1BRLPfbwSlA3y9ZkEzlcYMEdZ007FByt6ElZwuPRCOsUOWlChVm7Zega2NHUtrH+3U
VPUWHj5UAVD7YuYrfL5K7s9KOTbzIRIhBFo5COqx6ZTLm90ioEwyFRF+mC50lwZPRRj43lj6uW/8
gsPifPJlNiT+MYGHedZTsXB3L61b/9BFyx2MKFlhXv9aEi0pA9YSBVX34TUHrXYNN6p+iO7uXd+/
S9TCrTzElVol777DAco2kmSqP36U/xFW8buN+QgGa65y9pF+4XtAp87Szxd9cSqT/E68IlrwI0V2
otCpxsvbrpWPt1zqNocz2Bz5Cubbn5Wj073Jhr/xOGQCHIFMN7X9C5oJOqMhWLOBbd2pWIYWE6JD
wTlnt44AAsZGFelvT2J6nUhjuDQKm5vaFILBMqJitS05T1vGtOVJEstCzLZgwDOEU0RELlLez7Ua
Gx151tv/1VVF1uWx8xNz0FtmgpItfZCapSSdcqocMaq3lbf0/X/+vimXXmjP5QCjkOlKyg0ht3pr
iYRyEd84hvfLL/G/IUzhV24GmBgqb+8nkD0EqSnjeBIj/HuKFDPVxLlDlYoWnI5cGkrnmghcD5/N
hTQqz7qzJkvmEhjkDFzcS46SUbJwUO8g9WeYg4FdPLL1f2unXX4MwfjHHzmRuJj/R9lAlesqCpJa
rl3A8AC/dtp9n31rSxIvtSNmhmXfcQSB05k4WJ9N4Ho5NLquYiPMUyZfsusQkEU7w9kxtKq24ctD
dCXtpcZN5HxGmq5Rdy2HbF7NcNS9WOiSEPT2nEjhBaCLhYLkRaUV5CyH19yUCLRf9NXoq/AfI8DS
szaWrwVftW2ptS80xOObQfUQ+fo3O1UgMfP1egwJbeGwEprST1f3+Mt8R1RUlKhU1Hut8lNVayok
PeHLkBU3+kycLx+kCw1nqvz8LNKHontr6F2GtNAHaVnQHHqRzTHDl3ARTDiTxMy8Hv7//9ogGgZL
8ueM+jmY+MA/ewkdgsc8dmcxfHHac/ZQtpBKhQ2ws3Py+CLWvlrYfCRcFHI9h0NKboFywpj0IIyZ
mOu+q9j6ApfwhX9c1TRIOjOtSHPFmeDgpgTC7+WEIq/Ks270Y8lL/1zadLkmA9W7qjwybzZV/DgI
5WBn6P73WmMOTKU6ipV3ckPr+kULIvwXWgGIcRvz6fGRUhGq5JupL4TzOht9oyP1MOgbT5hMx2Jq
QjTQMzS5uuGZ4Bp4CSW2atmffOpW9ycIZV77vJa+MSU2lgbFmuqRJjEgT6DnjmPJDAt7sM+nZm9J
E7BHZiGjxr7NBuNHfw7tv2ad/OYlKBKvYv6TQt5yY1y+N3mSexkpXGZGadlxpQY991tQHRQoCVJG
kVmPU3w2lYeFpI51t6DZIhb5Swn+1fmb874lZVp8JEbT60wdAvToCitqAbRWSBuz1OqIFxUVnUcw
1nzo4Y6DzLWcB7DBQrtcTTHlxoeLnA+srs7SZw0PCstCRwnAu9jyL4xDKIOqR783EAPh0cycSxjh
UAsdMfZMYm3HIO9NDoiWmPxLmf6NCvA+RxxWyzUf00GOiJQ5JrpqX+nkUddjayuWKlTmMZYM84iI
jSUWcqxckATq+H2bL/jSJX+LaC7DHMc9HgnBgi3PhrnvtdDbzSDOL1lKuwGMpeV+ygW5DgveFM4y
yYrWV7GPOMo6GsGZgmlV8H1ZsEz8WEKqzpj/8ITB744pSpMLNmWWYFdGtqm7NkoP5DV3maOf5obQ
bbNSmlaq/9dv5ZJCJ04H4cyQl37m4J2bfTnsDSUsKqTbFyLvEEZ+CbPXMQSCnVtUgh8RVm2+GFZ6
hEVsL4gl9BBJyfc5xgE05wj+yZ+7fRbnD5D4RwDY3mjHOed6MK+n3OYXYuoMhJgifC9W5hY+lD3I
6NVZ/oOUXpRunJVuQ5+Wj0AR7RVLA09FzwaUzd7Tsv0+hKffBZeJS2d+usMh5jzvDdBlxdnNM058
0PmvOnqYYA5sT2wFrs4WJqSheC5SPCw0h535DM8XtBb50kXGkyWG01UPGFd/VjJNJmpMJyLiKnCH
6ao4y+7efh6fLgv7iz6Zhku31XXgbIPVcHVtG8opCU9nO8/weGYqk6AejWCWATXQNkSwo7VgKxmz
zJYd7exw89Vog9jtL2E9NuuA91DlusUBR3aEyeI5BzJ6u1qwopcYaZR3yfBv6DwhmddRuQmlIm6V
L0zXsgtpZzYcZLG5vwQK/lINiqYYfMzr3IQOORJLI3xH3w5otdok1FWT2WPK98FKBh0N30Zoyqe4
O0zlE8o9wKe4gm3FSUDODIoPyJlk7zwMfvlqqXNp0Q5dlmFOjXGWFRmoTo8qEu5rWdys0Z1XaQXI
7eBnq8Nc1MHPxQ+xmZiKq9QunrTE5WzBCo1XaHvN4oA/RMfnPUzAY6hr8UrfquiWuhWj8OmZ5JWa
Gv4tbHhFpwotMp9ntANgupxdPhHmHNjJFLQTcvQv4OLIXjnBtQF6GI4f/yNIVjzXNv+nHdfWX2Le
oVPDdHHpUnd4Mdc0sjQ8mBcBFvRrwPw/0QvYBBxn6B7mr6+pQYYPGfFRxB/7Jnlz+yhtyvGPc9eV
NLYodRnCK1MxOElgoLcgs29lrys8rVhu2n8mmEyfRYezDRKZCMzEwlQTR9E+4AXbQSaS67+7j427
it/UoUx2Fx01WWoIhGMkpEPIqxn2dtOwrLGGIzh7BvOlQYjoXEC1pmJLxyYV6BoflyLod3SN3ss3
bcYxJReIQ7aDRH0ZtV84ZVghKjUVb/bBYszgQmEG63EJCo4SdqmW8T+gqdH8obPfi/Nu9WtYgx3L
aZsHeRNyhP9Sfdi33431Wobqqic6e3oAeygHVX1j/IsbQxO+hZirDqL/4/zV2mVJmsUvCwTk+GWc
sW3jjjfGs5hO5D6nXYMkhfpPwvpCYGjGsG8ivTk1rWTid4BLZ0DgXgd414MnW++qGASw0U8iLdGW
yirsYPevr9uIDujU1ImfxSWUN/BtVus/05zo9LeaiqFKeTwKh06d22PWJiOmBJXBigVGs6SGYS2C
gGv1QgybZXJi3nuiqfciuVf+UkGmVflGE/3V8STksVGSXrcog0OwBTJguD2Ccw8rHhXmFdjN5IjP
F9vvUHTgXnUn2SpN8qO86In8B2hro0vezJQiKUcHccAam+OV4pNxCdPtoPNyp9J53vPbh/pR3Axf
xgBHdQIQN9V0qzQEKxFsSwAwUnfa6RmlXV40scldklzHVqzcprXNnHkKIZ8LDbaZjzj9fQolUKPw
PZBoLsGZOVS3Ur5mLQtUhMuvqnloLU4JtC6xiY+n3QYGuPLhMk9wY/08gXyPy905+9fvYo4IUED6
TgK0VXj1jD+o2TP/tzoZy8ZbLGNequzVcOQigrQlUGZC3k3QvM+LZe0nIQL4/8yc8lg7XcJa0T5F
gosnSniEV4QH/xHfzLDS74bYonXzkjVCZwuqYEWpwb3SrUIqckqRpXXTIguCwzyAiiUw/YoH8ouT
oILOPbkKoDEBTfHK3Juivh8bTJ6F0MN9gsXWef3OSW7/2mFSo3m2686P4uhrfoTRKYg6z5dgTaoZ
v+SElrT3QbdUX8jkrYep+3dBw4JgJP7WcczY4RbOk7h4wwaCLPy/O8ln58utYy7dHGJyChWltGjC
EHFceBcTqmL/4ly1GGDWsL/njVsXHfsAgW+Bv/9F8N/Qd05kZpt4ne55TkDJA37vjOtXe1UC0rfe
RFChyDbdyvC3NBUqFYpYlc1QwgAWguPnwbBpmhzF+grBJ52+iwVuGLQ9AXa7DjAzugfRxWeyjjkd
eaQ0QYNXL0Wh9z2EqIIX+TM7fNbiJdsp7Oe/GlNeQC0m0YB5M9nEujRf9z4VHj9Kd+MUBcgU1dio
aWIeWJ8wf0wTdoyCXUbSiVJpgZNVMHVqUJCuvHdNreXM8dFlwm9fOaLNvQdUIbmZkXuk2aHU0GPZ
VoLSwisdvry4ox0UhNsRFEYl3dSz7iLEjUC3P65zosbFJwAC0IRzqbRpLqTBxObd0ZBqIVXHiQ5C
qsW4neyaJ0mizi20NjUGWYMRoFu2xtTLknI1qkVHocuBFDzCt5H4Rp/NUcJOYKD/JkXayY46b5JH
bhwJvHqCyB1jCj437m/yL7ngTaoWo8sUePxGmPAr8Jb6tPmAkzGQzu+D6dVKPAEAPY6Jfgt9kIpA
ryJzKFiEl2VLgsQeno9PfI/xQnPQYzQaDntgfZyGG1p862Ba1RSUGGK9TQ6Qx1eYNn0UXaa+itSz
eABfmp6vl/64GXDQDigqrxoMEiCVujaH4Sk7VeyBcKwme4MPWenvpY75WIPqJpeq7qUQODTG0QGi
sZPU0VYYhx+oMZgFaSM/DezdngRekKLompbxlGjZFBo5y5115GMbNU81TLz2zgrHQXJmUISD00Ra
YvEHspWQtoBK59hu4Vmtp5BAj1q3xtVwKiLQK85orKQu/HfGtl8H3ml7qPg99y5VgJKY+SOzOTkQ
EIY7IMh9iIQIe/GUoXMITHnUgaONipS1FRfLgJsXDLI0+PgIJGOxUWGLQc0GqPvhl7xBbiJYlxbS
WUslMa0MWeRJSk06Ay2fAfKSZWp//3vFCrqggjuItuDO/v8yJaV3MebhoVjdJw6IpYPmXqRRF+QQ
AlZhPR0wP1FFkFELJ4KPkaBBAc/hZGo7iZIGT5kneBmgguKakxIhGNen9p7Q9RLSXx2bqlXXzH1y
TLrvsUwoxYsbVh3S0RtR+4OMgwdIX3xS+fugO2rmrScnUs50Agsh1J86WcDa4/f9ujv3mkBWFWmA
BK5SMtlHJ3w7aKRvcbZxo6fLBcaRv+RwEcTSw9KvBhMTjiTiZCgMWL2CpM2LkVnh2y2+4oNSHVE7
hhxFGIhRGv+aRHLoEVVfRASF54Asgice+j11uPZ6KJvMjcvRKiGBGIu+EBXrNfNMAzGZwBjkHM9U
N5kA+XR6RTABQu8mzi/W21e14O625S3Ra3WKkYRJ9ENViIeB6yA85OafXMeVu6NyDJld4p0Ugy2l
Osm5IscWktH0RuIYFCz0sjJST5cyzGxARHfs8eQ5wdd2TTKcw9Egd05KPw5UgU/1Gy1sdFq6DdGO
G9gNy7bzDDW68UfZEkEJX1RLUVOtV3bMqiWSTKiAEoV6ayPWXimYw3Qk1to27sT4lD6prg6nf8GL
DGcTY9sUVU7t2SvRxSg5o3NAEEgG5S9SYo5CWKmVM3HEyOvT2WJHpY4siAiLIc8nkI1G9mTZRSL6
QbovS9kU9gxZvaQvpgkmzRr8Skolpqi7cZ+ZbrJwEQBZDJ1kYK9OCA+QrAmgSzR0E4EIAYv3WKuA
KgZS53cfv6QNl509IzutnJEgboxIdWyf9fdROz9PsukGTqCOrSgAT3Q5z6oL4TpkMErdw9QuTJVB
NGsiRfklGrQtCbpdKZOXTMwO7lGxOw+AHWajgP1Xf5+Pxj5QXmHfmcz4HivLqifQFN99o3tmV+0Q
EjJm24hD5guFq3JvSygisyXhqtB3mx/B18Uzy2ajxgTKtRAzXhFifvdZ1sJeqtmY8Izma9uBhuoL
F80bmRvOiW92dWsS3md4NjEbXi7wVNNqwQQbA+UMJ7AuH3x+EWftDs28sxF00sPKygEtgnvoMHn7
8QcdQFwil4T8rgKpBubgo/nv0Or9bcG+bxMGhzDfCzIU9WLoOIu/UD9PkgzIWAv5s/v/6Arlonjs
P8Lse9dTh/W82exnJfitfJLm9okH3pinh66gpSzN169Y5UyLc5+cL+wjFkj8Eu/3hFs7UFmglord
dJCnRHZAn1AR8v8DUoWRpjUWmd8/stUBeZ9Spkgz22ZnE/Avm7LNBQfP7G17OG6TFqY4Rx+fcook
El08DqBD4AKaMzU771/i3381Ct5pbdVZkZgyFgF8nJjS5dE269V1OHQZQlayu5kXn1+DM5JT8Jeu
++q8n6notk51rLJOLxjj2QKUGewagBvsanig+mh11Jrmallu/S/x37XxubeKPTwBmpVpa4Y5hrie
dn+tbLOX5Vxr+g6B8eZMEHiWBOL2L9bdv+AfRA9WiY1kQo1pRlGiJ2+FuTCsXbOMIhlCMUSs5BGq
E6nvUzPXcx/XQ6zFMtTkPHg4VyZtxiT2FWC2hgn2k7GaiLO8nzAXb0gTwzn0iqP4Kd6CIRVaNa7o
GHw6f6e9kFaDgIBW0WKZhHIvPUm5DZ32aAOPCK135ng5U10gHhHu3M/DEjecq8F/Fh/iig4IeUpy
Hho6zyf/CkrH0pY9pSA5TuupQfoi7V9OOdaG43BVEOlcp1Bwx/mHP8wNvlqec8BvRRfzhYr7QHjU
CWdNhAl/i8LvJ3Y+ZOSNE9ALFYBYJMQ9C7UPH0mHWk9NE9iIZG8JJU54MkFZEVp/hVabXB2I5PZP
ds1JNXm7CI14Zdev0NcL3mFUfHo0XQP8eVBwGf/hwDBDVaryvPtv5kV+JOQ0NSo4JyjLEeCimgTq
Wmp3TCcIkzv83+DeDjpkErRELAfwL63SuFHQfndXdZb8mjTHq2WABiwCYtsju2UdbPIxz4eErsWL
2SpWzuzAXkQCB1U2cEnPG8NrqxMNNaoLImOq5l5j+pxW7YdW8t1PunTIRahSdw9D5fBPsBxheWaZ
ut+hPB7jnPawmp1JQCHOLvAnB+xkWgnBr8ytib+bxAbYJHTmHpgS6Ycd8TujV/lwNDVBZD7YTW3L
7cUC7Pba17lFj8r2uvgcUTLKjb+MqR9pDBnuClQNbBtXkTcJ6AWdi6loaYuhF7aFAYdMVF6eEMSI
kZWB6vUB4GE5dfVdezpQpbySBdBE1k8eC7q5W1bcFb61yvCwJ/drq+xcJljAa8VhCExy6flW1Ftw
f6vtyMqRMG8C21DMrecO0NBO1EOuSkpHln/IH3nloQfRd8WTl/Jh27z+ZgFazVeJZ79k43S/ieIy
vDa7+kZFl/Y50+6cM6J+pVvHb1B1LFykNIwthk2jjOY/axM2BIH2e2SFxVdLB5aoVip2iHDRo+1f
QJiep1mdnbVeNG3xSzJ8ANllQbX0Qitxmwo2i9OVBr24b+KJgMYqamXmaGftCcPZGaPTCK4LsKl1
17jjP5oSXGaKSUYNayA5YANE2nvYgGw0tVe4Ad6omHSf980Wmv5CjGXb7e7uSqieYtuzqJSqtgse
X3Sx3OlqmEaj+TaOB3+coUWkFHAfmn79Y1/2sdFKIpNQYMLgw48dl5DygQxtZ+P6bRhCs74RNlWg
RuKKC1Noe8gcLMPiR7CjHFj8FCtJ6v8vFI90oFR2pE8+8hp+mxGF55CMbkzAEWARvNuNb+1tFABS
lreRg1rws41apWxP06BfaYGl0qAytA6u7gt9h0yKwSRUtgYmjuAyQv2Tj0nuIqYX29y7b4rlNNCh
NK6QJQxe14udtbfTnas75EISG9nEemoy1TndZYN0OJ4T9My8WcFwgQX8DvNUC5ZYwdSmVzSThfme
xpROA038rvwSdgMoNcOsDYrYt/0K/xwRX01T2lg2I92YUCBRO+qzFYOTjI0c4977S/3BTu3duOfS
9QJHdf6t0xWz1VzJkLdElAmhp/Vc6QlgBLZjez9SqAAosmq6HtIWWSvF9KzulPyvpVpffkY13pD4
QXdQi6swFNBE6YdAxhEig3whXryRyuOIJo9/8KV9ETE3ri6U1LSPP13FbKwsZkEPzhYaKdmo3uwA
bDZpceeSia75ReSgVA7FvWKrmhAQ9eGF/H8H1Gp31tr0v30wsSVp/KsUb83fbFRfXcZ7d3CLYqYn
RWLbc0pxZdNS4LIfb4f4RWPVLLREu3+DfjHewTJWZCteQ1vBy92Sb2VSx23NXASFZL2NIC6+os1j
yEmtdtc480i12RKMbeKC9aZTkuBPU3yfW9Xygln2nYm9HCEThXnGXf273RHG2MVUvn2wulS/AAvs
dbPrd8evk6Z3lKbnkgXPxaDMPdojXwlZoIPwvXHDj62QFnPJpDyrsSZ2Hh5wFqWenjqGPwCo0jK3
EPnpQ0nfjT8gXtSaod2eCRbEfGaaqbI/F0Dcie2n0CBLLGwoOLimPym6bbf1tJ7iRe5ZxsbAkv+U
Zi6MHjTqhXsNkQcqTJHX+H8jHIAOGmP90Z4ZM/NkZ9QpWaSQkXu7JEKObJOaqfg1gg/Yrp8tsSaU
fxpXmsfQWenrVH4Ez9uFMKeON+Jh8nwxY5XHxnu7CADv+gLIFIsxkNdVBgjxOYVdJx1nba4W9EB1
1pFT658EetFebAAuyuBvXktIFW/uAJumnZFdGcg1qg62c5a44dP4RFdyjd4qOWurvXJaONalX/ox
h3JXBdsrDaSB5jCu1//k7YnbaqPe+IVgY7mXZhBS/l6zgXe5G6HHIrxrsZYzLqZA0rveLKKUYSVL
45EDLNm3MaXjiDKeQ156Z2ipRXGEVoiLZ+2VFgLTnLcU9BduhyI0uHGjT9TOJhZamRqeLVUEJtj3
4oYYWhSGcLVAffQy8Ra9wwD7ZuM9CNPvODsXxeKSm97FdbxSjvTcJkBnsS/nArkjJnI/lh0y5J72
Oy5VE6vov00o4dPZ7YwRfY6xWYXBLY6x3vkEr/XXeN72SkokDws5lyaTDh4jB7yu474j2nLoYbd5
NU3uIUSJKmIDciJxPUZAldkh02Xma9KL1nowKYwqFeZyheFsL0d9VkhRck+osQlxeW7Z4xeRo1QK
cTZJG5qt9VwcPRgePaa8tKXvNbA3hOtWWu1eQ8gEMfxzJS48LeqjO9jfA0F32o3MaxoYYhAeJJ4+
5mBfY85b/LyVLyhUcujnHFOMO1Mivl306JvyJNpYX2rxT1u5RuA63pSMWuZb1ftKMGzMbU0gfJP9
hkHDVbC1Xp+7q4GdWRq1pESuD+g0h1HlVll0EiBP5O878AONVVD/Gxdznhj64d9Xb7x6sQh6kf3L
sjn1MQVc9sZl+JelAJhC/gn8KpZ6XwXDJkZOe739WaCVDyU6emGeJ+GrtVDE06D/MMKAsWUEMI28
N3Jv7HMpZohVLzsIqLhs/+P6v/3axmtgIWmmDufFdoDjari+NFwoJ9MKmVO1JhGyD/4BBbArG2rM
4w8iyh0lUN0eyjYtfTzXIxdVoGGt5PwhApp19USdZZdT4V6YDDGOXzuJit4TrrRPHXZoYpDiCZk6
VFl/eWUt+qqhmsvpeK7SKYxLv7pbbBSWm88bfWMkYzU0wGmApmt+WYUYpU4YvGTcRhHVSgPeK39j
6xFB3kb6kKKsqO4Cu8QAdgYunQQtSi67+xFHiZshJM2/CDzc/awC+V9qk5FGbNuj+wlPlVwXcqmK
xM++arz2HqxjfHULWbjQzdpS36dM3PtH2dUClBlRpt4EUtMttxvYDuBE7LPUAEPoZeEYByP4JdtX
HQIwwpPHwN19CqFpPLP8MSZdj8K2izDxFzHCG7qAQ8xbm1V/wUNgA2tflfanOvkossjfWJzgetxz
aGksO/RB+xRKyjscANe4HNPMkBKoFLLYWWzX2wuYhM3bzeRPufxO1CuTJ28RUjRPIJnv8k2k4PYU
5KW4wT2ylo1qMw+wsRoqpstHB2rIaD8Y7YOH/F9OwSDOIT0ug4huqdI4q4kmH2ZIFVKhFLqdP4PD
qzid9PaAqT3fq47A3PnRNdd3c7nF7XUJ0GIT5ttzPmSFEOBM/eBw9Bqrt+OPVXDrW80c4O0Wa0X5
THSOwT3cg7AzhFVeALdtt19DbyssrgAvBt1cEJrZjMSaZ2zGZMik2Pm41HjKEzam0SjwOw/78dZ5
yTJIvchWrIwIAQfzjc2SBLdjENsXPGmbjHIWglpPZNhDcTR+54sf3l653PU8921/mo455nUnN2r6
W9wXF7Cx79UUkWo66SLQHQvhvUnO4TKkMoUYvgS7TW1dRewSw4kMJxmeZNgHccwBmsMEH+MxCuAr
JNtIiqTynMj4WKLflEwHVIJzM3LIA2zttT7hSV2z5ZFoW3sQgiAaZpTTyPnCAG64yTBd8BhiUpa0
cKiPGJk0qQx6aXKLZTjeCjz6PuwdaaV4I9ZIa65l82yRken/a2ccCACuZyPaMJghHx/hucc6mlMV
iu+SGbTXo4YtwUR3UIcLnaXrCANU27JRB4FjkGbtBvuQUxwRrBve8G8pTiaLmiZ4n/TR697GAOO/
pTznj5KUeI1ygWVyHPJfniKDx9l/VxNkSPVfFTFvRYwW6P5dwCbMDPsBW6B5JtY6I7Dcyg+aAVrH
woj4xUvI3tn/PnTKhTAa30IQv5StPoY8+1TzmlwIE0BR+/8ovn/Xzjq6YGNRa2T2EHT7higCvA+a
TSKfHuDUIQsyOXNknk5c0FdGXaui4qdM2s+SsIhWHK8bZQWXRui2f6pJBtSxKqNb6FeXpLb97CpC
1q3sGxwURDMW25u6Srjc97eEe1nMsJoJ6KY8vTG2Bj2iHiyIIBpmWH4mbDfO+endIlioiGCrEa0G
+S2lvVY3mkJKvZRnTmYWXrN7rz8LuD+o1XJvMJQkr/YbFE3L0Z4Yt3YKpPw+lDME32+usXraGIjO
DzZUoPZGrqm+1Wc816VOynDwSLTE1Chm6+z5YFwp3FJYQ0mFJ8icKxfScFEtojtobduDWyDWb+Jd
yGVYEleTO+RMF7poolFz7IwcZUFTkFBkcN4ws+Xf6HryhSLiG/ILZe7oimwORKbkhpxeJdqH6b4g
7+5MlogbXfP1AviMnHsJjzO4Wrb2dL4gCzDm66BAMCl0zRmvzrMidHuiS/OZ+6LzdV+xGBRhO7DO
ceOSnL9lgyZThc9YmcmgLfTC+a42iz7EfP/bu785L3TypI7wKYgbaMAwbFZvUSA0Jo/AoUaknsM/
brjMGl1bhjFuexMxmll27KD4d5PNMIaaXqv7+bACxamKfyCm71NTCNl2x60pLJVkquxgOnuYgfk4
CNcYN6P6hYPMCIV/WWW2z1dOkhwxEPEnpCtJSOgXRxIom8y+n61cGj2lcCrf7ZinDiWvLa0BXls3
kZ4bMWSQHe7+ztow2v/3M63XKzCUjyrIWcofL1InI08OWU6jIWRp00doU8NvaeJ+ae9AEo6y2i4A
z9mLqdLJ77ec/JAnBserCx5vNJ+3fokzlpl/DCV5t1XbnHxz7V2BufJDWfbOo05BkVhwOReU2EPW
G9gquZp9hpH0sPc2/cTI5LNvd8LsDUCl59NH7LLQ6HExKhrqqV2x1xgWvroX5XWSBSv4LM5Plmu7
GXw8zR1x6T9RKpNZ61G2xG1IM66wo2DPBb8x2U9wcaPle2ZEqVscgl5prev/0qyuqxeI6D2bfxcm
VpsD9SHak8P+xfFoQhfx7ni0zALggC6G+rX2xtGbK5Jg8keLKL1QX8QS5VBSGukxdW1oJEBiQGHY
f+xodYfttlw9TkmIX2N2LDssOGU/9w+stxf+kNUkcs7aHyZADQSF15RUgQif5auhIdae9iAwmAYp
XzUGvEVqiVzsy7DiEzE5YNYZqhHvLojEbjUTone98ERweh2i0pbryPXLPf3S6m+hJNeFNce7AWFJ
RDMuqxM2tbO9pi+fYCtRQEVDNUqVBDU4eYVX5FhIk47eFdWXTB3vgVCPBt3b1j3BnM7EC0qlqhQ6
sxSH7YoxnM0tXvRdCjE67MhqN/qgX/Rw8Ey8MrW3mTm3v4oQiv3RVlExN8hJ+/j49JuJdxbfGche
NMfocaZVkO3xa4RdynUbyvL5Bmt4OW2pY4UMBW58DngNJBMk/T1A+pyBiTGavl9Z1kAiIPyg0CRK
+FkgG3zjB02nEavDOs4iqRzQOADd65YWBchZFMA6nIEwnJ559H+e4HjXMqx9+Ta5OiHSKqj+FncO
y/Y0nAMHRUC9dk99L1bwbMUHPmJsTheBXDDzLoTFvH6MjKdyqCN20QmFdFXhMrno7nf7RGrVY4lH
vi0EreNKO2x0qmNJG5uaTELcMapVF2Zc+xmH5EHfO275pTPvTt6N1TqIFyLRufcu/ygIEGv3bf1h
/UbiKyWli7NuD7QJR2ISPgKpY6dD+cy6l/R/1ZwnMRXILjuvxQlt588GWr3wWSX4DrPBQ6QQvLbU
2BWFGY2MZNckQ7xkldf955zdW0tI2Nsu0ihEOo0JutgGkwfkYqf8yYAIWXpjRET1HZi2OmfpUxu3
FoKTBkNNpswg+Nw4mN/aydq02R0VJosV80jE4pKfQjCHR57JXycj8KGfAK31zl6ZJos5y30VABxJ
CHKPtU9Hdd8a4Yr2WLRPkerPi5kbHuOQbNoqrD/Vm5Bu8fkFcXon5DrditOZRj+6lLSUFp7Ax7dR
HIV+WpafbIezryQZXHNIVGcwm8NxDFfUsfYUxyevCfyN4dIWSaKXj8CJbIBEdcdwBwlXa1p6P6U8
yxOGdnhCR+vO4RuPZcvpPENTGVyt7oYYhwJThdfIlvPLVqda3Z8kNp2RZbomzV30bOQq7OcaSung
sh+M/m4GsJvQbXOkId7m1IOpfUieFhzc4E5n03H1a8FCMuo+xYdsdMEgopcIBGCuOOmMc9ddEaAT
RTa6XTiKTqKkm2vQLey00brpJ7Aq685o7kc7gmqEmcsZ0aTadNffAbkEJvbVaNn09JPxfB9LsWkv
sh2Pc9lb1/Ob5v7E7o15dMeM8ktUdmGZY5SPYiyfTH2l8KLZhVCBcQwndxQv89v4XJdMut0k9D+g
lkOmE5AxKTKWxINUfaJkZAbU8YN0fVwW0bj+Ajf1bNTj+1MPJP/s3CkKpGCDwlRurYh1Ks9PA6Ur
1vP6WM0AodAxnUhJ6F+9yRaideSKIdoP2Nk3+jIVC7yZIwmfY9MFSozfqCzX1XRa+ax7lMW3cTI7
l60ltZS744UcBa1rdcFSh02BBWhgzzmKhh3Qj47NKzyFj79b+waxXPXn4XYWkhTp80HCiayF4EBA
WahiJYePyT9S7Al7r5bJiM93YjqTcddbhJ2rnSJ6M1WCS7RecJ9oKXdr5r6RxKCVBNARwe0kepvS
+kHn74sZp7l1yEQYG7QPYCufeU9Dypc2eNvkU5WGTcIjkmbR6prSEOc+rygUFhwcUOsN4ot9Twh+
lR1/qgBsJ/O54xTYoAfIJ3pfS9PABMSUJk8GNjOqCpCnlTjgxPiyOYb7PhMIED562+/W9TRYN552
ZZcjJx7UdRutBTqShUIVigR4RdsbLKiHG4vMFAD0F+61cKfCJjW7U8FyL9A4IGFdmmLB5r5jpcAN
Eb0wdqqzPlsK2/+kEFt6YjvsvjwU4piFYplPcWZqN3ogj8yIUA/I/DFKCCTpDVpugwMKaQtt4L96
7up5JzbEPL8sZDLeEj3vl05rwVm5Q2E3tuebM1wXqrX4qSOu8Fdl1QGtZQr+hBr8UIqzzT964nsQ
TU3G+/+0HbB+YzRW6T6N5t1Zl7K/c1URIaMKU8zOgq0SbLo0xFupBuYs1It2z7weGewZqs0Ya2U+
SQiZlqwbjr7FtldKdbBrXX107kInY5UfsDOW+cQJjXzGR2aVCZeL8vVE3aWpo0yxNXNqw/F4IWfa
cIEUxK2Yj4NxnG+/r28HgWrMEjLMmQdP/N7jgVsLQp9SZ6NqnAWBeXG/0IUD01t0bUWTcs+7z/hz
KhzbsbpsVwsIqUNYOt92alkVuQhGZo9iAIgufmueq+lDjAx/AuWEiL4zE40t62TGDre4cTD7vKVA
LNlZsURVu1wg8RwK6bFLgG8Qw/8m83rfsKtj7x48cheFuPw67zRl5B33WOifhuJi50XH5sviUeqx
nWHw8s8dPoTSx/aYmULPrXx9NzwNlryfw480ifEbwK3oP7DPFurML5cekdry9MB0xosHbjSSuce1
h8AXSNNfAKSZPW7Sj9WqnMMq1/PAa0+BYgkS3MO17aDYMC2TjNLGpS2BJsB2JnLAAqwetbCRhkqi
1WQPhfrQOOcWyTxBiqG1VxubOy4/YA4aiPi+igDA7aw5mlrN+uTV1RuBV9jhuwUus4qq3UXUHcdx
iIAZB6q+80by4Yum14uy6Uf8xmSZWFPvWQ1SapXutQAWNfaSLqZbp4Mad9t1MYv0Crh0LVZn4Tc4
SytDtCjKszz8lQehd1WGRJrCzMtQ25uTJvWSEjKBPKIBese16rbn5VnvxMgHHpz5SbESuzqQQakK
36YNP0JL2SPEV/ft44Dh8xe2D72rMfZHRc9EDlBQf4c1GodVjer3jOynCRG4MRWlX9eO6FQkNW9V
301Z2CdyxWLqRwQb8qAA2cO4qSn7ocuRQURg7EYQLytp858i63rPHORNQl2b0arib+UcKGUzJrOP
547dakwP5nfNyXtV8XBQWqDY+k7ATw1n1GHKIP3e9qJ4TH4hzFRoXdwjkqxxpr4aot3C5nyFRD+y
GA48NYYwz61Bil4fgQpa1vhfpbEagHQtSDwDfUyek2xK95P3vFQJtPXy+rp91S//D08mxQLD+lef
frVjJw6rgm4YV3DRtvUcV0fJqxwXzHaI4+9XDOcrtY67NmseJMeU4QrNWPJP1zHt1o3/NTnWXazQ
M2ZsmjsfXpaF+236bsOfvLAnlS40V0VVWqQax+wcTFm0IAMxT20e5f9MtAS0IecmxCqwEOsKBEFy
s18121hIkm1iYiUMDXof1YJMG2vAhi03NmdPHpWLF+bsZzUBd86C/4u8WHwByuQkP8Jpp0fzApkk
UjZWAJDYhZQas+Q85bFMnNZ5pKRoFmNhEOcf5RbFMpTvcugcs/A8QJGoMiYjCY4ISRNzGvBKuf9V
6JD3XoToAU9F4xwqhRn70MojPf9JzjT/SzmlmcAPwpAxXNypZfqkbjKV0/lLnkfmMD5EtAY580B/
OUK9Igk03hR/9VSOP7gYGKdCMPocojndho6eya92U9cVK23jGfT7GiOzQRQQO3GPt7zCmtIC/4dR
ld2C/4tn20cZqJ1utsFQaw1ouGCzGcRhlbQ9l/PXNW/LCU5KUKLw8bRr1BAz1rJiFpevLWaEsa6K
oRtz8AOWcRrfo9Fy+eOcnPeVSfqozp8Y+W+S39OZD/oAR0PVsleA4+NqcRT5YkIok2LmUABFjs4W
oIB/sn7nxjRc7X8poqFnsbQj/AQSoid/05U5uyHzpSa98fSQ/wh7CwFsoazpkcqSj95P2fp2rRlT
kCdX83TrhOAqGS1rQ+w/T6HRima1OchrOBswnmfwlhHIUtnoCzn1BLXB4Q5ByA/evSbFzmRRTDgI
IjbwWLp/TrFkBXIZ6Ob22hxdQgHeLmLVLxkEixt2F3faCXs0i6MCXxK2YYDRBaIBlAizj6VDAXdw
lhDYYE65RhNv/wbHNsdjOG0PLxIzx2PtNDg9akeEFpeF9sGISTKyxRSer/zxVmfGZtqxY+O1OAmM
ql9kFRNj0Jee338OFEjH23WxZW3POwl8kZIDlTb/fk7TTexcx3ld3B0afLaetwJTT0TbiqUddJRA
BaUJDulx3Nb9TQ4GKYKTUR4qlx7J8rTbgvhyALW92hNZQTA38YdJvGCXF5usMUA5bWGXwfhOFcSK
OOVld2FjzG61kdo12YAcYS015FMNTYsI89+rntxuKRjGCxSaxVQCVM7CnRuLEIQy8/Gp+CJ11hec
jo4l/7xn8o5uy7uIVUP8DnlfBDJxLstwKCzdn6WwkpGEGVjZsd5ofi0pjqbJjCQzBcQfb+g1I/g1
0yZoT/oPlJ/X0TpgilZb1dqpemzfU9PpUHjDrQ/Ym7bYMrIN73E7ynl7RoD8z65BkqOyDDmYPWHw
iybMYyqgxJ4GiVB1AhUOBIiNg5Ub9caEQMq1hq8oWg/DHCsPwL4dpdFDFHHKwWd7CTcVVuWgd7bN
d+0gs/NO23SBSRo3cyOYTZVSw6vWjlKy3gF4cHQfMfMxJ5nkSFUVHTvtgFxxoUBmkJtJcnWJGfhi
JT+F+dOV9MbdUh+Cv3AWvEfisbMpi9RfSe9yREer8pfIXutoM9rmqPED7p+d9csY7Tl2XWJtuDHV
olq0b2fqfKeSA64c6gPFSNrnIJR39OmEndVRS2zvmbzBVRe6HpNisGup6eHdtFrYgaB3QO8jO10f
dUsTzuDX/zJ3WwQ3olA0SCngYywbKb3qU9oWW//tVgFv3VZfYuqzL2ltY/W+GZUx9d5SDshBlsWX
MOjMB5s+3t9EOJjoe0hJ+xTcUuu50FSaScIadiB1bjZ6Mr90Zrqk74jutCbcTdFlhhfboWGU5Cmk
6lJxC802/Q6dmhK85hQOkynj5tqNCtd85ZQdzht73KnmCJqfXNePj/cFTAlTsHIvvONWcDaW/U7p
QnTC5bNgNBqN9m1fTPBkj+ohncS99JRk072povLyC6o65x+x0N2D26pRlLtCDnb39hILjUuZ+BJK
AN1MNCwK/9yGQe8ckHb5TOmulEFXHbGg85fdhZIOE1D/FOZMBTdZavE1gbxUmpCnFsPuQg6SYPe4
rq7aAzqw9JEyqR/gYFie/IjJCS671Oko0GdaUHSLIU4QT9vywC225zgB+cYim4wnZavX2+GkWUJw
yWcqsavo9sSmcEmb56YSVq/dOB84bdUNKQU6OnBstgwfczObH+LfZk8+ZZ864y8c9fPd0I2FsFa4
StwnrirA8VcsK7wrmodRGZChWJG41Tzy84iQ8qtnYkQ2iIGKWg3z8Pi3HgpDVsC+podiLEnVCteo
/mFV+A5fHm70wdgefLV3qtNSnFnWWfV0uI6ezc6+hENdwKf6jm0OKud6h8596npCY/bGsww0Cloz
uetRnKlNvTMzB10UpyslnNaWrPg+eqQ641aYccPSu0gBtSOQHAOJu9/ImYl4RPJ67CVU/KK5J9ky
hN/iZDVfkz3pGKCR2YPAsiZZcFyYcgj2W5ELb1flyp4wsnomskbzMpoInW4S8Jzuq/MvtQNepasn
bJ/+hLROTYTZgXxO8EMqrUebFCT3bKaaUQzH9BCnlq2g1iwe+clMz17EDpN3+/JPm6nRb8FOWwxa
+QcTKE/iHdnYGDubVZb8qQYWyJhJXP0CL5+38Dx4c5Famz9bnnxs+63O1ksv+mdN5Fp3lSreQ1YQ
U35NPUOob500Ar8kMCsBpxqZv3ImCFAwq3sF46jKk2zf/OM3uYdMkYqSZ4ch2Qm7wmMFe3BfQh6u
QnSAbCatTRfzVCdqjnpLpHG34MbZt6wsc7DtwxCVFx5YRLluR0D2PUI6qK++iXjoTndgr0Bk6lGj
B22CjJ6UFv4bT95svQhZ4ZB2DfUmDWf88uHB5msGnnVAneYAOfjX4a2fDfMuiP5BZvrFh7nOiPbs
JSo2UkIIyIOWH9GUyL7OEaoIuKY0d7JCK/JkoC1kPkL77zkXN/cuVfwQdpiLtqDC1GqPR77BmMp1
1dNVct3/kHPRaqfXyhmFWAZvpxAZ9rUbSQDjg2rmJ+jj6d2SZC+HbupfI6n1lZyrmnsOrB+XWfC7
SSYZ76AhTNu1O6AHe+G8WnopUMtgSM/5Jrjb5WkEL4alWdyrefB7r5k6n91OQOjZeML97mv/Gck6
W/0Q5vI+Bda1ODGeIUvFBC/BKgGG/e9ClA0SHiGMjJb6XGd0JSU1xNqxrnfxxIUVo/Cw+I0AxyNg
4MT/PpbDutpgRBQ9we/T/pZqXM/m4rFtLRdrywHyzxBy8SV8MbVNyEUWdr8Azpy4BZ9K1bFvXle4
FhaFh1qeleMcapXeX/a739YKT70cwRkvfeHWNVlBH+12OOqOgsRON6m6QcRc7yaisRiG3lktfU1r
UWcTcRnD+0nWxOkrV5bRtIqo95dZnQ9HUD6k4Oq76uPSWgj5oYyYxh6pzBSDBM+i9UeOQpQVZjEM
aqW1Nak2BY7ssraKbg0PmAtti0XXOFAe8s8jYJPwkjR+1wUTdNvh1tIB/xNSzYG317B/basvjdkX
0C7zIJpxJkTG2+ivk8RKLWUmMyEyaQPyKsNZlNFdbpCZQigOgBVUx8s4gvQCqdPJMk6uTVcX9rBR
qTk3WUaTPx/H0+aUTLnKmi32BeVZESSRN3/v3QFrBf4jnWU008YyuQ/DfIkbKXnmp1Rlwx1jx/XU
9EboEWNWdgMH/okJCbupXGzI06DFceac3QBpaXQtmegX27MRVeni8FNnRPfcYgKxz3g5CxiecQq+
mpzoLFfGgJvFGGEqG4e0KoPRwMQK5qcKAWfRex3g3QFj2Y/AD+tuA6HLUj8jW8hx1phAh8QMQEYD
RKoICr6P9LBjz6TG/cYbvCf7M0uZeQl7yCpFkYs4QSmPDA26VWezowXQuylOV5C7MVAIDVYkaDDE
7mnriR7W5jPvwZXFakajpBIqakqrF49RgC/ynjy+lPmU7/KYv3PKWczFlfpp/k3xNYqndiPQLpHM
c1h6P87CQ/DpYMLlu9AEiJAo3ixYWJ1d++gbksjmiyhLFFPSQXyRu4X2lepnv66vg+M/h5G/k2Bq
GUmMzr2K5IL/qizRqb+oF7sbSrmnZrci5a/+NjpnKuRJIbKQWqxC/EmO5L9IOdLJrLETB90uXxKp
e3XlsmDgqlaI6v7vih/GgC0osiRlKma8qL2SbXzhEerIZNkU9TK+QQVWg5ahm4yjzXh0GeQdrA7v
UJROc01jB8K9iK2YjpXjmRwSyHgGwxHeHA5iNnDhtRtcOjHgwvsTfy/8H9m+R65qAe5I197482VJ
IG1QCW43WGfumaPBTQ/o/Qkkz24lFg/wmC1nKyH14Tn+6zIEg8tETZbYeuuhWcVl95Z/F4pc5Usq
NKigoEN9akOLgT+QXXgsLsAQtbiU4ug1zP6zVL3z5ivU+RZd4Wu4BdvqLZCBXTMjkOHLKezMMxF3
MUGL4v/Lf9s+2N+Nb8Kq/aOYgODbgGRCxUW2hvPeMOKh6GMFRLTiiLxFvVVxE1XTWd0Xb1w955S6
LzQuWwR/f22YDsCzPM6OXJgni+S02A0lm9Ky7eY+2lRtuUJUGLcUCniXYR5lOiH40NGfH9OAEfI9
h3hKlRF5h6a9mPrD2nDkC/zjqJfbeMYVl/3Yhb0wfxMML3OEqk8SePRDzq6uBWT4KsS7izCqDh9V
fFmKQp1ZscZMJhxrm8+r810/aIKMU3CL3NODi7y13S7HcWi3r+Wr9bUGL9UJrD4S41ZDTyeQ2MiY
dnHKLP1bleaCl2l7faTbhoBGqLl3C5y2swBjmaIbL3X9Bfc+SOP5cSuGtZsnLb8zuybRTpFT2t48
eaGCSmCi/UA1l9plZU3o1+1WRSFCsOH9BpdHeCJ0q75V/KOe6VNFCFnBYz+BedeKu4wMF+Eg1l37
9PfzxYnD8UBIjNIGzJ8Sja+df6sgEYBPDhiiABqj/scFv9aXfcQSwRraTyfcBsWFDkxhVrh9THaz
pWY6RYhBRalrNOmQwt1J5vBWUDZmGZ2LScLHkMlScj3njUqE395PwP9FmRiaYmf5ADbDtcyYckCR
QZWPr0w8PVnf5m+Wiz+bggKrp+KubFGNYe+PQQfGMyeRkuiP/taxdspegNmTrsieKqoICWFvCqhk
qapVCSs3A5oQ56DGLKXD0ge0PKe1QnNfH6coSx/S4gKu/p/WQncPISe7bJu8TypKounMnIONiDOS
D1YQthTR2eQbOCZ/NsDu7EBAQGDTX5dUk7z02yW+6Vl7M8Opjk4Kh4uYYtYaekxikNMQnRzvD/3R
hSOAwPxpRAi+OWe5HuSt0b06hFjAbB/mALaZ98poXyEV7Jlxy4k5kwpS7s+KXAuDEqP9y5aHa9kD
o4wh/wV5D8wSPSWMoeD8q4KpZgOWa3gT4kQAz6E0OrPXWuQCC+8zRhL50F/bWZRDBg5cCSyEynD6
HlNrT13c8qV7cYRsEbbn6hgbmp/fv/Wr6hKBw7pphuD5+SCUjCS4mEasXl1+MugFKYa1mmiphZYd
w167OtGM0cGJgbCnrru5+pSs1uNPDW6wn1KFBa7Mr1/dBwsKf7FV9WD5sMx+zTx99/5/ipx/A4zJ
lox6zR7sJp8fXLGiGdVJZUIYGeGY6luez4LnE0w09t/S00sBoFehS/elYPqLTanZ81rz6EDKpYMu
RMNJc6mhdgKcbpdv5uDzWAnRUJtXoYvD982nMkxv4/yyX5QfAkepYi0ZaIopZxlfg1MfpNkMjvDk
dkl9NKF7u+dlOzk+GKQkI1vReU6dE/6jfXEw0aaEoIu3eF4EQ8gvmnyZ/itiUmZ5mns5HlnrDT2v
6yPjH8WlUGhGMvuJjRy2fBEQciXVBQiYaLoC5AHeixP+La1EtEN9zzORTSJururVWs7RHadkyd5n
xMD7Oo+pGpSAWrjGOxdBbu97PQfq1woGR1g6QTaHLbU6w6N3EmKoMrimzbQ6T5FapCIZjowRPE9S
Lhll0DNxT0sLcF/qvWXti1m0xOW8tZnLby/CRiBd45vgRcazntLT9WaN6kqCGJEzc7MC4SoY7ESM
c8J2n3LEzQJRspinALMDXsFnfgPvhaV801ZyrRrCOTXweAIeipPT/IVERwM+q/daM5HzT+Td/mFR
ianrACzjfr3QpZvG5fzQRPI74Ha7Bhz4UBHMMQb/fWjle5nSaNKVBv86J8xsmExLt9q72CytLyZK
OUUAMC5Y/Gt7RfG6oQWGYIT6Z0GNejAfMxZOqN0aDUOA56pCTPutw7QIZ5IQP7wYRZCldSLoLfUd
nOPEYdLGp60OkkH9P0KJcpDzx9W8FYjtpZlj1SeGY8/jNT241wxfjZAKbwAse3H5+FCMbgbDmPj6
dWYI7VbXP4gIn/IG0n62bW+t3sXwB5nIH23/qm9U2627oBv4scEtu1+SuQoIorClRyYSyj0AWDtO
ecIJRykdgPhmhDzKWX8l3hd5JY4WWqpO5jHT+X/wqYzAObpVaWCWryNqt9AZlgRJqJqtrfqwItEs
ykRVScJvJStXqP1ey23npIMHnrJ0ElXTi9B0yiFvx8s6upNP+iqF/BBvtScWHGUlw29BjnLnN40h
xXIHpmBl+DWKmFpfsU5g+JuxkMfs/aJn/44/O7JHGoyEyO8Pa/yi6zIo0Ud6Brv9QzRuhncozTTD
BjDkvUDHDEe8nYDEEthe1sWhbnN8LmYBdiyf5HQDMPRdk7WIcCaRe9KUPYzwyT7oyWjngqbaA3op
/2cwgjrWX5Y1NlBR9C9sydXscHWOgcX8f0g/P1/DzghSQfTgr9RFLVIqj9m4sZB9acmCwHZSEuD/
YH6b+khAKli6bJrNXknmw7+BbnNEIZ32wLyPeKCmOkuCSmHnuzs9NQM0BRYJ1G0vky6l+Ccp2qhG
/D9oSC02B13MtC5GzBcLBmtvzzla1YuRc8rcALOvXDX7s83oLoLov4XF3O1sTKpt+PDhLlq4PSRp
xNZkYevO2yEAw5Yf+71/oyUnNs2ccTUSznCCVc8h49xGWXqTHUoHz70QTiSjhUniK565svj+FlrS
kqUS5RTcx/DFPXP/WONLdHFJfpRCdsNZcH7V4FUXCK1cYxU66dza1K/ZydGrHKmyeN7pvGeHYjBM
xwPz9UOnnJZWjRNEUCu5idmizg4hQyq9XGcPM6b2XuetcbWv0r1V2FzRGEfjuIY9xFnC4DltyznJ
vntBhhcxQTtTvV+vA8dRgT8O0+WZ3Vin2LGWHsOWQ0Fe+ISAcqqzeH2fWFh1friC6AwCOgWedSb0
FAZ5u7rtfvrPF8SVYl6eYU2M6hHIITIWn36BODfO4DDyZmr2iO7RJLLMezhBJEzqoWyS1LV/3gM0
0fylWvHCg2qRVT978HINHPid8z2T3Dy9FvZawKY/Be0zti8MnZSI4DUqnQttC0Nf5jPaQKzvG9B6
Dgs74NM4fqJt1WcZjeAK7Hd/U8ybf5K6/NZyAcWS2HUns/JzFUvK1HK7SIniWcXXsXMqdruGbSxX
WvdRV2W2hnk0HD35Frrxf8/Y6vINKRSiS+4NUl6Qn4M6C32XLoevi+AwfePRUf4ckKWBMIt3i//h
eNLZnCFwiEK3LIOIGrjSuP60omZiB1HrjDu1GmTqhRt08XFhwpMs2X3Agkf1X4sLJ0AkWLa4ByRO
GTInQ7Yc4BKF/l7kSFl+wuJwWCEyZQEUEnh+z0LHHZ4TvM0YM9upx7YHlIppWz8gx7sKcLd6vOgs
vOes+lq/GKhgRWF5CumGqKlMGkIpoOWhjkOj9tWiBW58yaipUY2fL+KY2aZyyN8X7DAK5snNatUm
yMj13gSnDEorOqYZNK0vE2IxZMC0efprVBliomDuqZ9xWDqlUvbCbneyrzjPh8LpW/sKbOktUjik
xl6V4Zh9VEvlIWv/ekuyDwWcqK8KROTcl0xVd0dHl1DqVulwAkpiPKJzkCBOkiT/hBFuKm1NdAYy
bo8MUjzjuRTxFLuUtW7rqyU9w2DfwQex3RFV3z4idPhbhhYjNK26atZ1SOzG5eliLjaDMvi0Y9la
noYOcVfankmTe98PoapcrCnLYGCT+97gju1V/TMRBpiWQPXpcycYQt74+z5FL6di4uo9RgAAHev6
GmhxkuDULGf2DjsbXwlqwSV/FKdvD6VaatgVYiMa1nCRnnolBYZVrcjM4ljeA15FAltUezrMq8Q5
yPv8ZbzjoBKtNWIe6nbwsIGzh4RbNlmHZmiF6xzyb3lgYzKqS5uiEY+x+J/6p+D6NnPtnJwiCNgY
Qi5hrpiaU8T3oVS/wswkGgeTuCA9o+SiEmNe//cEV1B2OZZP6vxb5phfjab08uY76J/ou9R5R1Ts
8qS1gW9cG7FD7CJd8kgXbltR6q6g6Mp2ZU3EZC1mT/qjWIn06RrOPjHTFQmwvkys5Cp4xdbkEaMD
aE8mE1MsnIjpNpCKjKxaUwl4WxMhCwi9Q2FYNL2z7RtLwpfgAAhjUIiZ8gz2vjC+U9S/LCDH4w97
z57fiYk47bBg2Ze99V/PhXszEGnuG0c08VfiKOA1nT1kds4WU4mV0LgSHMZFLb3IJfuOjedJDuIb
8wKW+6+VFjOc7CvPmd40UdysgszVkczuG2VjnBTNW+YIc8A8lqJHC3gdNhCRzGHREltE/tsMOFIN
pfsiPkNoWZXmgzi9pnmmbvfoJ6KptbW/UUTDAY/nTsw7ley79cV8weFRm7/vjBlGnYKuQKm96diI
7Sc8ZZn4jLVdHtV8xYcxuWyPnsslNwtq914a0peEBkP4p9iV0ToU5X1F2wUFfRMEmS91fpy6yTdc
mERBf9ORW93WHxkZ9sunLpelfWaD0HVCBP5YpT9yqmtKkV9RNDgsG83bQn1tahmiS3Xi/GVkZx1N
CSTjrkGV/I7xbY8Ww4yfcvyEjcBDcXYzP8DnVSJYdBmkQf0knUXutYvxxmE4ET7sVVr7RTQ9o7yq
2BDO9ExyZpyzx/gfzy5fmsm85UpDnRaLuEw3s/ZbYQRDZ4I5G6tRD2H8U/ROx1KLslNSs69VHL3u
O7A+k3P/N5LTimzoDIiWCXBXYZUumMPmACpp98AW7wcrzRF6UNvBbvSZ1kEmigCislINc7NqUzD2
l6dggyBoU3AsG1KR8F+9Fa9KsGnPZvEbTASAbPBo4r+VkgmzUrseqBLciGQuvDwe/MaOVEKPk4/i
Iv+Gti1WjrVRegfFnvRzs4DR1S3uCBSGDzdedHERP+nBahp0uZviSupzhtMfxWSXCKU5Kd7vNlck
mrKUWGcvjfxIHsl2nLccPTJswBJDXMnvOXU1SpU5rmnvZXRpLRMnmaSPr1GfgCBsni4J7SJCC9kF
VO9hqC3uki2/BurD9C7BAA46b4Jjbq1zFweOEQF91T1Uh/gcJhnqU9iawt7YfXFBH4hPOrOvMlol
XtOAuxlGVPQKSUGrBoBvTt3gjN+A9KlTmzUT3V3oDlZr2ENPvxfFG2lgqRqz1IKyX6S+KInx5L0D
FJdMyM5e1MTJweeNLw9zJXMvZ/KGNsruJv0lNK5tEXYQds4mnfpqZ3PYkxjRdrJ9v+855QGfbQFp
0UuTzb7I5zKowMkSZt0wkAbWU7llzlVYeFRet+h0mHMLJ8gWzV/J6XcPGvwLSWA/ROMZzq1mZJQn
MN3cl2Isi9/JNm4u/sSGzVqvs7vyFYuuJy+TSOlAwx689mpQKRatpuXVUgwppNukT74n9Eh7glGF
HmVDWh2IkYmXPKe+gd+biyk025Bn1+8bIYZRun4UBUNJ+9xDk1xxmBibpCjIDv+vUmRu2QoiMu09
RH6y5WVOaSykDVMiCaJqJUw0OsjkQh/47yVlQp21D65gjQJ+tuYBOKQYOKA60PMpPMbB/m1fM6dK
3gidu+gDYKsx7d3Cio4sXbaWuJkCZmNDNGnRDzTCVxfsPMm47SyLr5oGUwUhBmsv1DPacvhSUTW/
tHOFIJfBWLQ/MLgWzxb66YYJ0HkE77wnEimfJXNtM7VBkRzRUrPl9T2kybhIB2v8FD9RU2Nf5HJu
YjKjwP1IqgbPmBn+1OYmcDNjaBBRIoQgo0mPq0Ifo4ogsuKa1oV4cFe6Rla7GR90Kuh/iHjMVNRr
bn2QmoFOp/HtsZBjFZjeEqStxMmOnnURHM/Suz562/9MBhgtozAjLeXKdYgqSvsry8qYKYoqfd8B
Ap9s5tkjKSvEPjbwcJ5h12MisBfyJ0Nkpk4ejqOrY2iCV8jklOxUU+VlxpeJ0/qxOP53J2viMi+A
pvh1f+7wFzMI6r9mV3GP/H6QzdghbAkNprAU+i9uWQ/ontQKej+3kg4ug0/p/mgUlDIkv2Oj/SQA
newTlRghPQy7zrBRCB76kkxA5s02VQ3AT+ZwI/hl1G62ZfvBS2yLTBWvz6JKd8Lxb2JrP026vJbr
p10Pi1PUWyAfBWa72teu8Ia5Gramc8MUDLXylE7st8d8IcCC80453IBZJnziZx7NZxg2QWgfcZYY
J82cMz4zAYyfmA6TgQEGT6Zm8m8s9IkPK87HMH99glzXAKcHtg/aOl3cPUtMMJakETIlFGyf2rur
RISGMV+jVs8L4/O11ymAQlbGwsds/Cw24aqDLpMXIECV8NFgh3DT9yG+GD3b3TL8c8Yn/nheMOF7
PiRhonhEKJKlVA4pIv632qdbfO5o/ogZNrgLGYoo18yPMJkfADW+TsjK7WVaV7QmNjHx7xVLY/BQ
5eA5gjUQ/ncEh+uN2I+Hi9XdHpUDOg1n3grJ/lrt1O8/gMiOV09+NZUl7zWH2WEM0eCrysKkgdGA
dhaw8LaZdg4nS09l+Fcp6gbcRnw8PApUXndyMT6g9rfjDpbeFKcuei5NqyWfvq/0Ex184rxHfjd6
SaYXPwXlNAQnxFMzJF22cteWfruM9XeRdqJL8pDLTCJAvSh+IMz9OLZ5AhPiTAvKJyxklBFRnUW9
Cp4GIibEAmbh1F3gOJhdJM2EyDrk605eUmTHbiTrfPBfPtzuYBztwZNAlxp4QqOxlJpIjrMu871P
jT29/lai/laClf+phcfTVoecBIDIvTjP8JFOlulht6lc3EqoF7P9ynyhcZaEYCz/b/nijg+k8WUk
oDX0eNLzBCBd0UEAEmLljjX4G5BkBIgNfo976e25xMSPRc6nQ2JHC3UJ0yT/JTegX3g1TI09McM9
y39wQ6Up+kS+GvqKiBn4foc0DIG8OPzRXMqVIz5AKya/1apL7nfQ9NpgsL+wxPYfb5kv6Rc9M/5j
crtm5RWVTaZltODL8pX+L3cXtec2So1xvpD98uPEUXIhQYv3BmB362kT9FqLGd85DAjOW+/pwoSU
6I56dBpWtE5YftNwpMZXUlcjX5wkXs/4KNRBv1xBciEV/BpBBhv9jf7J0Y6o0uSwsSK43BCZY+hM
LCas0vZrz6KM8UX2hAW0kbeG/z8KVS7VA3xgyn7CSunWvaAd0HrcRDMVMmWi39VQWYiTd3HgIsM4
Zsq2QSzZaEVWIG5T00B0226jYGLVo5Dn+5OqH1Qox2TJpEZ6xVKAupy+J8xq9XLIrAnXZfnDdGAc
PcGjCfnGVzlbMJ+oJcmzeyjzJmAmZoEN2p6Hpft08ep6Ft89m1drHOF/Yt3za7GB1AjU4uxmsdFf
6dKBUPmujfrLDscsKjqa81mqYl+5vp2X/LSjZi4CEbp0TyGMDcCA3LfCtBMWAYU4KEjz2Jdg/dzd
Ht06qSBeKb6ocMXgMFoGppXaVJNu6Ux6JD6X9if3iRu40XwQb5+WZHNabHE6M6wIgcIbecnBRMwv
+wz/NV2kX7rIChcXsL1hwmta9Y71exLSt0eptjkIR5e+cHIrvcVGH28ryW6AK23iieV1NqSjy5MB
zF7HtPO4gr7bKe5gPbK2jgrxXYlVgwrCaTF1ec/aSnk9XaNP4CVDTY0O9KGhqUoLmuckGrpVVxzz
w/ZpIhzvMAOwzcGY4ZiYz1QqgMUNXmGnE0RLjuMPlmpaOzRyRYZlRMlp5TKDyJlz8l5Ay/YxcJD4
2BuPvGaagDh0ZJuhuqQYAiJI0IIGijT3kmyfEZzPEsg5JFMSx4VSW9CQw2UP98xnOzknpHLXd3oT
6PYKaAmA5lALVtO2yj7t3ydFZafZ8YnI2Vqpbe9Iu4yTyGcuZBwEJYxa0cgvjWoJJGFYw7ZSsYuV
U32Sl2gVnYK/KmSYhYHYwfxStespS/9ecf5TNI2Cit7AlVyWXWJxPrPrcxK+2usrkMxVU4Eo3SSB
MS4sQJpOjy+f7tqiwuhHAoeaep4/KYMxEXgW/lLBKr5gmAbeG0Qsg2HPNzVxXPUrCls8C4miN5V6
AXzetxbxp4bFLY7ui2RaCOTP13cpwsfPandv3Va5/KQ5s4H8Mbl9ufIaFJ//crZdI6m6kRLpxVZl
Xxjbx7raj8lBYpoyq5A/FEXDb2VRsUf40qDZ9wpyWGdRH/ltY6fJhTv9bUYF1VgkRGL/O/56reLU
t/LhHg80J9w1rr67sYt9H1dCkHYA7i0hVQmZeR6Voo4Ml7iZKQ/XjyaVLtYu9/TDExeFpH9Ac0dY
GIKa6Neh84WlXxT4Y3ZMyGaMQl6tiyWI97vdVh0HSEKCN/a8Ojm4sg4rb0ikf+t2OcgrHn0uSo00
D5Jj6p60BQQWFSMFJ4khu9PO8bCGw+qX3ttddY54JbA8PEJS1lhCHXULbMZM3TMZTPheSsT8ORSZ
7VHj3CeCCYNWjoldjXYzpckDrU2kpbaBCE6Cm3VisZJBPUxFhr6o5Te+joI1SPS3PQi744b089YD
QzH9M7QmB7jf7PZ5fSIINklsBrUlkCpqSTDxAMOlDpKN3CQKNwmceD63CJb48k3uPz5xeHYU0j62
x0HBNSja9kcbWfi5cCsfq3zezvGCuDw8Q3IOMeeOqs0BK/o59+xZUuU4Wzdyky8VHMo+VlKL/f74
0ASbkcicTV5OqQ2d1Q6JhcI7OcRsoU1Q1JagjwnfmopayvRHxpdXITeUbdssWiWqSLDPIkLXo8eA
DoKMnLMNHlB0AeQEwXlNQA2SUN7r0sHLCkpCFhHh1MKkToDfpAkX38Yk6FcaTF/shZjPmYobZF3w
cRo5/au4mXKkoumi4jAOiPKhxozZoUlzQg9aO6T2iDYdairiO99yMESHtMD8OSlvmelgyf7e4QKD
VM1lZnsHhLCcawlZFfXu+vxTXnM5uTtWryjAoE0WYyyyLgsUoyKe6M+iOh6KM29rog44Bwv7ZT71
fQH92GUEOh3tz6aOOjHLmBMwAqq/OR5P/wMCWuy+CfhMQx8U/yFxtSW858OR3L0pqNrDwybHeXZm
u4f9zyVwAQYbFhbixriYVpOvyj4vurMp8xdXI4cIyYgXVOfKJzTf08a8woY27RbK9NsKZd1fSkt3
q5tkn7Tmq0tk7TBt41xxQ4EQ6Yw4LNLNi2Fqo+LVllzvqEV2Botstg9kmdkCh8f/pGHwjrGsxQPh
/TmFSnEYWgDd4GIhfqG4KtebK2fMVgQVT1fmEIZHkxsDq/r/Ophjh0sEzym4F8HXqO+vVal2lbX6
iRbLiiPChdZ/GLneOPHvW7fnoANEsNhMEgi2f+NYkTOTn4cInJLVg121SSBlBrt3BfebuuDjl1D4
bH10Kl/ieRJQq9JqA68oHcPwrLZ7vZnVb69QjHwM1zH+AC2CJId2dd1knvRWNYb506zEGPP2KR1x
IXOc6LzvIYH5EZ6ZCImUjrcoQzmBlxHw0UOzsgF5qVs8nXxBTLPFvH0DBLm21Uv0n6e4shbqX0+m
lviKyulOFQDbtzJcRHaiBt2+7N14QECjXOSQtE0QgRgMT75LaopXE39VadstLgMwPtaw2SadAicr
/Uhs2dlai6pptrdfbcBQS/YTojhpile2QIjRzExawEjZGF8GeQ9LZcK2RyP4WG+6ZHpAqSGmsfxa
0UNuOWq/XV7V+hixWhcJO6UaiDzQE+Ur97jG3Hw7k8BNw769KpZGKcLl7LbdW/BEeyo4d0ZZqP2Z
rq9ToLah5tD9q2Z+b2n0IJRVELFSAuVeIUU7ph+3YWHut2ghNifP9yNip95UqlIBrKcoXQiZNqA5
31pBNUH4/VayL8aAcHixzuhtku5wIWdswv61+EA1U+gqsjMvWFBq5QZvz1n7/SY1+TDpauuMW/Ak
lKSydDy4CQcgoRlSQSf0f9EXaK/ZPrS7jEK8aV5X4Gmm2EP86YyE1Pn3ezq153tU3WKT0W0yySHY
xIgVpI32sFee6V4ei9MkYVRKq6wxB/YEygh2OMXUqcwmvk2XULzxnWqo1b1Y4eV5fRc1QQGiRTYF
ph/nYBxrL3GDx/VH20JWPVw0wogn/jsGmzsn/dC91HZx8oJHiGpMPy+xlqq2rOYvA0VeBrymdukl
r0TzOzvip6lOB6nZlxuL+cAHX+Lg7upi7IhT04jFc0FqWnXoaGPusdjGpDn22jgq3qa8vXEnJ4Bc
+H2drB7vAOso7/HY6Ucj/aVr/Y+UPPB62C5Vd2hSLjTveK1HGsGlm43IIGMRq1SoIzL5NOncNh++
Josyeu4y03dv/9LScLJj0zAbDZ8jvjpEThagNvYKy9XeCpmaojGVGzaYqoe0I2HWMnG1AYdGpC5v
woM2jW6SozsRn+jL+fR9aVKJcfdtvU3BqOjNYghioU+fPachEls81AO0FGTWCRN9AV5/46+U4CUP
09bEdhHWOdkIh6aPM8FxOZ1a5C+81RLw3+LqLdZOjLVw6ax8XBY9DTNYlhuAITau+c1gKGmio+Cn
X/pqw4JOCWNUA511bVZtLpcx64B0oZRE4mYdTDaxxjI9t2Ykul4I8pQNrvKEFEw8bKv7XKzaREWz
7JpULXgubZ1bJ8PQesqHIoYODZ3eblkuULqVfTMTXoapwbR0R72tPIjiIh4vXe11VhGOIGCzuv11
BBauAaNwWyE6c5i37vXflXVyG2z0VxvQ3TQyn8sfZ26S+a/UnuoeAAa/5B7yWTMEbsKOE9ELe832
Z5LcdybcuML+VVwt3SGy3HbvMyLgY6UL16v5zbRJ5aPjagdqG3Pdgec9/o7gdQXC44xUYvY7CK/4
NsQK22DRqp2iozyEpJ4yU7duWgD+dYdnVyvbm0ixO21woQqHOUTIFWz5EPSd4ZB+bX4oRWSjzfqL
sfpg3aSI89XcZY0asJozJKeGmtp6K3VIGjAPr6LJHxvMoQZroh3stGPtHqFikl/OnW4UGhhgrGqL
RMe/gkjYQiDSwlcfplql3QCeC2b2Pg5lvb7B4zQHOr3v8mOZdKleTg+bumpxCA0e+R9wtwiwHFGz
z1hbHqUox36spn97ukDIVbqit6m7dWJQtgOvrXABlGmFcTYbNkXMjNjYgyEjjLIljZAKobmm/F7h
EMJSKyqNiLSkqpyez4ITSIF6nY2dpx4aXTc1DzP220I24feTw+29kbeyI+nadUTcPkYugdgljMjU
iIGBSfrC1DsBoTNrmYoimWz50yKV0/1qvl1M6j4x0ft5/2CL4RAXBOE7EHhYrjyZrJODSiTH8mHQ
0V43qQBJVqF+qhRlOjBYIrnZL8c+bCO9qYLQ5vXPkEAjeN38bfxKPrMyLUyu7JC1aNbeFHkoR0WI
T/q+pQvjBiKPLyvDpp/1mDDjNtzjP9GPpPi0KwFlCgd0THoZFzY1YBBuI7eH+QeKZ8lAxj/ChcEn
y3MVvhOWLk2b5dBHjH1Gyxk7SZQsUAfRBls8wS7QoqQnlm5EWi3NfGusobuo1d4dB/ncxcg7Bhki
4FKC3WGuIP6TBdHNIxzBugh+elMWWybJwSXRkSLCAejNpBdjGaW5Ju5HEO2QBU3I/NzzBpLe3xzf
06w/NbVKSuHou9CaZnod1/UUH+AlQK5drgug0q/fLm0nK0H6pHI2YldYNCFkNwvE+2D20dRx7KYG
tNT9qyR3Vw2WNVROHlAkxrGF25nrhLhEs7junEwG2Ks+wPlaLlGCrn7nuNCS5f6CiBVKe0Y9TbU1
GDhrFS1jJc6x7ATJSY7HTW4jdSI9ytZQXb2O0Rih3XNgNn64YTyyMTYQcTEqSW7TFIUS1/S9J9vg
gSb1jNEomCawSFLQU0pH0vGgmXrWo9vEa/iZwvkQzpRtfIjWV9Znhk9JeD7XtzO2fhguqh46AJJN
MPioDGhVyGVxhattoy4UZXi3YhRBvLi0AnCYD0NIc/HUbpknvB8B2qF94ChAe9VXH+HOx6ltgUY/
/vgr1jpgR7Oy1JFfclnwHeeqlfGgyMsddx05EDlxvzQA9wm7U89LOUZxdx1FOch+HyRZmOMi/VAL
EEzacQZVoGTq5ydn0KBJZF+7BHv/5JgrWaQkKvEAD1qD0T9vbwxCZHGNI1XrgiY06dN+pOzGZ0i8
+F9lbARScao5iT9ua+dSwrJ3Y5/ErpiGkElbeSnOU0HvTbE97jMhH0QJc75soajn8xnMCyGBPN4b
A6BRnCJEj6ThMITA/7xXwc/n5CDEVS0TH531JSh5LwCJ5HxqgKqmzaCwh3WdEMQiW3d3aSSitrqb
2U3GhW+uW4wuX6UOnsr2U/VO8SaX3NNYbOyL811p6L3ukXoX4PzeHQZ8x8uvhkrQaB9eOH0YUSk1
bDWHCRJgw5BZyiSOHlZt4/Frhtdg+H6MhKx/gpTeiGZIt7zcnxRQWyVDmMH7Ti4oo//8Fqefsvdp
7U0O3TLe7OMcprMXpIdN8gf/3PGcRelYihFci3CPqY+A+ieFaMyMvsakLqYc5lT42Iix/UbL4y8o
JpAZS78/pkkYLEIqYUXL//04Mz8nt5He58xA6IKuFfc9xjerBA0y29yCqgaHnXqgoQaKRnXvp6xQ
LbvP/uzoxbYrGAjx6f6h7dwJy0ktjqn5rkvCs31aHnnf/WHnARGj+D3m7xqyETZxU2xS9gG1bhY5
8vTb+aisM0BMVs9EIBR8UFTR3rO0CpyB7A59KRNoGMt+sx/zoBLMhZq21VQKJdNK6aDMjyxlSGJz
54gngVTjXK5g0GxVs8PIRqUmd822Upkw33qO0O9AJM+VSP/rO+HuRuoeI01GrHCgqmSLnPdZ/Fht
2xNZeMZf0oQOEyMoW0zYYYomDbYPBzMD8AaUI4CCRdL0VqXWkWVEKjR21fEe0iMccywuXDV22CFI
xg0+3j3yUQZTLypYF5l/+BKslgWL9q+BW+udnH9RI7NXiUtLz8ihJsYxGHMfQI6StaRjiPRTBkqG
9jTyY647FtC7YdWjjWbEvEnQChS17xfkLRiPGZpuHXeam3cGcBIMgX9lEf18GImsNu3nbp5m58jU
T60DctGgS8DoUXJDj6DmgNlXQE7U8wLQ4onGLD866BaGCGoQNUU+uKkm/rkQOEEm5fam6IDCRhU4
jFPdsJGgumrmYSdrctsfDb6dcoAUxRNoQuhAnStxaLq7/6jTg7/0YzL4Q5ZHIgn6j8wd83wYu5aL
GBFDHGH3UgxEWAEKiL+mTtIEAMqRBSlDLR+Mw1pz8LsGpZBnfYxfzTZPS22pEBUEuvve4jvaWsZo
p2GEzP5TdAeOlLdFBBeg/q9W/ppQgxxt/sSflpWj3Xk1VdFGiMw9TLlX7IoEAbU7k1HQO95oVA8v
nYWeAhtNnyvUVS9mdRKLLWRe0aSjlvQd/sg53zRKG1t4V0SLNhOcGfSHYnOfYXxbG9/ZhHZAB9F/
6+bOT/OkW1uiDQHGEzy9RgQGqEY26pVjqBQ2e8r6C/GPIiJUwVvTB/dmm7vOJ8WgADG5P1CeuLdo
Pr/hZYVfPDLbpqJ9t/9fGJKvivJ4vzW0z+7tGDwc+Sz7+XqR/JH1Msme8R3gDxttqofMQWiotlZ2
pzQ6rqjaOt55XQrZwza+CB3TLl5dZ+av6IG8rOIFcfPAjtxP+xM6e3YQTXmAV7Dd96e7v4ixjDzd
WqSdqRh3vJuZl09DGyigfUGVKRRz0a17jBD+u/YviPQZoNEvxOFKLwrDMF0xThb2YWMJNhIbvfJa
2fwRXE4luhMoosh/ZID5NKZeqBZ+ua/JMty3+eOIiAYp9ubA51eo8LvjmkiRgfccv4sS3w0QpfbU
KVbPJlBfoxLiWqWNs2nFusaRGTqRKCQmQ9r7FnWq0AD64k0aM/QIx0uAuRqFePtLEnQVnOeSxFev
jneHawaIJn6JxnEuuvf+Zf5sKj1RURF6MA4MOjbxYy/jXthXH0Cj6wA5xqw8BzqjpTUYOv4rINEY
sBZPpsGYoc8fk2bad/i1q7P3k0dfo/+p4aPKWCZQpXC+r/GlF71m3Azs8qNNPNqlumngvlqf+q2K
KwEY7etBuKd6pnv2dzfTrr7KIAV4b8ov5edSnH3q2l+g00U5w2G/9W7Q0HQd+tFs6XEhDYqddN3d
JoXX/0VW6gs5clVL5kFyFGAX8YVyyU+yBqppe2V2ZvJkUTRga64Ow7L8mrnetkzpvPeKpDyEXe3s
PwAKBtZ6y0Rk5+W3a6+wTy4v+FRGEv13UzRI32+C0lLgR2jMuO7ziTw9My/qTDrUJDqAMGXKcV/w
9u7gA3hzRD5F5dYdLbY6lWFb5ksFdX5cH2mEYZDtWKhtf5FcX8pM4mSqbr9J/Zk3AXzE8xfN4yxT
7WEVyDV5qStH5Ty6kPS4IoifYQymbQs1HQFh1WWX2vm+hX2woKJ2MwNG5AbseBRUxNg7g9bZ6Vna
W0pIHdRj7OhIyIk+9w03KP0c7Vq40CnUWIpxy84fQ0qYUUBs07jDHtv2lU3XP0MdTQVIlJnKGVJH
0AdDZ3VbLO3vt8dekdTy21+KWkrPjUhKTICauYCySGfE9KbZuQAFwKya1BhgRpSq0QjzLx9LIBhh
j+usxjbUleZOneO7uh8bH/Tj0R3JQ+H9nW3sBTDWzEyoJi14PLbb0NbvNwuZ3uMxaK5Lo0o4XkD2
c9a3zTIOmRmAgd7p19rZ2+uKQlx/W6b/5k4pB47LZUw0OfRI3h42HeZxqeYXiyBEJZiQDWpLMAwQ
wA/eV+I/iOR/ciEG3P8cxwdnntKr7KVx1Y6c/jlxLB5/eTX7A1Rnz0y20oRnqqgQmYVCLQUh/EsU
70mTM7QaIiWcKZwItrlw1sWAm/xTqvuzR1IqaY7avRhynNBT2SWjp/xYrAtUURukKeyKdtFrQACH
t1+jDIxHOP6XQ5h/44RSP5yDIaSO3rKhVq1VBshuVIz5ilDJitoPcUgH4cj0KfPWR5IlO0wptRns
Kwm3hP6tVRx/LvccToLA+rel4PoH/KXMenXM9wkdaodhbyqpfWZC/mZ9uuyHVtopDk4Q6BXBfpL9
c9thacrc9/I3rP+gyfilbgY7OMIK7+a2/1iWvQ+d5Njal+C4cej3xOwQn41YUyfZU0LXtOysdV0Z
D9RQ3GzHxOSTFhSqNCioRtQLQOjHvM63xP5ve4IPwmGcbBvcCASGOuIbZ/PaYTDaEIe5oKcACaed
z5l9z9hKhl6nOMV/ay9XWVKBUjRVk7K73Iwr9ADCgT9fES/ISDFsz958qrnqh3MgG3IZPJ3HkhRh
N5xBnBL9zP5KAC+hmTRv7JZbHqfBbhLvxIYqxhhiTSfqOA2NZ6HANmuZ77wupQnUMkIKvYUaHTom
fanXHf3oPkTTkPUKcO97PKO6MT3Ohyq+hoS6R5hG2LI3/W9nUREE125b/FSXO/jSPeRVUI8wmhbA
4RBeu/fKUIa8TKsv8U1Bj+QFfwWTlEphrpfQBACag1xm0Y4hlZ/4jK1da8GG9nqbAj1GX8kXLE3n
WrVXgQQGkfeYYyRUQSKMiS5PG6nbaG6RHyiYapM0p/mcRH6SoZeve/07prA5H+6yd6TOpD8/XyA5
YJfEeWQeqYczKTGBNBMvx6uIIUdS4bhFvhiFud+Kd9AAXu1Dex46zRRdKAZqVQxy1CYeKjVXiCVd
21OBKHMkqFvnHDnRYkCChJvksqUF8A5zdpBcjtk5Va53rdU2OMqp+2I7tJuwvszz9UOp8DExJ4H8
1j6mMsqK4MmhOTb24heWZzIt0560H1gMBJ8dOR0Hj/ldkIhGDb/GhrWjJBPvSFqO0slLmTDruZK0
kCtSIMf+aQTpsLoVb5X8l0GAx5AWXm4+Q+gK09DlqwjoemlTPsAR/coR0QxoDuXije3Wem/OIVW3
x6KgMdzwFoxoPB5N4J9X/8aGf64q6/jNH6Rz83iS9aTDpQlE8gcLDRsKfIAtGuiOx0V2gpVlXo7b
aBeKLBnhfefGvnHTxDmj07cxvS+ZO4ILe00cbHP8LBx3WCC1a4+PtF2W9SrcM71B/GpF8Q0npRmk
MN5esUjqLeu2Hf592Lw/IIBS2eFVwxANSOY8L1nLCGprmgAjLUAROivmIrcJWbSCQios6xCkONaQ
rT9ybdDlqr7VVFaS/ASeNL6r/NTTJHpnnFtMlbM8iAEWmSF++4Z/ijkFZEtReMOehlbxjOzwGkn1
ejJaZRD9TA7fGO6tH2Q8RNwDlgdZ9xXRhKRKlJlMmFOtWf+iS/2soiwlh8QBDYcaQ/uHyRAHHwKf
5hKyu6fc7KDBAVPKdEMIEQbpcZwIxZ+7/puWowbziThsCB77UlChQl82pZiu+NmeybVdlHCwBSew
l0iWF3QI7rk9wxPbtJ6jHR75Hsp5j0Kha0j0U0TUW/EjUMFuzYbIHkV0cUdiPmP8pHLH1foyaEAr
+wts735srRkQ/xOlcQGyDCEJCK/Tx21Hl7BvDVcblU0VcSuFvmirfNg4/AxVc/iNG7TklpDn42f+
P35iM1L7ja6qjUVsWSJoet834wWl7SJj0LTce6pOpAuORjdiWS0Lrh4fMy+ceo4n/cbpoSpcL+/1
kTHwy37SvvjgyGQsUBCnlc1HhkZstv2ZV3PSKkdXexXBG8hpBw7CwNMu4QsMvEgXnMGwDV8kU/Ke
1spNGcsFH+0/LxPXQ+ZC92hX1udWu0XPXPn/ZlVJiyetFoD7Wvwr90nMUAS9f8seu3y229GMnMM8
96DIwMkX48Wm9VlznlmCG9IY+TZJpCn9k8xLZuuuj8ftiyTx81rCyLfSCa83TpIc6yLGmktDQGTL
yyAgWw+FAYdnbZ/karwLnS3hHuZh9+HOFTeBmaANRjsk+tmu0D1RNzlgaLsA/Nlb1CxZNzQhrKiF
TAIMVSTT/YPGznI8z8e78jEG14klUB7xZilz20Bco5Z9cmOmHAbXFybvRwBVvYEzhZjCPajjUWdF
SVVkaDJ7A77Ccp/S/9RilReYgPTCczH9LfObRtIoc1wm69PTrQ7LU3T4mq63bVqffl6OfwQBYiO9
uB7ngN4YwF+dexwjoovTHLehLCWiVL6bnphZzpKpHT+5q2bUXK+ZyYBYdTyg6BePVKG4SHEpONAC
0O5DHW+pIG0JKYhr2xxfTNnBaZrVD2ilF8S/Iy43gk49wog6Jc80ZBYpvPriIItd2i1DM4aNvihN
53sehoWfT8RHcYy9SHC3Ll4+mUucbNC2xP3WuuukrLWbegPCSAD8DpbBjhCN5kKUzW5Nak08mPdc
dXFcPvHpnUy+Yk/cktWEMrScgj2/Dt6BrqfvNu2JIKVxo+DO4LhEbtXuLDL1obuVqUMU2RtOeVuf
8mGjTwQEajinQZhGBMFUvrn7syhBCc8SqketjJ6qjKi8FhYm6Hdf8aJkHNN/ZcL4OO68hSibPNDF
p/Mlwxa7LwKbR62gS5AsxttpUMnB6Tb5OxnJ0LO+mOC6/yCTdd0bdS1e+nDOjI6r6hjGdxYl9+F/
/rC5WFmN0K1roSEe1VSyNDsXH4CwjBQ7JP20rRCBEq/aZW6B3s9s2tdhUXgguyZewUr0uLedX9cu
neD+xDTQYpJ73LAyEYkUK7QmAvJU5JAC7aQ9iBnKlygsU6Hw0VrHN88yaIviPYZdgkifibuv0A5G
9O7deWMbMgdOoC/nKzF479K7NqzVkhB9z5Z6eIrwd+DIPVCv0UGNbBDVnD1wt1fMu+uxkTk601pf
fMUgua8Im7zFPJMTdHvNx2iI3ctXCtRhOuvkNSSMYe6+z5dd+qY0bLRxQKIA4l6Bsh0chTY/Ev2G
5Z2ZSEkxKLnCRgDoZI9dmN9ypKFGVAkMPjBbOFl1tDhzmhevw5Inz9xU7YDx4LJm5cA4C7nkS35g
BPmnpvmskk0uwOWP42NVYXQr7C4K6gU5CsObYApr5JSwT3m1TbHw4N5qpQqGDeIRUXG2653tW5aY
fWQq3rXDgV6cbbcOfhs6rP3uxiBU5kKkk4XseYXf4mfLIgIFTYcizl+oIRxHXijIteYtQ3Jkl00S
EkN+/EQuBlttYHKhOGgSxIlvB+9CiEWm8BEZUJWX00CUqVOoFXlRas5qqo4YPhxn5z9+BKNNGbOG
2Se8TmN3M8ZUVKZE7FJlp4Xf+boqx0eblq/B0Dqk+kPDMvpmftmDfW9hJBIAkURlm7iiuvwmwHcV
huHLg0jzux8nACgkFyEMRzJdcEhnR22qkSiBG9DpePk5GHicASLhApLf3UoedwIPs9GemzkR/HSg
PtU7F2eFEY5f8j7TDcusvy5X83CUI0pGFctUGrmWXYLX0lsFHyzNdtN7aQQ1fHFaK13MA6hVG4Ms
/vrSMKg4Yk8AoCSUWbO02yL605PCg7H7GrX6B8cjjXrwgDFhOapZd1b2dBdxJN73VrhBTv3Zmo5I
ENXBkrrA4Nws+cA1cMSdUsUQ8s+ydz9STYqo461+4mmWY3ozuI+bfofygTRUEEg6Adr0j3c3gyPj
88A5UEzT8b6UWlN8Llhz6XN/xiZd5/rZJderf8XhPVrQfrcItNPnOlJsMosQ0vjKtEBPsxvETc8+
YwJfdoxgiluQLdNb4GTA6wHRMk7+0PBkhPDAsMd4JA+xMMgdST7KThXvx3TiEFC25f3ZbLVtH6dU
zOEMv+ni6zKkRqHUPhsYJFJBuc+WpZjTM4D8upijgh4/0GGmEQaurQyjs538sLYjVd6icTSKI680
aRZ3sam3fBwFMPyAi5x3D+8NoJgb5/+4oz7LAEsMlobg773uHSlzj/mIMviN5UJjJ5IMALBbrZx6
a4RI3vZZzlWlMVJWdAgWK67o4ofRogvQUmQ6cMSVHVcOkbxVn7iWhc5Vmv2QzgTx2nsT1W0G//UD
zQ4gJCTmKk3PN5uOcU2vKP9Th2ju+mY3TFe6ahm0oAa64S2sLAbq9l907o1EkRQCspPz7qZOpYCa
OYtbaKCS0Ap+RhsH2xtDFTp8gNPymJlXuG1bhrcNLspXGDgN8l2fPyYVOVqIXLq/jtmtex650sap
VnNeQkMlwSZrA1elmi4zPeqZgysGjNPruZPxTbQYBtujZWtOA6MQmSy21kecPDbvMLx7DNnRT+/L
waAaThByeaTmsMzePdTmX5zSiBvt9k91CcZIA7nb58kSM+Y0Ao02EaWkgoHONH6C4VRDZQpBYVHH
uFOb9ZLhnTssZHZxi71CrdSRqdQlmpmjLNdGK14Pp51aKd5mxdG3hRlYoYy58vw17oVwLaq2EMjn
/ynIne4c1pF415pqZv9sO8BP91y9QyQTFvsqvT+KV/ix8QfJr3smd63UqB5ys4dZtJn2sro32QrY
ag75t6XOu0D4PoUOtXuiP4dg0p4S7rIiOJ4b/2HT1avfKmZUROsmO+purY6R3N+gI/H92cT2RuRI
SzbGnusY8Nw9UyztwoWMs20jzhzL3XHSzo++SNz4ooY4h+BaeoZtnVRhIWi12uoFiX2ueObeL7y8
wz60mPJxInCkg18dyf18nOHu9Vv8MOLYBXojRmhExsjiXCkws0T6x0ouDvMzsqVlx5kHbdSn2cTA
Hg8LcWK7g7BDLHfqgP2VBMfy2eJVTOX9sn8IIP4FL/+dBkGPXjjw4yii6JaBZb0+O/hk0oEuB/AA
jyyVjntkrivFgkQMOlpyvLd8qYzcDq6IyF3PvzhhR70G+KIY+Qv7//4SDt/dOi1uJRIj4T8kMy9k
n6uF3mwkaNH//1QWDEbObt8KTLsaGgJqZOwB9xZFL5CFiFf6qwH3Q1tkEjMnbmbkCZk5DQir+37a
QzeQ5vnTaHRHtnIZNxxT4ZdIl5nSO7nQT65iALQEk7iwGkZLkGwTEBMyeOIfVabk++4yqqPqdgIo
8bMb48mFWwI3KuN53QE7aTRY6/rcOwJ1mRlpKETwu9OYuuaBaFBcE7j+2hvGZn4Ix7TP6opk26NL
JN7fb9oFxJBCO/jQLwTePpmz5OjbvSYijYuIX56xBEC4P5xKKsHrNyS8pCEBljt0lpFFFp3Gsk8I
KKTOBOHDrDQc2hSq5ZjHEC/Rjrk5UgfvMgiJZZf37w5rW9FYETjF/Et23TEBLk0jO+9WVhDOWZAP
eXuOS9vOWJP7SCHwIcNCwoMiRSSaX7+q4T8o3OlOaKR1UnRCgxTg1WO07l/SaQFFcFenRaHluDfn
Vf+/N4SP1xJv0sAwQCtuzt7J3J4x0Y7HSQnPRPQbDUGLRgu4qXYbplzVH5iGZHqZlFuxYnzSd4Bl
hm48ubbzX1C2TmAAJLr2pDu6CgQeDTASNV8aoEgDm70YhdsW3zUPrX+G0+5w02SeJ0nNXybkjbhB
EW6vuLemCsDCi6a8mK1tIoA5HV+fOdvnM3AnR21FsaBzlCLzGhzUsrdFNVVLojyt95Z91dJb4lcD
DVWJM5f7hqTTmnBk82WEZzhzANGCIchFkMxIT5oxWDshWJNN8IP/FC9fGWBWdIO11wMJmIOQCl2R
IS6WXo9oau7Uw7NP93SJMVCaJBQWu81B1b4Y7goddWzcJGEg/uADnnszY0P9SN3jzugUPabLxdih
DH+2ERBGRgzmmGnYNzPhxDzbMV3qOyhsqG0NK26SIzEdRxvs9IW9MGCAjEVG6Ko9G4C0P9pPrXyN
lqyxtEE0NDbWoB451VzxTaieA/F+CzdqT+32ElSRt1rjTeHC66bvO5UP4QiNIcVn3viqNu6nl06I
guorwSoEMXkkDIkWgN6O2pxIbbppzE3/Q1IDHNrVpCM/Afo5bkasU20IsmNs8TnNnh38W8i2ovm4
SzkChNul0X4h8pdvL1uOcqERFarw4vS+8RiW5jKEWOdDvLoqdNikBuvxmexDfVW20HrmNVg/LsSm
EVsFs2SW+zMk6whDgADT5Zt/ETdKnQz9P+fP72v3xwj5rSRaKEl+PqRufKBqHQ5VqxynxOZ6gJRY
aS57AsqLurkMV58PpbG32pDE2pQK74RXfsDhm3vrl8fzyniwfSkxwslS/I+STb+fuY2Sb9Hlb05E
XtKePLuYV5+11QVdIRuCJBtupVe3qUajoILHxi85dh6ELLzRZTq4gsxXl8gwhuSVPtdX0k5t6I6c
Etd6AXHIpbD5E6ZcEiDaKHPd0m+nq11GJ6DkblK5mXvJTOqvYL93+7rHwrTE8Wko7cnYBrYi8rqL
SxNU2LWRyPYUnS791Nwi+YWp+8m602WaGkERZS+RQcm3nb2UxTjcJzvw7J+T+Xu4e6pGLPLDBKki
S2KcmAd0on7+TM8nQT80a7x4QSzLa7vzUNm8swrj2/qA6SJQ2zp7fg7/NtnBJ3JtnmYl0oXz7eHd
a0gd8LHuIWuXn7qqbxzqgzV2si28eDWEfSjc2Np+7+iqtsNNChsXSUFkJ5bixgmKDAEU1bcPnVFM
5QxlB2J+qVvrNwKg7Pg+BmOYagOuHjSf1jrOAynzpIqbP672K/C78P6FeVFMVWiw7KOKqYJmwLqN
QCeyOOLPjcaQu8ka7KXw5QJr7HKvmLEU59vp9mjO4UgmhV+nLKZDmg5DCyAnx3eN8SUdthDHe5qD
HB3cu4/0wHqg01yCAjiVKe2PlOmz9vXGH4vUt5a7pMMlPCEHNe4JCrykkus3+IQ4yKvj1VPAI3Mx
+brZVom6VBe6M7WsXyTfiVAQxirZ525nilIqi2DIKBVDnoAhhESSDRxbvEc8RpBzocUeXCShySVW
91wvrzMSBHev3vv1yOuRhmG71X1ITJBYw5e8nKh+h4Jn6jLkp2VTopxYG9plVLE3VB18LkGfOAOZ
ntdcPek+M+S1hy31d+rEl97t9azFvoq3ll2SAAP/sBGWlki726QnT7lEmGU+SJeFgQ72n1aHFHyI
Cdarpus6/+Jnrheo7vLmEy/nejoQqrRki77v7bDGExADiQX1EFV4hlfsZVyI6RzpJlAR2YBn1WnO
0YC+Ln5VZaawJC7IAGW67rnM3IrZEN4AkCtD+/Eoundpbrxz7TjgIzICMwNcB+1BJBaaTRi+fENo
/PeHi9DZCESDQgBDkdCC8tmNq7H+o7e5qMe2UlXBhmP5Paz+C3SjmKL/8VZq9fE87UZqM6/AYmAd
V7q1bJTvkiDE0YYKM76bfvYhy8eDxYLjjufFSiv3uS1DEJ/zriWMB8TddekTeGiEcclQUPWBDfKa
lbIu8QjfaPYb7wBne9mXfBLEYiis/hQc/7h+A4z6KwOkdtwIix6reXtwQYjUAVX2oZ5EswSDxBGR
ccsDB3H1mfYo4LIp77L1tk7AEqrez3V7J3VxYUCvnwDFAXEjsf/+VwCusDnkLevt3BmM3MPQ5RS/
hDtNChu4xN0NXYF5vvc9tsCsOg8MHWzX6HA3woZ5DQc+LY+q/aK9tXB1cm1JCooljZsbUzkDRDVy
/tBpdElgsis9vZm7ty3fc5Nqwnx3zBGlfyiFXCiRKjW9XNsolF+gi2EPFvUPOUyRIwg16PmTP7LE
bx1vvGXuvdIeskgbuoDYyX3EvVYN1fyf9FvCvxM1OPj9W2wTxV4YyQoJ0KEySAnICWyVRdOb1EwQ
SbrSnmzmyP6vsS4oJJFUBok1vsJx39DNSjDKUfwF8fNY/aV5zWV6FBOSTplLTzWca3JuBNSjk7QB
v8mxznXCfPH0QwFLvMvJrnjbJrCrS7DjV0cqDo9dVFWgnh540dTXlJ2F5MXhCq2z4qofF8Q4oPgu
b0uK4BmXxM7yt3bw8c4BFtKuMM8SVPqMP3wleWlOaPfGytV0EXfKmZZsAY0dnAXAZW6lVXtPk1FW
t5ArkdVk8EcL1OJOG2TffUiBd72czH6p+UOaKcUeBnaTFjr6DF/RMl+2JU2hK3M7Q+LWVYzmn6yG
Wd+qBO476K7lOOSt67oOKJJbD0qzNumQ5WXk/0L7OAVv2XhQ1JFrtLNvMrGBrkjZPSNO/G0HTvwD
mwkwdR0AGdS3/pH9Huen/CeE5ZoiM/2IrRX90+/BiRib2tIQOIwfVNcHIuziaVNMp5u1YBTysHp6
yqtYXq1s26Wjb0apN5cBlAIIgUN28iGJ5oPbTzbWOsIk/REmTP7zn8STSx1brqaT8G77AyNwvMVF
4IY7An1JOgSesQRcCpMNuLZ7KdX4lmt/89bcbAiLVdkFsPawbHZx/ZJLKDSfwXHJuZlhpqt6MY0d
2ImbXiDMKOmvRz/Yu9JFWh9dKX/fxgsBb2s7cr5fk5n0T3P0Vj8NJHQ79Ad9UAlrnn9OPR0m8Urf
jGsgDMjCfzOkKADfBwVWLfbXk5X5iBWMSaRHL4WQpjdmC0uQH+skLMWIdTNZs5vbSJQL9TP7cXIk
Vh0j81cWwpWtKPHEyt0LPRAvWETtWBpfs7Nrl+qyOPMGQ4EEO8LVCzyYKZPgSsv2QUFMnoeh6J1Y
CjsRnperXPtsdkY2dH/uWa12bqkFxdtp1WABQgf8Tgmh9vAPUY6igQX+X43RGfDWSHRBYplycSM+
DJ/6pZdcwKjKHiXUyBsWDQqarj9w2Bnp7yCu1yX+pW+P+t2Lf0zRK7Bi9bsKGTpLPqhwYeNZmjKj
bEkHTgnDL78kmEAutnjR25cUIAi7FIHS01/owY4pJbNfy6ZuR4SyCShgvF8GVzVaJDHC6Z3mFrB9
YULl4NsB+ruqbxZ2due4+0qCtZ759Pokvxd7NKp+2gLQj1pN1fbkCugutwZmbLhyYpymI070NgZv
H5a3IwMbQeADQ1VTzXDBlACkt8tt5mZ/6Nbg7GBcRqC7ES/kJRX3e75/ZTX6bK+TbWJjGsIrBqYg
azQ2aEtaRp1JnyRGVrUUWPVEEkJi8+ubuhiroZR89pjuLCoTnp88oyvnktKBVKxhCwGzCZs8mlLk
ev8uGTjmOH0bFb6Gz4htHzn4+TZbXlald9i6nDraHtBFLgTAjpF6T9IRk55dk15TPsdE7Y+o2rZN
C8iD08X2H247rdEIKkxLfGr0S/KkQdVaybXs1LsIgcENPCoJ7T8gZk/3Nf3XDxB2xQ+SW7Fwgtay
3hxcOJ/kAGbPc68vTBT+6Bcor1/96Z+es59jkJXFjqgiaBju86YWhTNGA+zVt4NWp4CjHrqK2mMX
/NgYzNNaYXANAQmFlxaXH0GyybfOnYOr6drsmlHNwOTqHAaZIqf/w6dBQ4Urc1nYfiv6mmElUXXy
N0xpqusZcpl7FRUhExUEQTwQhXpwSeDtW+XqjISmvKrrWDmOOHL5weVzUBDOndl1lKZrWn9xriQO
1ljC2JP89rJmcpCaQ5KkxNE8AvZ70XK/xDlHwQ9CRCel71TYG2zSJKTRbnHlzGYbL9QYROjZT/G4
20Fh9X98Zoembe/C/Ii3vQwWNRo/ty9P7iV6HvFT+NpjF62PW8HX1I3sktlcKjBSGOABGgcxO9HL
PeGTAoubTWbvlEuYFWEuyyqty/hdzFIGX2gbC42HSdhpzDNuWryd6aMvEmIMx3Jl5OP7nZaFImJS
ffePuQgnxTZZCmcdHMWU+jCMiVOBvv108CM60lHCOnhI+B11CoeJX57cWO0RDoEuXdh6RQUWcN1O
uGXWd8PKcN7yhv4gdjAFSZaP5uToB4FPP0dFhMBgAem/CNiU1nHBo13xrmP2G8VQhdZF1MfmL6CV
CCoE6PEdgdewOudSxvJxU82Nr5B/N+ZDkgoNv95eJF9+E7rtAQ0nA8cOitukby2kIv30BFHuIYsa
+SF11GSJ1b+hHofSMsEGBFeRGiVd0Ywr/EobckqSo1wBx+43/kEjLajc7DsIFWPUdjop9fuzgPX4
Ctd9AdnCuY6Ne99ps5AqINmDl0z2ysgl83k8QkptoXPYhM0XZlDCg0KTNeP2bH5WrnXR1vbDl8Yi
zca8cyvES1bOOy1ykkpiuhONLDl8kZjTDeUkFDJNX8IEmr0obC/4eki3R0oxf5CbAgVWa1nOnwEq
8D2oNCQe3dktVGP7026rv/dp+3vVhyiXDRmNKgrM20J44G1Py5ghCZ6b5jikql0+KcER+wFy6PK5
FpbM1o0B+pAYKZQ5F76qBDc1D7EpkYv3l5w1pU7mKus/E+I0RGkjW9ERk9yMQcXXo5Z4dc+GWhVc
k/A6WD2DTWZ6uT+goBwalkuWui7NVGwYt+FqKONi9kRz1d3RxOyvAHHD3n4KSag/qcof/pr6s4FA
f9b/lSxRa/YKSn9UEbg6BP14Rw8fDxYMADl+zTBzYAEY/cqyvX2hXfxqFAe03V0L0urIDDCyF+wp
CP9+V7E4mUbovGQTz9m6CYnCBGGc5JK6qAbnCzXZVTp89gxRp+PkGec4Q0bRQQY92aSGXmHw42tO
+d1kgNwBrQOuNO5CM0Pxe9/eBBKq0h3C0CnZ+tfGwfutr9ogj2PS9fwFTnIoDz0xO1eyP1a0SDt+
91fsXuUYfoG7SjHmxLOg1TKANqqFUdyBr7hwWy8Jdd63dXv+h5N6VYHw/QVv1HV+tn5LXbykuijr
qJamld8zk/igMFMewkg86jZ3Q0WjMccykGa94+il5AsWcJ5q2tTM7KEJ0Wr0fihlkaiv1Mbd4r74
JHTGx4guOMdvj05+xaSeaAtwF7wNBYbcv+c1zJWcKbzdnsia6iBuGL6p6v+ZgcPFbio9AAJIrfS3
6XhMhEqcvjFUBrrNSv8C4JF6xGVSFTu4KoNo2kYUTwEEYI4s1gp6wBl8B3lXpRc5mNQqu2vE2OTM
BC7kLghpi8qjb7+Ew15NfIGwJZw3g7Pd5xYfP+PGEitcLqA8M3Lxb4lT2S0nZXad8XesN7IZHTjn
h6vlwQzBp+zq+C29n7WwedJRobzKOmwTJfy4bdMtSCxzO+6OIryGBW8S+tIedSOp/atR/GiVLK5c
7m+iTT2JyIrFjN1tpRIKZ9k+S/xYkDwNQBe6QQIl+4SsqqMZly5alWzZXoha/3njT5hDHBdp2Mvu
ajcRRk9QmdqbuGcyFicOyc1E+EloolVeY08KbEAKCuPw/AZU3bCQZVjHnzVraACf3V4L+qLQmGGl
7hzTg7l72lmxyAlDbH6mllxeg+OtQa9q2l/zUBur+IBDT6rQ8op78YooH7TUOiPYJoA5tsbcgW0M
YesMXMwtDTeBw3scoQXY7QSlhKiICTFPtD77pVu7sj15HsZcJF8E4TPhP0xL1Jj/1nItgnfMhB3A
9sRANDAM0a0errCX1NZVdUyrQyG3km8vn8wMDk9flxVUspbmC/kZS2hzzxn1As82ItrrPQm0RXMJ
89NWJa7h7yqdldNMZbisyIi9i2ETwo1OulaP4yYd3bpddUHBbvW7nIaWTk3FvQ6D6+fb0rCVxrbJ
o3uSxjabn6E+/hq/2xVGVg0QnUitJmUVTH5O8/6JQCTjHyNY/XmPJMUpAmn7LTaxPdmU9ykFWBLV
7NObKUkd7ZDO2qVdUczBXXMSRxAS4gg9GNAeCNz70pXgXOQs1CkKHoFdBnbDDAhNvw1dal3aqNTT
TeUwFJKnnVT8ucKouzm6RQqpOTvwj1OAwncgKQ/oSwU4m3flASHzk06o/wW7MQpmc/UUEhN/vLcG
GwB/s1qgp7ZVv+DrReQu0J643GL1+SEA0Rj7klXl2gu+hdfKv6vgXfvGOaE1cHVlpHdKX5yfLtAm
sa89JlPhi8DZJJER/AYiq/yvpswxl7y94wyOJVc0MRtuSqknguUBXUFkZlCI+ilbpQcS8i2qxpRw
RBRQGrfe4GIOeIPPZQWcBqK7VqkA5GILwVrkwWKGxMSd2UBKzXF5rrVhfK4WOGyU5CR2oesqRrrv
mSGbaf1phHzoQNzxSzjJfygUjNe8OKrTaNQ4mkHHn+RtwKwkrO6WR4vgU95cqdlWVX0j9QQ0slwU
xOlVzO01UO8xdFBV62y0vsd1EnPXkbJaqqMVIJj4MKQK+MMAUy+eur1yrDjOtX39WLRx2yczXz7Y
K91hyxUpFVSJ3S3tNqR4ARQFiJLaKvRmQiRkSHV6Dl2rk6N3WC6MhWHw7tOEMdQqnSz/cxlWqjib
0y53bsVP6bA5BGMdWLYnGSuqw2roleqKruAl1TuQu7ZZiOfMeuPwpRT+LOXOUaxuSwsdFgEsZ3H5
S/s5kd3ZZiIz2sOy1QVqNY8e/30yKt3mxnK3wZvAKMRCvNMcuOuZbaBex73HsCtJMSojyrSDoI/p
rVAu7InXGerEafTy3kts5CzQxFQgXwl40cQ9m75PuqLFxeu38RKp8KaBdmlfqa5SL1YrdfiFGFHp
YZVjt8POIo6bRrvUAmYvVObL5+9+zK+/8AnAloZ9wAAmHsqgUc6vXNyix7MdVoFKQLBQ/0V4Blcp
rFjr1VQmMSKNR4WysyuaFHRjIhRl7I1b1J7pfPZpYiRbzaqBfU204cTPieJc3vuyqDZQDeyfdPb9
Px4IXryLaKu8Ac8PziltW6NCS2hP8QEAdvIhJ2/dvcXkLdyCT9fxIdhnIhyy/5lMJ46ybry1HTyO
zer4n18yHvzFhS8KwW3szEzk15I5882ZuCt6N4HaJk05Ue8CyVvYYd+odvzVsiTUpxx/A1xVOIrO
bpDl7+KAJo40sRWrupVtTDg8Wuoyhf2/4pXiqNj899rn4Ve6C9+0oGbjkyc3P1s3RbL1bfnjmtRX
GgokGjWVWBIexES611TR5aXH8cHukDpEytYEjMJA14QZpNwCVJyR9vNSdoRxYNVFrBI1BwHmOnPZ
o50m6s40dMGuqYEOVgM/2/fwgPxguOZZFUIgTqa+ntpVFDkwpLxzOIAR5TRryqLHuYarqg6VSZxi
Ky7LlQdD1Vcnw8JX1JwUJTvKPg1OqnimyidtmkJHlpywGEK7OTGdWeKRbmNQ9PeFGhDg/ipDh5/I
kz07Z6mtFTjq/+7KEMRy4pS3joBrNtnioaepErCavFPBtKf5c+c4aVv74ODpkEVjm+oXegde2Z0/
A3oqzg/xAwP/Jt+cKsPakXJJIAj1iq1SqxPCBbEqtmcjr6A/vaID8DwHeiu4OikevLwJfTV9kXaM
lTrsIXrS1FvUAxo7em/BPL9Is53mwnpIO9OVS2Di2I5gvXnQvxIZHrbJKV2e6MmPhzel22h7k0sb
nZZoHqGIHAEJ1EIKLOY9sHQSr2+qxDh3HrW368oJlVBCocPlkbavz3IZUPxiFhOUAk6EvET+AjKv
0mhy4rRWeAzknTlk1A/ddzOolUI6gARRDj9AHWisSanLaqnGZNTH+CyB9bvGba5da1b1e5fDU9du
TjPr81bZfxg6MhvMKdPCm7HIE2I0dsPtCVviyoxIIxAck1pr2YZtlji5faA+J4y29SjPlVVMWogS
NJ5O32l3mOb9KC5G7AyOFkgH2hIjCym8ursKrHC6cJedU2nTKxNo3TIeVQMwufnpbnfTxVXJuaYH
NNt1ceCjweXXVKcxK0+hHPrB7ifqGlHid7OiZ4XU0ALTNaUW77CWbKPFBvkZqhKUXXMkmWxKPBLZ
ayv3h89Q2hxZp7y2rrEJO7i562NE5ZyVWnXUBN7MJW/czxtOckxEclo9if0k7yAUqd9zL4KQAmim
mn3uGnU8eni0bhFLQ2QwMMQQcMKhnpz0g5G+FNL66aUs+me5br88bJ6ZGGIIcGI8pB/coaG06d31
v4OIY58rvVv6zuJnX1mK7h8PEmdTbkWmDfecAx3ktpBJUzzI4QuWbebDXDMt9LUZjsQ5+piknjqL
DFcoSrt3vcOWs5P2KTNzvPFnRd5gO4EWILtrF1fcOeCWQmYPYAi4mlu2JioJ2I6uHABHJhhLADIJ
LyyJ+zNmlOIt9J9jlh9HCySEOEHf5EilhcElp1qnDynKSx99nXU7VlYNoKnlhCQCSbr1lWSiIXCL
ikRkTR/2Hh4m6E9jqPQHdUm/MkTT4XQ77VuKhxmoWwRajKvh5g18wC8JhGud1pWPmRa2EYvFIM2n
j+/yuMpZfdDo53BE7qr5p+wH6L0USvGe6lG7eyzXJ+Qt3SwpbUBPYwjjDTpV3AhzWJI71bN4Z2Z4
2qmOvCpFvyKneuE9UHgD/UhAyPE1RTsZM26jZQIXTTBfh1o+ve4xv+CDffBzOX+LPWnp93H15XQK
eg2Z00GWolfuF1shR5D85ePo76Uwgo4tMUuwTDMAB1v2F43v9gnvhW0WCUsjaQM1rXsYxp3uVsoP
QtSIU1INaK7cszUB6NH9xE5KK9L/Mpsg8Zz5PuHr4IW2Ky3VZuXY+ZdI1/iTnEzuMBrnR6l5B/+t
v5n+N7wp5/8Zj1vitlLpncGXlQa4y4b2Gj/O9liD/6CXF5kuhw8kO1tNp9M82VD1II8Xu58wKGPe
Kt1e63HFzPu894UT9pVjFDIlz34Odw5M8TQ3UfGQwckbxrqVn8eRjtbFK27aFXVRxSV5G3Ufjc7z
odutAu/5dUqnRjWJZAAmK+CfF8W+zsDNtJ2KwVCFna1re8+Y92HZ9D6hA7LMtwGe+F07dIQZgh/T
IyuNe3trGeeKZ5ssW5oKyZbaWeVGHbpEz+cruo4Byc+5MtA80ktd/i+ToIZB2Y9DiyRDw/MthciG
0QwoMFO1sj659E1Oh7FVRGxZIHhenVosxQ0zcoLzikTspTUP0ut5B7/onoWXIeWgvfkhYJApp0SA
FNozcS9N8XmkmT1VVbxlMYDmP/yDBuXGzAsyl72ORX3huUnwJHAu7l1d6Bp2IffcCuklPMFQYr7m
Eh0rV1twsXmU9Y3vQh/r7G6JKb1Pr3U9bH+zT0wHP7LTM2C+udk7VPBnBi580VVtrgM1W1aLCWVO
zIhMW92U5fBa2Vu0kvB9QmjlaIrv+rEULQbrpnWig3fRuUlKBWoPfkITw1Fh8GYboa/QEIZMWCDQ
eC4mTH1NloV0jernVLXHNTD2WfpZ+j1ALFAvXAmpGobWCZr4czsq+/sGGzMWlmvxtw7TdL1Lv9An
mG9aE5EdSA4rtymrQIt2h4gJicrHY3lReTuBsak6dMQjZM7tW5/5I4D50jYSYGSstMzL6E94zeWC
co2+ATyvVUYFkJo6SinRgeSvbbxvz0o3HMTbUEktCoUdCDrQnJKKSYM6F6brP0isODpMQMoGn21p
TgFUF+UDqzVOiiF4PIikYp6MS6+kF+kHPJ5KCFKXKmPdjM2PjUW/B0KUQqK1IrkQw9zHskerIjFy
r0Fh0VqNYRNsb5a68xO92ODdiiSwOsF5MTRF6ZWbDVlQCloaFAYouEMRBesBL7iO9gcRX0g0Pn/a
908TCf8qY/N+LUg1FqLzDnVGqQK1F2qEEN08jjp+6qsHWYq7cgUvQT0ylLFloNaPTFCvfYCMX+AU
fjTThnCcPAD7GyJqyJU4GIWYiQEJtICXSvPh8yo9ZU4MGY75fW6uANjvHM3aPv7Ih0RBhGL3Y/Jm
dETh7QJOWPbzbVSYucumSybAJoz9ZPY6K6c5gAIU/VFIVMninYDnCF0QbI03yrKVY5YRw3RODElF
lUspIVwWpKq97TWnUbmO0NL5i/1cMyOjdqtrxfd6aKu9EZDxegVi/n1K48WaAq+4BJE+1HR//fW+
2FuGK63HIUOD1FvhKzQNiocUOjZPAQrARQHwwN6xnByIbdFLJA942OqeeE5/hm+R+Hu7yG3dLkOP
78+rIBmxFkdHbahphLxj1eWqWVt9uvxR3mXla5HwrHl2t/XjqfnlGy1iY1f6ezCHdfFNMrZk2nMJ
XoarMZWpEj23yfWkmItbvp4FamJgEl501OHmHp0RgBBp9QIn8nkk+2rrhdAvY4LM8Fm85MkgzvVH
Nah9WF0v5RgxqMPrrJjGJPdn1tqgQ98irCMkuDWwa7vWM0tXcO9yU/1WrDbAbsnK5fXwySE8S6DJ
S5eAWVSTl/JERYFJUc+liKLaBHUKwj8kF+KEbZ8cemgFzi8AD9ZmRPq2jguGflnsaNaMTfBlB2yD
zpDFfbjX8ie6AP4Egca7GgCpqSIOxHndDAJmVU7g+5JNTBGHjYuRtaFA48X0Wkh7oURWUGxbsv4a
nJhZn+FYRA2peyJC2K9R7Xh7KZ2nlOaifSxXDWXcIVmctXN56Kg8FcO0P8DSdexlcnhWo4gPd5R+
nBKICEYPCOBrQjIQcXeqSke06BdXGJAhSrxbSObb1pF6I8HO5pWoJ9sQQ3MxYhlr3C3h7Gykrbmu
+cFIJ6Vplr5MAmZrYrXx6MWDhFf2jtWDuhqAOmXgTppxBKO0KIsNtXxLFyQtta/lyBxcsL4a4A6x
AkanZn28EC3LmAEmq6FZmLzOaC9lQhgjgb9IQ7sJgZnfnt2DcrHXGlsQfqIYABnql1fPaetJvyqU
w0w9uB/nl10/BZnRudwEdT34L2FGnsl3LpE0BV1aDN5+FYzUpn4PuzzCDPWBr7EKVL0veHmuAdRE
foGoqOOUiXaDQa4HZnDK7Fm/JdjXv+Pcj1MBkSnhUoBGXlCwMjyKOmgB5tSdAL3yjZm+i2xI7zDn
eMx6Ytrg45XbM/ttNLk/YqOJnYzIv82ALVI460cZz/dQD/qqb7CqtrPbGArN3+Ess7zYwKhcp0Tc
n/1UWhCsTqGKEKVuQmUDsswIt9DxZ/NXVahIffBUCuziDjPzltOgHH2sDeYE2F0AngiYVuuxseqR
r6hKVU//ubjYk0B6DFL4h6nQi9cdm6FJSVzGiot5UbEYo6nyClazJvuP0xXLwGofu0fm2HF7z/pI
6OyjrtkUgdUEnYuHxjTIayP7QFFpVJk3d/VHiZe/GRm+Qstutbt9ZEvYiceuD+w2geIh6/c7zGsW
awGlbzsgV1ZCkz8W/U9RNmJdOlChCIGX6wbMLDToLtoOSnN9Vx/TTNvnnUxs8Pwpnf6secLORpqH
ZT1pUZnnQyIutY/evEMsBlVlP/bOKB5gYs/Z9MLx8qcyenPkyUzQbuvULHxe41yZFpO2ZM5vGPNs
G3jQUrC28ypc2K4afTSlaGtfn7uXiKTDeji0rt9z1c4fS1imkQOmGWAJnJG3gTEJLhN4jOYrQvns
2G5vZn1u9kNYXn5OSuGZ/WEhSw1Ok+ntn7BBqIwoJq+UBRKDnctllbJNw0Zi2+EAWgI0KUa75rk4
6crW7CaNajiNaZaalIwedS6fn/qPPS4PUZEInDEP+cLZPboRA/HZQCR1LLMnPmbPozJqGw1jVhwi
vsoY6VX8gMni0zkj9y9KZhxu/im97Pnb2sS0/HH0d0zRsi4FocDFVIZKFylzwHf+ptzxzcA1Snd7
FUqITUalZhSHskhEwXAbOu5OlxHWjsrr70/HaSbebpadICb9b/q+RlE6MkGVAU+PEGf9kI0srJvC
HVumQDFle0Y6t74QNH2qZ25++ciC61TEkjJLdaij1n7EQzB6KEWL9PhA9SdN1zd53IV6bvK88tD1
Mo8e26qJ+lSrqEtE8NKYQMCQ39a7jZy85hDpnC9qQ7ttx2RDkh7hrkb3Ywu4gSQ/anp4m8rtA3TW
34ymH7YtqfXmpF5XF/pNtoSo7wl369PdMClkatB8QvcG/YJjKPcOLP9InUqLPFN2NF/kmjli0OUp
Di8HPlnRdf5YRdBm/AHUDlE/aN2qxPdrbImgaQp/UiCoHfWAf7ojv8PUZ6TLyi9e2YLtK9Rje0KA
S/df7arPO9kpNwrqn2WYKZ+zLnwrGL5AlHBxHeCAo5GZhd17Zc0AESthOOqQHlrlwWExb8626p9o
qoXfd8MwGUwlXW+Ab0VG17bOG4ifxazteyqUGsdsQ/aBUqXS34Sl9IW4axCF9G0lMk4uFtSOXmfe
dqp4sGohl9s7APswaK7Cm3VDCq71jf24xX/oTe504kPrL7ESTUa0nOtbg8565d88i/b9Mz+pGSAP
qkArT1a3ffdnTydgXvYnawPZ00WxRHgjOLGYD/SS9DL7SXXu6EhZbSHic+EW46AVmWlUcDK7QqOP
101X2WRc34bDAUqfY1069YXnt9hexKCyp7dTKEunw1gm2wsbd2W9tHV12DFotMV/VtUIq17rvMTy
4lXJUiA3BWry8JTx5kxpvPLBIHkFp9Z5YYYkLbKMdrf9jWk6yvlaL8hp5m0ul7W1IUHAroHJf9Pg
ixvSzMfUoQRkB3PCyrLhLzfYsmyaOqfBwg0uMRtI+BGiKNi9Pl8IJl57E2Q7YO+M8kZMWrG0vsE/
tutHS47vzfmOmItfT0xYYUnC3NNDp5MfEBUl3BwBhr6q17krB7UY96jmIcQLkT6X3CiGH9zJ/df/
sU+6MsUsdNNynH4TzP9EztUWXdIUJ58WjgK4bMb/gkRU4QSFHQ8+7Q0Z2Dr8PaXmPdzn6Mb3xt+S
9CN40YXj3+clNrnP5wgC2w/RUGXJ3njRTQLPR/dN0p5rT/nLcArLqwBeauM31De/DYh73ovBqtgz
ylLX2gjFRP6fv7pn4yfzVBcnz7mPuXUAR8pl/NAK6WT277yljTzil9uUPBpVTAZO5PIe/8xVr/TY
g6PVByOt5murQPb8twihlfSrBDKVzx+CyCcQ4Fn4svWxUHbJ8fyuZ9pvNraJmGLEc+cTU5J7c9b6
5tMOcH1seitBCyQSU1HqNthR1JegMt04IeGIBdKsi240Q8iwcQ5GTjL7d3ejtvAv8AnAyim0Brxf
sbu+mU4J7/2950VjP6KQU8mcVS82yzYWe/ZZ3hH8l3sE1lrWuefWwIk8jDWp76IeGxAH6Whmb04f
w9WnJLq2MIk68347U6mersrKam5RQtQNXUMhnWEYyTbj4QB8F6b198xYuBtVpqC0EiIJAZvaoUB4
sroarHsKDXTk56QbWqOAqT0PK0CgQ58PP/9mo/pW/02jAbNror89kh9ueTP4M6oWHeov8Ai75cf7
O3SKDEqES+qbLyD3QatDtOtqc26PlR6iKW51ym2o9JLi2IEqR941tH877s/3kAlbfUCZPzNzHETP
Lges9Y9dBUycUey+gheMVCFzG6pCwYtOWOzBdb6PrSvCrmdo8hBrQe4T8re3FflknJI5sQw3aeiB
em0g4MX/OZ0rKYIHEQ1aV3WujAtNnbQlGNn2u481V+jRr/XANOG+fb6ic7q+snqul72vC2m/qRHR
wjh6P+uPiB7kWsYJ/EVdtrTlIZjc1v2laR0YVmRk6NbvwFN71y/GIIwmMx0N5ewZeiIE+r4dq6zu
Td2R7J/z6lCJK0CrTFv/9GchBi8vqvtFXL7FxWcBtpOexDtpmcHEmBRW6IQTNpaILsOndkqNaagW
LJ7jMh1pGxo2B+mOrTti3K7pCAfZNC43Hw+X08lptHYYda59d3PFNrjXf2sS+rJS7vlZN0xNkcXV
xQXlwrRMLVB5ilZXM/AWUoaXpayGGW1texzFg1JJ7A6Xg3T5sMY1AqbPcbTe/wqFTlEnVNLBEOtB
5UkEc6GfA2N2BoeJj4X/NujLAcNd466Rp+za4nA3zmqTdfmbnypIxr/CNWGgOEwDo3Pna7PXPk0T
35XFn/pbQGhAquQWkAH1by3H2UmHOuQynsi2BrAZ1R0tDUJDYgZAJSxY9JoYZUvoQnT0KXe6diQQ
kAyXKUoDctBNkvoHpNVQ9GQE94Y/ccUBb6d13MSo3XwGqArXLJ1sfN5ioLxmFt6QLkoVIAPjC8y5
n7mMBZrNUuJRGQmAp8zilCovuB3+x2f9Bdy+O84i2PQyQAOSKu/+s+Y52odFq6ucC53JdCmOF3vE
1uUjAxXqyHZTCoWPwxH3a5eErnmVGZD5rhoSuNlBfDguLatnfzZXETLSVKQRvEABWP6ffa8lu984
0ZqiPY84hS+VhTg/b6EPWPsPEaP5WjB5zkzzNKbmgly3ZvmtpGI87a0YNLX5dlBCVrkhFDbmG1m/
tRBUCKsNophjRHGOmCv+mb0Yd2NOmBm+uUORy+nXvMvJowm/mmBiv8E66Z4zNuih2auaoib1tEO2
AL7/Y+r0qNO6WXxe1gmA2OGvvXFNtETYUtHNFg7mYlMQBPYawJ0s0/txwEl27OLT2kedKonQtAAA
nY/0cb+C61gqMgrjeBK91hZnOVywSL5B26YNJyLhTHd00YALvRKvtauR8qgPdATmZoH5uLY4XrZy
jKsEdrJs024YUGHtM/Dxf/Z1gOQls1YGJNW8sBiUm/Dq1V2SgHLwLcd8EX4+LVIgs8SoSTYqIGIh
1sOWgkEIZbsE/GxzfwK9hVw3wDFDdc151+etrKQeg/R7cPS5ten6jXMS6lrTW6EGaI3B1ZdycU6y
wIQs+pwr4eb7Ws8ju7gNRr7PKbVNxPYU+Cd2YhN5iRNyKlUFHXnCZkkxvxRiG0fid/TjADyvK/uq
qLWXmQW2966Bx3G4ZCtwjgpEaV6UebS/Zuc18br7lWBIHOux9ge3Hpa4EumfhrQaXiEPeo93cRum
o494u2Hk2rdbuzK37kw49WsBBcr7RXbKlYiEA+PQ8WS/rZHI1JC+s6PTKfVjJw6Z+BU6mOhHFweO
1UE7Intmgm/livmv8pflIYE6mbSpa0HmhhfF/Ghw5uCO6hIeIAOt6GK41vTRDZsq0gUAB0zZ3ebu
WqXQCjsmad0WBOKs6rQDVeDGvQav/0xuOTS3emaeEBsg7pkpm65bo1PSE3DgF2MzWIO8bEV2puhM
+z5dWd3tfIg8FtN6sMPKBywhg6uQlGm8mN0Nhtfq6zE9Y+kZ7Zx1fjyM0dTqUIY92L8rTI06regz
CD2/O6S4ll8KGUrmjJK2BcsPfKHSGjtGVpxZz3W7rTmefas9P7WjegSAgD0JOe74s5od/Tz1vVnq
6WQiuEr+vxafq2eQGI/WjcU/vnATgSKcL7NLN2zFjNkZq/G6aClgNyltsAKIWc6m37klA/CTS/r4
zqt6ITud6fBi2Px84/RPMLVXvtSQhpxF0VcD71kBDKAnikLTCshG/0k5lcm5MkJ5PVXMxHGJWpuc
3S/OquzUOTc33/YEb2t6YzjttlmeIoIimlqB0HRzuSj/6lP89TyZ+vUZQhAgNUdBIPLe3Ua+7fVn
GfHXPKGjJbOUw3yo8efvi1jFWojHgX85jTx5JW0dFFun0LUZBZ7bZJdn2BBsO71B631oCYMpvoWJ
d+6hHvRSXu6lvU/YPDJuGPhXSHrZ0HUFE6mMLBL1WsP1cclrGMguU6CtBKv9Zr/53Lq2rmnEzhVU
VMkpRLuiwlO6u37929mECbhmYenizwy1k8P6zI1zTHXymLtqemZvg4J7I4xm3Ua/IxVJhUtdiQs2
rqcEZ83POi5CUREbOk8osZxjRB+MAaB+D5G1FfxhsWiJHoRrDNOsu2atxNQ23HuyfZ8P0wvq43Hl
jlk29otIX1jrJkW8NLSo83eok3gcB4a42COy6USDYUj8cYiwFinEur0/DSceMKMChEQZQ4v7x4Yh
I9MCRYuCPkCcbvTibPJZC7GXHUWrIff42sbLLvCIUkNF1jbvnuL/bl/xqRXgx4wd6c2X4gBUirtD
x+UK2HsrkWLTpSoearGB5ozwcPvrPGzLm8JwjEPsixIGDjdghznfvU8xO2/jYR2s+pUlpWGjZWek
57ipTlbJS8/Lxw59+MQCe1mz0ubsU9htFkC8+uKDL3eo07goRzp38Mzud/Kw84qTV4A5Y0vftfPS
0XTX1J7eM9T7oJpAm8DFwHHsmMPaF8TFnW6qLel83OdJppj1pmw5FVTIFGnAe4J4UkCSwnUpdxTJ
KUREmfLPBRE6Oi3BH35PKdBIvEpXRugtQ8dscgVnLQR8HROz3FhufaIKdZwYOLYXTabXnJHUwLcI
bVOh5GAwu0aw9KrRtHD5bOvGrvdvDihomqcn1S1pdVhZqZh+3E1jnRDFMmIGQz4cPfyLjxQ9vyWD
O7A70PKND1jtf7cPK18muNv+/ZB63hKUtwM1cGyJJqTW3OOJJulE37nNHWllBvMngpyf8H1Ar2ep
zkWog3cuodbwXvc0k3RfiYZbN0MgEltqxcTP2IRL+iSRIgmsi8w3EViPGbvescYQCrTLTPz7zDIG
hTSKCXAS3khcYfgJB6zOlVIs0veTnj/MYgzWz1NP0nYYM7YVDgXPvifve/LYgrIVwy+TNBaLSQv/
NeW36dX9cJdl/IYxjx6AJdZP9CjK0BPQuhcALmYZhKLekDFLzv+wGWuP3g3GRVBwhh5ByBqjClIM
KMC7BJ36WOhlHaNsLGQ0rFqbQuObAobeTCzBPY/g682FzrlYcUlFT3q0RyNxMges27geMWh1pGXM
dJ2LUzNNY0zzDhD7Fs+YuiJ9/ViM554ZhHA/7ewB02ozIl8g4rsZLw2EEaLQ+k44TtZYh86HIeHW
qglIlFt10F4IfeJ2H342m/hwc95R/f6B7cxpkfaqrmAsV+Yt7vvsvHEQW0mGlFUnXexC/f2urqWx
KN2D5WZlSth8wJo6cvUzY5RpKXtJfjL83K2+gKBhc+0rXvLlWYgMWZgydZSXYrS1KKW0ojZCavei
RU1AyMLCnt80/4j0v00zHQUMY0yMFrkKq57pVfx4CUdKzP9l4c0HDoHJCQSgxUys8Ii1KeBcOi25
YGLzs48Y9JESjnqiKHrmLzZgZ0VXKg2ZIIJCj+g1ZB+3eohA7WlNPr4fQhBcl1rlHB7lflz0xqh2
aYc9jVydicAdVi5xVbLQupEsozXKpFSOLBBMhZ+w0UkdXScG6gzwRfZGBOR6GCvoTEDOiE0k/JQ/
uvnYx3VStPomgIUEFf9Zh9V/LIX5eE5K1n5uIZDXee86ptrKjT4sz9O+0BCwMEdxp/+8M8U5Qq5Q
HM9NPdEjIMZwQd/0b63N91MWpLQ8w4AGteHq6M8bb6iyNuK7DeD6A+BNbXk4uob1NyuA5PjpgacN
N+s5Pc7x4xydtV86sJsY7dQTkTstQAztoEAEUev/uAUSpw9VX2hR09lBylATrkZg2gvmDJJF1MqC
PRjIvOdSkep2QYljrnTc+OAdk1428CV2fkN84LHe+w1tiP26ym1ewGONnCEKu5LFw0/o5w5I03yW
4Tfw13E32yJ5swtA1xEmETqFdw7/6aSh4DFlJkHbYjtECH2xCs557Fpwne0A6MGka+/TZaBpL4Hg
Kv/l7Gkh0X1yuDz9qoOXrOoS48ZELQQt7rSfoFLfKd4Pov1Mj0Eb4hkELfZWHJoXW/FNm4hy4hS2
LD0Di9xNwLL2AdGnabwz47J2DJ3+aUqItuiEUfHDWFColqSmNVUc4EMWPfTA0kXxyxKADtOyex9A
EET4wJAZXZGm/8TUyvR/RDs5y0euhskNVYtMtDmP9ZXIM8SwGCD9AEKiKDaQ3dz6S+4bBlazSvk+
ib5xsntYLmc/hGev0QnrxYYeHu7RxWp94TAwILO2Sn/Et3tdsWdv7BEoviiUIEvAidZ7/IxGqVyN
q8AJS+vzt2r5G4ajYYj0m4s5Jx2VNuaR5j+lxL+16jkSLvEyKxnKwfv5kPgOMK9M9Zcdr2H1AOgl
eiUvdt1dVtxIU/MU67ooR1kNfqF3OKF3THpOpYPHkeOASjy/dvVmsI8Kv0Hh6d9TGn9fQQsohXKw
S4fSenmbQNXrJNci5zlJRPAA8YpJKF1qm3cGznCXpCn7GMgaZZsSthcDS9lsmfog3g1w3tu/G0BM
NzBesXktSecvZZAB40rSxu01FsmwEQ1puP9ZZEOUT94qGuzL5y6tPOsJO7JAuYXrUKrQHHQMN7YZ
9cfnCUI2x5pfOKgo6xv53JIBlWpcPmwaxnAeBagy4tNAWEZ9NNFkHvnpu4uGQJVjBumLFR4Ftvis
XqvBNN39GjFtaUezpBxMXjFBv+HjU2RmiNsMXCmfMicHeQu2jeyyc4TobPyKI8ccyk8hcyKLsajY
IUDea3+ThdslwKNfVBs2As898YW3iKMHI93ovZl6I4Mhk5j9l8nrKmJH1CfpTvF5nXEaq+CqJATR
2Fu4EIuvuo9dMf6OttgqukYqqLVwSpnBa22ZImicu/+PZQydp+SoUtjqUAi/E8QRb51UodZXfGcK
Sk5Xysblsq4VY6WjvziJvf1ZmjSc1TmjpQ/nN+qX7pXQunf92MfczChGvEVLFQ3emKHGuWHHB2iU
C9oZyzekgUjZ1SBV3bHfafz1/98wjXEfz4g/q3HudSuzn7eN84dV/2LkF7LzPtEBFhHilCFXUYD7
l8B0s/2qKCY5DApEA5WmHzP/hVOoqbPdaEA5mlA4gKkcEOfncjmAKsQiyRQ3ZaT2oV6fDn9oxuu7
ehzZnLvkJKpoiIuvtGuAt5gnd9Igdhb3lQFBaOA1aDlLdIk4oGrn9XrruDJvNA0VpjfY+SQG+ubt
glA56GoA/pgSSN18dbYsTP552x7g1eTTl1tMrLEOc/+SokkoGoCJid4quGm4/SUfg33b3LDCTZoq
kCyQW2a+CQjgC3NnUjEgIVLjM9giZeOpOnC57W5kEDVt3nAcJ4UDtBHtG36uX72ogFiUJdx3wj8h
3oT/n1GjEMZF1S0DmdVQnw0sYx4UXtQPv7ILOPuEH1Y0Av0nHnlpNsH29Nq+4RukqQ4nrHSUZgqa
3vTxFITd011p6w7ULgkZO+tR+PTyONIng62xmK2VahycR5qIjTeSj4Oql9Hv7u6dA3WR0wOoYa36
HKcfiyh/BKPfbOXbPX7aEb5Kt76lL5C9Oyk4sLcYJaML/p6ohK67RNM3fQnzkMrJwuUcJEGoGwt1
0heitQCDg53x8ZRmRbdvL3mJfq8A1x3ZohR05sGXFr26AlApIwlrNLWm31mh9xfIt1n8jB1rU43s
pVBuVAUd+eTvrO8LklscIBVzFy6WrVq5/24ynXGWoL3P1cJColDUieyBjjAe+GvGSIRtgkmdObhY
itPpRqr4rIMEkIo2tf7qqTtqwEim4rgMCDJSMmmS/rQs6tMpUrYfuzChhNo2RglN21GRK8wiV1GQ
TchEZRgt6X+WDKZN97ihHRum6pOojh7TRHah08xffAlZRJPZpvALrYjOab5Cy2GOwUsh+bS6yd5j
XAcAcw62BTORjfJjqHHU6se7Vd8QijfZgHUUHeBTFR3WfmouRz8NM9lzwtVyZKkWEgHyJHCkifzx
Qgg6KpoDep7HtyAcZ6TXJ7NmWQU6qEKiZD42jYgX0ev0GRMgJT6Fb7qvt+nrnDvtLNetg1u3Dpp7
Sy3qYWrVIktD2ZR3qyOvkt9Y6r/7x99lI3VL66BjZK8F4I8L+qtXrIXcDkNn4abPv8rb9Km8m3kQ
3Ofb/E3HW9V80cIP3cO120ZTgRIUBDk0nLNnrodcHCYxuPUwUvJloBbbsykXj8T3PBRt8NISorEu
Aw/iD5PoxWM7jPY+1MrOpqhDSBiZqYIw6lOxLFtHYRQpdCR/ax5TcUlNZNJSajQ/qTxneTCTE0ug
O4Sln4lHJRckXlk8Ot5uO8DIiV1xRL2jBN76zVfZJNyPP+6LWKFL+n92BtZtG7XMyoLPB9P+pJFE
8CcLaspPWFGaFmifRWIUPA3fwAMc3dY30pbiHXOZU1Zamp/yMxNM0SIeCtTR192nkXt62Aw5Y2wI
U2bkMclt22VkuxPkly8TYwNHbtO7T7V4o10FlBdCsHqVu3VdtsLCYyBSPYGbrHBzdw+BTf1IDTqt
8/BRDQV+RqJYwWDl1XWJjMgUum7d1MF1vpkGeugoz8LuLAMHTR8BiVl8FkSPuNeShqKDTtXSVYk0
o6KVfth5FufglfAAkW3O/4yS7IRxfcTYKTGGIdIPIxvGzQAmlIHBfDMGxnx4R5XVRTayBIaF+NlL
Ia0ppFIZi/0JnOJ5kJsm9+AAtyxya9NC3NwLb6WknFty/s0HDEWkw6VfPx2ucwd4V3Hes3dQ2As/
oKgMDsMtxOd/PYEUABqUnuYrzKhn1PbhARHdMmtyTbuFVLjGMLm2ps3pINJZ0n1FMtJmxl97UPfr
VY5H7FNNUjXrIjzfJa7iz1Kg9AvR2s4Rh4YzYs0wRY3OUhD9dnYhXlUhWiyIKW3UzBdZvaYzREEY
q2ErWYGds7cr0KKimwOr0eIXjCbQMndogWK1SUOPc3pgNQxobUGA2JvxNf/8j5bNC4KqnxHc7qrI
ibBtCqShTi43HntxWl8MvonB8vsUXtv177N5ODu+YmavgXbEaUEvDUmL9ONpqVous0Ri7r3ZnmIX
w5Newa16yQ0WpYJt6In4H2GIzhozmkDlKlk7EVyqoTU3WOfiGVdM7GE8PaUFUr6nQ3j2Jl6IUKtc
Xwvru4t1UvgcZ0Jn/2LRfpTwPjizNz+apynTxvjlyEF7DTvRp4cWItwkdHH5oB8ygw74ptfuWp9l
CbRJ/o/nKd6fJT25ia6xcUFzF6ydOfegyFBDaYKoCiooxB7Q6FB9iIgBvEFPmSqPEMN2OFcbtf2j
bCnAuZ68rvxQ4mnka9Rkg9U5yksl/xBdmxstekS2siJIxtI1HYqRhNL2wZF3gzQEYmBF43f4MEAE
/tCNPM5GsiDP7vvYrxshDNFLgQR6vLXy2OO3/el1J6g8Xx+WP3HAS9CkWsIBs75XyOJdacppvN4m
Z8Cv0Q0PgFNM1I1s7CND3h634/1U17DCUEmQABgZkKdAun/+l2BnPr8tJ8CEGvQDxZd+BAGOOkmX
YrzmGbR+eoBXXGXwOA3VHganMeyTjq5WQoy4q2icbO4lw3EdEDNbcoe3p1dEixDcN+ms5V2KpqyW
w08UL/7JpmiNSEkJBGxF6WHeKagRCdSUelQrl5qdKhl23eHy8v0Y+j9WjBSOekR/9uRdhzdMDuIx
TyRq//9nMuOqM1sP4AFnPMIa6PaVznhw1DpiEpGdSmDFRN5RV5MTaPgvi85Rhm+LkMHFlJZFB5hE
13KMXSNqRql3Mgrc/CWVSAtesW4yzAKdt02Zrtt9iSBUK5RpUpI3LmdVtTbNnPs2S7Jrl/xZgxXy
qvseBAgQy49Jo6Ju1q0uHDtyS44wF/c6jGzR3p19Pr7hfoGPY3y666P7zmRkms+89+HGOUCAT0Zk
MmPHSGgU5Vph+mmjqqM/3ACT45i7huRm0LBYud4pvd3Nkg7zlDyW4/I19SKiIYR91Kzkdiet/UAJ
mf6TN1pV6gYw6dAtUqYfCuwDlIZcLkdY119nhuwspKgLOd5Hhn6URUONO/YXmsqjGbtHuWlXooJN
sjJQns5ZMkeR4dFvYtdHkyQ1BitsY31IuJxOzrSBIFH3K9fXtKK1u/OBouEFFIffnrNv2+92H9+u
8EmE+TDhMmiwGyyxVKlHKP9d+7Q9GIknuTrKBt5jxritYT/blO4awudwFNxkI1XLPjip2EbpdSyk
xtRqY/07YHQO4ECVNxC8SDgQzrbWkJ45ts2dvk2q3AxwCd7Br6ex+r7nASFr+k4iPnas+wIvSreL
AQJK01cS3k/T1UEsR+voAfNu4mtMhsmoZ84WXiiwa/IKIPNVruYdJnjI9TwfqPF07pTLe+9q7cSn
ljZpPvybUYqRgFjGwVCBDIPr1ty9ImGNnmOQ/YDx1fV/Ap2TysBAj7tftwQUcinkqbN6fV41vhYP
1HayMSFSIrwHDxIRPPAoOLL8b2Ovwx6HOfKUPS0O7T/DsaN2yCd/v5G9xEypDnQRUggpYbTe99/e
aVl+QyW527idZpZJk3MVcNTvyau30pVHCrJfkewmyWWWvbx3EwlMYTYls+TqP1Kdo27zPd49fYX+
YrnhfHN9k43mRRK0iWTQj3zk4ILByXDw80cDzYFGW5o4bL5mQtsvdvMoUAFEcXWlcENXAet7IOVp
vwiaERR84yqWm05q2hQQTZecNiqwUJ9Tgi3TML7BhHMBOxwKQbpDhYIgjeJFPdGtQvMhSzjKpPzn
zvlHC/u0QPmkTefMQd2g7UCHhKKVm+HFUTFImLedWoYxFvXb9CU3vwS82pGgYt5PiKU5nSFPtd8Z
vFA0oZvsZruNOAt9+ATUFHwei37bmuEfGy0VRQG9ZEwTWw/eaGzpHkRQN3lUgCMkyM8WTzY/jPju
y+LzyWxgXp6aIolYFG5KC+k01YLOv76IX0Pw+NFEeNDVU9i+4Jap1HbcHMWcZJHU7a99FrEetl9T
HJx9dUtpR01GNBZ3SLQrNU35HJ+Z/Iakv39abba18dOsyxk9X+gAyeRoW0Xzm0dWhVUq+zmAEUlY
cul2aTzAayIV/e47nZglPGjTMjOtys1iv6FKsBgm9tmcJCNtmpkqaegaSoozPoVR/m1xWpVzMQw1
EZz+dvXzs4xV48n7bJ2SszDpOzmcL20I79+zu4QYneE3CFPP4m9Y39PnebxODGtul327UeR4PPoq
kJvc4fTv+aO/tMr8wiZclFgilSSPGGP9GsammpTejj27Wz2aSSdSMzeooy8v+Mm/KO2bldT19G82
c52xuVgUKHgaZJuYx4OeokKWpf170b+1p5GOUQNds/4ktZMlk1RPDK2vYsW5dKAVSw7B/PVGsjfz
C1ZVesxBDqXZ88Ag1SzGmyGgjjNGGUl3jn8oZSW64Cw+mVh++ajlze6yOmPZDYL64VI0huOxXXsr
aG/RUHC0bQLxNey9DEazLWzHb2A05mvOwK0iPqfrSMfu5hf1zbbeBKlNAjlynkp+bOXeobVZYzHt
wMWTnz1sTd3p1SUDUqu0XWC4lkipxq7QQlxG+ErHHr/dfArA3TCZc88OQg7A4M7tyRIiUeSMfHlR
n/ZDwSIQ7xjIK5th76484f9iSk0oYZjMUGdapZ4dKc6SNa6discQwKYYLs/iNRNV7pKbQbM3p5V9
B1WOxRewmXslDKUSk8xO+RuPNcVelPPFFfOlakkLqaXXwPER6oDwOr5LUxiwymS7MpVYF1lDz4tH
F6TEU8JZCTno+o9mlVPAJFTURQ6EN7KVtqFRZ6J/F+avjDLdiJbDdqejNAQUUVgZTE3I5XDEqV42
OJichtZBTpCXTNs2lQjisgijmwqBrup3Vc6lzbdnSQUoMyhdyUE+OF8oQkqbGKX0oDehvSsovdqd
30Mjxpk8TruUL19J/RyOnXosOwh7DKC7RXJvLkQuq573dtPyeNk+ymsdd4YG3XmGw7f2m8tq3u44
9Fg45XcFWcOLqSEDlote7EfWbSqZrzHSUzK7RnJHn0+RpDKwcCmq/l+7ZeI8zQj0csWJh5JExCkS
eH7eTKyp5p5PsA8gukhBu8Zhg3SbWFrhZGbfLqqc/aQuHR3c65BCHywxmZ16quOmVu7lw+jI56TY
oLXELYngZZ24s05VyZ15LTFTKqhgU9RJSE5PQhqbhud8m9LRL1I63wM2Uuvprnc5vh8I2rVid1Gh
OTq1+cPv8ZxS3YXpjoL8sjPfiLRCLVd9hAPDDGkn6SgClqWo7gLXl21UYL4+Fkt4UZv6qvQrHqr6
LqHAvI0nOI8BdhjCmdxaL0r23WFNB2hhh1GQ7dJ+tFE9W2b0agdLR7A9/Tbj84HrxsXVBn51PITq
QbD4T89WrBpCdZ0NyCABN+qITuRANVf+gCZEWQyUK8Potv7sP91bi98lG3IE9QNvAnuN56bp8tzO
9DsrrU1mlKZQmwkZdAGT6xm5IhoLgU/KuRcPEF6PND+Lf24f8VHwpCsN/3gH9mEbLKVGdOZ4oiHX
KxdK2e8Q447JoFmwjt0b+IilqPxMyBLIEp3tkyOex+/Vh8p07Cqp0d6P2q9vr08+AzFX+jHekuO5
U4EDSuWDfnzpT/RnIneaKmOUHCgYYiuvwWmSY1xo6Pg+nO7B9IUefAJCo4gNYs3ufPSGMJxGTizK
T1+fxepTV8D3aNIhDSVxW/EUnuzjvsuDHJeHUT9Uq4Zrn2Z0rRwqjaBgXxw+y2ok2NOVENhGMqOA
0ptSxxXpWPttrM6vmWtB+FwlTFAe9Iur/+xLT20tn7tJrKPf9ci0E0VxfdmOnF/EwUwyT1P2EPS7
JfHItZF+t9OxDY0VFvnn3KPgqxYW93rgBcxXTHsEf7im9ggwEMHqOHh/nQEN/vJaNjlsMTPQ52vk
NKMvyCZgQ9QlPZKujZ+zwj3YY8uFWzX0GHwRFgf0Pj3N1XEXKNrjXHjgIMDSPJr4Y9KqNSacGD8x
cQmqN/zHsZQhovLGYnJ+mANxD7787OeOI/xe1QGcWf4zuZSDsSH91J+Ozx0NYWjh9w0sO3mS2eu3
/RfSpeFHQRQo9VTaLizRGgFR52HHZ0lC2C9jKgKxvATlKe/+t5cRiCxf+bQyNQ4HmDpRZLm8ucrF
7xFbhsA3VgCZehjA3BlUiApDH/akYUfkBIBGIjeMwpLlHEyAlenQwAMruIyHwv+Il1ks2kgI505c
Xp5SAUd5FtnPEUI6OFhtoyMrachQn/QNZKeDyv6y9pJPNkPqc0cUteSQeyRqnEx6rfrJvJXC8q88
E+d/KSMfpxdcVQ0erWBEJ5N5ZVlpEALo+tZF8JaHLh2z837fd3sjH9BhvmcVEobdfdatZ0LC13to
A5/1grSiad0gjnzUaTJXbgDryQZ/07X/wMxfEDinG3lT+OOuCY3+VFqeiR+DAOeVb4D9CeB+cYnL
ApKnv4vZmPMdgwXWDI8ZI4llQtwrXfw9di52Tvw261IM6Ed82nWjYi4GjBTy5tQbyfzhSPGWsxAn
VodaynKKpFPnD4fuIsrHu5GHSx1f1XZ4ljMdhu+VquCg5//3k9Wyxah32D1Xbz9KT9FtEtatZI/s
dKVlc4frP9C8W3CIiWuSStHgnnZj7y2w/xzRiCmT1KeacSu6hkG72/WvoFtZRv1R64kX59vefNPT
RUQWpCgBHYeTEFvX6liJ+7zF24QX6hDySNrygGAnRrBzRID8MVsQYETJTSOZinygOGIJl/4hBzOn
0RinCrS+9dTl0rGekKPvbCKPe4nQ8xaX9dvVQm1JbIF1vN9+fBwidfKvqVJVl4zr5EZf8W4DrIaP
Ef00W57xkCxFIZBXBuM5R7ktxipZG1/3IvwzG16OSWmAlD8JcY/T4qV8AuXvCoHFYOD5Z2MWUigP
+Z10LVw79gvZ4zr5OVGno7tzhdIOa3YVWtEFqERX6mraP7u8QwYlzzqvl9exFb1RL800Rh4jabBS
Rvpf/7Yshe+tHshab9uXffgo1clRodFXNJ2SjUUrZlChrD67JSTVV1pLWhQ88W3RKKQvlfLKmq0c
YOmboBIKNAJEXIy5mh2pczQQC17r22fWkZmxa0Vuz2+jhBV0aHuuk3S1ChLcHyyxmEYWNpvvT7pu
ug5RfTInEEZoXpi4PrXYCdCvjvVsPmbQNCBSis+k6jYNonpWeQCagnOlK+qbJW3Qnn6GK4C1qSBP
z9w/sFzUc+JCNaXm/uQRcVTnlsjdTtP1BttRRIGlJZeEttNlSkGAEC8kA16StLm68HEPiFwLHz6N
ki6jt5cn3GPA5JfG4X1pcuZCfWsjJiH9Lw4cQVTe4GM8mFq0UBTOhBVMWezs6c4IKUH47/ThxEpt
ulX3nmfIZp1DKe1zwv4vhmyKB40AURB1D92nVTIQ5+Poaze9JHIs+4fIBiwQxkImZsN1RpY4mnU0
fgrSAn215v0sFeJIdzmFhmQh/GbCshIjZCqmTXrw/FIVtB8Q0KTSzHvSIFJXiWEts4C8cs80R7Ig
0OvhyPErojf0GqArrabXI9PhNgT4WPknUR/0wgylOpdfGRsbSo/v0nRL77OsLpkxJv5qKespeoO2
lButlLohpwCRz84TgTYqIK2yOtsdsJ6O3AiuDxNLx2xP16pP9EKOyLS9cd5+RSlqzT3m6H/eAURw
poCy8r9xfe7HRauwaczP0vE5J3GeYGHIB4JEmc6sCKdIO0ADqHmA5/PXNsCZKmUVTNFLw9rGdCGJ
ZwQDoONO+WZY2wgG63ANLDCEim/8F/VCp6eMJjFhKWeigUxFW9kLU0IrRAFz6I9K+on+P1RtRcq4
oWFxZ48sfdE6Gg2qWk3UgGk78nu4ADmRT6CiiIQTEmCctvXSfXgXx2mKPr7/6spTiITAk5sGHOvQ
apHgqdZdHwkDdII7W6yh68JxwnFhmVl8lo7Jsie/L3rdTljZpmCew3APFFmpeGDNcNiCdVgq9U3Y
5Dpq9bUZLUlllV6TCoN6CO6YAyUl6saosdSnTb4ijPJJIetQ2PnIZilpDUJUwzX69FOT32/WbpcU
4/bEwGuhObycs//k/qlSdMp9kOx3E6/e1AFNAUoG/PAqEtPPMtx0LIDq3+lBe2k2v5n5R0C5XePl
eOfI6dhrsZqqBKBfxPDlmy55tyCXxcx1rt38ksjFresAylfiYhApkR+ruTIyOqYJ/Kl52+Gp8SdK
ORJlWGl+1Xv998MxsHRVRIvUSkV/ntM2C0f9dlXscMiKGYtbQDll7IvT3pRpO2uLuYpYx0ejwLgW
2lvipjrHe/eux99yjZoIYMh/zuxXh5p/MNpV2qLhQGJxYGSsO12QyjTeKaumphW8lt2ibbubfE5e
p1Z+2U8HcZavZ2qrbVyO7MGQ6Ip7Ar7dJd8Bf0/MFyzVc7htLuZyuA7X2xShcYjJdRAclt0Ci88Y
uy/HP+yVOS4y5nGWlfH0fD7eJHe4ytUYG3QV694fZVKjf5CSRFVFK2nUPX4kHnUzOUkxOXFZDdTx
KOlfwAKX8gYpmQeME76dtn3zDVa2p4YJyzy0JQ3CuDlfqrmO4a27rl8OPX0rngGdp5W0rxX9qTT1
BOOhfS4KBHMHYypD4h0zQapmbf7tQG21V0cTNmEtEFZHSzRUOfx26XqS60J8dxwjCuwIBhJn/N72
DKDf9hKXnVKLTrDLgV+ubjlcZPsur+rMhZYrJy3IvxdEzGtShBMjVwP1vrBkX3Q5POJr35eNRX+N
oOinJqr+nm8cMqWMpSdkCPw+Oaijn8Uhlq7nezofFQMt0ZcU1Jy9UAvkQBnZsWJxQ01iTzXHjjzX
wLtsVx+r7v7WVNSJRyE/U0v4gvt+Dc5YWrY+kifELuaV5XfW6hS8gd5VSxhRcCgMWXys4mOB03lN
/7ddQAHOmMxv/TldlE3j78Ubo346FWJZXgyeqgyNJlNQPYtUhoDlhq6rlVJQMUXfZ2IDIH+VKh3G
KcOUnR3UAuAM4J+cGLIxyL0AtaXXFFO9EoEkXooT58e+46wxU25Lj6kxhn+azW+4NxSFe2azuON+
gA78hYf7DE2vfAlkz5rnA8kFqH4KQROpD998x6jf6RsjAPlf98yy/JUWpfZN7TUmyZM4a4ibwJmg
ghDkAxuPAEWkckZ/BpihZprwiakJ02uFfzITEdk0Li7zlkZ5ihGoEwQq0xfBm0fCiGGQ5cu+JQjs
fnAc3VlTSgqrcnLq0iglvhYf5DGU4A/akpjcPVjp/3bp0o4SGurmXoSBpCyXj//1Qf0OzGvOQZ1U
A4Jv4y9oFXQO4PZQfN6OAfAIQIs7s1UBm9NXIMlHEE/5kTfFhF/us45ZImFVITMYwYjJh1iQ6WvQ
F3xe5CsBERaYPuMllD/0Hi50IhbzbYGD06fC6pvQ3huePHeOSBUn06+6QlGxtJLQjLIzhr1a0S7V
4lGu+M+tJ8nS3WhkeBMUNAFLAOfOicWpr1AcC3Ab6QFMUcb4X8tuCPfe811qBDfg7o2cHAFxCA9K
8kPdd67+EY5qsVJZfTEjjNUhWrP0V6nhG8MZV9Sq6uV7G6Vi65cLGlxKkyq/YaHQWcyEmACTlGa2
63jQ69GhtJ7+LfKXWFREdTrv7A8GJwoTOGphpDTt+Z5hs/HOqQecELOe+XaxXquiq9KcFq6A6MFu
AKjSBmlBIKxwAlKTnStEP3M83CJAgy/+ihvciK7EsMEWjmIZtgXoGZnLcIX7X3t7gzNqdPeyLlM+
ouXkh/WBHyLYGH4EowGNC01l0iPYa9GISQqA64cJcbxpBNOubf+x7+nz8e9UY/5ONLjVWgg2GPNz
rNWZL+cJhQmNecF/Deu5RW3/4Vnx6MYcVq9E8oFlt3ceNY8+/wDc0EoVFLBAFGPwxt4VTVDIimZy
Jhu3TkI5ye/7/oS93Jrx7jTPIEzfjL78KAWDOE5u43pzJwnCdf49nezwZCQuWdy04TDCLGYLa3/R
umevuQsAGIurUWIXyoqEKFIkpikNU9xrA+Ykef2eP9SHVRbRrWb9zWa6YaVJcGNlz0Tx1b5x1Ylw
0aJzXgd1zxdYZKghpUN6nHhqOmvkSxc50aEzSCvAXCukH+sKgi+IlYZiF/75/JrAA0r/Oul7ZrQf
pahc3y8nzp8DLAeYE1U5y1rMjbPpa5PMsbQMXawCvrhr1g8mbWIngfteqaFDaqioS4Yv07XacJBy
V8drYYMXJoEuqqXi8k4/9E821PTqYRLE40Gj7jrh63pM6bbcTJoQ0opVAxXPjGMfJyLSgg5q2KOr
OBw5i37t96SA19gSM/vHoDvI7poJSnvLl296YVufg0x2HinGjMC4+FMM7XfqEpf7B5MVnxK1s92c
61R8vuxmCoYjNmd6K5YPgRevvcDyxSEyrX/fHD4QeEuy7ZaTA0r58v/5kDv8mfiYsSrJhUbY+rQ1
RC8811pzgd37T0kLaJPMX+yF5gne2SicPzZJFM6veno1qjAQZ4HMvcOSwn2Fu1aZu+0n8YeoKW1z
K0xFOVkDFbiruabCBUtlwX0mQHPpY2+/SCq1DlrxqdM+1IgB7hN5F6noRU60z8DsY3S7g7IpODLE
Saj3qiTq5fgTFrEgu/GVj7ypo+IGaOFRXJkpYWD0K0/nHa/vogzOJoug73T3x2LVRYKXflUdC636
4I1BQ/rMNk0AQ0kXR+uhL1wQPRKUX7d1rl5cYa1z4hVSylZ3OXZTPMABEbug3g6OYU6jT6sBs78a
Cb1wZpHUDgWgt9H0ER945cVgQL4tZPL8cB4dR6OmOiQsgbl1MWA/yqZi8muhkQbwAg/1HQhug6aL
Jkpg+GPnCzuo8HWbRQ+e+e/oMkPBXCkHhlyI/rL2s/X5ytnj4pphbkgsTAyQt6QnxOyvTKGCjMsj
gkqu+Wfkev/+JExV2nUCG4UEdhcVCV4KKwX5V5bd/lVac/nhXjr3i0qGOEuPoRPXEhUYL6AL249c
ruLCs+niw+qrJY8h7sL8TMaF78XyUZDImNhE/ayIUYWb8MIwR2tAMyFiUU2HYUfVOglOWj76eowU
SbS5725YmgWbpD0qg8lBJ4AU1yyR0MErDJYyFd0k1qPT5zoqQKE4ZUA2UMCO7ARz1SzcsdyjNW0a
lUs8cGSFyxP5A+ABSamAzMVEseqRWlhV6OEOvHH5G2MsXbM4FmcyhDHIfeDdgx1sYp1qTSA3CKgV
F1qbuNRxtYN/H9mCXKnZ95ERL1cFL7DMxt0Q8miTyKhiPicCiVXwXKrca/AH1ahqlGU2WaaKSlx/
T0ZyDSvqh/DLqvb9VTkHwNhx36r0WrS1hBUlZoQLjB2FFO7c/OQB9OixvuIZrUdI8TNKFQhQwjgA
8ekSzg6K2cbZjDIxHUCWlnTcgWDkYUtk2qZxE5R9/XN7OvbZqsrAa9zm9EQkm/gbXKdClW2sZO1o
NfNzrWRwlLcLYeCfRAhLmQJk5RoRvFsBl17INtvFKKC8yknusT45y1e1DeJ13EcjmkHKlA/jEuia
FbIBdwqMtoP5OfgJm40GyB294Ss5/EElwJgfLdJcnN6TjtosoUboGhPZGibj4ncz+VUNu0geORpy
sny5ceI2+XzLrTvtpKYzgrP/wC2BPjzaW1hXvYdXb7crGcvXPBPHny8wOO7moxx+uJd7cm/ic9zR
q/qvZHjv8e6bjv/Zqvwq2sSOYt4uB2i+OUae4wrDvHMJv5zQnplKiYN23YtsCtjbTJqMFf3yBeGB
9Lw613HnnpzaSIkUh00ZcTUzIFDm2ukdeZFbWcjL3HIyGO2blUqaZ+0knGe3Zk9opeNZ6r/OqBPs
DetHGMfDisehHR7h7o8HLAqx1xwxHdmOgqwpOLgaEfue6Q62qVXRnYWdVgmNLkye8fAx97wC9ucP
T1Nms9mEqRUrUWHyzD8PmS+7GVA4ajXy63U7cGf7bvxinrgpRdzAar2Ypd8BMHPc7xLsFneqQOTo
54ls3HWVg8N2cH2abJnx+01VvQfXn+xWvJ17VF/BBnbzySh5wxc2dQldMUMRJPMvfRqMvvQonQMv
yck2WA1vDswAPIUiU5jrYd27mbJNlEsumBPPhLV3amQvxzOZU+KvVyunXFlTfnFioXRRu8DIwTpZ
Tj9kMrTpj9zWjwrAz9qcA0YYpwLXGklOns3/P/UaqVoREJ/1owOfEB09WsHUqm1y4QlaZI3kZ9Lc
S4yhPzhMcxYX+HoXLWphucUdujELi8BaeWZ4gUsvmeub+3ZNsDtM00YaSaGA2RbQ5zKHGXcnkrmD
aICi6smgvZryxeFXBjIdGodqqwkFOFamzr/g5c7maAkL5oOlQfrRsgn+nLlzj8rPlTxTInXY6ENF
/fW377lpbX3QUKg3vqvlmQv5CJXztZGUImO6n28nN0H1FNROKEhKAB2FFc8WRkNn9mf2CmwG4T8H
DpEtiwaMvAHlaeZhssvMAW3dIl5b/pXqvTju/OSpRsEScxZ6aCc43XR20BH6Eyp77KrtQipZmKdJ
E2eqiXqL0qr/0clz6J5gIQXLcHStzqv4ooW2/rpKrIOikeyAKVo8pyK6drJVcb2kjkf2Y71Qw/Pp
JkDyDpKeuJQ8aGdcVCLBkx9vTlTiTk90Umnus+vo0wGYtlvNCbbJMziTntFDjm9fBIfGXX1lksAP
kXn7znwjAHb4QBU0svdKp5FS1ufOPL39kEf/2wWKWQ0SUi0Q0PSg7r8tiueigJAG07FZds0ve93q
i/Jx37wi5VUASm0S2n7lKPyLvIaQ7J7SBSFIU3B+mT5giKFu6gh3XuMzSc7vBS2Fu1d17VPgaPeB
5gbVDRbSUvCLcC2LDgRvvHlXJF6m2B98x1uf4eBtQugx3dyCStorAB7tmNeDqjZ8M4uvfh9ogwow
+GIz9TEtl85Oe6Z/7XvwBVpPxHAEeKOX+zidjtZQfZqFrQPTYEy2bHeZZwx10CSMDVKdHIZnMuTt
vvH0mG2VA7uoSDJWReC6+pXJ+/toDFLSihH/4IB1iwUr80Rtgv8FTWoKZx9PVsy5srhLN4UfudUJ
iUwFkg3F69JSCGAJHX6B5y+A/pQOhfIjyl0pp4T9WhtFRazjBDnSCnX0IfqfLpCVUePkeJiWwvTj
xiI8qvVY7N0aW6/2JJYjhTKs+Jfb2QmHO3RlwuCDYBvcAR5LCeZ3WQHnFctu+ISX4Y1IO+UXTpMo
WiaaQmg36UrreorhDbsiWOin+mnwiPEfbWY2s5Cf2fwSOqeJNeNvRwpa9Z5QO9kqu4eOj2azvCtN
KhIP+zSTVs1D2BdbzcdezhpYVkcvq8DjUgO2dR7n/HZ2d8z1YvClLUovharkFByPPHH6x1A8+SRg
fGLUmXDzO26IOYquW9i4pJiTPg1KGNtTJs1vJEn0fTYeNTJP3OnkWsKl0Pyd3PkhkV2E+GTmsTEY
vfhlx6x2SLXqH4Dda/kV+ONfVgrSU/Dhhlehjie42YuIhRGiC9R9z9nR3oZZBR2M0/JHZmcQK49q
q1HNZs5U+cSYKZSF+0ypmsfllzdN7V52ZhT+diN00P6xsiMBDiPL8Y/6MyOkoTKbS+5DU847EPMa
HA97QjoONSGIX4FWHKk7g1odLHHn1kPmN1Kiu35HAYgTEXn4Bya+7BRUWmP32fO4+F9Ec8VtvGDp
o2mx3c3Xmr9UK93lJJMMBr+KmBCA1qreV31M34htEyNU3PPM/VLF2dzsqiFitbdsJPQPy0Utxx84
VTbNxpDvJuuiyUyriWdpDImcsXN9ZkCNc5pMGy/0LtM2A/PhoKC3EZ4bvrFPd3KNiL6t1uwhmYaz
sRczStIyg87paan3ziYOE0JO0heNYym9lca1tGB8dQyAiJPugzuy0+Vp+RxPZLk9m/siHIO7OSlB
WRTaQZlcUgsZNnYii5SsYlGzVMl4IeS9eO7AXu5pI0CETBpxtZpBb+zOo0YkLtRS72UMYmlcrPoT
7HkuFBvHucT5NbXthUFyyPhOeDXXXmVK+mV7lNOo+aXvpMzW0jKmWtcqXYRlB++eo+QWYAFSKZmx
nEtwARAduAztIyJ3FumgtTED1CHAf7NBOoMnUAM118lHZGEkZC5noHPVRkEqx8d1O6ZMErurhL6H
HC4RSBVTq8FMNzYd7U71F2FBb4z1ygt1vL9L3HL4GTpectogq1Crxsh7O97Kkj/STZOJWHVQaGvx
3xPfGtmwCxcKv8X7+uhR8nUKim7GW+g7NuRHl8i0CMda5hjpVskF0r4zSMaqEAzv6Ow76TXqHiHd
5v9xLUbrDxCa8TsER0sLFb3rFsezfLDvL2y1qgEeL9Ps4/2Aijfmhic+q49FrGUnxlpEMDcWWh/P
GVLw/MckOJ8X8m2ehJVWeTyoRrsp8g3AgfRFnhiZ9CHbURQfvPQr88nx8kKIjO5s+VpLNqA/ix6h
wqVcwLyh3WuEKMbnuNL2lUKhpd5EOblDyEZcSkj+ewk27xUvPoEpD59XgX4tlgMkqq4qNG5O89f8
2udhVZqhuwh8Y5DRZf1Of9UpAAP/hrTDu8QvtTVF8XqD46GuCXlQBeWlibzUndFsE8m1HaIdXRzS
rJGZKX3DNL0oGqAtcULwdHOQIcqO/7JhzXnJervQLmTGYQ6+CZCsM60MnXNQCyWibU948atlQUjl
AQM5e40XrRAPmLRghLZEg5RtMzZCz9qhDKX/i8j2JPiLdHC39J9rRm84cm3e2mEerryk3NffTAMS
abtdefMJdz6Ofi3b448vxZEQ394aTL1LF5JN60GZ04iNfsi412L8IPgrv5Fam1KOTFagSMTwQX/B
3+7WFwdf0VY1VManXJSzfBtKlAGjOhsE5tcs3Ivnftmz0kI66Y25n55I2hJdBfJbt00k3sJbUz+D
ljTynX1ra1WOSWJnCNfnLUcy9JiOG2jJLRr8OTJ6yRzB2xP9b7PLJ5XG5zOwC3ycRnLDhnYdW8gX
extLUZdv7LI8lh22AEuu4JLxfi5CVHMz0eJMDuGfGyuia/rz3JKkaqHuxsYY9ElO954cXX0QHBhM
K7PywfdnIo0ybcMc80E9uPPRJsoXxL9v4Q0Z15Kty/yehaMHXh99esAAEgmKq6YLGO7h293vWGWw
hPpk2axjP4TpU5LP9WNytogbxghd1+71ey/xGcy5VmO+YFpwq6GYu2/+xEuCmid1xM7raMKJczNa
Nd9iRYQgucCn5yc8FSGjO2br6QEHwRSZw7FFaGFasYsbOXByutfIQfcLp509UtITSguxlInkQuMl
jWFUiAeqdsYNIY+q6It4RtBn5QsTtFhLXQavynnqbfwyCXRkRcfVj1Wa8+2ZVUbk8+To44rW9dSZ
hPYjiwvRhH+VrwSU9NoAVYBda5RiHfA6r90S4u0vLgxa8GAbWx7XJgVkG4P8lY9beTGrsm5d+spm
u5bvD/fRj2MbRzo/PSl7nyic6nKyRKfgNQHvWfWHTVuGKWgLeyAPEYUPAYMmHLOed91+VK3T6a1N
2+7n6RZQaDqYVcaxjSVKYBUtgzDgMfVBQOVab1S/59lQdOwYQ9jTIurAA5tsxkO1oxADF1nrNRpE
NtOXvMvCpTC5QoVISlHypsEcaD5nn/B7LyMRaU+V1sFfQvHmGtIoeQaqPMrnVHp1ze47XovH5k8k
++RU727zYWfEkdGlox+53uvsY+eoTqSGs7q2BXDtLEEsxPkGRnX6W84gj1l0YFqMMTgT4l9fd1lB
f27uJ7mOvCgFwiA/1Lgi40f0nmYvmglxaQGmbxBT+VERN8z/FcjIuWSY+uR5pAQgn9iaPMM5KhuG
KVt13U4yQKTWlXNDfFLSkIWsXSyB1WFrvury2MHvgyhB0g/rspPDu/gP+pIOKO4jJ4iK8np4byK2
c/fVSCpIH7ReF3KPNOwvrd7cvDpI1HvkK9jnVbmoWMyrZMT3206WZKbA9Gv4HSBSRaLmH4G4TF+6
udmU373Iax6QgRYOswIkm/FeMVzDMWJTOtcH9MURkRBUpZVkI7HQdukzUh9t36tjCgiyXDvOCGNq
AmMtRn5kcIXuJQRqeNG0q32BpqD8XWLmDJs3ACjuDp5k5XI5n8YRBt03zZh42SjIpFmLiVyFgHji
W2aQmGEmWe4quhEl33S0lh3u8bDCYxSQWJ2PGf01N/1Yt8iUxT+OpSj1Phrb2nKCSro7IkzM1fbE
8GE9TNA6MQoOJECb4po+RozjvicVC7xnlcfBwGJr1PpN6klI+coHBZsmM4CzTCYeUGgGTxKLxtei
FaJwPAhtRUa3bYBALNlEdtZ2tbQzH9v+os6FRoSlLYoiP84ltEBDt38jDdSUO/T1wPvNY4kkNzi+
lMznWfetewAeS1rSHE+SZbgFpZ1Z6AvipPXYAtmKQA2y54+s69O3ftmHXEjCnFHUs1dhIZI5QKpV
P78UyP4ALh8cO/YSxKNYaOJvGfqI3uUfScOBJ39mtD0MkNo3UwchKkEQSd2uCz3tBY5yC1OF+nBN
8DaHW6r4ZawzjXu8Jl1Z+x6yVBSo+CgYDQPX830DDy1DS9B4Un30ZLO0CRuCx//1LrsfUVRDgN2i
QATkM7/AYKIX1LAdKrFxk5WYC5fn2YUvMocCU65mUhdMDI9ZHmUgeFFOBPiCl+2Rp9KmGr2NkTZn
OUqKrW8dvvr58J4tSCCudIyAaILmOt2zEzRCtpkhGRyXOUWHM60GcyDo6gWpEFKKb8jQ8YoMkNpI
1ylHMjjZDr1r8vEJ7S8zwwsWvuLpVJLRwGPH5fs0nZC+8s1wHj1IK0UwEGOYiHEPBTVAwQhceg+4
1PGxO6iO+qEesYI7/lG9QhRUZ6/xk7IvZEq8RGo8kSxq+bf2BW/e+GmXYmxCRvgDFVimRbIAKZ3j
zM0HYSdGUtr3dY6Hufi/FzwH+YvIxgjr2saGcadW5Ab2BEkp6g4FBxy3Fbf2RWZm4YZCKqKxxzW7
T/QyOaQYVz6joAml87FrToDAyXzOFdkn7SLqehZSY87c/GO4hYvrtmNUq0HYjdMm7kk3hUQ1KrCr
JNIBLxR57emLtswjhreLy/XQb5m9+ZhDjFoJyHafZwhn8eUJKh8e0LJ2j8yGxIRp0AaJgbYxCbzz
MBKqdf3j5Is9FBXhwsXItq53A+al92aDtYXmklbdGRJf8Pk3BfSrEocZ4u9fP2qh+hXTvJ04NMpb
hKpNKctkZiB3JyBdQ57onkI5DmHItbYZSzJ29XIPZBj8+H7GWa/vqB2P29PGXudwocS1ZuBsvo93
Lou0kA04QJ/j1oPWZFFFq/vTOiUa/DkyxgUrcbouQpi87Nj46zi6ZQtTlVrjUM8YozidFFDVjwoA
EmwNM4OT8s0kwU8OBnGOKbGLomHywAEEbfEg9SM7NLm161D15SPnAMjpaHip/snswsz67dZTViWx
1dWzRXFeJEm5S9Bngo4TveZ+I7jJMypEM0BzWNWnXV1gfuBXUQgyFyd5imu2VXoW91h+fl0pPGAL
tdYb+bpmXclu/i9t7Zn1qr9rwLhGeK0s8gwc3OWi0GOW1PP0HRJWWGOjFTp+cm+ROebQZFFyUgn7
6SXktv0Sw6ncnjo9R61aSNMiwCDd32iSfYCPylReQKMfWYeeFaJ0B2TCGKdfOQxTnN3lTu9P3wd8
NzKUk3sR59bM0/EPUCzUBj54NvAWnNfhZhmm+yU68ftP0EB98WtavAaEwFv3Snr7Z/zfbQ9qmvxH
Ag9erqNVrJwt7csv5U2r4PvSrGVwbE88aCp9Vq7bvm7oPvDZquKW0kzA6Pks7Kgc9UMot2fQwAko
hz2stjBDkyX51mNrQeGqxAUOQsLHLNDvkCN3lGqSj+d/2nabCjqsbh8I54oI/h9Us0N+JZr+Ixd8
oY2zbBGqJCV0liKOAi7jZ0ffXAyZrZDv29oteYEYXgHk4whOCLeCVbM/DZ0hYN/txGH3g8oOQFAe
72vG6JCzyBOeEbe5FITGtfypMEminrNpkfj43948H93QpuHpFzas7+dQn+AmgiLouRxurbCOKUJg
NFr6pO9WhbL19Vnmys7geCeJJMXkwMx+mqs2xsdUKZ+dH4DvyRk6j93VxcsMG0moPwUnhUp6vIm2
FarlD3jd4scbWIQqdrFNwPCXJ5csLDvryGa/gRHQ8Mi+OSI38ORNGi7bVfycTKxY17yWb5Sn8rgN
M17P23u+EZY9RIxs7MDOG8I59P4PMEA5DAL+tLUa1HoQJFZW9IC1lrirM2x/O6tykj0in9iuQwfO
SRDqx8o4V8KM+C0h+1FmBv5e0PfWbF1m34RLZF+GjSsXnsG+KXxsanqOhBXI3IS/UlNuYobyk1Jw
fN4SFNTLPyjBkhHyXVYUOIsbqM2yDGt6IDD7toch2kR5ZIX4QDudtEBpE9vGUEEtIZY54IvnSEFZ
uV1o6GH577s9d5oTrrOapaKKxPITMYpc82OqTyCpcFVPTTEZUc4zGRkBaETu0AEijbGEYke39Ex4
yDCjA7p7SxFM9uN4oaXo15XN2K6Yp5NL7E5hK619o8ABg2h5Fin0Jr+SL67U4ck7zgIYeDaE4LCQ
mfWZrDViziCUJyG1+zbrqUH+NtMGV9a3CKhOTXnCq4XWMmZq2tIKWPooQhSm2LQn/CfLR+kIzRkx
lD9UCr74U5nsxUcWl7pcFW5Q8pVK34xOOOR+P/ZBip0ebnhxnJIvbs5v0UT+Wt9/ITL6tcsHO5SP
aASpJw+o1GFEUJPnwQyCoHyRc62BRs5hXDT4K0Uv+olepD2Tu2ydXzDy6hBYU/Gi78hlU8zfTCVc
K0ixrxUT7LVnIyWxUbveDD6jg0nz0bZTnq3dzJEPGYe2GAUDvY7AuRAIAUp6MRNV1FlfgILOyGIC
ZCNQPDke5rNQg+Yq8OjyxYcUT+LQiMokDUEI5jjDxFxS7Kn3df0DmUN1EiteU7U1QGS/dwUlPhzO
oF4HUxXHsgfyfwWnHGhYlJMYOpweLsLUnc61200+VsAd1XRegUyKfs2woJvfgq0cVnJbGVOm84Xq
5Yx5fgV7pJLGbN34LNpYoy/jHdSAD/jdfvYMRpKib+1J1arkj9px2o2tgXd433iilLojszeL42/f
8fRREfYUqK4FDyGNnr/R6jxfSo1Pvvah5VY+YY+HFtOeVArGZfBYW4ynB/1VHaot0Pt+s6XTEEUo
nhPvAWYBXROGG1cLTLDa5J4bWogbgO6FTuXNw80i8BeCosJ1ofO6K3skaI+GbBvv30gs7OVFML34
Bd6ZQ9oAGS6y0qOgf7JcsGMWevalKbGOFkf25rintvf4o14Sk8gDAPwQfptHfQfXdIPBFLP//jmb
yM8td5Kkmyn9+nkSaijm8FqD5lPGV+YpclWqC/KAl8fF4qIu0Gz3rhnT+IeTCdZ//2tSjVrVDoYW
MwPqRx/AY/clQnSZLx2xEAob/XcgbrVRsFxlE5tNdi/nzd8SFbnV9iFCPUNLLzXrQddCa/rOyieF
91fxwl97DbHipSc9GJppXOMpL2Q0IVQA3t2+SCpP5NcTTOc7Mpc2QDSQhB6//mUBAUCSIjvQMP6q
OqVw/uDjK2qNOxyfniUajQnDOxq1Hz6tyy8IcBDYZ2Pa6Gyys/fzBGGeQcFlsHelJLsSSXxCGgWm
ExQA5H9EP9DH5LMWWVfge5ikQTe7FXt6ELbMyMqY+jGY4b+xbZoMB1T4lGx7AEq8aZudXCgCj/sO
b43Z4JY+DWFQhg1+icq5d5penrRuMM+avKt/T3Na9kdajdL10x3Hdf3BghblEL7xw/4ef/5grwFp
Y1/St+jyx7UEGbdD9SnLhXS0WtXcaDd+kyFSRtZo93rrY/JPcgQT89M5kDy1mvrrpxiNWRns37OU
CtFvS0qr+xxeEA2PLv/9Oo9edQ9/fUfQZHpW8z9BGDr5NGiRlUuWkyax7nbxpslAR2gBaGE+D7hl
ocqhUW78SpQhjLLOxRzc+xveITScnfjtK36wRVI794WzpoCiVuHzemPB/32BCWXQ1Kz6JBvTsNgo
E6uSJ8MjS5nr9BYJiE9e8KTmjmZgFLh9S5+29r+9rzhpxVH1VMK1jl+BnzXKfeU2qstovbyrglAN
VrjZXqRJ00I6aI5SUzeyANZYCjlq8B3/Ylg3s7YSGlpiDpG0ulmTmNcWRwtr+8CMdvGOZpBMZXZm
59HjfxLOC4dVJqypAjgBISqvL+oLfrrykXiMvRW1BMMgH+8GJZKzt1h2KosRuEyChZvuh4Eq6Tux
A1Mg1CZ6xJPLpt1Z5kMzaSZn2xUEfM/cdC5cxO3YU8koDKClC37VqWBapBKWhkSGGw9ztfejDpyR
PO2Tq3DpU7EGPYHgtoQQwlCj39FZxVrOcPYu+CFmGNR9LGMJc7Ra7P8/vMGLQ0e3kP4ELixcYVuk
/xULck8JF5Rip7SQ6JqfjVBkNx26L6RigtEAhE3atWURjv6BMnYDNSEU38HlJBXVoD0mnX30nOKk
Z1SYjI56tY5ZwVV4iq5UfbpaPqrsYFybYYNu/SRd4FgEQPALR5zQGP/YA8bVLZiQma9tavXC/iEJ
l6upf1afgTaMKDFdjejFVbPxZmMq9B2n4kmq1dOMyjVmK1mtpE9qYZqfxzCF4D2pGPlWUOu4dZD1
1FnIFaIYRnH+cdvHGf38diyeAlaYMzEibCkBL/Aaq6SJ/oQ5iTjaMiFW5217pb+jvJ043rcS5iTa
rAoL6B8OhanIAT30ikl+gNZ4QRwh51dSiiI6mpvtnxpYn92HEPxcTZUYUKbNxllS/H9slU6D28Zp
OD+ztLwXZrE/58aszjJcfKYmAUlvyMUVLuEsDrNHZNzM7JO7Tr3G1TGDMYw+7rU0YAr2M2+q5dCl
PYNtR7e3YyrpU3ZpFh6VY9N8ipNeqLa1G211vKQjOMk8EZ34xcPBuEPdpfuBihHgKwRuN1//4jvK
gLAU1ygfO6S4bFZL46yJpyqTPaijZr6vMbA3SZzf4+w10Ug69CTpDBwGIuPu8KRfQTLBlMQVaDse
EmpENE2M6XX4PRAP2Epgx8Tz6RUzu/3WAfzYCU9jsHQS8V4FrDIbU0rP5zGuGFCv48grWb5Sw8Ge
1hKnt2eMwzI9rqLKQn65ua60dBG8hjD3ZEaPTxzSeUBWRS199feFw8vYQxWooPoMr9CQwKjiIKkc
7UhpfL4L4JGlz8Of1qRn7PomLXJfxs6DJByFPWvAxJH7IrV7NaLq8gOhibBumaTAxeuE3vu2tinl
Ue55gL8QTDDyL0ug+p1z5GcVDSfLLdKJNxIcC/bBciPBcdeABc+a02TMnwEjgmkaHZglhud56AfP
C9rUh1eYyrEi+z8etvb1Cgy4m9BRTkSClfgzKIOV98cFpFqFQ+brQYeaRDUBKxZsTlfgCCzE5p2j
G317KSFzxR9KzP+Kru5xYTdUiYYSRkmXYD/U+TOnmAOqnOogXMYjdVPLIEHb708Yur8WIxQMzCcK
EqXJ8jMdqIsM6fr96qP3cECPiqC4QqLv459w44IPUqEFg8IIVAoXGghCdZTnTRXDT05i25YW7XyJ
QlZ4cmy+sCMzh3RWi1EKI/3HyNnk89Oh3nS9bf16874wjvI9EVjgEozG8J3LffI+1eFRtUbbfSr9
tNDJZ802Q9fVmqaA+uvwjGo05XFM+ebVnoA+/Vvxqrgcmuu80/2D9fjgbwxOgJCHrS6f1y79IYJX
K253L5aXyGM2ZK9qZmB+CDtS0vJCLyD7Oya9W5mfCoByB/i3THHNccn6aiNOY/TEgAkPqKeHbjWG
LkwpcGCg80kmjBXFXEBQOuMEYJtA5IJlJSh5Chxkm5PR/A68Bdl4D/JcnBmlUfaE3Kck5ek/nXL6
JBjr2mlmfmOu+MABK/2G3XxjuVHD0iM4nBXKbL+tkfy5JaXb+G3A0XSWpO9RdDt3MhQJGrvv6pY4
EMvUAV37eqe3Wmk7eviUX1pGDY9BtpLHQeeTqEHAgm26T0tNTKmYUF2jzSlolTRuD2M1zpoQFf8V
z1teJ4PuOF5BRAI8fcZd5ghM+KkMMnmtvAL8uiGaAFLGQDQDecfWagxSK44DAxgKE07/YFG9yNmP
92rF2vtYi4T/Naz81G6CIpcGdO3tTr9Dd+DjBcuA0QU3xCrcm/TnkleKoMR9EiwfYtiTNB/7Hpj4
HnlmAKaB0VkkUgXYyT06UyN+NV7NnXafujJF9KDPks6Pf5bKKoEaGfd3A0XzNZSHkiXw5o75H3ar
mE5tQbNfvnXwFaLgCgVqZesw/nFO5rTDaCtPrSynalg+8h0F9Gv8Q260jjUgu2jadQUEH8+VBzZi
HV5butzjwgAy5RfVQJKGV10zB7KhOp4DmJcaiZKC+yAcV5CAJl4VVfDrwNnHEPziyvwyPdnUfG/r
aC8FWzkUh9Q5mltnM9kuwYGj9PMkhJZuBXWPAcswNXi5la+5S2UHxvOGle6Z8eyLO9mEDehMyNXe
BbGT9OhF8gLHjam+s2rHOfjVUanRm0GeJ1mwbQ08EwXLByb7UhWFGpONj5YYIeV32YOVno9Z3eHx
K2pJ+yhCBHeADaQnSoUdDbDVNLA9zymbl8V3erDyefN/gde27d059pyNjGY2TnTs2XGXhOBKgaaw
nBU3iipSxFeA9TMdY0TM7gYqdvSMwBA+WKHUJrDyMDf+LoyVMAv1jhx6aFr/8zKAEPHNl4dO/SDJ
TSpti85PIAdNl3IY5jcGW1EqQStrDoTyfDaTC/1rJSnqWixpcsgrqdZxOAvC/FQGgbsFRCl1hrO/
e8X7/uoWmS+hGgktGI9G7/dVwNcdSIkRVm3wbQySMfzBuRIoHvtD2WQHwb4r3H1eSHNajvzuwGKT
uMGeGERLTlT8B3wbUw3SqHGOJN+wE+Z/TOWO9zaMbrm9tqpmuS8RaiSFBAh8X0mnGn7MtMuoEHMU
tuah7exRoRC740jzfgTY6pm3FOBG68epiqLew2GfBcvqs16lBNSwTu5DiDifCUCpyVksc+RYOMfl
TKc9i5HN+6bptmJa6DqGGY/xcbF/wEIj4tv9/iddQ46FXEyGepro/36XoiuZWOVNnE0G4HnsJT5x
UVKFOtWs2+wummILeVho41w/ciboaO2NIZAoTixetB9r1JySblrdnAW8jDhNUQpAmDxG2o+DhsSk
ILZe2NaeBNBoh85etnGl7yW9c0Jg0g2AwkILVF7AxpRfD/kqV4UH/4WjNiPgTQ8aHMm640ThIiqg
2PKNspfz0xHjz7CstMUDV6/32Lh0s3DUjbp0b6HxzVw/WUbcwfWS810nBaDqyEEOaFoNkogjtYnu
S9VMbAy7fEZ0cLJU/BabDkZOgSEO8cVJ3nhNm4MzsSXHM62aJw7uREA3m5NiwOpvlIUn4gEp5BiH
SyVhmg8aVPBTdDkFOTzcICvNRq/qy4mj228X6Hruqj8O0ktHqwsLymO2U+Y77U9akCGJx9HIcpdx
0bwbhQGlLwpjl/Xz4S2A8+u5sxCJdP1HI4slrkEBzacNWEhXD8IhsmsQq9RMVjgMnht4dyA369PY
hA4TMmIMnPOjySkiSJTaN45jHDj2x+3heyf6xfMmUE50/4w4zZEauoAHTecIvZxJ07hwLPkvyaBY
DfpU4gSmQPLmwg5/zgexy49dK68yXUnFAEuWrxSpog8nUAb3RYWvVXjLYgLHQ8t2W2g6QLCtWdjC
0NJpiNnB5GOh4URVEaTNW5jIPMKFRCMrlp+pW8vP9h49eFVyyDsYt8ZWJgxAPODXllgXMsHIFBps
OKYQ+vIJFss/6xT+0CA/tYf730bA+H39EFZmT/h685QufwL/7HWyM90vP0sAli/OdH4KrI0eOhTy
IUjPsyCIR5/OiZz5T/3fj0bYYmidXDwrM5sRjW9FAm73TJ+ZNnfefrGKpAaTjSjEcnUEwqL3Ly4K
obpbmCeBW3cGRI7k5v2k9EY71+q72IIKmuf+/mkUFZBf5vyFG33rIn1vnv8MbtA4HURv5pbwCG0I
AG3Q+P4v+stwsINNsRis1lOrrPXEBubXV428ktIjRFNGBoHhro/0SjhcOK8PgOAeiaEFAoXGcRs6
7jglol3G8FYmepgGzqTunP0Mvo5OaNYLvdlcLKsrBmMGWX36lIe7azDFVNmA1Uun14DQPI30bujm
zVdVrCgrZEAdxhcL61S6ZP+7FirKIUAoM+n41jw7I+iMu0Zk3B3QdcPEa5a9HbQJxXVWWmTRSLEu
nNiMrxfIq7vweudpbCFf0sIcq6A7MtefXLMH8TAbBaq9gLxWWPx+J54SNWzQxW7rKjkTrXx8Oqif
z/fIyYIKLO/Iiw+hkRTvMqzEHtpU0se+tNgTQJs0aiR1rNIK2xw83B2zVF1+Q2yZObJMH5qzzR50
sbA1tN7tejL2Wb2hkgLuGp+GNY5oAXkHL6T8Ev0/oL5VPXKfo7nFkJHI0l/ZO6hvVppTYBx1FYR3
sHdpLcqMu1iTOZJ3d9G44RXiXC5gKSDzNiW2Mvl5I9i1WawybFZsHlkg5DUWSLlGfqXJPyCTW3I8
YkVpmPKleNxw3X1aSil1Olq+gcwUaIV3F6FL/4odf/qWrsQgfMsObIIf9g3pjrwbfOL754tNKtP0
5kw4OUoxVF2zF+i5ZNHT7saQ/mtZ8AJb7MIYTaom9hmEHdmBWSjVb+IBP6Sg9uLbAvP/OEIEsQyw
emmjWpLqLLkfNA4KXF1SeFx0BYrIFMxC8x4LIkhpsVpLtyBmkfJfnKdGuqZkJETWMdDshUHNp2VM
MHHj6DMRalD5ZScikE0fj8ZufRtxLd//nYGgx0RLERIAeMELakUvjmkYesAzz4XRhpR1qn6eMgq8
ISqqQYHxMrS2WVBRYzBWI9AK9HwfM8R2xCDzXVOjeY0cu2uNIYmn2HsyXXXbNRDrek2w2xoKRKsW
XEMI/pRafOhrdYQuShCkqmvsSgLTcbRTEcMn4lGSxiQHRdJ8d7XUiFE1JEN9oVgWdz58CZh7hjDu
pgG2vnKyNx8p/FcF5UjHN3r0rewMAl2oeDuZ3vuU/BvPA5ues+seWdcsnD0aNll6wNR0KaTmmJyP
0Rm2L1F1mFmQODJiZ4qZkBDzs438JIXZE4hi1sUuXjn6vuo4oGFNN7DODfvfgq5serfhUiEiESId
9tbUeHrKOUMv+lsrMlPaY4BQFe7KpU5z3Zspk/uute44s+63HoFTXb4BDAEPDDJZrw76rVti42zl
ITCGdNdixrRVk7qzyABtdaFSUMXNKsqTs2alr/oY/eH2d+1kiBDEbI8qHVfAk/a+iv/Z7iQY+i7C
033Qbd/iPgFJ7NZOBtjxXlXGGlQ1fZhC+UOYPGV9ilmXEqbFHQNlWN85Eye8d1PLmXkzGJfSk0Qs
tIHo7HdqjtxMwD6OxU/qmIeQbr0pz2hG1bDuAyWPnnR4+nivwYepVd6zZ7XrdRkOXASvbq8AOOR8
dblSk2bw8g4khYYVMK6KWF4W2v72/RistE/sSi3HFM/yqg3M7RWa3QX+dxk+s5NYiiGqqiOUXiqg
emaQnexmh077NUej5R5MuW+POEc7f57C60h+rnCBiJEHJ++mZlhzxMY8oHpI6MJpoHn2ck2Kc55L
1mPt3VjE689ZojPlqGWPf1tey9jgil/AHmoGWS9BPbMXsZ6MTc114gKp9g615/jr5xhOgTmWfd4x
Ir43ca97wubAywufAkwNBxoPBy6abQ0FocVeoJ/Xxi+uJglwje8yCxorBit+DxOBRek8BThnYY8b
JBTjh0y67vDwPEwckAJGxCZJrj9J9SSBQHJfWstHMQRb5nDF+Um6+5pyGyL43N5b5SUyMLQwiKKP
sw3GBKmTpOfu/hArvFIA8bejOJnpZ54RxvO9LPHp+ByKggljrxtIn5ARYI4nEYQGMkOzatJ7qtDn
QFehJ5zL4hrjfYzngn8O7qwQIn/pRH6yI/1HUGR9HPxQqUQeDukNR4cGI83lNX4I9u/ATwgfSu1N
3mn5ckFWcf51Jyi5YQxnQOhy8f1FNnNyWjmFYglFlOWgkAe4w/pBnfvsGDQ7nqstekoOLo50aEq+
lpCpYshXzsdsB7qYxOGRecj1Ze0g2T7TTayOLi1oyrpHqJwilL96Rhn/xYVhSr7F7enQ6gpoBUwx
ucVbth0J/1DF8ynWAuO5z5aL49+AyXBgN2M8CWc1U0KfASBongsSHilsD62RzudGBVXbW3REjwBk
x12nyO4WNi1wYTRYco6z/wUNcE2Ub+RUbfPXsuE5jiJse9fJd9Uni5GiWg8zRcSgB1v8IRdXD1lf
ttMBEcLVgZ4LB25WJkkDRkBxaxaR01H06uDlNh3T9sljv6Gj6tgxP58vpVvZIFpJqRvgbAr6wIlh
IOuUL6DMvYF0vIstlHbIC+GXu8RaPYde463K9+JyiQJYDP22i4aSdlg34huehCmaRLVth7iEjTea
vJuXYtt7mNmQ/EmQmITOAIYrDQS231invOmpne0/km+NI76p9xgmI1CN+B4SODDYffL7JTGLU8PH
zWJhH/fYrfoDWGyqEOhJW1/tymcIhj5kQAOV797iOrNjRBxxcmHhtjFi0hs3/7Wa5jeYgxVlsMCq
zT2ZxI6svTXnywiz5eJLrtlmZRuoWbOo//AxAIFbruVfRdnj2ru5GzZCay2ISLlyJrOaEZa9ECCz
lpTLtn3joxjIixJ3UMG8SV+Gbh1qond5VLFDtBxocYVhNMFpaOQh3x7Xost0EUp5OAJUO9Nn41qn
tsxI5zAs0cb4N4N+TXKZHWpYEtK02eDnflHJO43f8G36cQtktXzQUGbZcTKKy3xl5a5egfmn1Uxg
jPua88oVvs2p4XPevN/cWzYHiAj/scZ6UKq83pGhTStjmXQ96Nd+SzN+lCMh60RgKf1JtMzWyw8U
f7WYvvBVlIr71uSyFJIvtmkRkTWrGwEO3BaMcPKWIrJqlL/EVEHuGmOh3hpN1RVK1tVW52sbBhR7
lHra3CYZMM515Ct2TubL0i1NX2zhSgyRWG6c8JRtrNDZ3O0nk316+Rm9aXXFCd54tQ6sUbmZFqiK
N6iFX1pse7/TfPprn2IuFpIFkHRneS4jqAJsk2UVgY5G0geEnZXQAFYXvkC8X/rI6BWBvi/7gc+H
J+/ZDgjnZuAj8euWWZlS39ZbVqh929l197Bq3bfId0kgge180nteQBmptNfjcyQv5TkgrhqM3m42
cKElBBJhvgtTZKRjxlTvZckhgTCEnW+yEZLlhBZecU7poBv5GzOCGWGPDPYBWo9a4WA2ONsBDewl
orCH4/StGnbytLHixPy2pZk4kZIbOdHQxWjeWVPa3X30Oc847MkoOK40bt9tw457ZYmi7GYB4Z01
++npl5hd6rkvPJaokgWVFQ1vHRUP+cZ2Y6eYpj+sPSkXLzQEPcVuXW9pKAzd42Spt6LXGI329FWK
xvEqUgbGlrJIvQpRGR4EEMUTt3wRoy39PSLd262LF/moLPFBR8IrjkvXXV/mllQLC/dRdE/kSjgs
h1BZdEadN9kIz2wTTBPCTWnThoiQY0VVS/38ECgX2fesbiU5Jtp0a1bq4df2CfqGV7ixFQl2Y75U
P5n13xIeDb7OrbAAusQ5YtQw7og4U5hKjOnezgBTrGEZaxBiPRdkIqDN5S2EFAJxI+ObAAv96kbo
+kmzL+E8xzIIn0/gbY/gMQJk06qv72pcGdTMbQI3pnftC0uzUGrrcjIm9eqT+2zYzOoTy/wsF8kR
1H3eR417JzBNRATUi7zPphqS8eKbf5TeEge2/wQFyIP3NOanE4aIRQruiM7ITG6rlaI+Ejpll9ct
CZEJfYtkLdeR8gb/CiM/YXHwQqM5aJvnHPy7Ix4ZmwFD+iKuOL7X3tPjhSmNtTIh7B8qzmRgNRNI
nn+FOmWsmO9x2ifqorPvUjpDvmghKzXn2q00B9W40gsv8yGGEWs9LxFvMcGRENwvGTXBTVpvL1vP
qHM8ezR3bpWq+cHpDvePNv0vp2DjuwGF9l19+WJ9xvSVyQ/R33sJT2XcLLKbXUQQ/NgTZ7vWiXgo
rI/tHUKRStOPS6iwigm/0qIQLg4l+qn+sOBbpLdtR2j+IfL6iGt3ZUjjbgEWKShLrDzmNvr07VlO
hVjv4Y7Tc7Xw++9YAw6mF8ztMienbewNSgBoMvrblH6ABX2fCA9tpwJOt+PgtuKw+a1uhqB+D4mk
rr9viC912YiMbq7y+r4mbGEIFmizurI3UkrTYEPZ6ioHrNOj/roZeu8cxfwcHeKNwQEcZhyXxoAP
a0A8ULBhhqNAH+n5DTxRYcC0txoaoAKfJr1kJ9RL91KGi6XNC9+Bp2P5Dgug6vdbnZHLZonSagsI
3IWoKhu9gmTMZolpQ5UYneinDCMbuhJK25hmrBCunaG1ZaCaD44hFiqZ9a61hIBPumBaI3TdHGcP
RzWvojgOxdtJkGCYXZNsLdLHWPrFtCafg9751Bkf1Ln3U9WQ/8IXbbSn/DEB89JE9wx8Lgh7BAWL
r03SC4HG0rPrGNa+gHDn10v4KKXEOrkRFmHTuzdUySYFX7iRcBqwixafXkpNVH3DMn8CX7i7CJzn
AHHfwFEHm5XVrPZj5GRyBG9iseJNRBckLiOwAUiqWOxmfGLqeyDfYS6zjYA8fX4L9oR2nVEM60+q
H45DoTIBvna/L8pDRr5MS2nCyCPdkcOD2M04A+kNyuZFAP6n4MbIt1brKpR0V7hUgmAigc/4JQIX
pcXMG4AIvCkNdK6ZPVcuUbJ874BPbs8HBmJDkQLRc8orRVLCvNH1qnu11NeoJaTE+wrltk7BUd5C
29/AaqRakZbLItaUgHW0YGCTRsPa59GvX7VBx4/SxhLOFyJtZDse5dtlhUvqQYlJPI721eZ8b0ZX
NBTDcLr9PzWbNQ5kgP7CffsuHElSfgKUA1AasOOZ4nm8noB7w/cYpOHN/my0aFRNMjtwHbMvo73h
pZR092YvGdVuSEZN4txU8Ic+SaqXJWn9FR9neNKpyCozvT0rBOvaqZmcwwo1x+Ok41KYx3uT7OKf
bYkyBlnR9tdQhWm2zd400KbxoKu0s2/8y4zPZH3Pw9PSiOpPUDwtJ1Lap2PwpJBfLTW+W8XnSFtf
9N/5jdZLG/XBCbTnGS2pulnKkfw8TMjKbX3FkrEOiKkzFFp1RD2gn8erFybcRPV3ItHlrOF+f5j2
w8HB/o4N2DpUbSGvEP5NzbTCg8fUeA7ayEvxU64KX9YJ3Ja1kOrEYx4DlaeP6yhSJkGxHB+JYBIl
S2ocgu6C1pqJNXFSCVcyyLy3PLG0nw0z8W4eOmfGtfdoCP0w6VscvuptQvUWGlinwzPXi74LC/Hj
UafurH8DS9paGmZZNYTskL4eamR7jRsQhEqE5isG/RNmsQFNKLAeYQ94huUVbpIzUhs6I+czbJyr
EIJjlh+AFeUgUDZp2m+hqSScevkhXrDDKrtxblQTWFllCNL0JIBvzGE3Ojvo121UXhINNLRe0xp4
3raq6Xv2nPxGvSjKj/XAg0ZopiFqQzPenGUu/8j8VGiaRWKPwOczCYMUh15hoPFCpzQ8XLbnaUPV
C2GynjdXAdN+sYHhUSFjV1GONV72bdrftGk0e5TJ4f+v/Og0Fy70Yc4DMVKEDXSr/D9JI10/bv3X
x/hTQsTRi4RdMsrZL14UN6DZMyKUJCVV0RYWpGw2mnm9PDTF416Hs2rWUeJueFHyPTBuRlqCdJnc
XAdBNmjZir0YPYJyys1LxseDMi5tuKaRKT2GG2+CtZDV77vdCqGIBt8fBQWPnf68LEgtHiootWiG
z/Sz27mOCT4zW2+ce8WNRxTGRzOivkSbDJ6oU9cIuwi8dhKUWEY0ER5hbU8IElhuPEmKJaJ4V69L
PgPncJiwGN99MfCQ7KXz/ERI/0uYswDvYYB86/mSqAm5Bz02DEvQ7OVTD4z8tHuoeFOJh2hwsPjN
BryB5pzWQCAc+NbqvoTjoG7+EySqOnclhJgIeBmDYm0L4ykoJrb3nzeVBuQ/884+dv9pHBz6Gf5i
uQ63xWcFNG+z8LHeP0Q7KqpCXuFW6BnRRM1UTkFAfiuU31lD9xmzef/lW1ARGWIHOx4wkv8wQ7N8
yxfPVwx0YPUFWygSfIJoBABH034HEo2SyrVETnPXh0uP9F76gWBKSYrsoFSpbwcVsYFjcv/A7q0V
g/kEt/lgjVfNzmYIK38AbZFPuZJhQpOF22A0ihHJzwpEu33h1NznMtarckLft13PU/NXYyyZX5iq
T94P6S2XILpeizT/KUG5AfHsNo7C2/H6+MBlwYFa5/kyfVdgC+dED0AH76cZaHlN1cBohY/6EtMk
4Y0jygJz7hRcIrNeVHRhXvTrxZihn8IRiedSpE/7gYjgyqXi0LEmzsIyyAmrvwKoQiI/S8IJrZW7
Jn29G+DdqCViG4LT+QoyJw9jHcFRbnLnnYs3hItqsIBRmBnxBHSnbzQej+dobgZoAPpVK45SE6gQ
dkP8vnhD1/zB05mEEm3JaxuMVIC1hyzOs59YmxRXXu3MnS368fjbt0Q3ow49C2JInwyIDIQY4NVZ
CiobJtLdlBeOaG/OQFEDD7Bcg3j5wj6/w1uNEcIXEKvnQromLzlbYXtv/YCOdP8E/U2FZPY2o3+w
pjxcNzpYA9PZcuGIQVn1tgvMy7tdkEF5RyQsG9/chSJYs5IejNtHlXGMWqczeiNMQbSkHiKZPwKr
hk5ClttAxtklR5oMk4IzUaupn+ZDwX8Ji1QeRieJ7gFTCD5+Fj33j+79eNX0IGCJvIIbHmpN4DY0
yvyzRvylaflc66w2DFaPi/20I7bRM63OGlQDvNi5IyedtCQSBOt01SxdEh0bEJh8LTgQbI29a/Y6
/6xmFcDhgGFVJ3ALNIMxqW92XEq10WbpDo6O4HoX/Xpr8M5MW5iaQVC7DQain7keAjMX17Grvf7Q
I7fvlCqtBnO3fEoO1Cd8SH8+rGs+NHLX4z8b4BXLtYvW57BSZoHTX5NkNUh2EIVx8Dvocu/4XPwe
n/PCItDP2x8gDLAjU8FisLbstot16nuzYfZzm5GioTsrDu/DcF+qMyhRr7CVJVIuRUNuB986kBQh
cWuaElh4l5SfsVWi7VjPJEeMgxWNEcnKGVwOCkV9kodCbyEMpLUeiRDUdYO3drlT3pPa2nkKlg8P
v+LrvfGJQrctUG91yZhSdDOqvGOoGWLahYSflcSZ8zj2kFOoxsujMP6E/EoHTPua17VhGOlR2IgK
Oz0rzAuHXQKbAVuQGMSlNNsXAN5JVAdMgcsjGoTCDvm+sbwY8e+VeK8jLstmS0L1YtRQiLF0GMkk
vJEWL7iphOd1LXmflSuAc9Kw1Ctjj08U2ThEuORqfFl+nbotK/3DL4MQfZ6k0r5gwqlt3zGdKzBy
s3aW2f+Dfpq9i0EykGl5wM8SQPc9vTBZJA9+zRo/nyL5llLa8cadkKK3qO/AzBE437yLwGQw288h
cHjjyEazlJCQvSNHLYo9Z4h2/ecb/hnthj6+h54uakq+/EthkVZRHwBwRGIV5XLLUVV/EKMORpYk
75KfOJumIEthSaoaMV56A9mqYo2pJY8f6Lje75Et7va/+Thnm3+1Fj6Ex4BhF5Shp9jI1ndbj/dB
XyPUOQfjQgskSSrTdsl8w1ZFAwNTQln9faioFEunh8H2Z77yEPog0qu1i/L0eoLAoJQinGv59nYt
sMfIItTJG5XVKACgHfhi82yyYMQlMWkX6cFOcCPE8VJC39LJfIG8NrNCh8uPrN5lyYzm5OYM4FVv
tbLqjux14sQg8u7bD27Xza731dQ3eCew5J7tZZNkZc8WBSfge3XiG6QbftiDR4QbMhjtfVTafzRI
aNN5bveJCIlTYZNu+J994rcM6zIpv0+OkmviPNbZCY60VH6Xgyqq0WLC9hfzGnzAJBjirGIhVv7X
lJAU7E3C0uhYC3FpdCyiJekIY5gru60bSSOQ/5pAUp0SC0+MOA6xs2ViWyG9olGVSz92/I7k1Eab
MWfM8ob28jxa9TAXwKdvFB+mC+XyNa80/827sekph3a8zo5v86fp0jR9s7ZT0y4MNS8GVULP5I9Q
vBuvSIQ0UmNMORsuhG/YL7rdY9oR47vZw6qAy6BQqmoh0hPQ2P2BaL6eQJlz4rwIjfNq3Vy+96dg
Gdj6ldpgosy9X0ArcM0OCdjVhr5QxYW17wO8yzcp+TRYKhaKCC760CDSxBuBP/J7ePknmABoj5xg
xFRrclzIF2OdWTCAUymqujrGvLl5Oy4vPCkkK0GDESWUlSemMC/7Pyd3t7TCsdix0SentDYVPLmn
KOxp2TVYsL85ykj30R4aZTHeFnKmPaLorJLWDsChUDFaE+OJ9SlzFqaCkZXl4vuraZni2lAG2l8+
95abnOoriT3yx3JkCs1lWGOvBJUeJX/uiMddNL64EFPQuS/grPo31X8cTxz6ZErVlOA9bebhfSLP
+AUbny1HDKJQqeoQGx5eUerbJP90GCLoO7By/30b6Hml57J//AJ7GKLz6og/+90flk2/cVdVkhHv
zfQ2bSMcZAs3Bd/NdZKdyhaA9+fxdz3Rh+NzvHI8Tn9/MenQhkDLzCrJXAR/oHBrpBFbpsW5YOEb
kBAzV+tEuAjNhqUQ6rKj2yoySG6chB+0YaaI8VGTa/ia0koG1TfDyR4NqdvbKKhUyJKkLDCowUpN
aZUbnkYpFLtUsKXOBzbNxTR8xNNBmdSWp9Ifq1mK/WlOO7/Eq3MmOh3AH+hQ2SrDSjPRl7sidHtY
mxsp/KPoQ+Xn9+5MXsXs62thDfW+i4sk5QCrSJuHFA2kp4Y+KSOXE7nsGph9RtmB9YweiqJX5o20
odN4HpuoK/OIGtuAN4XzuvgwKhwasfg0Qd8THT4+Qt20HFOepqWbJABkH96nExfDhy37PZVlGknN
b5SYdxCW/+CJghub2OdOXNYNB/H5IeQkHgGIbQWyzspQMyGn3NRm9YChZXTaj+PjE/Srn//hhAjd
nq6CnZ3zkaAjJKyNMxnclzyHDz27BUp4T8HWpvBFbXpVtNaldyS7aEzhNrjQyROej3TnJhX76Oqi
LB7cVU8Ux1Fr/9qGnG3h3PhOAGNhSKEw1ZdnNoUDaS/eyRk6Gy/MqlcdmQsgMlY/cyE/V7qke4QO
fN5OyOoDWWE5ksydXTR+9MEPan+GbYc3dDfFuekWCRcBCZ22LZ8yrXr/5Cboo9WFSk0u4OaVyXjM
hNoI7jugSRqllOw5HyuWFcG061J3Kw/Q8hNzkXjQZoCTY5kA0isk8JprfRT7ekkTLFVSNVkfPG+4
65YPkfhxJwMxROoKdbrbfAQVovYoFiGocdra3Ex3T2TUyCboZiyzc6DOgnTI08Uh824Kb3jjVa5t
oYelQ8zGRc2IgH/4Z+VMzOg/RuPpEiGwbKw0pQVcslVu2b+DNhQQkanNBaW4p/r2bbOPIz29P4pE
rEyh7vvo504uui5KDc4ztf6KRB9jrVbgVFnqDiCcZ3hSbSwbt2ZOKgdN0O9pxiRYeLVdNexYhfv9
rujh+oOSWOR7C3QxaNUBqfYoaKlS0znNuZJrKZXx1DyWRSxjJtdMeCEW/QUPlnnJTRefpWos/L1r
fqU7pKJbOPpOLAdmpd6zU6Ud13XF6GdtHjvzlryWSkhYShEpFsrsFeZZEvQ7WMHLAYBUO/ZGuGpM
5Vb+etYQ/CM3nzVIWYzvPEtdqg1DSc7Ttql305taV4wLPej5AybQAP+8bad3LDCvNBF7RiTztGuu
kb1WjHePswMp8QlSdaNPDP3VoSCuAL6fjfqvyyHvlvvnSWsee7MaxO5rfACbxsobGSE96SQxjaaF
ZSxXPFHp3XmiWlZun8u7r+Q/Ekq5n/iTvsUL9yPObMOgGvtG8/i5j1IN+SuxjYEuE9kT4ajNgbXO
woPWOceCKh71i7kW6UlYuRGNTMwjMGS50cTkCd+evc5zfx3K/EkRFxjiu6/RY7bQpR9NQONh16ET
fE8IqhsAaxTdz6HvlzN5dqLsnpKh+VSxi+MWvWYO54WsjQBsHUxd40F7GNmVS2byNTjUturpsDT1
KCWLYgdlIGgLxWtgfCJkSK3da7k+53gZywgEFrpdd/SI4w0ZG8oJLF/uNm1q1RQ1u3oWC6gNw2a9
uliOrXMRNKlbs7AvvpSinm7tcQo84qpXyuzSWJQPEH2YiRq0RKc3yuAX5cQGkkG/FPxoZXy4tmsw
nLcIDZbm0ro8+dL/9mf7vJ+wB433ejEsJQhEuMAqxekhK9E3ZptpVAif9hjIxw44CKAY0SldAowo
a+eg8hAegtWkTNFawPLOrUO3KLyx9c/0reE2Kebx7qHaOrxjZBm4Fgh0WtxupLUb+tOE0fj8Wf0d
z9HhL+Y1/46Z7/uidTCcfGA89+1OAADcXm4uK2e+KjL6WWFywpueiHPpPluicFHFJwGzagsKTXwa
L+/OvYgAp4jRIS+twb2GbDs7EYEmrRa7Aej4MiVri7ShGCGcMF/WfyTYthHgUY04+oXLOgqB9bnK
l0BUdJEOZJLWXBlzSQO49Ei1a3G0MAhdgZEBxIzp5ZeH/jRlWs1Yjo7FLehdlW7d8KpmUOCUon8v
BZE0d3h0M6AW7L8XommMm74Pc5gOK6k7lKWq+duVt7BZgwzEbCD82muAWLA15hTyOMqQWvmjFbKw
rkkgFjb39FQoqFuv1dayWI7XSpRw2FbBY73qc804HkBNQJwYTpmgpmkEL+2/1hCz3vTp8m5a/IAv
FM4P8IrvyATW1xx+EH75JTmvAAFsEuhKIU7vunqMIgPuq3c1gyJ+Tpds3LyXUrQg2byCZNaHMffr
NXq2LCcDQlhFeae+uXTsuC74nH+YuMroEsawctM6dz6EvCFJVEge8EUgHzKlcd3xaPRptbTd+xPd
VIlgsOixn1caworILmmAvOevkByQgfpClpvgQLtIZFed9XXR4yAm3N72xvu0fWaP2kv4XXRMGYp9
tMpZKjrBIiC/L6ww7xHtLABY/Fj3VNhnkJNWOE/rtbZlJKsuv4BFU4Eh0a64wQ/hkONVTYwjUQo/
0mgLrqVt9LbiRqkDzR6SkOh+R73+YNNNa9HYKTQ2I42SKznIliI5g45Il7CPZSuHqINSRxispLJg
3aUh9yLUDP2Mxlu9ghdqamm7uO3RmIB7E+J/KzxCsVdV+SiFc+nhbbl5yqIsGOP1p7bhXc6ZX3gr
ArHhTPXEWLYFbz2bksjsi7KNi5YehQL6wd83z8oezTOO8ZJT/ZbSGAo6mHUuQKgoczwt6F2+hItN
clEZGrLIv/7dEUKkikvLXatkY74brpF7E9LH+QmIL3/wZK5ezsfYBm2TYng/zEXdVIYeOEtJn/9W
vddMh4fxJEDmHBLa3jTicfNDQ2z79bnSnEX+qqSQLJp4c/sL1LjMKSdIe8CkparogWLTtyWtctGO
Ay9urfUyMURFCqxRfb6r6B7xzI05n/A5pDksbm5oUiyLtPLhGBnBrWJAM2ABz25P2T1GceRHvb+7
NSUsvM1jIGGYLUmcVRYlUi4bjhtoUBirH7PLW4oyRV9wXfOMn8DlSNliYnM4dp/leIDm0YFV6v27
Vk1AIURUapOj/yfRjEPef3xtUMLSFXOIDP0R64oEgaSvr+XWZoXmnuAoqxJLu656FJqHa7A70hpv
1PMEtKly+BFr7p/l3jgK4azVq9wKTJiUaI5XRAAdaqlLEjkBqgK2TFRTv7YYVbAlyEuSH/rSLFO6
/TfyaNHmaqq0YpJKbHFR+3Vg95NleV/1B3hJyLetOpePAsnh32QoAa9EpPr5/mzkcvx7XuG7FElI
f+nL9rovXWpwaUHPqo7J0ivK0LDhrSsxjSQ1qgAp1Of+h4H/F3bK+A18PlOaiskBXlo+KQ8IV8K0
KcThFUEGEPLcNTNO7AFZG5e/rgwjcoUXMIiqEPg8G5gbv/AnncW9HvA2k27DPeb0OO9+UqzBdTUI
AaTJwl7/bYuHozOPV+EPchDGBSwvO6Ztt+SWHHQnn5yZDWytuZA/xflhmthohwpMrsuSwQjxi4tZ
NgevvxzNzgS/JI3pKeyncurtaycWU+rS29Hb0lDjNBv2Co55iHO+AwVaXALEasmoqe+jBoZWI1/F
FI21KuFP/80/VpDK0aTTjVQdnEOZEP7++nfdpCE9Sf6I8wujeLLVH452qTvd9ypOn0myMsO3rIOl
Z/Syg37d1mQt892oW02DuJ0fKjnDB/9vi3eATh8Acx+s1hNnnlqBcK5xwKJAvOkRPHm9B6OVG76U
CSTehV2/tGZh3PX8ZbTQX2oNSZsHbxxkC6Zyu5n0HB2xXobQquxiNsFOQDq/yI7LiPuVhYBwqETT
o1M0jAbhx1bGT5X/NmWbmnP1wqbUSzQLgCRuCnJYkrMaL3J49bhYj16puNwcH6PWXezc1gGI+mAQ
iMHI6H2jdo5hwZXlu0R6aiHt8/wejTkDEbFbsNCF8saIgM+s0MaysZHPunxugpH+UzWXw7GkuZmX
sduk083j7DLFzjqBEiusSfaeD5WomBzne+73sHWDxgpt3p29DnJdbAOR6aBgV0a5lMnVPmjq9Fls
+Cm1T6vXtzLXkOqejMb5K9qE/PgFSikYiboC6ouptAjrC7vBiHwNIyOFhjGmOBfNmktc+bMgycKi
J3oxBgXo5FRbIHBnz66fmg+lLgXQi4kBXw2MZaCkDbXwWwfMUzQ+rjdDniNwwBYR+i1c7TobOzxo
C0ts67vdfaPLO5uk5iqVNJ3cODd/lVzcSdKWsfn1/C6DKeMCLX1Ay+dRB7Gfz5uvju7RTMlh/i1X
lXydRuVDmx0DEH7jfFL/jyNR6d/IA408+wQAzfun6kYb2yzS8yePPaZjtNh4d+5bORmBL6WFvgna
/6FGopDIrk2DkQvw9pCx+uDuNGAkhesQQlYpQYILPwljmJtNyN7Zx6As7MUBvl/nwaJz3m43EpOt
/eihlg37WaIfUokFSXvUSqb1BgLWIEOtntjLfmR6MZmMQUhnahdOLXWjyYf2uylNU+GdMfZVg23R
aolD+qpgdpGM1aifH8kLlo8q4YdC2qI54fegHJIrpcodtd87YK1pyBR4omHliOb9Lba8g7MGrOZM
YEm10gqhomc5uKKvY9jy3gCdHksUCnbmhvwNSLBw5WfWrO8HqZFw2T+lqsh7vKHiHGyWjViEc/gF
006e60XGlZmROk8GJRgSYPabLctjtrm4UlExlJnYzaM88CZ8zwdnbql98qRQs0WjZ0HN6bBQGDOs
potHHm8MtbLQGTW9V26qXMudzNUx7tmDCpYuDAF1BXVQ/1llmnQmmbXxjv56jXuTDWyX9BDgz10M
KewhkzS3fXyWztIeVOUKcf0lRN6C7gal7xuCwP6OuGWWqbVESmo0zJvX0xljOu/06W290f8amVqz
0TmeNN+bEWGRo0lX+T+WJgnQONTiDvMA5AyOew1SFsh7hSqZeog7ycliGTrpJ34ITZUtVEfCwT+y
fgM4J5sgpDoXh1jydykWSHTckaHYDCoiLscTuo4XvPbyjl9f6gbTvcEhvRb3XyXfiNgUHQGiROdB
sjDa9VTrJZQ2YpocMn1xtxBFMGpi+WxbysKgC6GUAQKuXJfEJe9+ebjO87XEsTZpWEIEKDYKtKoo
CHNaNL5o/kxcKmvC0rtGkPoE5FSs9YcMucKvrqQU90LeLM4plL9IhHwa7tjRC0pstHCEHZ9O+C2Z
fzXiF9RcuWGIosWSSBvN3VtavQIpw8n4UVTtSBlPmiie0VVRqbVQzFfuz1W5msN4/kA+bNFnyUR/
lsCwHK+arzlMaqyocgbGMY6vI8iJ4G5sAJSf+vB5w5n/tWvG10SFcvEgX1KAAZv0WPCd2d8VNTmN
R5LzrgYAEcwukG6u7VED0UipEDZwYr8vQCe4+pDjMjrJKNJTFHyh3M1a8AN6Ecw39XBAKCmOjeyo
bFv1FXZEpJj6cTu8yHoMgU6qkMN3TNVhpfFT84/cXrtgewz2QLX0Nu6dDFFYdhMgFsDjk63xGBmm
sRvhPAi0xVsAhNCVOvccE6OLc4TUrbDx0lFr2x+FcN0A6yHVPCn6f/v+BVsUhkI+2GoBo+oXxL/W
zNj69kcPa+/kG94U/dxIxn8Sacxj4boANuL4uidcC6Kg/hX1ekgCx8exBKQjXBr5CvqqoZne7FrI
T5PVEDz4VfP8XG5alZxOCruSnfq6nJZQsuX7h8pQlPhOXeN6JoMIkohkW7EI/BvGCtBylfpz/yal
QCtznutpjMrGK68L4zgL3Kc5Q96ghp8vTZl9n2o6LrUtgfxnMZyhDCoL5oNWotnD5h2+dJueh/Fo
XOdJ9IQHUcSzB17/ehIQlML6IEAOT5MHN21rx0ZnOsnDtCVGThzuboE7LnJQ9xFysv5zJgNhWK9f
f8uClV7+zU+lNHgTccSeHI9HsvgBz5iMG70ATcPL13aINYoAG6maL9ahGGOWujLPWJdtb/oMd9nJ
CuMszFpTRd4pYvGPMlv/IvU4Cf46KG+gmA4DefF7NtCVEnYnMPDebUF3JwK2OKGLYFCTxu8r76Pi
uJOrwcBrhbfxBTGADrr468DCk9AyTIR3QsAEbgz3zXWWBq/QhABXMvWyRCTGzD9IMLEq2yIf8r24
80B0d3kVs6b7OXvF9QcGgB+pWv2xKWK5F59GhJ1x4gS6pL7iJGvnP2/Vd08R0IKfHp22Iom74OJR
NgwbwjQ9zMyxOdlJKoa9j/xkvu3NWs0hhW+kjiV24EGlUBdz7RUIkJ27G7qME3W5Zc6lCCmOPe/f
NMqNOdVXujBM90ddFMT8FzjQ/PBSGy5nKo4eSmmLXGyfUBnd+dFaaWx12ZoS4IMPmKROM9TSz5pH
uCxDOVqeK0NS/wEAw7rYTNjYwJgvELoK+RBEprdrRifzS1s6wwDbhlVgONv2QNw9HnGLzK5R6lsz
zCbFk9MbV3fkVgzvvfbpa6jq25TXaCiGdFtb7H9/4hdfyU2FUCG/vYPbn95L0ojq2nYz3TNkpYN4
N659C/fmEDib8+4rozxZ9sY6Ox/+31cBZ6usfnX1oB3ipr2AmiKmIoTe730SDQtPhGQi7pBlDY1f
p9I79q3LmnpCSvYh3T74p2yHXf75C+Oj3BbJcsM2gsJ1TmQhz72ickhN/dbDFSVW6aCRgEQPunwF
fhF8bkz2L5+HF+8DzixEoJIFx1R7rolzCAyXfwN5coorvdIBGQHsfAt0pJ3zOnZH/Az98ii+mNuo
OxaBfVAHQUXEKgjc2sLUmVG8FI+cm0jvlKS89xHu+rZt3PWpwPR13i9ou9Nwth3xeSmJkX92rXh4
u+23qgZKYDDMDxJBP8fJhlN2dM+bhECrDWOXn9DgaxJAXVNsFA/f9ctUbN6B49mSFei15gH1Xp1t
fnYIPs42wQS1oBY3S/PrugMCvBUAEZjFAz4pg42t9we61nmGF2yAY03mRfuOZkbR/qe0WOjubBSL
qu7NCto3eg2Gy3LfmUBXcrSQgi+CP2sZ0x1FwHue0rCVWZO9EXjxQiXMt2a7ItDM7cHdqU8Fbhfu
PifWqiHtwlTkQHbb83l3TBnb7FuZetSRR2ewKO628DC0C1bBMgJ2TghJWzPYD71C8mQE2PeEDxYc
hknu0h8/Ie4/ATGgSwq9G5ShoNLtawrMBtXC7FIk0x+ueQz1hfuLCN2Ro3glNB4Zly4SxLkW2nnd
d4j6yyphdEN8StXcTXVJTdWvIZJ+gQpu0rlxsrDPkeCG7RHOafZN5unQG9hMCM4k0JU0ilqnqGmc
b0zilAlveqtQhe/58vdArflU9KlBgyxLnObbbNTiHTZb53H+aSlwKqe5XSDK0pgJMCUFAKPko1cu
WsQyFcw4cVZ7+aPIl1ZPSHPCg2Bx9a3/xsjXBuL3w1NUtI/5HEyudEzciou6WCX5J1+0RJl+ktAS
gBDWsW1x68fjcQUY1JGDNZnza/1XZoacnZDFK7msh4pMZ4DUcbvEVEFXLUvQnlVMSCCpisczygh0
Vf6Clu7I+NCwMWTzsZ8nqosAFazqfXsJE1++UT1/q03UBsq6EHwtLDI0iOe6iC9a+pp4Pyg/9gK0
JRt0xaqkITn7UN3xuRwZGvCv/PbtaC+5NBVv1FGPqXgdjTP/TdPTg18qnoqqiV8WTDStec48IMjW
M82OkWZZAXGd0/PhtmXi6rExdczQQ6DtyQmb7BwWcLm3Wi0e66S+3inztz1XJp6boAwq7yLiFmxm
YPlTakv2xzpWsGvRbJAQw8WwmKaF0o6r5lVwyjV/kPQJvo3BABaI1/f+3kZhooAP4RxInX64+fIi
fGVLREc3Z3Y957QuurgcX/xI1A4UdYzMzAz1GDGZ6fTm+vvrAYJmDWYTcptJiFxoGhEyy8DJsCL2
OrvTUDkz6vH7oEhDF7hEZPIUfBK0rXAA6oF9Vp3l33cXJzJ4H7bxmXhugtzpDSbMLyHpWtmqAWhx
MdS3D1QB1veMxoP6TX7bgzTab15/aMTW6VALy+tGCrZkxB78wXcJNrgblRoj96RPNPFzC+Q+5qE1
WKAjsoj7mj88Q1j6QtMjveggEuraYdCh6xjZo/RAD4QaFf7UbhGhp2pPXhB6KTlPMRb3+kaAHW7D
V3eMqfFzwU/Zt0uewyVQxUQ0zpFUlcYKM3+s+9cqcemCw2PuguHVuSufC6mNA5N8xIxUnXyLmcB0
BUMPjVBSSbdGA2Z2L7ZnFMipNia+my4C5rwtdCooeGHnN0vLkeZ2W8eiALXGINYZTcdYhjlY2fah
kJFAHzTOfkFn1LepNoL2T8vAL67LGsA2Wcqhsk2Bwpy+X+LxaChyD8h2UdhRr6bfm+Clu4GxfbSR
Lsyje2Vmw+319XzhT0h026kCeS0/dqRcA6HYw2kRT19hUzhbpUbAs7S2rNl+SdtH6D8QhsOX+CuI
ISP9o+tpT1wKMF4tqcC+3rUzBRH/zoLoiEA0zegzAugR7fFZZ4mJxRaYlumKIkGc5b8wYhp8lBRR
MCNLoS3F7LhkyJql2J8vg+0WmgPw5SRzKaX4l5Pnoh7b3m9r7k68vPq32FgHF28Cf9+Tn6pAQucx
F9FsAVeLF5uzPnU/jPjmk5+hqamKxMMD7WN50zLvLlNB3THIgyhOaeu29osAJCQxo0LT/s2lM8Nf
GJ7RbxenZeZwPBOmHEMz9OA0IldHA/tY6QGyZueH30A89WhIlJvlGL/gO6fYer4jR2WyvrhXz4z2
z0GnanPypWjMv6pYRP4q8nWlug4M22dYOdkw+c6NNCwBPdLtZr2iouoF9p0zkA4WMnhKWF56Ou67
A1Or3Sf7PHz7DDAnXZlEIGkawTilUwDWY+bqYzrsO50T7SKNf/Xx9e4WgO26uFInAllFz+PM03dC
hhbaLbhkuJHAKrGfswiGse8hToGvEpNY7GuuDVj16+7JBEx86aiiXcXk60SUKRAjz4j1bHWPBfwd
QoNjlLvexVUn5cbYYk4yCG9yjBnWac3JRYQJqF5fnLDqBW3yZLjpBr5xxdF2HdVkpipwwpXAjZ4p
+LIgv+tu2KNlBq/4xM9K6Bl6epzsyAyK1he3BYn4vi2i1ZNc68i9WkUClrwCGLpTMr/1c90dIr9C
W2rc7aOsF9bCHC+kdOuQykr5S9FmfqqxBpjJM+CpMIWwaCZgo2x5HOo/cW58C/+khU0dei6WaGP1
yS26JgpPOSRQCmnOq8c53uEIcxaPMrJuNuyCR3sbwurmSzpPi8w9+wjc28Nx71YJEV7RuwzIzKME
SGbz6lOk+BvSJoaC8FkzbQ4+5qY7LnIttWe+PsrJQ1u/PFbtq8li7C5LpmomeStSTqX24+vf8vDP
R7ocLES7s3j46c/GoPfdGmBmoXX/YShISlxpgrPTGI/NQHW8yL/5LSFaxl1h1T5P3kY4gjKKaekO
60kac6SvfV9aPAUmgl4pGUfy9ajVqgbBR/xr60NfArLllhVnEqHNdMwujNQb9xmtp4GeBKJtV4Vs
edwEbXBRfTGGHIPBCXjnV9qmvfokn7vKNk+TaeeYtwGjPNEvvtfD7Z7zoabH5zsr5Wa+oW/YAjCk
uYp0G2nW4BPqmM7fXF48fBjCmaEce/zr0jCg3qHQow3ate3PjYKti83shBom3iG7bgbkUgu898Fi
ngktELnt4yw51hFRNH6IWvNQBG42TmEI0ByHJ84sVxHxem1eGeSUCzFHlFvsmLG5cAujWEAbAXgV
aXcdcNbSgPM0n1zOm24R7EmEHt1AAyEMrcbaY0x3+w1ZhaXzNfyqBBQ4U2ZbFb2c66j2cMlW+JgM
ESkUj9FbUJFNZIZVMnwC4KU2FGwsOhHwGublmc0C+21xXbqIu6/4eYlp8T/gTNlskmdU8HUKcSmv
KwltHM/DxD4pTcaK/G3Uv9/AOLkdwPNMK0rTt389LtaNLS9h2Ri05BLanid5LknPwl05lT0emqyi
HYgauQv7l0WaEfzKavAmLvBCQ1KQnsUlA7/543+6zbb0Q6wx0OUpgqNFjaBgRZfhhsn41AJl7sYR
HeY6vc+U2RP40AWvEyYRvoqAJ/P1dNwk4511BzuS9DtN3ahBJ9Om3o3gEF3sVp4JmGUiwq4Cf+tu
Op+pMqMJUDfVPmIDZkA5Vvh4rinKTOTspFJRo5Tgn+BcsOu7mdEW9ZA9C+EMdct6pJtp/UuiPbWq
0n1lmDSJbSduXpY1v0Qkfl0+fvmr9Ba+/yJHcgLuCGcxLzXfpCUbBWsT88ULt7SBOmv8yQRdiWbL
ErasqD4GWD4d4Jr97CDWZxtcbrCsOWT2CuesmqSGOd991bZPRehRWC6aoZ6kR+fCjmQkX0ZwV+F8
ef6AkewxiNPyFOG+GN3E62hsP4qs1+UgdAMfnQCXecpV3F/Eqo5a8+/97sNgisV3uDJk8nHc7OL4
+vnbq3HaNhzZskvDy+2OXgUqmBsuUTlyPoX1xKxZ5x5geuCgwqSvVJerEO/JtvhNtZcpOilEvHMx
K0RoBBF7sePRsBRn02AW38DPryXV2Qzg2TPV7LoboRacVz2xfo7oZOA0YF3WX/bOGNayPmUa8q1Z
EoPULLjXkOZ2Rjz3UKLltbZ+zchxVmfZmTnrfBgRGxLDoM5bxrqkU2BwQ5P5ydnWb+N2WLmDyzi7
h9fVzCg3WUtyFvWtEI9RtBhAA0eD4zfOYVQDgc9aunzKvw+TDydfBCR+M9GEgq9E/1HMQvGbWmpc
8dzXN3TX9XNBLXAUz+eWdYJhaVdubzFG4MA3LuKMVP9r+857ClBKW+0/gpt8sLMetVk1weimffHV
NBhKpsaRMlx/j65yaHMQUN90aLuV1coJxJPhREgHFxAyT6vxujT5Svqla9UtjVXik4j6eVz5jL8Y
YEXxpSVAt08/6wUXDwutb7VFD9x3ADW3b784briJ1oeivMe3D5NBzgY+00+9lDFZZamzlQtR9Mf9
eTMOw4TTC0NLnXNCx4C8elG2w1qII6g2PRTrpptCiVKm4GOMdV8IUTpEj7GbHxY+au0mEzXJUcW0
yIYO0KlpQeJrDzNm/K9zQCaENNLG3z4DLoFjJIIgNQSHXMzfuFmV/THmhK2UDN/GY5GHHxaFU5j1
8Fwy5XeaT3FbAKkYCzJUzgFH/lXx/MAIwGe9AfK2PfWfIIGrqIxuFrfd+vDjKF9RuG4n4i3KR3t6
g/I/UwsZnB8IOmaLpYKonk+/U03xzYniBYCt/Gv7RhlKbaEOOJxlzoODYjABWJWaQEjNrw4f70yb
Am8itf1e3TLmn2o/e55kfS0/nV0Nl5iH8olVkE17K8jKWlmKIzfFlVpRg2lpuZiOuqRr8w5iWYNO
mElGrAijwm5K4PqpwhU91Z6v8byeX0DB5Dq2rgrzUFGI1TzHoUcrulIwTupjrT0JriUcXBLBp92d
s+eqxAI5+l1xWHOfJTJ+TyIphrAxjV3OL5yGFKU8DIBF8Yh9nBd+zTLiSQT/NtM0Oj4N/7qeA55f
vYH8OSKt+dVBEGrPyiIVtYOrHuIbIa4qBXp19H5lzdxZPY1ARqsJgquAEdlHBnMb94h7XFByJ/ZD
MsrorISxwRKxHT0Namko8AmJW5Qftf4ov5cHiJSNGG7bFEJmK02J2CbmvOzjeheCuKk2HETDOQpN
D2111NcJt6gXCOKaEzQTH2qxUCMoRkwdKwRzgckSZd4GRMu4yvaf+W6vLzu6cTillfNT6aglUPEA
xjvKwH2d1H/RPB6HLwRhuwAmEweCwScXsTmNHNyo3fRx5pa+3i4lkiEHTWnqfMLUMNvefpxd53Bf
pLJiDgkc4rTR0WAIpnCDGzSaO+8mXl704ojRrZgC/nAOxKUXtdAjng+UX8Mgt746Aryq6wTojsdx
MC/0ly2tjMONxDvy32Sn6e0FnEnBfUtl1wAUajwNNIJaRGgA6l8NQ6kDGzslGFWZ2813j06B96u4
djWHSeJKn0v4SPU1Jsz+4E6nKiNPeB++KMYwcf0wRloBzd9nXY6iR4bnITWd6P8L1AL791Kt3Wl1
sIOKEvr60FsB27pE5Kpx56lPokzXjXzdPV1Xu8jkEhSjviwB2armb2GXLcoiEuG+Os72C0Pyr8EX
Ir6Wx3FyCpllbfrNH0bFzYsKHUuS6dVMIQ0qe40A1UE5bb9A099TkGjSNUSLnAuFHhnTUj8isRvS
v8JocfpD296JFxOEarl+QMdcPUS60xkbJHP33qCs829d998NbMjjmKkeEs+XxLZOnqtx+Y9kHfV6
HdFtMaGLTrFiMfLXGDq4YFzmZ5vifNvvvgonrDOLSWHKf6EtHQf/RYEqRyv5u4NlAYL3MwlE0Xs1
osMtgvbbp1HbVErJ8q+K9bWj5uQZxfkEdbPc8VyxnZKQOgDvKZiIjTa6YLExp+zCXJb/9lKmiEuH
QQAJXlJ36sWwBMHCO/wyeuNanyhpJHqCkFHbWqELIGrPasII4QPXpbtAWnW678bTGK39YemmUnTa
N+j3PQH22UPLOfTPR089C0ySKQ1xkzmzqzfmi0lXqww951Wj4YyhDr8tS2pBy2qaltvXYL4HeUO+
WsjSL8YwxqA2uw/kuNsZHeRrm/UI3MvhocLzrHIeBgHUtecfw4Yf+mwsq8c1g1DBQH+E+ckw+Qjh
tO/6f0xrSYtVqVBxMgVl0Ndq/fJJmAP0jMg6dl0QGQH80PuueCZMsc5vSTVciVNqeu/x3eyr4Xhy
H56a51pO8SFqrEDXV59EbWs4P1aIR07ixf3fpiby/9Ve034r+feYOiFupAc8IphlV19qgMCX4Fyc
QqGUfuUIO6TgGBo943GDIFjYOa0IFQsE2MBLXDlSfQpmYy3mees7cgbbgtBg8sdpLnXudVYIKI84
YwQ7xeCTIwjVv2MwCWUeHTE2jODUgXTEVxBOqZJSNOTuEnNv8A9gFn8ggzqRUnzg+IeY9xxlUCPN
34aISE3knQybOIJ4zo9gbdSfa9JqD2leE6/4rfdX2NHCku2ckbkFaKDyLEHrkQQ8pIKWp96okywC
q8AmcUXfRWdbEFZWHBvYDECW3glnUoy1gWDU+gq5fcQwInaCMSnrowqHisX7gd+2XsNpCkrtPc64
H6PdJpgv7VPt7LGSd1H6VY+/q0sbqYDUZXrTpDV7ppQqjuH0D+bYZv8avcTAzCB1Iq6q05i8Z0Uh
yNDZBR/LBKSBsCipPnSsA5mNros6ewoSkQgM6LUALdiyml6nbNvCwQu/3bubIFlUUdqOqfkR5Jps
JN//NuS17JLisoRShBLZFrg6AqRs0chPBxNgZ9amQxTUXpz9Y+4p14FzhiOM9ninG/KsbUjftzVc
Jy4Ub/q/Ea1IuYkbpSDNSWlq1LpUB9g2nIX3qXsPhrvKn9SkzViGgLUrYeXgYBU+uSNpFzMIDk8E
zjyS5tmq+lx2PgmeEosdFtS3K8CTULEPCCK6U9RyBhIuhzO3t19MiVKx4VC/O7Ee1aMl4vnUou9g
9XGsBYT42xz4+MDeyGnB4mzjZWN4AvnRk4FA9BTAy0ouH87ttmKT+rtF6NXiKnZGQ6CDL/G08mEm
yWECJGnTsALjoQNbTfjAtJjRSOAnvilNQHJHmELS8/AnZXJgxVHG6AeMO7xZ/YxL/LWB5Qgcl1vb
fcjdVYdq4Z8k4+79+hEAszCR+8skyDc4T7xmanCuDnBZiWjylO2Mzda8fZwxL4yPd9rWgv37Lnuf
C6eI9Cua/g2PoXYYCxi5G38Wv6uX4Ka/LvAhUHlUVBLSS/Y13X/pWc4Qucu5mYkQIlil3ZHf8E8c
4gL2b6gI0iSN9rHzvmKSiXB712wiyufuqLoOgKW7rOqT1dl7BuT0KX71VWlDSfu3yQ5a0jnAQO/o
9dN9Ath/6zvRRuldXxfvulA7+KoxDLhidZYJ0sITEymphtMthqp96gFAN7m6KzLDk+/I62X/R+hP
gVannp6WLH5SxcAPQeo6aYaNDPMjlWUFu/E2qjEiQK5T2ccX0j+/xg1CFd7GFOJxWqESHqqRRUrP
g9RwdDLEfSc9ipnLQt+zxy/PfMZTk6U4MswxsvCDIRJQXpbX4azuoRkmu7f6pUD4V5PEPBfNHmyS
9qzXrXMIGcKeW6CaQv3s11hlbjGrIxvbumbx8RyqNL/FE9YVn8X5FUZmPNuYYbtWQ2OVLguNz5Db
2QlIvaqsaSEI5pt3O1QF8fsbRKiuDsJio3rlrjUhkxJ0AraSS57pKlCvDEUCXLTusn9yslcAEKkd
ykLeZxCwemwEuL1DV02+G2bdIDtk1f1jWChcNVngGDEKumPZE6uweIle/BFluBXSDM3730sYbKCV
u6pjuy5Ff4E6P+Md2nmDY8zh5p2pXn/kvci1YeAKB3UFVcB/x0ce2IiI/uYpZXIjQltbn1/t3+3d
ssY1sfgCxUd8T1ZLge3AMIAjdZ8jc7yvTvqYj4KnMDKSplkToBAXrtmo+QU3XLXnbXXgaM8/xLkF
YW8fOatSRieTmaAzEh/R/rpkpY9L8sWKMjmbeCjsSNcOJ6gXInUjjrt4t9AkgffuKDe+3JMphmkB
/5CN4ZK/s+wC0Tdz8Q9BdyC4MeCALsCEzHOSwlq0ZX2874vwuNABLvdvHF37YtpVdpEU97eB+MsX
UDrwSR5ORiQg1HcnJEiJM/vqx9Hky4qV//tREe+m63gBDiTb2Fs7PtZ9lO1X9414btrZnfCUTUrE
GraX0RCXO59qR9bdcjKbQ40dhhxVlk2cbn2kiCrRw4MdurlfIkx1MHTa05w7rH6yEtk21ZR9Ypi4
4g1xHRBUgsf1TKNsp3PZvPuYuuICYnhcYmglYl9OQQuqIr89AwVeNcsp4UbBXScLI/++YbU6jCOU
pfIQ0QRU9PCK22RHNmffMSkT6IFLWiDziBUObsVdssR+xqezvR8AVEQnbVgD1X1cgZ8BWpCDmGnR
Dda7H4ct0hza2aFNSMDHU0uONXx2tC5G7E94ajsnIxM1uVF/1+Dt4bwWXK8zSqRhrO3IBfn+grtQ
qyH2fs4cp7qsfSXugryoeWK4auW826vBxEsVrFxKl07x0NnTZwT/Syn2qAvg1yYIdjYiOOIxAOtJ
lP0X9zsZXKzmGwXrEZfydr3iSG7dsqmpDFHRkOUr2ZIzl+rIqYr1DjplFnaPb1nTj3lmFGKoe/dU
RYrDv6m9IhFrJrabnwELMxy2PstNgWciPKWO8uoB96evmFP0gYaHMD7i25LeLdy6NPmTrKS3lUBw
SAYrC6m63exRaZ4Z/vwd7OL2ehOo1OTtm0o+BIUqGXJtxAnFGvxcUDNkxK6EK3me53SEmM7/5gaG
G6UFxbUi5k9C3mR2gPEX2csQiQxHIHAvbTvoXO7pbgeUcXUNo+63UyYiAeU+/SvOrbE+QCL81MyP
dRgFKww96uJIwClrSBzZGyVwdAyc0TspgLEfYXh8uaeZgY6zmKrQrvgrB/k4ucqaQ0GD0IMyq5g4
iHmgwTF21I7v9ih4UlK4VcGOrvDTLIGZtBDkk9F4Cr3wtg/KxyusYXe0927kk2CcaZJlxsVZidwM
3rzvlkDbjFjHuS4njtFfFnVGsm/VSd3hZ4gOuVuJ+Yd3M4lIBUcqBDYUjj3Df5YCHI1UyVL3ZZTN
tNMKhuXVE8jHLo56OR1VmrC/nebW5fqy/wlSv81KU/XyT7O8AnlaQJVmnC/rGwGTlfR74Hggh06/
S2ShTdNzBg1dFrLMjLM6hq5NJD0JsTtzyLiycKxTJoqpW3mNrssQn3QF8iKrraGXrYRodZuh9a0J
ePsYy/Z3upxMB9yUbRDswm2PE2Ex/DG7NOjnOp34xg+v8/XO0AYnovO+23ilTktmcQ4waho7BEAD
iqWxGFQxDUhGhGS79UBA7mQ8xLyawTdy1LNeycuZsZUGvKCqLnwOYxauOnQneswZaI/uJocolwiC
1p7wzgWkTfyLBjw1BxqEUvX5NrYKmPhxJzNqtwnl8hDmVYrDm2209V1uvfu33yb82ay9bT/5fnXd
lRS5k1sRvQOkkEbUY/z9vmBWAtQApoa9TOSOz0BS/S35FqUuxyZFf/fUB6kRXSk43myJERSUWMWB
Hiizhen/4gOo7nfWazC+Q3jwJXB9/kxVY4lg41Lr9mr0wq1h0OGPHOQUSALLT3UDlX3yMsdc2kUB
mJOT2he5+85e7CbgpynlAhltb7TGscCH7h/MVqoIwSwkdfKBHABT68aPf9brwWFGhogPUEOXzwHr
zzPRpXTMcHoLdiU7Xsm/fvzQot0eBh6xHA0zCsmq8tMHPMyAXEO64zut5B0ZQUSxmKFKqZOof2HN
51Cc6Cq5M92G5rkyM6lhlvZnPPqY+e/fBqv88OPOC9fsfF4Ys92Cp+54dq8To8fR3ykRivbS0qvp
CuynCRgC3m8YmnNyD3oTsAzzNGm/UDdR+PMuv3RTn9Nj61auQCv7DQmP/2xRgB7VQC69DcpJdEXX
PEu3xiLKjbjCzuz6W3VaUVnnX8+d1TVJoqLfhZa6bC5b9DLXamAW/g4wckqHn/HYCYg5Fy+IDawr
ETXDWD/GGhWsFgTdvLRryhtBwSJCmg+9NmMgtwS/7tQBOtFNadbdit86kRZQsUBTLHtujRu6LiOZ
lZNBe2hPXKpMm6t6jUaYQbn8BcOEBy0MS+Dfsdw3bOPUyHWoVkqiIsO4kbldJDJtmeeU2JHIiUFT
nX4mkHGcvQEaU/SfPekCC3IU4At7IU1sDhNxJ62+HWK8tgslLAvblztgY+bX6BL4BCLeCwa4bNEz
hRFNIz8b+G2u5VhgHqRmOiLKn2PbURxtdrnAzRevBl6EIVrDLTKa0J9DFwyqzl6RYXEs9qjfqGBs
xdlMzJRAv1AVF6AwhOBFuO9rWnyOqrFBi2jj1PHjbjM6uv+x9EvkraIs3ITIFGoKx9CBkO7tJRYn
yOQaSSDvIdkGBMicgi0at0kmCH+r3CzcZbN/bs3HlZmvm0lCMZgZZZ07D5wM/PpGm44tg0itV/KV
5wL5eHipH8lPYbc5Gtx0t0cCJSLwJ0vfv9yvySnWtakqt1tMg93xFmlE/pPO1kw6sAS0EfCzfE68
SO2KhbCu4MmqhdTaBsjl6yRABzdX5o06uJeasgfv97e+p2EmOleKZew+FmUNFlNSMzCbsk7S7FVO
dIqlqVVwZFzp2UO8uUXUmRXcGPGDC4P+BcJrRdW0gspHdOic6jXKPJaAurmP9TIZP0FS6wuuDGdy
4NUZsXxZtk6uJWhecgJEAinDAhNBresyFZUjNP3VJ3/HRrTut4FScM6qmlW3qlAp0p33QNlE6/L+
YGvCDEd0zYqpqZ/EH+yAqppnbf68hrHrG99sQ6fG4aT1PhG6KLUUNKjjuB17v+gxCPqc4fKK5QHL
AEPK5XhlLn2/KGgfvZt8W00N6ubhebwvo5DUbYofwgyXxeXJ9vz8CN7Bp1PyX4jbBIcvlmeLotyV
bLuhwRD1+NW0d9/0a3z3vcr/ooYAwplQTMfqwq3zCXyXSKNIG1xfZUMWMOdG/gry5a5lOUdq6dci
n9unCCzT5M13BMX98+iFVNTV7BaVROFDB8wOkUDRr0dz4oahtt3hhzaxekFetYbEjhXJIfP6ktI6
FZZ7IDWpeTtwZPk5JXa9dHywLlvEav3diriG8AWNpm/cvIEkuo74cx30NpcBO5lVvv6NMM5gevOk
7qodSNCAdzi/eNWCDm02f3s5SRqD8R1zRUdj70FgSGQVhs1Sx+Leqw48QrfAnO15BIOF/pog/Vdf
eFhpQfDcIr/algzXzDhG0EoVsMzMvg+tKfjM2i7MvEgoM25/TzhH4Cv1ddRJ9YmNGOYJZepFM2rq
g8HSXch69ibmpBdQvpxz7/OzZvGAkin95YVIQJF9zrLPcpAYxYL6WYffqwvqDRzWCe4H/eJNDYou
RZ0LjeTfvrCeGPqQAtJcKIT1n/ThDbTVLUtQZVMvwHRpCyJbyAcCKnZm/pWS67/yk/ioRh1KCZE7
LilXH7RHLUa++mb6z9oydW76m2njBxNQIZKsdXciDxzJKIvuVfmepivK0eQ1DnIgZTuZlbx7p7B4
L16u2Js5Cr1yUw6SrUY45REAXC9Qdq5XGF6LMNTTtqaGDfKeb5FYxt+LVjijrDXufp1a9IV6tzti
y7+NWxGQt9fu8TCtuVxYNuuU+k7UdcOw1Ug6KZneFJCJUJEI39eGS6eDodbftlPagTWfYV16HI2M
ph8vmQfyImii6/FX+1ZSP+rJLPCiBdY9XKlFIpxxTfe4g1lJsY2fMU4xjeff6YFPcu5q7TOBQng5
JJONvvoVgQIRkJ6K7eMKATytPNJ12LHOQAVLGOXYUQjNpKE9wUT1aQ6Og8ohE+ipSIZm2XReRawo
fTYpD4C98q8SjKXWHMLMyWdl0D7nUxyTpDvWPyZLb3hXHcx2wPLv9O0HJHygNdcY1F7KUVEXrXuw
iN2U4bMkzFH4G7IyDOqI3ZutPIL6Ev6FdjG3aRXVs6oo4Fdu9mWCVuAuZklmX71nBm5SZLBKa1Tz
H6pKC8hyZlftM5wUS6DPXNhdDUrNvtogtrXmEw4T3O8R2VBQoEw2qUWQuKYe36ICu5BISbL2eqJc
FNC7QPpVnKZqRAslwDNK+xGOo9fVn9wHFa+vcCHAcpb8kQivs7tf+TwS9krnzwKnfRPanEstadz4
ZVEv2klu7P0CQt51l1rm8SJb8gmEfGSbP5Jsk2dG/yRgg+L26YdxdQcxhJV+GnTYb41pT2Okq5Zm
z7DltY7047uEJt2yEmR/LwjOZ8CnB/boktQfGFDf/uzKUG8CEao6hq3S6stFoeUW7JnENQUiJC6N
ehtKoTOhso65OraSYEOEO6AWXkKWP2iNBtTuIt2p04dkK221UMi3HU/YoQzx6yDQAAvjBsfe9VUy
BCIHP+SP8z/KQC7ThuWakER5cfeJLiVs/g3BsITINsi9kLUOGYhpvnBm7gg5E1Mvo5TsFTFk8vjs
dk2DqY/Qp4UlI4N+XMlOrEuxwUNp3v8pderCheK1e3b1dkqzJbTtLPj1YI4RJm9V13svf9jPIkVV
tciB+icQ/wGRV7gKjNgYHsSUNrLidHRTFt+c9vUn+wfj/E8C13uG4EYXLvx9MHktyS6wuIElvpEY
VcAvujE53+vLzOsTzXTOOwdHVLCCq4NMpAcNL8FIzrI4GZxdJZ/Joj6d9oX+MyamYHaxlk90smQ0
DbH73e5D2Uch3kymHyjA31Eg/ZcyrYTyFlzadIP/aed6OWeoWY1AG1LAGZhUfAih8DZEzckd26yX
8iqT3Lim7D3BuIkn2PP688U0e4bMbW5uAAluaCgR+DmLi0x7Npi/8wYWD460a3lfqyXbEuOM2wDt
ZyZiDylZvqKQNFbCnLZJn117JsztiZkfUPAjjJTyOqasVcAii+wQHsXxcSLIhY4BdMo4pZo/eFXD
Dq+p/8jvihpRM2YAjTxT3vIwAcFtSCcSS1yd3xl4iTiK99C8fn+U95hieBYAqNNgTCwFofN8R1nP
YMPmVTRGj66DLK9uHUJ0zeSvFJOFZHq827VAypjJqiDiBZlfAkYWIM40ZymseQeEAHprPdrx8o7n
XxO6zqcoj4y9s/JsBGuS3RQxTDYvf4l149BxN14p4oZnfje+Op8UbHXQTV2DpT1/iFVhYcG4ts/D
o0GUK68jpBd/WIwMeRbg5LBm29Bto4WJvrbfw11x1AO8jVKqqf0DIQpkoEXV3SG7V0fS/Ndilw42
x8ac6dfdgfDnXU3D3DmwZ5HxO4vAvTvVhTa7kSQiRc/e2PuArKWfWctL/fnuQ/U352TpdkI1On2Y
5YHOvOniux83twbnnMXH9fghmxTOIL9uNvGnRStaCmnL86fzINvPm/D/f7EsdmFeSR2ZU9Tq9pME
ZXbe0a9mfWge3ShqeFBHDMYRNboqpB1Phw5kQ5ofEAuIH3AGBfKUMOp/vAS5aYJc5DipxG84VUS/
3T2GlXWGPSO3Qn+0LoVvRL+tfjNJdaQero+hFoYAroedn4PyMdXyHRIvCwMgdtWkGX6qPjsF6mej
+FGoY6g+OcjDilEAv1+xFTbwE2DT6BScv5PiStHlgpRlWP8ZK88txTp1QuakqfHxvRVeQrZIVy3W
Hde4B/q4IIBHbSJqw4O1UdD8ng9anLC7T9nknlGEd+HW/zXI096btX2UbsMXxqIdebNep4Yv1MuC
Ku3pWSJUruUGEzSvIb5fg1Ao5njBX2nYl0nzwDV+rya4HajEBvpVSlEYHGy+BCxiAp8Hh6oaE4Kq
9VQmjp3VrTWoc5MI6rCCIzw+F5CY6FJVDsxta5mURXxJK6cmkq6wbKo1GUGB4lxkGnh3iD1uNn6+
PsiUFIq6H/X+gEB1UgQM2y45HwDabU7sti0iJ2lBeL72jhbZdLA4fPC5e9MQK/PucCxd8nWwFkFl
YnbNQmWaKg09sVleJVmzy5ZVFzTVmfcEpfG3BPyiu/me2M8MT6OYjYk2NMRUZ+k1XU1Q9LhkARl/
ngcJ0dYEW9nFBMYwpWOVVH4kb4GWW9joP7gv5+t4ga23A1M4/k9MWZWBsxXKVy1IGy80M122GWBg
eZQv+X+hxt+UVXFt8W9B4iutyP7IWA+qwGrW+4HPNh7yojGeBtNJ9PWRh4+eovYeFr8Q+ys2ZFVx
4XpATOJZVXYanHDWnObsdr4xR7MEbAR7b+mOWlF1swsmShnOpIf/92Fr4dE3Nhziz7kY+mq0PQXW
c/KjxIFscMTmh+VqYxG9QFHtte7+s4iilAi7eDopqMdlNfNZmFkh9S2lFIG474yzWb3okSPNxdM6
Nmwlwyp6/znzZtRx2vgtbUUxH27+uwJo8pDnQQCm2oN61zmZetf8XWMpBVFeZDK34xTmSUISFOaA
yhcXXT2oi4M8vaGdlRoql0ryIwesV3ba8Ai6NbO+8yCU0yEQhe/oNPGA0p4MjGlcvds9Y2iF7lBb
lLfGlIajqcuV8Ftz0YfNrsn8qAyhg0U71rjvsUFX8yu1qjnUOmCFhUhwyAPYOlRQ+TmxSEvpKOZR
gRvcws1hqMVweERbxhSM3DAjUdPjBwZ0oADnv4upqxpZiqpEnsoOMxZekM+ZsPHLdH1dIRLe2eKP
+UKXbVC/8zQxvtYTNdGIqaDmNV/e2JNlLwxN7J1rVaIRchqTCnY+NwkBpYnQQt32fsPNogVWtOEb
hfg7aIA0ntS+e8p34sHAH5WflAByJm01EtGh/LkTUGEGmp1xQQPsi5jS8ccc/0rP8bZoHiD7Ac5v
CRSMQ269J+VsNoDu37bylLulfAM6s4H6gYKY8bQ7qgdzEDHOzkZrxd7suXLz/ujBJyPWppSdM+Yz
WB9BMbzj8Q4B9nprNMFrQqxdbRgSUVZ12CmP69pv2W7cUJ6Re30ytw60c/5iez4hWHcn0KJzxSjk
sIsBMG2oieiLBv4gFx/KBCrfGjDvkMR0VKfoH2BZofvdcGCFWWUVu2fxYCZ68Pe791HXVUKqVdFm
2u4Te+/k8ajz67LNA2laACd3b4cpzGmBTZeGe+Zna2+/T6smlUzhQGIaZp3MPyTHKMY6HHLwF7yw
XGCDoQbjMKvosCjaKDA3ZkOnM6v5jtnIqIb7AnTXuvGvtNabnHMQ9cxQ+MdsY6yX2B0r19jl8mPT
65PUTPHd5UeUGNTy/Jyj54QYDUdjVPRjWvnQvEHFj3Q3hr3Fd0ahdrxTjJ9JCJmR8/PuuDxpFZaN
LK5LkuPcHgMLXqzFSsxrrZ/5cwIzXkmfBICsliJ3Whnh/M0UpiBzyOvsiOCaEGoPyLlmOMq7Yb/I
ZqjU4lQWmcHp+IgvhlpjXTb1Xxmw/6xcWMsrN1W/JGLpU3QhGws+kwyIreSqOZswj+Wy7sQwHS/C
s7ZYhbcmf5781IBxjiNSt61IFASBY5KHSy1EMf9NAo3QutCvAtalrBX/9EhOSmF0hKDEbz95hF19
cDhhHKqO3+bk01hGJNu0WrV3BtbX12vW4LwygO8iJW3LF9PFtnhGbSEGljRnD0iwdcKoxLiw/LKI
dRa2VDRsowWo1vYXz+ViBCXrOH55hVdzEn9qnFjfRGbsuqcwlbF5CJ4J/U4BUq39NRBTwDqavBVJ
SvCMhbFZR5IBt3Fu0s100r+MaLehcgi6mN0Y5lpTyJh/zcGgo6VsQmmFHQEvx5wozlvK/n0I7E0r
czu9NanER814qSIOYN1a0T0tmLCWHOQbZf+SS6MAF3aNDNYLYAJhAfhQIp+itKKdtAIGWJvhBg4R
rxxjyIT0DvknQ20W9ekgiPbVvAjXS8nqcrDadVg6DupW2efA+3ewZ5U7HKNYDBy2i79igOCkgKhC
rftEX4IWw9N6vD0KjSyI47Mz/KQqlh+YRYH2bgrTP15XX/eC9bdJxFkWfIVoz8LTCroeM3dny6bj
LEObw1rUCT5hfr8WgO3teuqAa5pZPJ/MJdXuodrw1R4teWO5xLpc2ejDRsYfvwJsvDNrvYGKepIo
2gHyEzp83w3H9Hx8GrHGnoebgXMExUYcxW5CfKuvzkw8dQ2LtB+929M5rMY9psKKc0qIvUkuCw5+
SAD4nwxF/49q8IJzKU9jifVQ6EDk1WjJz+qzKxhZvDEk8pm4k7Rk2CW3DkOVbleifGPn9sZti78V
96C+weK+jUXmXPWuVCxS8Ax/cAE28o1dPNMb0MAlJCeU9VlVuyYEpYBX7aBWZ6uk0j1g9+eayzpV
sjRP5UZY3W+IsKHtKZ4ueKDETwLqJL1t1oS65lXOpjBKMlxlGXGGrqBzL8evzCVvyH5ApKOllR/+
ATWng+xBeNKhbrdokoyQ+9C6GxRN1kFC1KdLXHADNgT+gpvbEFzkLT8Q1aY5j00hEIBJ2t72OxSZ
zxP2kuiMEckU/aombL4KicEdz5synwxeiwVwE9ysLYbcuZvCz1gDII7kIkPPJxZu/YEdfIOG90uF
B8DDOKkWB0orj8De5Ndat+eJZPcfMk2YlJVlWEGu/C5NxCw+rKzxWWrZoJ6qgH3vq81NbTQbwsTf
vlBrnkae52c6hbMBg2aM7nj7Mc1OhAi9WmiLprt6gG5001LjB9inPTT9PKBp0Uz591bf8BIUXD3C
GeHqThCFbk1tSp0VvEYDgVIyBWIVdHU0DVKdONw+JNWBYFncU7O0RYZCK0ZjqXFub4s8TYZWf/qw
oukyJbRG+RWtTe066+3v8dJBqWhbDCAhbT9Ww0Tg8MfQI0gWMy7r7nGU3NJqj0wBylDTHVyfweJL
q47bqVrPfOGf2+g/UPGHZj69FA0Ak1MwO2yQSsRD9SMvH4VFtZDLMI52145l9SJWXnXiclK4V9Jm
EseIKROOyGYYIXak4v3f79ESh5Cs/EZ/HkLb8cU/Z10b0YrtFbIp1Sg2ypdFL090eNrRBIOW44uS
ElSGRbCq/3W65V1mRdSKBqNM+WfI5JjWhMXfcwXeMGVCsflq7pM+Laqv2NFv4l3xiyUz87iFdvME
iOYp8ocYv8i0QjL3PG0HAF1ty7odQ4wCKkM1s/adf70+GbD/OBlbSYI198rlmkH9YnPCzL/JFMps
0gRPaqhHKIhnAmabCWmUbhuFmHb8vKzv5uGZTHHQkMmm6z/yIry6DoQkOarLbxW2TZkdPjSffy2o
TbvzuMMFoQK1wXuGUnGSs7ASreA6AUckoyHSZ6U+2tDNDO8c4do29a/NOq8P2gj3KWFyMaEDwmYv
fWaftMaUzguzOeB5tZ41ED+/inrN625CiiFGMhuP8zKVWLn3vE7YGFFwVDVG7Z7+rWAN1jRSDOgX
oP0xjAzH2mqJ+ZAiIoZVmP7uiEumyAyABiJWXagqC+c8bmkiWv5PoCym4ouMzftzX1SAuoJJFdvp
O+RK+WuVqbKNaZATB47nqH7KH/CREztXLjDLmvaLStgbPaWX0cW2p9W1wOV/YyDvuLxuj6RuDd/U
51e3p5rCrQ9QHcp94Q7nTkf3A+FtAgHg6Oy4W/e/A6POoCiD84DM+EqwCBq3ojgtDnJ4BQCNT/m8
ZHfR62C9pIl7tUseuGzKvtm7WWEXx02RFHOVr0teuYYyIuqqKMKe30KyBo64a61hDAyQEDniAZ53
81QobvmDgYArFJ5N6hHNLLCGb0eO+TEWmGv7TZCq2wRAR2pNXEc8Bmm9lFM333BfZ/EBiJi3sGEi
RuJGxm8ORqkL3en6cReA4PVeZ8HkDmBrvQwH1eyQ6ms1aoPtKZxMwoPB5kMEP2SEZxx3zbQ+ApfN
sZDiXh8VPDBaLuEEnakJGmItdqMRdpERfiNpMruNEvc8n2+MK9k87Q3k621AD/m6F7HuUEPnqzSZ
X0kQ5jzL5chWyp7A0gS1DD4F9P/6ItQ8cCqiYWvKBKJbHoqv3KsLEh2rZVGSuH20aGRMN7S0GqZW
OHbhBP+9lHQTXJg6XTicm9xIXNHgaIXp0zpU9b84/eBnHqrC1EIJfHliGo6ea5GUwg75iQkZk9nW
wZnjIaB9/PXrYSUJoXdY2djwCsfiuTXOCo89O90dbQoJA9YDJ+sJYzF87rG/YOa7DKUV71w0jiCa
36BX//aYqa1EuB9ifczmyy56UiJZp5Y4+0dMuI7uFFATgeSuDnqkLRaf6Ly+4SpoaOqhb+MPO8CT
Qy3tZqOnFTGwvgMSXhWtyaiFpDDq1dn7vP8y4CE9SwdS4IExTLHfiwIE4NDuq7VGF3hor8vGc4RD
u7Hk0miWg1gquYBc1uXxAw193YlEanNhRXmG9lY4rm8SK95wNb93ld5VPF7ITVXjtzxqWyN5t8CW
gWrvB9lyu70+JUMCDBIXq815c3N+rr9rgLbD6ogBw32bcMK1/xMPh05WoOgRoT2H6fyfmpiKTZ/S
8MwE8AOxKPF4ReEjgO07KKXEty7DCCXQLYUjQR1p8NQe1VFvesm23jZx8CbiF+vdijlxx6Eni1sY
wdLFFis5j7ezVUW+JZj4qbpCGNrXmREI/ZKvL2nnBQG5C54rnu7v35bf65UtOTb3xiEAt/Ivv5Mc
DPp6dmzHpHQG8OFjEFfG+8fOPfqkDkD0k7vnbJU0D+U2RC7L0AZGh7veP5qd7VI6Wr945s2t4ByJ
s2v/e6HYTYk1SSQ/9N0RByzyoB8saBKzDe+elGZQUvnPrFnplj8IiAJLyg1dnkTb/NGMLahtJ65W
DMx+UK1MnFBzB4FTXDS3re/J9vUb6M0BoKiOVuVZu9BmPZdPAhCzwkhw4StTwxG6MDKGKCnMT8g6
mVjPAfaNk45iTGOjrWBP4JMg3WTGME391B04JI4Mb8JohF6uwcHwAp/Y4o6iq8f/aUsb7eYryhte
D3/FoEpqja9aDaleGT8LQ1c/wMJ6brZdmltoAxe7Lr6mfHMdDay5bil2L6BzXkNvlVh6EoQrldy8
x/yQbq9eVt/GuaR/1h4apolE3QwQaboXmF/TBHUCNMq5fMX7hK8L7PYhyg33LGuQZJNOli6BVyNI
2Ya3PJvOUP276ZokoXB3iXIVDpq9QHj2cBqrjK7NiVlTpLyorYpvyaOVsKSYXCfKrrNWM/dj1sYh
r8zPic/xXTyPDOE53YyKmqtD2ym2lQ0VSAQ0ryu9JEOwoR70nwvqYsjHiujRgD5awWtcGSMKrGhC
xfry10ClJwoh8mx0kyWV8Y2BDO/b9TO2YeLhtCVtSI3BFLGLCHeGMf0YIUOmMwEOrbw1GherWTL4
n+v5WOe+qQwrL6ZXAEq9/Y5OOlkTq77MxG8klTaUz0u4J/5MXjEy3tstngoYDmH2mMkfegcf2osh
eKmSLImum1w6tXqigh5oEGMkjpZsdPM91e1nairlZnySge13zBHm/bT9mb/nD7Bg56QfHrzSF8wB
G9JnoIbHUIPKel0PLoXwqr3xMJLpvgUMrSDzVLbX6p826inn0zzNXQg6jnM0m2mJ9GEN5RBiSvRD
hc9eSlcTakdy1jB90ffeuM5lEYhek49Y/ggbZ4mmU60BGfmINeA91Ll5Q7RKt2kw7VaW6saZV9T3
G8JmCAnpjn263q9zfvJMWfqrYpxNhE5A4WXWXb7fx/AA3u7SHZ+JoPlJDUdKSe778QvL/9zWx/zx
e6pQTA3QOaxdFUhJHm2x8JARVjZNlw9zuHVoawnBqvOChpw/wqd7OOs8CcPbQIfaEIOzGIjZBWYU
QJPUEerxS0jWj7vtBHdViYhOfZGFEooCZ2Dy3iHZkFYgQI92LTrtjfVetXhJSANA9Gu5Bp7HrOLR
wpHXXvaFTLG3hEtNSBC2wuTLl7gi40m4HQtoAp6fmktrS7T4rEEJYphBhV6TI63UUucjk6cLYGJj
IVOJf+X6BkKmgI/DTz2Y+B2zCZwbm11oPfrfgODT1hcPe1MaKt0zkX5wQe9RzZCo6LoQ6q83ZhH8
/SDH9uumEaQtQSMPSEkVPCiOC/WLcu7okQURzY042TTrZXV0lLWPF1pZEGbwBFXUKcazUjB3MQip
vx22ZMj+2mjZhVnHBrhTeOsaf2i5JPP1gWXO222e432gX7i5oo/56PwzBa1znbmYsCD5/BtK4HqX
Xf5ddlLXhz1E1bNh8kBkiWHJmldBHZ0aVFbTteb+UQ8RfqJuVbGWWNdQdmDs7ffuXGP5uJlGNYno
Rp5s3EmgprLPsQLmNSpM2cdTWA07mD3bfqC7+SmQet3O7l51MvOKgHY83jHeJ56nfDXpCAAoXqM/
6EzcPwEK26MAp7yzzBgWx+3nJ61Sc3R3j3BvQdD2D/G1Lvj+LR3rSaS6Ia0ooU6W+UoqM2nT3OsN
dWjnU2TUeL9oP4G6iczMlTIjVC+ozU5f1qi3v3u1iE/mxozegcINLLHFdxvgWRYX4abgf/H14WDM
eTv9h+i0v4MuJjZSQx51Tm+eG4ZMA8zdW8cjgXTd/Gmr4oscF3MnIBWi9R0kYZ+BdfcO/9AAp5wo
sNOBQgex7GPM4/PVOTfRTpB0Fk9R8m2tGP7jeMHgGluHdBrTtLrKK4i2i+4fW9NiXYVzlmgGICUt
4L7HrDi6iRfglRT8TpjwViTvUcqH2KFShgD8FBnLeipDBNlNAI/pQzCYvGxOnavn+KPa3N9KDHua
p90FbIkkw8hnt7DDM9Yv4A+u5q0XR7+kfZwM7yk1jX3HBab0/Om4mvPxc0g+z3YumIGxt2u4mjqg
VE9yTjdkdSpEb+iWsOuDb09jyqz4ucuOQeeHeWz+nqXa50fwHc9eVkNE6ONl3taafgIj6aOqJaM6
dcklXbZqG8CnBgrvliijee/iCNtsD66dRkMXP2P7CWI75yxb05ne27VNq8++PVr1SLXdKV9TElH/
YCuY/w1qNSlGwW59+5Q9rppma3VG+R1WnDdHVZIbCmRyMFJ844G0YfLKyZNvvG8Sf+UInDsyxEOP
Uje+Fmj1gBupChoIykIYVFL3lq+XdyU8WeOy967qW4B91lD0M5Grbtyyug4zh1z0SoE/IsCoedui
J/HHBpIi+ughard7aZGAPbi7GM8HQJ/GWNpfgmJiRLb9A4vOmzurTxsK8YtTox2zzrDmqWigwbeP
ZXJ3PmFpr4UPaxd1gSSzblRPs+0NoHHV+Z5g6HhNcWhFJTh58dgU+uUcYjYKsy8o+81nz+jexj5w
Fo9ud+CUSIilbkr5lPSU1bzOpjNE1TgQ911x/LegKBytTWn0nDFIsS7GYFvRo1Hb8WGUM83ApTWH
9/8Lp/yz0yLiTxWz8LaDlUeaYabG0g8W/0wkiR9etxY21D1jWihyVXFQLFKebOUqn4iPRR72szlp
JlBd7wTgXgJ9c9rmHeix0WyznHXqgDdhaSb3gPAjwoZc1NCFkS6nUyv+568edjkjh1bXDr4gtfAG
keGMg57YmbPJwFrzAFHnNAO0jo8o/56Hl+j6sLcSf91pLHFCkAywnW2YpPG1a3nr5FTbJb+VR0io
pskmPTH9DsVUTcjRjE8LNEi/YeJES+/RuhZ1fvFNXw55okXDaQXkLZLBzdGP0GUc7N/XYSczck49
qfQTPjFNLz4Hm2Br9ke0QF9PfgsHq7HbPRjiiyPD2FI4IZCOn684rLM0gZnKtR1QXW6Y1AREsHbA
66z6NSWHfLuUGwOhhf9dWHKyz2DBU9DIw1fOr8SpfWLOYTJT7arlafizilZOUickeEHKSKtHJ4no
58oxuFflj2AaEgk7dH6INJu6I1+z+WpMDDzubQ0xOSTZbU9N5SvsTtEVa0DaOlY8zgcJ/KZEMbCk
X1mOJrjoevG8+K4npgj1UhJjDSX01htalBdxx2KhklLcBf2QLRg5ai1EEHM9LkXn0ojpobAg9OJq
3r9cKqrvzvVDDda66YUdEUZ1mhh8JFRc52Dg82iWR/9zCNfQF+nwdNhkfZOy8m/8NZ/Qy0Q4F2Z9
YmVPFRvHMkbJULCujbXggnxrcnjdQFyvPcfG2KrS+LAZ+vJdXNA+4cVwyUIG5lirI+Do1hR34cuN
rf/+K2vZ8z6IsWEH1GOFKTbdW93r/OexMrBlMGQSABUUFkJcAPFvNYltriIGfrXuxaertFrJe/1k
yXoA05spcB8MhdqwYmlmISoNHh+gvGTGT2YdE5L9iy5q7MdiQcq73RGxZ32rv5mhCXhbp3kBavPk
wU2CXbIh5Tit0j1xt4EKm24ZIrM47phRuZ16Wms/EqfUekb+lcKuaBgvUcf/k0pP26zw7RnBwxJF
K/+TKxykZfxats12YUGVAjpKki/AxxAz6IaIVjv4MBVD/6c/rirYY6pCHZz/I1YbWMRMJ9GHP7lx
BECCsldOM+q8VDQoZk2cCAO/Edlkb4jnzagqUjhbwrQcK+IkU7ZAUYwTOGfuNwaWySfA72l9qqer
i7phC3ZT69dNQ7YiScw7cW2KMzL+Q73yLrJsbfq0txRFeqZ4eqrDy1CT+mG5I4+pGvn7oojfbrEG
Sav2PZNpE+d+5gxq0EGYwJQzZcGgqaL20qsc3uIEOEnB9uWoT43b1Gnbo6Os8I/wN3JYbQgLpedT
bEe5XOP4C0EbGkrsc0i4tkxZCEaKN0Hejyn9WmP9oQjdrH7ardlpgbh+Gk4uVr1cjOWFRQYZuA+N
zpGWElcWLSsIBufW+W66KxpEvTU6LTy+cBChF/6dkTek9u07iV84mqk7iLzy6FcWnEiS1DcD1Dgh
W2kkx565IouETWENMcpbvNU4U39U3S04yWsAArCNsWWj1rVW2VO2elYKynKG5Yu0omLilpm+aLL8
XOpL+BGQmJ2fncJ0ZMiZi7EtW7Rsdu5/KiccT4MaetZiDot8WvWO49Z8DF4cs1pT+h1gkWejru9c
73orduyvwW2aJEhJT2QfH0JdgtPpWig7vVgYQltkX2EWFHkPRQb0Hfgr3TWryyUho67lHMJjeRF2
kn8jDedVrSqLk9tlYpH+WlBBmsIYhqRVef+ymyxWun+ycB1gVch5zWMhq7ZB4FnYqNHr7dC3Z8QT
LfXLoash3OmkDwKppbeJ4mbYzGxjBwPUxbFJCCbQl8wXjTMh0wV/K+KO3Oj8Kwg9X3veNf5wCMsS
E1+P7+NrZFKZAFpLfI3yuqpvmnnxdqtvUqQgL0I6qEmI6f9Nb5AhIa0e65FE3rxQgleMGJ/rizjW
y1L++c/ubO5Q+dgbDNCQB044ikUdoj4Zbz4eeX0hQLts7H6DK5tmeM89YF+5srvAmbGreRKmEGeo
F0ZqfRJxhkSWha0EkLizt+GnWHE+yDw08s4jJ6mtzsS0FHKIOMusQA4sVpOAt7cUr9xf1T4TUXEu
UttQKyl5EMmspMNNj+r5E87KO77SQvHTVYhBfWW70zmOQaPTvEvFSuCKafmzKMLj+jb/MzKIZOF2
aFcpu6tYgVuyDmr1al+cnpqf7GiSVcO9vPKIFuQS7OXCyQZEllP10+fZHeJpwnWUfRlRxoljckXK
AF5N6ux50Of7MK+UKblOaEcVuSjerqVkkuQAdiE1jQSNRxjQPcsN5uy1ohGOgBg2wEnyrUGx/QCU
I5Ul0wBy3bicjoxtfxZ/1VL3aIBlxo0zlnejKNwKKLKWLvPJlgKeEkHenQI0D4WH7J+3YD8EP+gZ
lcvKWXKEhHMqRq4w+k2IMZImxrDba/W9jN9ALCYHVlUeMKT8eQTbCl7SDrLhjbagLxMsCddQH/63
727xwMKdlqQlqpJHZaSLmK999v+tqKf21Jk+2Ap6DG8t2BzLN4eqRKuP27ki5xES16BWHU/EC4mv
NkSbER6CKc++vOTJCREtyaX6+qMoYHJJoe/CEqB0WJlqcHnXIac+UimW0PwnmCRvdjrRUbPjYTF6
sBJSP8f1h1POfwfNZ/yKFgvA9IAmZi76nlB7Fl+6raTztqXmAMFEdrfm4kW4XfF6CR1Uo69Hedcv
j54oog7/i67ZBBEW2fL128weQ1gL7CIXQMoiDrzG2bX4EjNZfel1oiTBVWFs5dkDdVM/DxiUFz03
NmXe49mrl/pjQ8ZaWc/UDQkJV7vPrnJp3RJfr9Q/+8C+8le1MFs12EYQu6bngzlzVtjtowPT9UiD
Yeg1f7JfoKcum8ESSwAbvH7mXeivulbJfka3cPcz+bFgceqpaYrj5hP2NzaMdXZJFhm6+Td+QcQ4
oZQkwE+ZHPdgV4jtKF/nNHhhbCiKI1Hj8sSb5YY+4jSBsk8KyGWZxZp+RVDi9p0hLjq8OAyxQljF
k/thLOe6KvuWBKJt85XnL9nvp71mW0oS1JAc+ntHwiHL9rHA++QVRqXcccmNpyOXZdokcsEkYI2Z
JScJAx16ita4ZmVEv3Rqf7IMZalqxMGRNirzCsJHRdPdNQo+5k9v1UaXIBVoKj052NG9Smaoc8PI
N5OumapZEHv3oxkMVF0GZbRbeSRXV5LhR4kVYIpRnWGFLZOsVHwuFcElawN9mcgFPXs3JKzRlD6R
XjrYmJSU0NOUPVIqvSbjEi+V4n1to9PW+nVPLFK1u83P8Ao96Hvw8nUdEvs55AJkEEKbRoKSuMMI
u43sb4UMAOUXWC1AWCSNjlD4aKV0cVX2Ok4N2xB78/l3/yUd4efnVN3K9py8ZwqqcsCcznSVt80i
I8E+Eo6J3APG8usoCKzCCzjoAE2ve7264ihQWHdcqq+W1GKHUaBCz26FI6qRo1WXwHaCvenjy8jI
3/igieEdDNlANX2VX2AYbpm0oZH+HA0QF5YWi279zZETTbV1GF7ocvzdfKfxNOGCORX5Gma/iJlv
fZh24mFL3VyX0jq7zs19GDmCfTUYy8mzJPLtB5847pBmu5v9Et7rS1fXF/TvnAbR/GjUcyAVaJMX
NjY33hg/rdfFqzUvRULTJSjQk+q8l6WsgrSS8fW+xcnreFKltt8jozaz7Vv2WKfG5Tk/RxW5GbO7
VvbrYo42AgMym0fo/EMHxV8nBJ7jdNhpEHVinRuYtyLpl/zTAQPH5dUifAjrMvCO4sMW82RfInHq
nWX6us2CxbyNyBwng3S39zCmtKtVpKNCFHgMuweTbfhM3IraXddNfo2vfdEAafhMR4Q4WJ7OxL/u
jgxgB6RJ94yx2sfdgfwqouRTKwGiF678fVsxHmggUl2e6VYmzpIAC9mu6SyeqYuC4W+vay6APvRY
59YmnZhBtHG4GSHPmKS1TUEBekL4zYmo9dfUKU39ZipLYzUzOOVZdJS+BwHG9uvHl/EKAUVTKT6r
iaDxUxE7Rj6CwNuiDOQKW0CKb5lR/uJByzvel/ybf22PU7Afh6x4sZdg0pYChhoUkkSzQ+KHXimC
GfR2XyePJjK1jZ7SCkg964mq2ysvB8j6mSONkvnkOsmKvYfmrk17AQDapIH72kZ1BCBH1t7mwQ8X
zw0ZVgxelCJEilghyulGc2nIioGP4zoNVHUgZMlxgqNemeIC7Zu1IgHaycAHY+sd0NWUwEiT1vvk
ntdu3T73EJiyS7nJkb3er/QbbQO0ws/KLPNBmg78QXFWKTwDDegX7r0Vyuh4jjv6N0K1cDPGzIcu
TrWdj7qno5oDCHBOB77R9g/F2jEEyTmdlb7+AOMFevK/ijqU7gRa71CZ4xm7udK+63z3dcUqSnMK
DAPdXuBFXK9DElqOxylU4Gx3xgFwfRAvytrOpJKexRP4DtFOOzbgIU42yHVSlbtfIRGg3bWwW1dd
iZ2j+agaGlV3sOH7hLjsV2nWs88blrXDNFP8tGPUrnFaO/AmZU/RzdnY1OPmf8eTU8oZ3tsiixxn
aTPya/dhg5cawSU0I/E7lCKzFMvj0/G2/u20ZP3Nl66gZn5a/M1aKcUAOJAlxTdx3WJ7tBaHfIy4
+/XI8mT303hsV+5eF7IPy15MQeCXobzFk/k5wI8zZX7sy62930GB0DSIlA6gsru5hZHfY0GNvXBm
VJu9gf0OwPX9tTu5TVEk47+vq4T8NMB7JXd3pHIRz7BzooWZFkc8SztdERc6hhkVORcl5TDqj+hk
jufXhcQciphOIennF68dBbkRyEd3GrOx27Q3B+B7SHkLxCUiMaqL8iPyMKzPF7buAYAZSChnqUmm
dhZDoyB98gKG9f7el6ESt3qd4LLkVaCqYv4a/HsJYlg0nQs+HCaYaLx2TTY69KvNN7L/yKQXZcau
fBLPJFex9dSHmQ9+t84xJV3x86kUixm9IWVLcHT0JYPxUB/bYTUEeEWCk/Qicd6POekBsHOngoBD
zTEnJADJS6h10TBJYAWtNwqP9GwKaj0bMaNLp/AGr3PeTwhyfjn+ttwRwZ5BjoFhUWGUs4Id3dWJ
PTjLZd98DgmRb3oLoCER/XWNyJX2cGGl1rN6wW170jsBO/CPaAs9imoJGhy4ptw7IMR0/re7cIVj
9LScJ7l1SIOj5e9mt44C0CGNCOKho7nN6KFvywL3a9PGPO2lsOH4aZ3R7ocmU/JB0WWgTRn13TBq
XBztn0t8zQeOXFNtc8rbTjM5voL2nRpRnX5a7issLZm7/k8moDOBMpjiKmHu2+xDhvp2Wf4MbeIN
C2+ZGbk8a2WypkmJKNjk4mzGsuK2jx2c+f6YuAHfVRj589VMw18plrmXpe8mTYmnxzqR8UJtqpRV
5nzrySJXpuLuhC0VP6+8NIR9Trm1hRrjyT+gO0voX862mR8fH1qSUJ8z4Tt9sKG4HudT1ESrPvAi
19ghmSI9ti9qPhLpkkzx2W+OpG6+5T5+AjkAedXfU7RiIH8I0jEleD9pWdBEgZK0copH032doZyr
sxFY8cl4FuzOgMh82udyX3TFfMsijTjYy55C8J7OHQQAXhmO7356+ZcqWBPpgsHLivw7ZjWMIClg
JTWqaObt1ppEiyE3LD6/BZ56tLKLTzqS7PaDaiwqQjbvSvtsfuHwY4XzHghb42ghH+gVYdhmZixb
uv8E3IGrkKa/QUkEpOSb1I9zaIJM5JjJcR57NH05v1p1y0xjmT4tIAZCDOrfqO3fTFcCrGIBFXiQ
5SPJaV0rppWvk2m6KOEvCiwUsGEZaaBSLE/Sj6BOwnY4/TkiH27ob7mub6cP6Q9QTdf+WekNH2B3
55IGqPUjnL8YnD5CuixbqW+VJ8EoctaRw4SKa1LgOPr/1C6mFBkh5lV5c7IrMkxPAh1RHDBf3ZVD
X8Y7CeDTsXpgbBkxvVzG0H24FKNulM82cZCTLbv2LEH2ocGzQnMv0oONlFiy9HrMgzx0RW/PdyYh
OiVDJa5BLWh/AGiJ11HBeJNzkmPYz6jEjoLnaFa7pcO7Ezr5Dbd+ZiyKHcgNo02m60r8XbkgrU1E
eNTs3XTZyL1wdAZ/IoxrJd4Fs0t2U0n0uqTSs0P7cs4Q+w7hqpQJrXob3lre9z7NZDCTltceSYUt
mJoudqdeFEy3vs0kkHa/QU+12+/M8LbKk5+8gW3xHlqv1D3LzrDHVZNSBbrXb3SVzunj2uoG8BYZ
0y/50mtDcgVShPOA9Akn1x7XgfDqUoIr5dWriwpHvMM4o7jh9GXOTQWn3nPrlM3oxRN0dDTKIeus
4pFrWM0gplYICfUqX3WKoF7dJEa1ThByAbt45kEKKydYcruIH+7ZzDweRJtRqa5svoRj5fLAwNDQ
4aCmPVFA8zGtqfBRZrCmRt4NmXnaZzF4HquemqWXQmnyxEprcm0V5PjzxpbtyRWAlZMOMr71+PDq
cOXLU1i8+Lr11Vb8AiDR1XDfSqi6ayd1JgSuzeIMVC7Lw2Xwwpocvrq5sGzhhiFOjKUIkw5aNKpA
I9sDmuQA71kVOTYd2hEJWp1tD6VN38rjQIuRef8Cm7nI+N65/q33lk3ysCvvnmodEHBDAZ+Sx2yQ
abKdttx01K+6bnX6N4b/nDmpIBn3XIK0qmp59XFRZckiuqMw+KQjHzUHXDvSE3Rdr/uZWbhQXd5s
fLnkDVb41+tUxmB2/diRVUkbBqFlvh94TE2QW6aYEljcDN4l2l6XtV1bEumEYaDO7oJlFJBxbGQk
nVUZVuxjGFzVS1Z9js55p58lCKw6lVg8fVn0XYxyJQb23LrRqu8kH2wynDXlplxwGbN6y2nJCij5
pa0l67xAi+9gAD2ee+Y0F2JY4F+zq1tWjYH8O7D9YJKNutgX9wKFfAdXDZs0LLBPhawvbOec0yxD
a0hpEB4xvT9cPxRJKUfPGSc69aJNdtnvV1B7yiTS8yeX01tKiAW1+AzS47dzS8GGmdElbcKTU/NA
RkzJv8MYPP+Fi4k21ReCqnxggyc0xGhTiLAdiRlLgs3wsiVPX1DJ4QFquiwfGpe+Nk3C/7/I80ym
wl38HRTjxwMi/JWPPbLaBzKpKzQXcMu5DhH2Xe6+fB2KC/V+E/ZKgVqjwXJJolSfxuPTG0ktEi3g
55mkHI2ldVKT5uag3tFPjicYNZSOy0UXqDCkUCSS0SfK822plozet1oxllQ3co7LvbBHsFUazH1S
RYKn3li/jvyow2Pt9JmQpWylv6lHgVPIj6YRMNjV88F6Y9uBB5z1GDXlH+ZbzE1fToxPJ61lxvXL
1RmBCLed51ZQ8R15JSeT5V7rhHEh/+XqE13GQXrqCN2ZP2gOUizvstGfY4vnAne00CshxcprS5Z9
NzzcB5S7KrH9u9OxnLgXMtqBNmrYzlAAWaztAkmtFm7ROHLn2pm9finQHPoHmtdjzHQoK6yTCReI
9n5rFVUdbT/FaM41FZDvEyUbE9epHvLKgE8oBlXHAueW4wOQ3dDK6eETtTsEQCHZ+eaiaC9dPDHa
H3jwqzRZFAdrkQLYj8W/BiOC1BG58FdnSSZ9t+8YeJEkNUjHSMabVYNjU+d0PMyJInWn8vRm2TUO
6WmiURwwdIMG8aAl4bBmtK6yYkEZIcDFNPgf7whqdiVrcoKK0+inIzgwDTEUC0PsVsBLWvwHqzJZ
Bi73fOzkrf6oipwQWCwPwxqLm0AsVF2nLz3psW6Axn9mL7sMD1lbJPidiP0QBM5C0n+WfNNjfwx8
CYxEVlguNE3MXXxgTfcpKaxiZ+GIG/aCgSd8D72LEej7HtG7e1TArkWbJAicTzq+YCB/DpvufbOC
CSRhSr8hCJIHKcsIrTRA/cReUWQ7moJt3kR37tscqU/0gpYOZPNoC1YBTvbDas3NVzE2Fc/SkBjw
HQG4W8iJDF4ZgpGWXyqs35CojpHeGcfWQ7sF4iJNilKnyd5IAxAab4U7NPiPrVyORz9OAKi7Fpi0
SfRv7WFCVzVbkflH0ChhrWOT9xMmYWdt63agMz7w3WrpCDqPRN7w5D0ioXVTLNkzKQdwHRW5epqO
huzeaEA8ew+62vXuPRIVA1UnCm+EmsA5kctVC5aqdlSQgR89vl8PdQMp1pl4ji/yaSAzBGg4BBvS
ICAeHMFDC7K2jvJbzkAZDv7HiQR/U8eNGrWNk8AJn7uspRQBQcCJBQJ09egvqtju0DXRe9WJKAK+
gASJfgfqcDkVni2K3BtgPi+oyZH+d2FIwLmz8qEOF376YEQrETUh7mvgnml29QoCo7787bxLk2y3
JAG0SdwxkhebvlKyX3CW8azQtrfMX70VhshU0Np3lpQMIyAOo7Cxg55JN/hYsmFH3117UwRL7Nnf
puY+iGMxNtw55RMALw28jccBLO9M7yQyV+8CqRs9BKEu67fsnN6kKBYoej0RdHLA0wnmQbABu2mL
Dt/8EvTIPBH5Wgv4qb9rN3yE+3WcSryDf/sU3GBVOml3quRR5+5R0tFSxdIqKKLUIcaf7AFNGALI
erZNMqBZPvOkHgMzHLE+lTh4q4SvknvpS/g/+lsTiiwAqfEHEm7fpTiye6Fv+2b3h0TBdAcUkCeu
vmB9YqM5lPEyIx4oeSxKVF9UCPIm1jG17E/g3odiNgA5Jh4Uxm8+rgDLlBbBmN4X8SWywxEXe4wt
xSw3Slrubqz1zf5ipGg0BQXt+vsU+CJkuI9NhxpklLHPIs/KkAgLvRonj5aYX5KBhpf+Z8UIgiQ4
S4kQtit+Olh74B340r3Y1WLup7udB9UMhWOdivE5f+jTsVjpu6mj66fqF39xtWxXa8zbVbrytcI6
lB7dnOProjXD7lAkBpNsch3DFCwzb1D7I3NnkBZVWytua7a5mBUZRCPUawQpEYorJfrKZL6eup5R
k2sIINdsFK0YsjV7sRjehkIr+8LxDpSIUX9ol2f37cWFMPIToAx4I/EveFeDBv0lyQyXrn6tvsPp
TYgTeIO7CB9sor/HurBleVGtQDZT0UQ3i5y0oEO/RA7LDZzIuzArcKPqqSLYK/g23Kc4x3FO9TOA
Lg+Aq8L4xKLHzfsAeLOBiLuLCmzIza9G9EvoX8NWjhrmjvY5n+E0XyB391aFkxoov+ZDwnmHwxfs
T4Olj8CSkGgtSKBp/fYTZoTC2Nkt2O9MRc+Lcb9lDdYIoUaFV6swlOLsPUQ0e6Iul2IV27V7Af/Y
oFsKJCNbzEFGuPClwLckZGM1vygd7apjV57k80YbF2YZCKUay//xsjTGo3WTPLRMndGzYIMQsHpo
J1mf4DSoC6AbvxePIAcb/WUXtEJuXN6F1ZysbKKHSN+oQNEHop4rErXGJvZ5M/vFz/WRGUAsBe59
IgoEedh7+1TyvfZd2UIsv0HVXzbTjXYj9WaeXTx3Yfdf4MWVdFJM/K2hRWNLck2RaD+Ef+5ykP8z
qfcQ0+1dvXw3P6H3LSpNyirj5dVM4Xhk697L+tKLLq0cF2J8uv3NPdE1EnWS7cBzkQbMxKNV8TE3
jqx4909HLZ+YqlXmuKUTZLIj061bj26vvBhQqTzVWy0s0gmRwLfGdAmZHNHEknVJA5LWGE0zxr+g
cNnOwUY9ITPt0t9zt9RUchEUoYU0hzq53QCWR/VrrtHhCXSH56lH1MwY4wHyCikFWZ+e8FknsMiT
pHTqGIi1uEo7bEd5rPrnajDNBvJSX85f7wpobz3ZOnESJf6Kzx2issOkh4In5CI2ytWvm8YBCNLK
UsFHmCa6CUXXs6IQkuFJq80bsDNe51UmP7idXsCPkCKCREFj7siogVTOHCk6InQY7cnn2SFA8LUK
rUubVdus6ZsRXuUrB9I0Eyy3OqsWWQ5UadD9pESzU5VWpjtgPCJyGDBWev2jBvpLrvSnoJbVTzqc
6HID17f8ggvpE30cMssCm+IlQivDu3TRUMU1f5HIfUy86bMgxpMSFP9HTPEqgJUtBoIqspmCQHc2
41FW+s41ViRZoi9syxD4kwgV/p9pvtwP0+WSm4kwfbSb9dylU2QiZYx6aVtoP/M1Cp2OnwI/Atd6
41vAHOR/UWEA0RW6+tutGo2ZHy8HZlJZOp/BUrrFDis+LwC7jANc7n5Gx500qXzEcSm+EMnTUfLD
TcfDHCmSblET/IhyXW/iLPRZ4Bn9HCLLkFq+MGi9PzXeivy2vcZP1xpmi3pv0g7MQsHaQzqyVKFK
/PSSyfZjDO+1SbEuWHcDD4aBQQVObAZqX4NNDj99J3gWfPhZ7xsva6itdDdCTDM1vm21eoef82ni
gzUv5E16d1EFBQl0NDg7/h0FWrPupsTRbE+XhjcelZCcUMe426m7YiS0huEu4Sb02usuNmYjpNgK
JULhl9R9nON3D2pUmtpsgFx/lvCbTnyyI31QLYCYEWYCfyxchmulbg6KAsWTsnGEYxhdgyl471qI
3T9ZUHGtF1zH0XF/hs7xSlI7jHAUPMHhiiVFCr6tWXOeMHFKhklt/wNhhRMAtvQbzTAEe7bWfTj9
x60rs2bPxF0unUekgaYf3krvEpcmexLn68vzkCn2SJh5FDvnOyfksuy0vvhAe+zjIsIDsOOMjoJ+
pr4amgo1hR+W1wfxy+esgp502bwO81UpRJ5OU60x7P/lEoMJfRIVj2EOMu8P2UNoUB9l0JJ6gAIo
5HcRjCK1UvL3iiq0iGb9WvW+o3W5KagdUwkLyCGXQfK3CxVsFlZkyOSWIaTBiSgoUmGLLIigJtQn
3JAIkoJm9t/xA6Sb0C6v1pG+HDydbyZi1sygZ52CfaGMS3sAbpKiHx78ZOkzxnG7kyfAzWe7BnEA
wTbmd7+OXXSfFp08P5+JRMX04HxOP8itT1pcdSk+x1HVQRDAkjKUaF8sxdLbzfofSE6n4HjFwHi9
6WEu6N/3ZElp6MGPtkLgDAHtBOUT4A/kDnMeo8YD1se+XhPquJsSB/VEVXJdIoBAZNOA/piTAaq/
mx5xZQK0L2ZZsvn/5jkFhDjIg5LM/iAF8tinrqwvGquj9wjzPf+442vxiBYMF39E2H+MAebD6/nM
5ZqpBhOVFRixz7akoMMbPdm2xzb6Y9eOSAxMbzJ5Q6opMiYmkdZBuEnCcGdH4bInTQhfYKBg7l3p
j8btAjRDRc8m/GSkaeo7NCrJ93jzc/tmg5hFn4+WvriUR0B/3k/oXJR8u12vgTuJqUybstUi/yuY
hy13M8/4ShMOoldxvOouP5yeMZR4fIf6zfBvbtf82mdCubppN1fN6wWfon6aUMtKiSCUdL7TQAzs
uLeT3P5QPDFd64N+hS/zygUW72Rvaoyj8BQf4aJ+SWvQNG14a1asM+GrEZUbXXZmZ/1B/f67H762
XTUj/4xwhXXQtJClkYNyqK1Hrts8rSggqXdcd/GvHrcJaFWgmeSDK0UQ/fLn0I0+S1yMXEcEUM5D
C1IhabRzj38tGFhgby40XmK/DTnh8desLvgiPdYK+DnmekY0oYbC/hMLtBvkRlRpS5zc49b0KzKg
bByLMzuwBmFAlnO2ehyUQzHj50in3tDF4bjKoKkvTN/fJSlwBHbVcKV6oihS5otA5J6AuD/gYq0S
Rjngrot+jNkLK63t2Ha0opjcLWre22ed6lS3Ehr7MIViS0iwQ/HplAAmYTR+QfVxlKdcuuuQbOoB
Wy/2FZBA8zNq+U/auc+jsdIx4dPceaM2v3Ph9rhfdDM0dzuHlKWyZgtlkzVTmNv7bFLoHAOPN7M1
UPJubTMjgVjUJmxWt6Crv4NQvZnIruWsoT2HyHwQfn9Y+FvJ7eVyNu5es3TU3eL/PYW82HSDQT+d
2hPjvr9loGhliKMoZY/ewKGVj0LX2HLNdnjIowAZmkJfMacte1jgaVZSke5CgKC1VFoF098iI9/y
vLv0bbX1z+4YaL6cTHak6LwWmd7Nb6rNNiNxdyW/74vj/ZBqyym+jYjfBa+udeLJg09Yidxj3cW5
ek54MU9OA5xgawUAstpVzAav32BJbzRdfCmmiCYJ5ny9ah6at9x+MqzXH2dDyAXlU4Dq2ZKUa6Wg
D+qadvsSfasBHPOzQMJLXwgr/mOpXqW7Q4UXV9EmxJh1jOHIsiOLghlc7pRX7SBGp2GmVier4Ipe
r70THWcofZFNYc7OYdGQrS3u2lnSqXWsdYGHZADczBDT3bY4qPS6ig0A0VpkJUSI1Bvyz1Agn5gw
sBsJQKzOFINy2eSunFCsyQDuNzs5SRy7U71GWIqgxXs+yYU4BDtfyp2vPlPAlucpUHKUQMOlPy6y
6rI8HS2RfgVN0Nsq8W5j+8Gc2zklOkfNJJT/wrjpOIjOIZb2b82MP9+u3cHVyL9VE3YZlhVNXD9w
6e2SLxYsebQzo7opbxyzXiODrccmdyCzaowbHFv12PGRNgx8Ho7dsL1ZsH93haJF/O5klDu7uzJr
a6EHE5gvNNrHcMHrRYQ6l39l2XpD/rY+rsRxtASj1eXjwTbNfqa4XQjsg1PxPMu272iYn8nmQT3v
zTt3OhIoOM8f0SDuIeRw9pGbjgAzqwgCYMoVyw5SSkjeh/rzwfDsIXnvsBcrjHqrHsJEhktkd+1M
nnXb8leVfdnXbO50F+aBv+Czd1aGhlX9GvflZhGPQSYkEsl2s1UxL02LlFSruDR6UFzlhTafS8Ie
7MrSVjmMky8foa4kAKBux8KOfrt+b9R2FJ4yjJ7twM5ri2hqvhRBFpwFeU9pyy464R64yAekrZyg
LW5IFaQXLTFl8azF80UBlRHPaVUVL2/W+jmiK73rKxnVK3BgmMXGJNtsxFgSMnV3Cb5nR3HoeDTC
QSH5YmyAP/8mex8dm4bamAr+vPs0RaGb4DI/g1ckXgXTD+iQQk/3IfuV/M/M3khiTvRneFB7uPrj
WqtEKPxlrRROlOxU6PAJl9UFqX2LKJLGQ18hYMQiK6yYkUnsOm8nPfk+nLHgB33rGhEqvenkE61a
Ah/jsy9ybLrh3/8Aj0d1id+3Cb9Mh+gHokZEwR1kRtjgVJjKhmOA3kfZJduMOQx6D3O8VT9i1z1/
m4/j1ZL26b0At+iTRaikC2giOyVhlpEboOyXvC4gXfR7i8r178Ypyw8tvxf5KRh6DyxxDNTExJN1
x7+b923tvssz8MfIbZOL7cJBzaYG77f0sgmNFBLjuzYrevzEkw2loCiCnfOkD+6FYyoRXh4JNlRW
qkcuUUIM5Fzpf1EcIuXpnAcloxxX0FU7FAKYtSbWqeHQYZYaO4d0kdq92fzjaNyaqQqzr4VB7ay/
Xal4jDIAZ8iNWCAgB62uI3LhYsVh8VIOhrym/ySmCj2sxTyYs7GI5Vha6xIVPexRg07TTWyYd5l9
3dleRVperlCRjx+zOleKbTL8CFbSfxZicehJnUQXrzTY09NlZh87I0LhinCkyr1OSHFZk2y2JclA
lnRo2Q0u7SDqZPxh7SJ1fNZgC8apLIFgqXVSuLxEuDb0c3BWHtzJ5+0k9rEop6z0aCqvcO6Tiy/d
rQ++SBqbnS5km+fh3YW6iV65KCoLgniZ1Chqr+ZC3ZIbp9HtsWaV1aIQc2CuLNdiofo9yQ9f8EmI
YgME8osCbnH+esNhIOJT/RQt/6RoygpkdHAL98BO/TU/6+NWSThpMyyuyFhngODLXLPhsFO8zjDu
tZk//PnKy8kxGNI+/SmFVdYKcE4kohB8s7PIBRdXq2FBEBpL8agFoniKcbpbj8JEWi+MimcUGu+t
obdH5x0oEqOPGB9kpeS5zrPjRIsnkfuClF719IEsGQ8eFf86CosSri575EI5zRw9psUBvmg5HvGr
5wOhdW6tPOfBK/TL4/m8oRUDUcyg/fxl9y0rlPK6TJyebPB+2LitGKikTfzAVhYCJZX9u1/7H6X0
tnZz1Uxrju+XdaGKI0Yy5eLfp419CNqohAXX2G3OOx+Nw1qyJOWjYvb5dscdkmmNE9+QRFq0PYI1
tRqBuG2VNDvE/5uhYBjZ+eeH1dvhoh1nZxwtLGWhNj5GnzbPH3M8WPB+B8i0sa1hNt2XJHdfSg6J
b2PITLLV3KQ2KVsygtcKkFG2E+WInrMHvcLbXRr9dopBi/qOfeZkPA52R/obt3qvMIU1dN7j4EtU
qQyuUUokxnpEsll8IskduFeUe3ZG9OQgnflbbzs/X/jM006Nv7nFZfDjH6GmDBn8jGPI1Geh+5hA
1bYNeAJ9jyc6CILD0O2a7KIOb3bKLYiE7AEpCRkoT7YwbWAGPcqf+QOgTW7r8gamxrpGBRpv+uP7
134/nU30Ars1UCh35Z7F6jPzsaDzO3Rmb8npQ6VdeyYqV9LGpA3iL126e9WcL4TmXnXDcogSK6Fq
LrQWn+KhsRxuggzbOiLDl6+HEdBZQ40cPXT1Esh42dU1+CqbMO11HHUX/2Vi2/ojwXmHD56z2ZUo
y1QiWe+NuN79MeVvLw8//a06oMWOK6yKlmtwYHQQFYnA6BwIrj0TVwpMKp2u5j6BsgvuJpndSoS9
6gpk0abr865oWU603b89mhHxuxBf28V76Bikb2gXHg0swkZxaxy+1IEgiHN5Ci6eSyTMWrSwTM7E
rnMmof/RM4zIhZHBXhEn9Es60Ua6lKjUoQi9NIg88blSRzu252NbZsPH7Z4JYLgoSVQATlxnm7ma
3hgKKeUjs7wSlejUm1j8/pAAp9czg9D+OMTTgKOt9PQNNyGvg3ofLPQmCZlMyb2gtRWhndOnVzbT
e9AWghFsU5fynuunHiTK0Qpptyw8GmHipSwqhDVbInMkVUJix5pNPZtJBIH61DlFg83pVFjl2mU0
A8EUHlbPzC6HFNBsIinBVFJAHaT9Gnr5gNSoUfPbbxPgpw9rTBPmC/YD2Ctvh+9/8viEL2aEAM8i
X4vl5FfS9BVIWJg9JoDWigc5GGROzqd9lxcm/cHII9TKOMP6zjSwugRAz/TM78lxAEuNm3um6n3C
IhP2QmPmQVBxDwtP1BN8+F0mwydQaOAET4vLUsVlkDRV3UTFZrcLlH3nYKlikwa+vAe/Y9c93kSn
d2vNr7owScJ6VTf436iARISO5K2tO3+CC0BrnaFji/I7Ul1zr+xHJMwIqy0XoVKBYFtsDtyct2Uc
v06OtyW0V2aJPqtYJJpiqTjhGHBaCADOFXzVyBwooVUguMeQ9Wo4fSbt5/naKsCCzL2XDbQrJrjU
kwk67QVo2eZPdwwj98lXMWzyySO3xBTvZT+86mc6pAqhCbsiH5ov7FL/HY9Ran4/Oi/wT0zAhwkU
QyME2qitEE9V9H8KDRhdByNRqliq0LIz8CWwLUA77Vk1YPuImwYwJ9coZHT7gSiPuGhIbfDqwuT4
nJ6GILgaoRQhx+DdhiOJAByrFxaGkWJUlKuotuVr38vmG2y0/iuA04k1/Q5rkh0COIpdxKajyGSk
y4F2P/dHh7TUgBXF3etggM62SHQL40sRTiPDFYZqLbn0eLe/0ov8V9GgfxJtPKKXEuXhEOuGfgT4
wI953EhPY18Gut5GYXg2jh6UQy4eqlLvQtDzjY4L4bILqAUutYrlGUXV1h37aDj/uBOahORdn3DL
zEjBlj7bNsq8sOPc/rK+UbEhBOzd4RVzuI1gIxHgSie/5JyDbwqcPW6wEVUZ/Evp/rwWkVk6pP2j
t6w5org6mspN7wWlIUrrjk3VTtFlFU6H/MhnAqhpKxP2bXKX5nsTywQtEkqO1RetSi9GO7wStRWY
H/k3uxCsTlfDazYWCNwBbgrJ5pXnAbJ2W0HG69nSx1dqKDvZagFy7RHcU1uaavjpsBC6DeUsM20V
drrZZr7p/A8bF0jcbMg1QQftXHoCcrsOBsUn3aOJlJ4xW3LG6EvBL7pfzqXKZgMMjss3YsJnwTed
5i7NugtQVUx/HkRC+J0LKpmCTrCJgzeHZsUdXW33dxT/cDVxjpp8GzsmIBM7iE/4I9pFqNJvY9mI
029XyXqbkTNnmfT2HFFAto/dDhlpLcS8zxYlADfyFcsKHrVWkbY5lu2omqACwre8EiWBIKmZWR+C
DDb4dy1JOBtHLHMPuiLqLgdJPnDDXkeKWPMqoXTxqoEgW1PfUf6k3vn+TY6/KjoQj5lLXhdGPix7
bh2UWeeuMZTq7SKM367KOWPQOVbcIxskMMf2eHKuZCGRQT3jb7KTXx5sP29/gHCGoNyEZLPAWiwb
f/dDwunen3kvOTSJDq9wregqfLLkA1p0tHG4MsnranDrpS0I5Oe9tjI9urwad7AcR/BcZtpP6LeE
l1NYTDfDcb+VIGxrdjY5ZBm5xKQKiAFF9rw5xaYN4mVT53pceT4mQCJuWK4l+XreKdF00hxdzxTV
poPV4f0uVSTN4E00YuC+fHaOTwAcPlrVGUc2v+BwlRjJUGKKi9DM24UYWKOob0hOuXDnwjTun9Hv
3iDPAwhbDDfQZrn/o0a9R5CDdnVghP78UmlB3M8IJFkG7AAfK1h9KfmQDOqkAWb5lX6SG/a1ml9K
6izYn32pm2vvcDt+PooJSfNkgQKdmAd9fC7twS/jhbKvObV0ehUJW9yHKEk9Ws8rqmwo/6EyhiHS
WBusiPw0VW93b2KyU60r1Dl1+rSdUa8hAp5cjocAxdsOiU76xJ41eWv0AphX85AH5HhEZDKgaOOA
CSgUN/w5GMppFlD96xWXrphrA98wSrDzjFHWpcoFYkZsyre5OgYCupGh6SMCI0+/6yGXz756Odsa
fMkF9VbPYPvFGoMj5SeZLlyNBhsvFN104qB4iCGF487BgEdwW6A9TP1xd5RFK2qwS2leVwLCQRRa
8U+NreA2inbSvkgQmCIKLN88VqQN/bOtPGoIme7HvN8qk6QMgNroq7TEISCDFXehMpnfREKr3d+H
dlnMcDi67VgLjTt6Wp6ACGbF/T99zO04AABUwGCaCCwZUL6E4XA0PLg9h1NdFsabUqDuIcyKaX4u
I8qVKNufxacX3bON1mFWicdNx5MNdGBbeb8Cr5wmhop234A0ZDLRkU8ghpxc2Sjtn7ktYCQQWFzk
RzG9/Hq6/vspFcLsL/KaAeOw9nlo1woejWnDU8KIwwUy8zWxW4Vp5sFJ85AdOJiBLns0y4yWrSfL
cI/Ji4ElN6mqyL1aKv9Pavnpc3EQlgckPj38LALcB8sfJ3q8p40HW0pMxmeCWWvu5TwxXs7UWJpv
mmaXt41W38us5DgdA8u8LcPyHVgKOchnW6YGJPLxeEUBjyAFy+63daS6XDmRrseuw8wWERUUzQP9
g98AkzjC0odbmQel7v4VOrJ4eyviL2mZkxX6nhrERWtCd7EVYjMuYCRvxyADfK0vVVs23OJboniQ
fEF66IzWih7SPdoykyqspHd7yyvHx1F+Q1JE7FyIAp0o6H2I+Z5UV5iX3Ygaatyy/nQXTw2Aj1LY
4P910T8qgq+5vDHxUmmTqMCDBqjzxK5X5gQJZqydjA5aBtp01QZI7xKIeN+exwnnELSQ5/oBznIs
3ARWF7yXSLLptGkQCgvgHtrPMAGqw6c3GxEqsauNAwOxF1qfoIGVBMcut/CAVVUD1kJEDwAzqK/E
UAaGw7fyy7d5IJhTb0YXuJrXeZldpk02eUNXN5rMT1eIZQoYv5f+FqMXXSPRfjieYwqzx1XGn5I2
d6W63/dX+RAtVqlKnI162qaYM8cpg0N8xrgIk4wacJT8Vwd0UOgZfgqo2L11lVyMdC1bughskyqx
Ja1XM+0+4Dd9kaHeJ3L+F5kdulR/W6R0cJg2sMXPrLcm2ouQEWBy9HsOvvyM26BEoq0UCMERD9j8
Vio85vcj4VJuXLD70apClr6PYPRuSPCeEAYKRH20leRMkNb2wcOF2BOUGdH3DD2fIcX5X61czECh
t5rUrqeQ6MWX3141yxb3iK4beeDgUCyHQyowTDEbbElux4Qugb0kS2gSCaTgL8tV2J4aUgrvjax1
X3qAMae+jXDOHX7EsjIkIxu/CTHWL6tRKReMB2NZiCP3hgpVoi3/HrK/pkN8mmSvzrjQmkddDZeN
Hvnq4FoY5aG5TK8tW3LYNsqfFAjv3ubo0WEtA5f8IwZ+tpioFK3z9QY9rJspBMZKWm/yPEx89oJ6
Olw6Yx0PfkX5iYBfT1l3Sjqx3buEVfQl0gAUIQUw14y2ouBNpde652gegMIB5HSmqfoT3vg8sZDF
sT/inDEFPMlmAG18A+cfd59YsYMPhgLMBInxA+8QvExrq/vHki3n65eOoGemkbgAnPvjhM7gpOkl
EmDdx9Rsf+IpUv1m7nDUfyh8ZMRdzAwxwkmoDx3KAeLWNKODDH/jteCwCasxez6ZdN1+iCxkvgj4
N0pFdYbd2xuJZt+FowG4tGbZG7kscBFtns78I29uyP+KP5gLEswQb7j7GlmtCbsBk4hZ0C62f2ul
3vrSK2F/VznzA59E7zOO1dQuGxuSsHnJ5GVIBNEZbk5faa44zQ2c4PVeK74vjZytFKswJmO7UtEF
pkszounzd8bRiUA+AYMkcAI64KTMjFFP7qu4R0i+ntY00OQA8miTkE8Kw1baI822bT/XZJJyybg/
DeGTOAS/ZheFCIYCWyrCwM2JsRDKKXihsZ9kqGPFuKiOYEC0/vwgKSpUukLShh6eBybd7Qe0SaL4
1e7+xD3Fd5s9dK2Hoa550WKxvfxTb96oM7tCeHykvJX02QQdyecLWYgws2n5GNv18Xl6NoafH/Xy
LVMSbigQH8+Te/ewEQ1ZuROFdyAqkBwZDq6sqfxTYPIhwo2Azq6V45d7widgxGI9oKJ2xUHULfwW
VMD24maX2yuD/UWwVi0cWg4GkHSrt4eMt0C3q5LnXp0NgOP4HgNeaddERDglOvEvL/D2FyXMcaGH
uRJb6PLTA+vyZw7JzHDSvNSt3IiKTpbpE5gwTlmRy36ZGRY97iM3DciQl53uqy0FsG7/wlVBmZvT
fb5zW8nXIeh1pjRRPiBJeRV7DO733W6VVUK8gwnq8HAKOWRIAeONAs1vtKKU/f1ceCxZMZfA9wRM
IO22ZtW/rifm3CS6amP4Axjz41BJaODnVQeV+rNdaMt+xFS256m0fSkiD6OidHw+IxZGm9M28/3J
Xp4me0ZCV4dQCqTpBgf/7Czut4OrSL3qdUgMHq6K7+mVWoS7PgzBFELxarfXW43jqTx88JFBabRf
84XZHdq/ngaPoS7LIPJBBBW+pYSR42f/2gU4ux9W7B4ILhLmaM1nAmWok5o3bRNHITsxkCRinakD
tFFuyphGRtVgRbkrtqC8ZHqxlgnj4cjq19j+DavL2Tz/b2HX+BhDpk+FNW6T7jaH4CLHbjpoB2B0
ZwHjU54KBukZuQs4sJwDMFbjjjeKziYkI1NUxUdXDwQMVqpdnHsPQ1kQifzcJoIlhzgwf8p91GFE
en8MlN7iXC+u4h6jyLNxMz5T6K5dPr4HSK4nwZx+Q3ogVgsVZIuWNDsD8akqdtSERtr9UqB7Enws
8YAGaxAh2QufkGPyeU2bf5w2c7y0WchiasB42w0Z5jC/usp7UfI7SXdPffhqZdOuUylBjVoQmV0g
SqQV9D8ISBEuP66+x+h332I9ByhEtA/+VXaJ+LBZ1Dgw+SZ7pm58F1/SjllCWcyppDXrZXvIqSnZ
6DECMJkdg1LMbuPfqcHa8wCTpHO33Yjmihu0baGitUZhgX3haI541fIeK1AL0oOjh6dz+b7l+oK6
sheQjRXEMgz9bi6zciXLmjKNMwEukUxuNUfrrfD/5yN8V1GtcGKwxwmQ15DwNaPLHCLuqcbPRqcU
v0NWIFQ7YUtLO26ZXx8iSnnBraKsZSNlYMIBcS78CJzTJBbFpXggVNjzfgiaL0ByCF8NR+Dg6ic8
alIWpdgkaABX7cjv3ZUmuvfuu8LEeBssQ5QyaEP5s5s6M0LPjCy6vyXWgFB3S+LlzVaoMa6Pjkux
dvZaGAsK9GS/sYtTc/MGvmG7v4H2R17MSOA76Pkrsa8RyIKOQpqN6g08C9P+/76mE2BoUqd5fixO
pavtjHNPrQ8cVdfAy9WwKZVQ3LwZ/8wmxYhasJKHMbp+CK1mCDgwkmtCMF36Xg+EwTbYjP38E+LD
poEBiqoYag4KCaKWTflBmKZVd74HTwEuev/kcXQIuJEAbVyVBaCG3Npb6XyGGGJLVEb0KpMCWgxq
VS3MPl/AmcjC8M4rOFirs37C/QMGQq4V5C1PSLm+qrLZi6JQ33hSuRWFvVzp6KvCotYOvNt6I/dt
WjVJP0jGke+Lhi+ayUdLvwYDYZl2pSgbd70+DWNeIJ9e65Edeo3hauKVw0WzZziT/nbcNodC41jp
lDtry0XRdF+OJD9zqTxhgx1a868tKZN0bU2PKSHAZ7X6ZQq3QfblVNVAbOouClVaM2CGr3IOiWco
sE6oN65dm0Qux6OAksocO+BbIDctYFEqQ/5nuhyLtqD3XIm75BMehM4Twex6Kg8QBfxClgYsaRHZ
Luh6Rc+luezN1FpmXl++RRHI9awL/RrhwDfi9yt6XKe1rT8Q5sreFe1MejKdbTzwIu0CG1TuBTYM
FG+/s+ZeYn/++r/l4l4Pm2AmzFtCLfotHsfCRx4PQFHkyQb4ROq/FItfq0rbzAyAujIFJKjFkMeb
MQmb3SgZmw3jDTjkChI2FwclOV7OD5FcjeU82kvvXWgR1j4NBu/Y0Xi4CCpZE7N388daPjhXrkX/
DVVWf8mnUdWmvl2JKNxgdhQtX3O0ttf6Pfqw9UDKpsMnosFpTVNkLUEh5iw6FrKxGliIRLfseDER
EaQJr/yTzfa77iKSFbV+zZcSQeKQgc9vvst03sFZ6fW59s0pDReMrUcGh4mcuw38K2MV4Nz2Td8p
bphOPSfn+TduifuOOeDTfizFbeaR3BlEdQdnIFZITfivJyT0vn6hdR/uxNKKox1Z4M4hxDWMucLm
7KzleFPTZ3pOLqKQeeTRbtAY1eNz9EBVZZhK1CemhEaBAZ+ITjT3WWzkT9NyAfnsZtStYMF7AirS
nHh1gW8GHGkJacCJ6uZjTzllFi6Wix3eUAihrS5eTDeaFGLgAwG2MJXHOLOgsSisrpLwWKizZeRZ
uc5rSoITgQvwbpvrl1ZKSaapiGwCp21rJrblTxjRb2G7JZIE6Ri+FnRGy3mawrWr5cXcvtE13XXF
XTMloc2MtP7CDIs4N0uxHG1JjiEzEYqBJBGm23SZw5lcCrWTjiee7GBWJLLKiXX8MOEyMW+4RCum
JuiJyaloW56WX+a0KASu438M9TUF6SXh/cgX9A7aw4KstvdWFcYTBzQLSSYg9UJOR0AFvtGxbpDv
1i9F3VZ1+2W4xiACdm7uzVBu/1qGxoq5v0MvRaykZrsLW7oJNJPar6QnRxvi+PwEXET+GwVH54EH
vWKJvdaLw05NZrbAr9N7LvQaFfT4QMf4OBqouguieBSBa4UsFY8uJfjcBXltrkwn6uMeXrZfsFRa
/ETxK9pJugPQjBoE9rXGtc5//uFswmYSdWx9z71917Pmswuw4K4tbeFGqsUxw0va86aH8BJ153rY
D4/6YagcPpxNN5P7YMcrQufobTZHIhMm732b4QJKHs2uiM/miPkjJqZHDchRyAVxNetVBEpgXXcG
Bp6dL/bsu2hWeNrnCe/Mahy4sTtWRMI7RtMJ17HQjIMOqGH+5yqrM5E9oFwgLDa00+id+WVYuxiu
jifJ4s5txODDSGeEBiDuVe9yxbHi+nzq4B2ORJEYtQ/6mk5e6sYLd0brd4q5dgSP17tJLuEN7a05
joJbaIyZ+M1tpjJ+VU2Dv7OitbYaa/jIsvcfFPtkxz1uJxQTcAinEzEy5ScMcRDxXAg0xzZfwG1i
N/NCEjBvZtorI4Z3MOaBe4f13x0chbV4c3WtCa3IYHG6J0APK6QEWkR83jpmzuReNRupsac3IHVy
36HfL/KZM18XA0IScx4N1cx7A/qfVdLyqQimfHQwR0xDz0GZRu6PAw7H7+6UGHBAImD9lMaPDR5I
9B121dhvGszDFXV+6gzvE0wjQhe1PE0pLm4BS6DrtgbXEolwBfGeRYJqvkXSw/FFhRlHElpucWT5
nuY/F2xEJXoNaqvhkBeMh7KkQF3sbdcEV4j+EwxO9tOeJXOeO9zgbU1Iq2v7lKO6ar+HpeF06zc8
Y6o7bJSKvALFXr45R1La52i7san1T/KVRrr7ZeA/LdlzXC3/++0m8simkr2/pWAzVwlWGTNubI6F
8lQs6uewOgUSjWxtysnCbq2uqIlC1rwcIfkd0Sw/QQ2Oq4wJDvKGTgByVbXoQuqzupGuMsH3B9+6
xO6BZDL0mv5MdiS2K7EuWtKgq16E266uuxRMXMzp1i/aT/vaDmLKiRRduNIREFSWCZIEMSFe6/O9
tFkBV6wzGX8/GIO8F0kzQMDKxnDkE9mMqYK+IXqFsF0aTIMD9avy/npsTmDkEckRv9G/S3/+YT1N
lEWpvsrBDAlgXmzYQCufG/nQpd7jEIg3qJ5JcbmAcYIzEgu54DFvvbGhAcoNpI1H308z9A+D2CwT
qQFm6alBFiQCSfBMuv8Up2OJD6YZzMeF7/OQbjXGujJhmE8UE8VMn/Aj81pc/SQaq5XUaJYQyliy
2uiNxgU4OnCDOfYbcAny+TEpQ1DFdg8b/8ZDji8QMSkT6PSdueece9ePi4nhmnDK/5p0XGgu9kbU
aYM2tCpoofuGjBXf2plQACMCp3VqyZE2NuhO2yobf/mrFnK44Ci2X+clMtJNw7IEV4c/yguCO+PY
5E+l7wkEZHI0WkECjKY46UVCryI0p2VUcDcioUoIRmxl882d+yNbnvj9POu+t7DWonKP0RqoXb2b
W/sjVC/cZj7jp/Jf7vWAFWba8d4hfhWp+K3Jwh1NH+11krtFSpfkgALdqp1hCDOo8+PT/tW1mPZy
ZMXhKUJzxTeMengEfM2iNMH/0r77SS2ql5Y7VNzBAGOSLApx2Zjs48bJ8qHcONia1FwWjwKvpqai
c589ASmEWQorl6mSTamV1xHm6UgLg0fbEpwRW/xDBYHwFvzrmgqjPTdkGqfye+tg6wOgzvqkrE1N
jxBwgFry05KdaDNG4cZpcjfuHv9mgaoVWbSrauD0QchTCoewxUgXmc9tJSYshuujGNfUnecFXspk
LrQfmVLNW1pqg6D67M6j8jjBp58eixtZhyYOUhIEpsaXa4G1wwGV07PpWFYATBTdK95o6JB6g6Ug
KVdXaAieLRa+qOe56MXFuCAYtyHOK9l+3lJ/CGopcbC2b6agra424gk4TkYgTyUUoOFdkWH43F3+
MKvVJKtyzajcv0mjpHuuf06h+wgXmWHuvGmpzqNCjpJS1c4NfO9/Mgkj0n6sKzqN/DiehxWHGos/
rmtbxdqamylI0g2QKz/qgyDu3aqhqIJmxCfprWXzvs2jLvJ+WEttZaxuqpqpwoSoNf9+Voeq0Xh0
AFpmfCfjJZR/xHHt+LlJimq70Dj1C72co1LTttpsFR/Tcz1bHPh9zEnwxQ4/MlMfY2EEioF6Sw0x
+RvnJwd5FCYN+Al0cb5L8xJXdVM9vnS3yAaNQqS1HJSPmaWNETH9X5ztHbo4LaWzsy/w48RH+QHF
IseQWorTSFKwSqjp31xKouSs/VhygRgn2GPAHoSkHDee6+nhRYtU4hoUmnMdq55IwmEisvHCbxCP
BWUCDgQm/s/A2Yu88LyeGQxNkEWDihr6RSM7GMfifQDWf69Jv/Z56RGuAak+Qjkqhm7c19Y4CVZD
/LD2WihB/d1hSKml/sUcc0H6ukFQ5HBGR0AzCEdbEBOnnMgy73NS0FZ+QfwIxGtvifw3+4YhqZNf
OOxreHxBgi7EQLdsUysQGnASiUea/Qu4apBDK4Ol0aQdX2PPwCIg/tBbeR3CZRjnyjDc3DU1NhmQ
uMQaBceTjnTl4c6PxLs1S2OF1mvqebJkH+oXjnVMqlpcgjpcUwZYORPicdIonfpCSckm19Exapgr
RPAsTZdgp8e6fexPS3ASK2dtwzUL+C6wml8hTsU0iZ2zqC1RSVfPz4qo6Fs0uTdoQ6D7RyjR9H2z
xErWKCtpwOUOR87KKHq/Mds/55sSk1bRkYjgSQaJsnpzvRx2AmzMKkTTA9FgOHYxLolBB5aaEkp5
dX22709/lxnSIod/EQFgigQrW9u5dTejJ5WftuGTRripi1bHjV5xrcD95nYypdsroQibHyypZ+8n
2bXMcbu7SVT5O7GYm6sqFQ8r1VzHcrgbWvm8ak33dLMpeAtFCO+7rjFVBmewt5yr1BzIItRhTUAu
xczcuCegB43n/pW0WEZlRZtozNDShtI7JbVVftOiFPbYVKnHaKC6tqHPPG4JFOzbJ/vgv+JyMckI
WY/IsIvhJ4ph74rcQ+UNUxHVx4dVTmVlulJQuN9s8cdbISl1f/SzWJ9gQMjzeJ5UfbLxbT5pRECR
f0MCDZIncvHcK6/eKQHmk4Kh/+0Z+weOm9VR4ilAE7jrMVRalS3Eh4t9fIuhebpWfSE3tgEApGmS
niQhdlerJ4Bv7Npy1lz0aqnf6Pn8qW2oIUGO0TMT6pDQ9V4rk0mYvp0qP1HS9lJ1ySu6Y8KV2Fp6
u7heuWVQ4CEIVV20Gt0luTZfHL5quf9qXJnuDJN8DnPWi7tztYxNRKvjQUG6c9+01NDxdFMEg73P
0ffEoCfo1Isxqwvnq2o7k8synpQJgOobEtDco49nYDz8VeAv2e02FyN5cOeBCXd9LGPLbSLJTyRf
0G17JhAIq80OkjwyQBnqGrUdX4OHAZs27tpgICZhylJ8saLEV+uGw8OaKgssdyYbKOCLxt3bqI/M
rRs5+2p6EjenLM5oHXSl8xNLMIAJp5nnOo7d94DjHzHphD5epDkE2dtHa0Osl82YcnzgEMGgjAI4
cdRgn2KmnFozMD8qTH+PYY0Xc7Jv4OExET1dmJa9NMU+/cDX0jN3JIofnElBHx8Mdb7hbvl5xjI/
pkZHfPfFiflYyZsn9VYEoH7f2uDV8gYlG6+MjtHHYpRbSsGjjb9+7GIZyfuC71jcZMvjrxQCWspI
6XPgqvxAIu8KIdpdatpeEtx0yTjs5BMu4EJMiOvlbp7MvAgDkPh1dCZI38nfE/tzN29ir/bA+PRK
HZI92VWNH1WeJeOK/Fw7GdniUpR/oZEvNvAAqe51O0qmBfdC6MdId41RRs80MOOY/UhOocpa1GQI
I7p0QoORJ4j9iBSVnsscMRApI+iEvYe6/P9b/PwmdvmUHz6ggxwcPGAjzBhz4iYDmFqtPmUJ33Dd
OhJtFSftuX0jDPSBGJ+2AQwIGc/gWAStZiDbQ97z86Ce/71RwO+kAlE3sfHMd6FPqK6veItvOLP4
CZ+j5I3dskUFqtcxIZZTJXrPSXcnlDL9he/2n1sU3daLGglfzFyxxSDAEPWbaaHj+KVKirMcu8uq
Bijr/V7B33VXKzmhDLUF9RIhKDWv11k3T4i18tTPalNCPesx8V3Il/+8zXaUtflCc2LVYLbxEk3i
JL6QOhxhWff8DFzznxScGMLQy4lD+C/VNugYw2GR/odFrn2tIBrWkibz7DixMkV+w4QEvVT6Q8VQ
FOcYzHNoD6HkiSvoyq9RkcrONtxT1S9wCz62f+Fa33KQlPu5WXTLFDD4qHOg5oy9h9mA3CSPBPPm
EOivzeTgCCxZXs+TI4T87gyP5h97VJst6lENywP8pDY/oOyPDdJECXSXsyxqbU+2px4Yc7HmoKMH
Cv5nP6PXSNWYyHORXCqGj6DIQhUZvutkZCxlmUwhjfa9Nz2KiDXSF/qTcFxx/0djfpNmKUPu+v/1
tJ5K80Q597K3NUHXlP8jqUw3xHlRmzHKIe5OVKYECUQ/YMTtyoVcevO8wJQVrhZ5whqRBleRJRdC
S5JGqxDtOza+5B/BUs1v2TwSF8j4kHQpLy+MRNCPopY/UHMRE+mGfMPD5Cg0n/MOp8mnObwpNj4F
5ptIT2AjB41fmjvE0LG7hp9IKoljf/RO0+z/WrckWCOk1PGT0lWS2vseT+KrMUZcLVwZ0/v0m+Rb
9Fp7nHBYohqpyrztha+LtvZLM/ze2z/cgtv2qnqdFh2C/LxoJqNWToRqOISjpC+3JC4KHjCIGpzV
7svAjFedTxdf4wBmnR+g9yuQJIEfnxEFwyvVti6n/ZwJu4iwgjCPUQZNjC2x4o2gAeOGjYdzccU1
Y4tCD9wKR2i7dTYYTPOF6tXTJfg9ADcjQnXwuzJWOjVdMzrmkIjlTn2nX92svC6dPYJDQ6KM2que
a4kdnj74Mi7L2AvbpJxI3nxHZmb0bC4fs1tRuACTjNh5QVWsQXgl0MrxigZ+akjQL91oHSknzXy8
fYGpV29Dv5OZ34+a3kRfd4OMnUoj+fw7t5yV274eDh2vexue4Xp1MYMxRxmAjkVul8DKn8WpTt/d
GFoySVdseiCxKWFIxASzDnk/YsSIBdzD8FKmB/QuQhhFcYyvQqd1zHXzN+z/oIx+bGU02xx+Sn4r
LRJ8IFPHeOwUgU9s0VX4dKgglG362lVtaHp3rQBE1gOXfPMPRQERVNHvkKoiZuTF/KV3aOwLGn31
P76S906CyveObbbzGrVOBCXr3RC5emBFB6C0HbRp4B93iLVz4rhOo7mIcOjfvEV+eEsYo/f375Lh
oMmwtlOaEz1iX/jwK0T7+PgeeHLQ6fvI7e5tpGBLaCFtYjuNd1Rt+NiU4vMlUI/i8ao4IMcDV2mM
G5pLrJPjtkR7Q32fPdShKwb+IHHccnL5XV6uGQ3s2hexKwcKRGEps0zzZDoR0nICDX/6p3vMblhZ
LdhHl3WT8MjGyWngFsxmVwNOyFx56OkXlMr3GWTNNrxN1CKEMPqpS6rlmHc+AulLZIHHfZQMjmmY
ebQ+FmAbj5ER/L8skEzOlyJ9Nejdgfayd/sVWap/9nm4m1vLOIKmasXcPCzf1iWn0bTKnl81dNNP
1SZgfxSvfZDfCPLGnRJ+FyXgdM2d5N7P4ykiV+5LVdUka2zSKDZaWJw/XW3q9WC/LUPv9Y18/oE4
z0epjeVyqsjuEZjhFUUExpdJZdENNAJk9yZ3DM8ZX3vste1x68ubbV2Btw+3j7RAxQYBrl4cq4Rb
C7tjpUmFZ7jfv9Dh87bZA1oVEEyVMAE64+yxvbaHa/XyahgAON9XSPkbiW0z9x1vMkz12R1xLbtB
5dZMtDgx2gRDslLzYtxyPGz25I4OwNI4a/TZVq0u+Bl5FV6TSuFHdeDcJC3VMB5Aq0TAFeT8Qjbz
5j16qQQOBCZAkY6cyMp3t7RmSWGvaqDrGtFdaANFFPED+vptqeGa1RiszcEzTQ5HDwGNewtJL4a3
WmxCa0d1VHitLOQLo/uM1B28E2mrJn16bxwi2dKmaBTkl9oMrfyyqbaV/r34cAmhYWofs/QzKqdg
wr/d8z6heQ5UcXZbAIlEbqW7XzcmVQJcwhrR2III6JYQ5im4A3JFUxLx2851ApafSFuyf5e5QoaU
J8nt6GQGednLESnXapXhtHUQGZ8XT6q/XI9JhcltAqJDSsr2uyO8J1evlAFDnQJWP86Sxrmm+Wdi
jcldodeoPWeKTnN33tXSOiueLuZ2eV/p4SIKovr8aAPcaKdsTRkDerVmSeb/nXfgekdlAgH7Z2LJ
1Kc68YY1Bi1T7jFMuT9CaHJNazB66uWvjfvVGhOGS7WB11mgb1I2n4dH+KsQCGzDx6JfKGU8LvGE
EcCcCvYLapO0InZHfd7GRZpZ42yIax7o4NFTJiducGFOmnuamPLh7S1APt7GbrUAzqFGLqEBllwF
LriDqdo18xV4t+ZvFGDxrWwQ7EnThjJhmgMvane6BZ/nMFmxVpzZYmBAlrwvvQhAVqcQxA18yecS
BagZspelLTUzPBzg5HDDhK3K40RuijVddUD+UDkHfRHnL4dJbRHOLI2j5oxar1tIcu2aU6hxO9Wl
KOoQMLDNNexCjSy7CCyDNYAw15qwIz1EGZwJCKeJDOdMnRtQa1aPIXnKMxXlG03pJ6GfdcGo8TFb
4hc8IlnJ18E3kQugatxcyPufRKG/tVuJW3+660J7DLjAC4jeawpIaoiQ4dwZF12CTgOAwEdrCQtR
iFUwmYa1UamRidZ7mCOpm94rL0ZHZBipORh3HN26wjnGlVy12ehsbPvwvfSDpMch+8F01NgU7uEm
cdNNg8X8PKexVAMAFSX0sbmIHyeuP37tXlrL4SVCf5wsnc/B4v6r8jIg2epBmKop/o/okz6lu09y
XZnp0mGc9EAXpsgZ0u9EWcWbFgXUVc8ITEBrJ8hYZg+5vp0tDikUYJuRbEKWEAppjySWOz2PKTx5
+pBda7VWBqkIvLA5QcucNYeolOAmxvSSUWgsdhKh/H5hfViKVuEQFbVWvFxePJ783Tvx6bsypvKU
M1nUS2T1t6qApWKAb/eNdFLs7Oz31rG0d9niXoXkJdV6sRGD3I9AT79tIzTbulsuLHv+1hfvSYsG
vLNL+c+p/y4CqELTWpY8Z8TyTL6sNB+74aAWztSDs2rj424KsAeom7/zsbLPiCjGgMvVstrxL7Q4
cFohAXH/lTSR2c6c/sfqjYxAMbdTtFr6wC8NwGl7L8tSHAG40lnEBd4qLjVe+Iyf/IygVAtAGVXx
ET27GoD62zuaRSLZECdRP325XlEJAFEQ3RWL5KBDc8+YfzARE8vYDvONXNV7N7BuX7ifIj+9hjtK
Zfs/x4sEK9m/KdB5Ui0vzYk3LXqSlQDP2FhpXgWJIqfdcfXOZGqVvYgey9WIFwkgAGTECe9M6aSL
t6bhtLpxXOHQu6RYJWYMGn7EISoA6lizAQSOap/iO9fGQnaGnd9DMUE7631xtwX3CLJ6hihbXki1
mnY+WIjHXntEMy6s9ATFhUkTEP5arl67ffT+ynn6tBQ1fGr/qjX4D+MjpaCMQUxBbgLs0lYaDazj
48AWc+DQmn8oSaBMY8sSlg5LTqa9SugLmB9opJjJyHDwy8ML7P8z5qMYhAb2gqkacaMoSbYrZusP
FVArTHAE4tI2fb1t+8IGTNmhmBYcKaI/Ady/LxiD1swsbD16ohABM8bhIqNGhnaf/ZrseVHbykk8
4JAuPAaDIVNGE0lBE/93xaiDX3Aec+4ghTHE+varywlNbv37SLDMBDIhp91f/1F3BX7SfnDB69CY
Z3eZMkBSHRnjgRE474c3pzPRC0s+0O/QUMv6g8y0qq8cwZsKyswpFppb1UPxd31W1ITx8meERSk7
lF98TXdU3IuE+TbnSFGe0FnlY+lQuS/wenB4vCAhTy6WA4qsj1QDs2ETeul1i5E9r9I2pgSWoJ+w
4L0uCgxuvB9q6OFH2XjsOBV77wJknqkA5hO6Dtlf4aqaGsmdDOb/CycFPz1yqXAsgV5XAS5AYFPI
xsBlL/lkeQVUzLOSxFdA4dk5uwqORPXN7iPNuLfqVpIpTaq6aWuAwwIO+yX4ydFGhazqb0dP9VxV
1yIt9JEn61IQf0kNpBdDNHwfaFcDn74495hiOOi53ownzad0Wa5vixwbJHwTn4bu4PZEOkM+whyN
91q3+XD5UZ4ZOp2p9T5MGftwVW00fSpckmFqNW28MP+aa9Qbf7bthI9fEoz0bdBjCrmzt9gm63aK
zILtMR+LBl6Hmr2f4U8OPMW/ZP3/NxFSiMm7A6cnk2L+jH3f7BPPy6ND9nuxveamxgrMYQgrOypL
v4D1O6Zxd5AqIvRjC2aVyPlz91h9QpSJryH0ZqAbv+XZf4rsA+zBTF3KWlzLLivG6JILisgqPaIw
GMjdQLLqKLpbHKNRpDCfn+n9TK5/kGMBncb/EsDXnci7yGHjS9NVaQRYQKDXkZ+ZlVuNsTFyw876
jNoEfN+hFWbYvthtToBjQ9Lwb0h2r3NQr+vWDrziRMKOwr4UH97TO+Eg//565KIyr2JWnA4fgAJ9
6a/XPKxqI2Z4yq6ixb4LpTpIxbWe0sVYa4M6jejpbzaG+BczEq8eOA93JLb5batdMdUsJdE+RzWJ
JQkf9rFB4lq6bH4DbDU9qxGvisJyoSkxhBJWyvliBhDA6jzuzSlpEM0Ja+6/teviaOUTEE675K7y
lC/ntyxOpoZCkrhFxkgdaYe6qgp5QyVwDnCRCyHvAT97XxdESoaOP9pxJY6dTQkWY27o3UFM+W3x
s6J+W3a+T1wmABOORfCkrdM8ZCIFUOJjh286kLXS+oTMzImfE2bMA6OK3bX+VYZ95K3OqoXUc7kc
gxHne26mwfnDcg8V1t/0oLsrg9QNZzYkKVsOlWRbhHYljzRAJr6xEf4MG98tJBiNTszTuT89cXQn
b4fum5UdSu2S5yuRI1sQeuCYypGnPRKCQPbF/rnvYM1lJAxFYvp1cLj5tyNsVv1MkBaH/ZGguPEH
skSU8SgXbsdjz+FpPd7pO4F//36+Fk8wSVJ4uu5Ucd+xBgdEGuyaUmTrIr98Tg+xVHOLSb5xQBwB
jgZxQFvKkESmeUj/LOr4dN9rDM7meX063gf/lQEmcsF5hlmHUJgWjcK5xQK8M4E9AUqXAUnhF7Sl
WQC24xT3mvimfF+vT+sCLNta4t4jyqjbVHVYMMEA1t1nxFMpW6ZIrfuCtJ4ufC6cOpS1M35DkfCh
gBRAJ/zkZMCvr19DGPdZnSQgr8zyWmB+K/2mjT6SQQV1BMmgdtfPVUsrtHPcVvutQs0vwVd48kZG
G+6okvrqeafmBHwKLOhoarSRyo/0lEWsgiulh1nP3TgcZ/8udhzo1JN6UD+r1ifL6eufOBnDYVdU
g8MDIHp7V5tUZpHnE6+Ogc18cEjDfxkqIs3y9rt2Xph3cGTAy7/t9ojzLcBlQcLTU9yWIF6RR5N1
O0cdgfctr4A5/LFL5khFQ8DflZoaRQA0CqEYGGI4gnTypKQ2X95TxJOF4gpE3jQwV7CVPb+qwOXq
pa8oBbgdJ4SHNHHtXsOUIw6Aa7nFyNsXDOcxK4OaeiUQtx+yfJza4zR6VQvnfVleYsQ2rceWaWel
1o7EUSvcuntJfn5PCHAAFmeoTBcKMRqPXSuPOGqtLDCugAhEjWx/S/SPnw+CBWtltCt0Ik91pm04
iSWTvju0uZ2WpCijemZ+yir6Kn2JJZoFxRT9V6UgWt48aAAO5p03TRWNLAX9wdG3bhbNDR0yOuJm
wGy47QnfPxwnBbHz+rje3fW2qx48AEqcbCneYDkx0f0apvmVA92hdrKJFsJHd7y7zYmcKTXXDlwM
cD9fh20RnKtVnV0IS9US/KxM1QGQzICExT5131alYMlYXjBthPCm0bvgjdoJiIKBjjgUsUSJ9Cd2
XIldhkotGFVFzhwPpfaaNJL9Q/D/hEuOtlzsiTA/scb4Z3hLoC88IhAVmMxcLQbHRJjaDb9awWyo
6ot3QvbIq32Vaf4DOjxAK4IHcpqy1W+JMlIsnhzF8ORfJNoAwrXv0zUMIPMVHYbUeh3rwoOKCFBj
Eq1wk31DvA2eeS20A2yWWxZmex8ZhLL1EvYOBsHRs/BrUQV35PzBb0QlrawWG4zFC4UuNADVftWS
iWzyxD6rN58pnjoAqFx/OyI8cA28Rp0V9I3oMXi+iWlEV6CPbj5d9BfM+YjT88WMXWGOY7tLGJRr
eRuXjgk4j4d1JjKvoJ16bf8cVYx0hB4O1KWZuKcIHud/IxweCzKFyc1Dfo9ACx2Oqwhg02fkN/84
IknlXRxoX+PNeU6GE//+Dm7yKMSqGsopq4f2kaC1SgJJrd01jHPVfwgut31X2FBRvSGc3wxfJivL
fHTWyIySpUVZUUA943wEENkqSR1KCDOwRjcyEKkZL5Sr+eBGzlfaWrsZy0x8gb0KIDXkTHJHdGCN
jPKnTnVxezA/01HqoMTkE2Xgu4iyBsIKVzMn3iKTo/HBsd/wUU4s0U7ZZFIAsCgCkEQBhGqfXgdQ
bKPDim/zSNYpXdeV6b5mzQ9FQaysW8+Mo18VUaf3DSMImGM+NufIPSnKQINEMeZnxiEi0cpLEg0D
/qdeoz6MV9Y+Ynl3E2zl89n6rdcxypH0KZIA8cnr0DPwq0Ficnb0IRjBk6wxvOcYVg4KrF5ju3pR
n2xjq/vHEz0CGLhAgwMzOZK2bktCguC7ClWT72Efv10HLMSTBohJMNrUm6NRRRA7kG9Ir9SQC9xa
vPQ5pNDmr9Nwo8xxr35Q2Tiv9+BJXDi9gnaOobd6hTBiN89Y0BvomIVMzzPFgXv+cUMqz8vD9kXD
pxJ5cDjAFiARYTmAT1gKogtgnZ2228Dq6QW8hr32Pafji1cJUTEwmXoeML3I5R4NYIJBVdwGnHSf
B9XAX7AjoU8odtQlx9r6DnnVLC82fnTI48Gb3/DwJ7gus2aPd7s1bGAQam84Vp3VcGgUW6loQBZS
cTFoQcRdxtApDnciQnHOUpNL6xdbUehz/8sKbrkXJSQw4wbFA8Lq182MOx74uA06EIXVuYje8uBa
cH1QjCD+YA55mIgBiUiZGqloffXwXTQ81VqWBvgV/Mb/TYhZk/SHSv93N1idXlRiIATeDuQRIdeT
42NIBUKbzVxWyHpipH/HF7kn5EVGWwILo2lXVGN1FurUmhQV9CUr9l7tPxnoOQpIxL/eNFJa15hc
gxl24DCw5gsTC8XKevbnrICl8xV+qYSIUUaPcwe3kfDx1gYcDQeHq3SeAWYqOcOtjmIFPcBKi2Ct
rZVO2dvwD7CBPUu9Nv4jqQxD47abcyZUqTx+85oAKNrTNob1qMZrP5pQigAxNZzPYffwq8/e37LJ
+8brgEaHtmGAlnMoYklLlUWukot58RK+gWnk/upl4194d6wBXYu7VJNc3s/rIz4Waj3PqpbK0UfV
wiR4TFnRSYjFR7OpeWcURicoWvuQ2NyKITw5uv7gIFnDew4l8BBjmqlFiWUh3nM7Y1qicSVXUXB1
dNAb9qvNZ8WkER5zFiE0sRwVXlZgeeKnWOX8eX/1UoSHchvWWb4rIB4CEAB/+cm7CKecoLEGPPhX
4+hMPlSNAv2dqfNpFQ9+p5CgEIINZhrs2WMiHhZVcYX8a77yAtDBBhG2V0GtbfCI/xShUlF86wPK
yaJDBBbDjaIUjGf2Icw9xbVXFbLolbN3eAzkBlChQHCHJtD4b7LFs9gHumBnAGJXutSC1X5YzMTv
gXvl9EEp6i1r3qKm1Gg0p7rnXwkDKsBlpyRu9onOl4JDUP0cIhLfiRAYenqS4H9BrlKYkks3PzVo
PJL+BFUltK3317hzDic4w377oV9G1CXklegpDX5QQXTrr1l0hHcYAXuvZ1F8j5QBWTqQAh94u2YP
817ZRYE+GZd7ez3Bwq0L01e52txJ4GUNim4lCH48eBBQFSOmtzg1dHaWuDi6eWoMsmAFRrpui0f1
txKouhnTDyLq7JrlhoG3FQQQB8KBjSphcyllUghaouef8x8u9pOS6FjX9TMhjKiXhFtzhTgMDMtq
bWxrJu6v/1jsC27k4MRPFr05hDU+fdyK/0CnXPVjyZD397nY4WPfMMg424Dt7dCE41PVZaKdx3sd
EYFhGjIq3x+lNDS76dQNlcTeOAEQl7E3/vKJrBkZRq+OgVKnmXWTTpytC5Codn+9u/JBLvywV6g5
nbLt6Coxx+7npytUmpzwF5jEZ0Zkw+CO1jBSRHhRFJ5kt8w0RzVXHE0Us0gNvk+DjIJ4+7yPG2rW
f4gBHOJiTdiKsA/0jVnEXFZJcxaRdIWN6ab1lZIRd08uHgFpjmRl3dD66hvFmpa+O0D/JS8gNByy
oOT8FO+SlIEF/03gh9f3wq/GVHyz91QdTUD9uzmyuUMviOoGBb4uLIZmYj9O3ef8LSekpc6mqfg0
OCZS9KulqR1vwVIPxpZz6eDPlwLvPLNlIhFitKuKTmP4gL1lMtCG3FeApZA0v30kyIpRHx33Ts2a
DRswMy4MzB/EG8mUe0XfDT+JUhxrZWIfXq9/9wjkRefoHyfqvxwwfR/N84ICnI4qdfw+Oki5Gcsn
H8pkVGItwqBJBqQGpZNq7bDaTCPtUsEp2oqmQkh8u/ULDqV9iJqMk4Mcdsux2MK6bY3xh7LrjmAk
4meCpZJGLRM6NNlWDx5d8MnN95CC1zqaKiNh4AIx2c1s9KaE8swu9XHtN2I8eNnmNAn0BGpA5zA+
9CYrl6dGonOwlDKJcoFelOg0kOcSGvnXpwBS3iRHeQvAc6Ms9x2Xdv0gvQYqbMiiiDLA8sYyUYaf
Jrvjy/GROOBA82HehVvrI51aDgLvvwQuci2V/xDvlXp5rMkm5syhSxqCptmhkATL5LRsDuRxI+2o
JrJKhWcWNKsrqinOwFvtX3csQmEbgnIeEPzuE5UFXynEpEKmycfS9AKfJb2Rh8/N61Zfdp7pWPIp
Vh2bYhvLdIk824ljX8Lmik4sSxNQsA0hWtYGqDkuzHeBVsXkpPBpM2PU7b5HQ2f8uBHHscyRcQq0
6SH1pKUj9tarkSL4dNnQpgMPbSp/fvngY2q7hplWX8YVXAPRZLpH3Mn1PIcbF5+ab4mSyLHaz7sJ
rxSqVASDDaOgugxt+b1t+6MbXdg2egx6fLSZ8/DIUxI0EiMgmnat4XsqXKrSlA2WVVJvJFBymQ0r
TLfJT/XTc0h62T15JZQbRJBeqNCZM0hzyH4jRqvOB/mUQNJw+x8pM98M6r7yQYBnU/91VkDuvqAO
FJSpFuk9qFl5m5kK0XALGrnJoC7S0oiHdf0C9FjQelEUilYz+SSuA7c3QJejgOvCKWtQaYCE8ap+
IY+vpmd3pQ2/PLIqN8V0xcorb8+uouZRH/8AjH/DupCYtHD/xoH8CkxA4uZStfPr42m4z5cIvTFz
lVKg5QZcPHCMDfyiQ/wuG34LTTFzFi/ZDsf303fJGBMT6mci9jbCQ6n9OCaCVQHvJF0cQDmsfMQ5
O8OKM26W6Pl+gUK1wqk2gnUkQ1lGq6RtCEir7bhDRgH4vvMoCgzodb2pJEBzut3iYdMShP0aVaGG
lnGrV4xsCfU0MSmAWlxfZgbPTOxB3rbMKxJRdn3WJlkZdMomaGJiNz9Fu/Ck/+G8e8WR6All/ri8
+hJwWdFVy14wFNLcDt0/svRbiiH1wZcfxA99Sra03wujiS5TrUyJtxLK/wpwVP+1ILyfBnM3+rbP
aykeE4YrWv510sD85d6bU/Iq8e8kTvcCBp6zm1vvtmho7YxKl4Tq3plwgPDLbq//nMbLqkLKjt1h
irpv0r6GMAOlx7qwN/TKQVAS4Usm+J3y2sfCzVAxNCtGpnyd63aF3dkD0FZJ1+BoF9OqVFV6DfB2
5Io0CLm3Zi9LDCQ2rE5OIjKBIa4+mXLCsDPt1LCFaiunF3KHJk2UFVfXHxrtj/kDyjZUyDa4I7+z
98/VUTwsQpDLFMEYIPatc3nPMcdomZZPJmjysXpf4mmt0jtL1DXZ9RjWE4azQ7aZu8L6gdofdZPH
hR9wBenc5bK+3LJL2OOTuS4bhLi3QKSBI12m5fNMgwk987vgE6j6p2/FUp6ls8e0S8aTBcQfVmWq
nmE3jhILjyr6K6TQNFewrXxeKMTvGvwf/2ly2yzNLJeeYvU14NVqfSTITY7jbS6euLsltscppwR/
F/9whmLcjcGrvmq5KUC3WktfgdNTomU9hHWKEtjbIu0ZVijYpqDgzXm7sO1nQD4sdgYj/s5L4HIE
ZAuLmLwC4TFmWnBan58gdRJnkFnHxFgoF4YTlefe0c8uYePZ8weOGutrN0nJif8uMHARTtxSI+gY
FQTRYfdUMzplM9ovHXjALL2kKdOPPutdGq0KU8r1qJIhM7kX9RWISNfIYbsgfVvmWP3oMoxq9971
bjIC8QNUKtM+Rac79bhiPKqWA6giZ3kUscAYWxYFEUo0zDVERimspa4mNc+K02n8Yf+LCTU0X6YJ
U7E+1r6IRsTd0Gx4nsN9BeLU4BkiNUs+9MZaYO6jS7CTChMIFsGMVk/9R4dzU5PoOWMLEeBBy//h
PK5QHl7T8r2BRhq9vQvucNIALCDWot0eqvLKzxC6JJ1aJ68/19cIEpqaw4vz3dUNRkM80ptNqU23
0gmVpPcxLV4Stji9JIKBy9aAPB4TjBBQWXRYocwH38MK9wH4BmohW5PfDYIniuJz2EOo4X6wdHVH
JZaLFIlQf81SB9XjHtbd7InV4zBDJkQ2tr9iR8HQJoleKZ+RcIVlRGU/07MLoLTEj4r33/Fqds5M
nfz7yGybS/ZVseMB2zgFV6mv6+5apNzI7gLkffUPKCHtRLMQQPvCdNFYJntOgR4aMQdxZXwWoRTR
z0FICtG+g17tW7nzh+EhKDZwKkMQy68Ke6Iv6Ozxk4jZX3zmlzwoffQBk1CPFX5AO1SLncdoNN2i
/J1JJXTgFExfE5dP5iy48cxV8RPm3OVuslQT1KntWI8RBYU+AIdVsl0Z0GLL6OuTyfVzdbthfl1y
ste42np0nXLQPrm2BhAZ85lKx/z93aedwIfll7IA71T3nxc7QpEl5TuKFF3Rx+c+z+c9J7CrxUIn
6rfuIgHgckkn5pCrPZPYj27duMztQZqjQMsam8gWdoEyLNQUXjRTrMq+JlHloCVheNRlQ9N8Wb7w
jbI6rkZv2UuTQqxq9OVIzccHHdxmxVvQ9i6T75531nGhR0sxkDi+j37iWcJ7k8e9lrCGIjwaox/Y
qE4x0mTRIoJP28pXxp3yOEEvP+XdLHnbnIJFAghploPGZrOdI0NFssS285z3YnFF5HteoDd1wFW1
J8mlpGzF6yGkv+u81NN40y3kuEUJXF1Huzj4x6HbW3ya+UEdyB0ylO3iJLSZaSqK1SrLoHuZ6Nje
lI+Yrq0Qv9JqrZ3d+XItt1RmUv8xAr5UzGdURUF/HiOi+CpmVEkbaRvtpc/EefuhTFaPtu41w3NI
Upqy0j3Ns6jQC23PUT6UYRiBT4pB8NW6iFQqgJTrZvkUhzir1k5jpF6mB7MPCsneKzYvJfWeYXjR
P9cxcg+7uJq1egVW7RoxGxtXtPmrosDUAASdoxlxKHOECaEgVZG+Dw90FLjlh+w0S5GPc0FAw61l
Tl4Itw+AiIGlIflQjWCPcskqZ+K+bdEi4vWvmq8vr6s8mMEzRCV+GzFLPXJ0+EvURlu872Yl8BJR
nAX3Bcp7XwRW+4/kTsBBe/GL5PuvyIPCCgf+5UDszmBF1to/HYXp9yICHdo+hUQyFfzoRUB/HLPo
lCrFd1J5RYwGbvxhqMKjGpYapZbO/cLf6Kuy1sTWlKZ6cpHFGnaF0sr1fA5qIvxtX7tQvCUsIKln
7THmvhaTQkRdlRzymZSzzI6roYSIRreJf3P670fQrtJwAXOugjoJuv/DcsU3nME1zUW7gTFlHfAJ
6FclNxGn+HGsZsIKRrUISQkcNhl82aUxAO4KG9MDFRdDOGB6pLXlaViOazkr6mI+6bEaUWbLvOz1
4Ah7Z5UklwTRrf0lHZwU/HpDNPHQly8u2ZSd1KHeqqWqZKybNLZ2VwqyF0nVpC4xCq2quv/R1Cqw
3NodV3qf4wNIMZN2Rs9zuUO0DA590+zgm88FPD+6fVyKjnYcW0qlT8jExY2xESrtvEEOjcU71QgB
zD/7i/K6qYxEJl92pCBFWQB3PIdMCLZjTYwgpO6nVtdxTfmh4PwyvfNMlCdFQSSaPdC3x842VAL0
RrkqJ0mQ4SjP5+fAu/LewMYZZtREYFZ73524MX5S78AngZeYdrY8iEMd9zaWoqPfX6ozg54cBAEE
k36WaWbVgquTqccy2IJ9EngLiqHzYOAVQVI0gFBjfpyRpvbNOdyi3TCCi8wmc3v+2oOi6dr9K4PQ
qRL14QbslemNWKqsgqj4SkLRLV+OMesB8rt0EQmlcSvba7FInPRBPSAF/YuLF60h0ui2KNdagQdI
7NLTHQKGyka5WCai2JtJVAIKaPGDyzW4pZqYBGnIYEcovtPK7jQJWvefLHzP6PhABdILETA77wC4
QQNY1hF+vvkJKLikdj0xWu6x12vraQIypACbdazfa2ExYeKaPb6GAFyyVvZ5ZSWSRZqGt8RHQWbm
uP5x8UedxE8G/px3o/F7+1v3xesoUYYPMbEkMDlqB8hHJa9NYeDaHjTpd9dZwcbU5aa0JvI8jmrV
x0S1a1eIhgNEu+7PLWI9KB5kY9rLKY3KioBpdxSJSKAT83I9DX+ff9am+aEabpU1b2HF9ul6BJD2
5VydMFh+eb745dowePyw5Vncw/QdtDTL45Y08thSHmRhw3/zjIMi8+CQqe3Wc1ajcpaxdY8T1+bs
NKVbHmdWgtO6mbKdnFof2Hu8x7MyWxsiV5aIo2T9TT9SS4JzuEyr3746JuH/a/C11tD+9z1nmN+U
t/DLdTZFKdkpkahitx9YPzi3LWtOg6cbKvUSBgFhtHXZnzfSvDI9qREAHMQ/MwKY0unQ4AJIAQfO
8+5ExLTehrcAKBHqgw42s4rSdA68gycYvfuL+FpRmWWWUUsSrt9xBTnY2ewsBytBehXfX/KLctdo
tjvkHFqEn53yc8Im1vHBLQgij6WCEU44f+R9AOvmdx+kJ0dDAA0hidCE7AGWmDCtjs9TiH0eqoHL
QF1nIjPnicEua1G7loIO20hI2v6SEx2bJQFqNT5o9bYVBqk+Gl0a5KAUhS49tvbvO1Y7740ANQTN
DJlHAQdLj4y2lOhiF9H/RCGqFqXKg3SOb4E3Xf24/sFPaG46zFb9Sff1Jz6tCs4TenR3CZUaH3m+
lQ/kt5skcqyA4ZCzPNCjKxFDWgh52rp3Te8YhVxcpew7dM8Z15HNDv/guh2NrArsDTmuPYvBr0mN
pxlK65OGQiCqiNDEH9curz0rDfKW6YgrHCRFv3056f16xotTiLH0gHMNDEM2fox4s/l7BAuJrAWM
o/43+1m3MtXMEmw74VqeSOnvvet8zXoGZtVhkGuNkNwYIBWQwwUgZABeV9ub2ptqfBzOsK2XieXc
mZfevNRXKifhvlZ3r2rDH5boQD3acfEPWOrOWqF/U/UisCWVDxIt7i0wkFomIKwmtAjNdHv1mvFh
FaQ+IUXix9EhSbHtpj5BxEaFmvq90/IeSoKk0JD77/4sUgExT4vWiT/1jO30Nn33q8AljMWt1oon
6FmyOEgjSwlSnrPfYuSJYOWXbM00AS00vTm5pX6VcP4MbjQLZS2RC59LDc3EgUCg/qE7oPsEPqCu
sCMQC/QfI7SZtWsQpOhOWmy5h5M5dtCdvR6jnzAOVtMOR8DjGAkjyWguZdPl39vD+v1CtgVnS6fN
loZvXfgDzLZBxdzvTpyZAb218jVMTl267wOuhfs1ocR4OqM9TGE61dbiaQPN8r29MbK/Nn+9ICYQ
alJWsMo2w3v/dYhXuf5qSPnHIE6NQqRykwcFTKKfXEPN+Z0PJw1pyr7oRh8N7PwdPKuLAYSeTZrZ
W/7Awm+C3Jg1kejkFkCKmcU7hUQZrGgbRs/DdVuign1/LU0YPVeUkT1S2PppMXS76Ui+ioJSJ0sP
pGnXtvJjjW6hxVQ2y3KoeZPH2j7ny1BY38UDjonLpWgI00/Jn8xZVOjM2wwpzgZPuX4NYYTsWYtQ
g23IXSHtp+bZONfV/jgnj5cPPKqHXQrA+Cw+2QcZevJ0Vj40M8xGzYdiq65dmljU/Ioj/DItM32+
yKJMw4YZT09eSO5WvkhDbRtUPI9VdcJxLx6Fh1XC+yzZfhKcbM8ArYSqshBvrTVCj7caoUpflxwi
lsbzJ8qc7GSN0W9677jwqvE5a+nWNEL4G98fWgbM4GyYV3GxDQvrKz4NZS4mM9qJN4K+7pA8l6zQ
kkOMeyy67wRMa/VqudKlVCpJzYqX6ZD0Nl1NlUgNbWODxrKh5i8D8kaRMlXwBeEjanPbPn7gTf22
QeZ2D9wTczJm/962PDMG5tk1dnXAbINJeR+i8jPrbINT48+SQE4wmsWbTpYVcbTk0Q8rke6Yfque
Eo6r6O64jl/+88zdNhnWyxhxH1db89mas4WKb2nq+69rheHEzg3KiQBeCABNi5uUiOOdywlzF5+c
Ig8cBw9KdKMFjWwVQhLeXhF7tJn8IIUvkk+vtTFD25InlBfRSZhGReVRcj5y+4iUBhYNCzoV8cdp
phekYAMrnMUWgT4drWaKfq/HhdIXOe29WXpyXW1ZFt4BCcPEZhfv/v3lYx24y7kyB1BQxx5ah9gb
2I24lGHb757LSnx4qjWMSaZXXZbxrta77XIwknl66pvmIIYlVwfkp0P9bsna1yey/X1kdXTKB5Zd
Y8NZmS06UNqOy0zEg+x9HifToX8VeqwBnRNLoRiRwxafiYNc147VLIOegviA33ZcNkzjsP3BGeYD
/8MVkiO+LUnT+ME4cWtcMr1vzaig8z9By1GjAciMHA2kDuLCmqnRIQ77laFaC0x+CqxPtB1UVX5/
0RLO5EO0AxbKJjdZYxRBDExEWD+2gPCW1y4Wbd9jN0c73xLTcZgcG4zqK58RpEGdwwAoehIXIHOt
bwFbtowj9BeyvY7X2uF8Mamx1Ypbo3+s8fYpS/NllfkoY9TQQ0LKkqPBqJslk2KSfJ1zvBs6kAPt
DD+AApgmF4H6StyGDi/BulcpdH6jdpmJUjU1awGtc6CXCV/eiadjrvb0fv5RDbG32o/7W7EM1JiC
rQbI2AGQY2Kjx3YyyRUWXrjji2qXRM39PrHYVtPkuZ/dcQOtU4YX7c2KfIv+FBI5wtrBjkckaNIV
qGtR0dPnUCfOBko2BtF+9F9j/NO0dXLqpIjsBpf9jrfyP1Xga2jjQWOKm1WpCROMzLRHpWQ17Vcg
JN4PymzrQACP2FihaDentV+jWKjY23biBPIE3uFhYmNWyoYz0OG6jR+kewju56D1G0YePl3u5+GO
JaZX7LixuvOU5RTs9fLSpXrzJiSzXmvZk3SuwY6H09Q5CXnzKIMUw/WayOOPIewu4OMy4KJ7qGwk
cYjWTTg++4RvzfucU0gJ4xc4ItVssT2gIcpMenEo8gmxqhtVTEZWt5yr26Xf9eukOxaBzp+hYnmm
GOuOGytV9pjf2HPPaXY8lNVIWNFk3d0ENSYpqtgBdyY+HugZ9e7USurchYUd3uZzsPeedcDR400P
TZvdtbxNAW0XtwV/7Jt9SPXPGqCJniMiq2pxaQJal4+tznQkvqjwdrv8ZFibuzn9c0HseTCnEoDi
czk90ZgIWEhA5CXBca0ibICjGYELf+1HkTV6jQ4V1e76LcfGfIgKh3jnyuKIWJ4INDH0ny4/EU1X
DLygsY875s9P5jj1ao8YgD7a8A7bl/9s/HXtdWT74HAgrk8eFso3mAx7SD6NvHneOK5yepBVazNm
x5OFiumGgXRsZcFE0jp7hxUuwYINGBPOdCiBdrZub73cIXalPRhuHhIXUwvwrhNqncWVjIOvze9/
xi5u5rTBb3SPs/GcGegH1ryOofnwWk32uY0kDN0x13ouestMjDjQQkkP42qFIlUXulO2YGv2N5/V
LINkC6Niue9Ku9OUjY04CXLA79EImJ1T7Jkgr/f+F7Xvej3o/GPPgs55dgg3yEnrjJPk1HAhFDY/
k/yPc867HOWL+f7Og7Snd6CiC7TslkPfqLYgeksTo8Ls46dN5mTnv11+EJDUtavItKCWR4nwP4vL
/kfGSyNaSnjO8pGUXNEmlN3Vr2nna3H0qAkMWvoqhcXrKeRzFX11hh3rlKI7WPMGCM0yl36Qd7Ns
LYzyInXsf3ctlka1L9NLnrKEZPv3rTwCH9hU6EdzC5CJKrHM7i4FjwMMsHo0PAwda2E7ujhkWKXT
sxfV3XW95A/UNAySQdBxLBZnK6HeeX/xz0kuBqdtqEMjeiEmpiFPBc3imynRzBnK6USspUfCM7fr
1WJgJ/lH8cJPlYprJBrOySciVZq8j0wfDGWUNrrHuwAXG9IefHyvfpbD4eB1VQUodaAr/jxXlzHm
jpM6kl8gDqOaI9qKpyGWITwDdu56m+qn+RiLLGiGXA39w3IK/7jS13nCz+bdTwIqPfqRzc6rPXPn
y/W6MX6aajoDk2UpioDJdq9h25eMYzwK8UhelTOcpWZMJ12/x/gD4SgDwdleAj5REIxOzYkV1XOu
IaCzEwFTNbAYTNtfdJGwwe8WBK6qChhEH3L3y4zbdrTY6hFPqjOECHaUR9K0E1SnveZCKTkcpMxR
8Vxhtc2pnrdBGdZzh0AYJgE7XA5ny1MXP2yMh9DQRtV2ogdVtXqQRIcqcQXs05EuGOpy5n8lLAXM
eumAdLYe5hu5dF0Df89QqF+06dwR/10c0EyZWTdyrJr0HjXrJjtXyoUqJZthIcFACfEwH/QZLriy
pl/EwpqyzVqGk8pHWXU6GFCeEnevG5voI+z5URWB0ZZOwGchGLtVg8xgui3pzSR2TIo2eKrWhlWW
GKq9BTWIfM0XtMYbUFk8PgEJ7mGToUedRewL/+VI/mxbfOJ281eplLfPMLag28ItWfC2sQJFAM7f
QtaRckm8Koyz0Pd8Gu9/UuegF2Ayp4kt8wVdXok7AD8194j71MQAL2TMBjJ0KbLGCQDEIHDfbvhi
4CngR2xyIum3BnTnQEFTRL0Fi6ZOCuJe1Y0r7NCTNWTGixyVosN0q8O4BYNDIdOo6wrw2dAlDyaY
wx/xdouoUcZsRenaxEv8EE/g7n60BVfrC//NwrDgFbo4+B+B0CSUx7xrVjGfXtR/GqAA4JnDIEGx
wO7DDvpy5bwgSxDIaOrhvQ45S4KXEMIEOuii0FZr4LjsRjFL884NExosqOUr9CFfYBwJuBONChAK
jndzc34LIqN1ouF4yCaTysCal6qCJOw9zpXBryD8B1woOVWuUaoj2MrfgVoO4eOXBOUJkiCLC2dB
5RQev83LsVfzJwyKIn77eZObA3HUnrE6BeEDqAEjTVsmj7hJjONoNxmD2MqJAmyTFtpKUHhVhIjd
KI3o1C9jsgfrghhttTETvbhwQeQ30wc/9ZoCs9nwLvNk2ElJUeCCsjsA5+RaOJv0nI1qvr2NHAT8
RNJGD/FYrLbXj6JGYPgMzcBXq9+fwcbUsWi1AEx8b0uugS2QHaMLAuzTK5rJAYwMeVpLLSRoSKFI
kwtBhKzGx/SjJESmTGBpEfu35ro1Dyi1AlJ7sRmTwZRPPjp3bO11MXmLVittm1whx4fv543oCMvU
JuqPNyf4QccopQp3IVVE/yysc/NnOnICuBE0NCrC+mImBf1tyu5qGvEOsBlJTibECvTxjn2+7JCU
Y43HotxSkgotFl4SwupCdqQjQEEk4+Op3E/IKt2iuDzTiLM/GyoYrQWkKlQZSGa1XssujK+USK6d
uvyNEhPpq0cdGrQ4+UH32kf2sRSTPu1YdWvT7x9Xo8LTIdwe+GUJHQbLuZYFaqFiyJaFJefs6HUw
2rC9X6m0U8p9B96VHyWGDDBrvikHNHmqGKb/FfjiQsW87n3qpwOwxrEi49WxpxlJ1UMPAp0XZrEE
xNYzHPzF6MPJJqmyIfgkDdQFFtFXJQ855cKpT8NIWpDmzzQKitBYlfKjyy74rFXw/8uMvyBEdoNQ
zSkbgF+5oS0hHJZSS93W/rmeELo2jOEkoLAmG7UJFVtNgqaGqDzXArVWfZI4i3SUi6MXN/A7ECty
PNkrjtjhaXOlQnJpQ2BzysbzHISkEaf6gxoyqlA+PEW0jksT5koISxiVEjcC+mTnIOE3fKJcE9GU
1+LiKDKpYO7zn/2PqAP3cG/78tZFWwew+qIFX2xwaAYzZB0ajc7no6S83t2HcGHSF7eFP9khTNNJ
UNceAJS2XL5Kzs+NKX+3wB/tAg1M5lf7LsyIgtT7c/Bvzh51inqZgJaSSNFrcBuXXvIkGR+aTfyk
JUgwyDHcoinYYITLiOC+AVGDpcdu/8IX8MqF3yt76FVirRB57z+Vh7m+4H29lkjSWZBWAWzpT0fB
QFHYPONHFv/FjJfFqWHBa+w8FvIpYBDJ6wGksLDRxP+a5wiEkYqH1Pj+QVuh3dfFk2Ekktt2RiIL
y8rzRr932CQ4wM6HbuhkgewvKvqmt+zIo/oRFXzdnNAOpw7476RPKEl5LlCtwlYCC0dvmGHgOSHG
pWemXVEPdCBKprotX6QGMJVhkXxBqzEzCF4PWyGdluM8NnN4rX+xm9an9hoZnRb8fzQTWd1Sl0TI
0kMp+wLh2WCi5PMMQft4kVZcfLpsT9+MIANSm0JYuqFrT10apkRygL6gR2QbZ23NEn3qe24WZ0AN
N4TvDAQB9xkOwQuETkFqDFMjri/fT8Ay6tq3wkaqe/PisB9x/xWEaQwKCZQaKt6Y+x9yLVaIkToL
X4npGUJBYeDw5KCEIsi9Ow74jjm6XsyN4cEfGaNstVt9r9A9dxZuOY61S7AMY+yjZT9UHf2nnDNq
cZod1C8DbGM9DTgvuhO+oXQlZFVPHhAQMNpJIVFdKoDPFRue3deSYEHRSS4P0TxO8LFAkLIlXez3
8DTaneAwzN/J3u739cronIfeLNT7M5skO24VBbLYXYMGdkfczFtgWHQejVucpiUCZKYQVpsAEKP1
RQ22k80qCNAGr+rNlkvZhMdEgUSEngbYCJjtiiCu7Zu3mIm0uQ5EY/gHXnpg5bqJeXhw7ejQpnpG
vhD3atHDcXKIRKOHY03slIojfvZVLfBYKN0MHLrxgTKxGYXWYOkK8CaLt9iccHwLnfW1LErxuTQu
8WB+uV/LT8x3WARCuJiauxFJlno4JhQ9CAcK5a3CR+tgu/m2VlimFuTA7CAtPK5/+LulbhZXDK5V
ekVt2BcEWYLL6hTsFE+Ipk/Oh2f2l29BcLZ5RkZItTSZ5uJ2E6IVSwnVnTlZXN7O2vMJoEhv0apf
+GEe4Kl14GKmSf34wHl8q8qw9FnGQmb//Z8sfKhwO5vsgIWH3dTHi3UYoN7ROUjYGQgX9WQmUWzi
3CimAMZ1NXH2j7KQ4iSyvLu7PbAJeDNX/P5XHtwBsMw8bICW1/jIxUWZ73p7wUmoRipPdYuJ8NVz
iUWzBC2yFfCH/4gvKHwzSaHrjS7jmfB3XYA4WxYk3jGmyPpOjXUHbDlNW74g59ytrDlvN9KBQrMn
9ilooN8R8ZpUqonstZDbhyDJY1dd4PiucbfQuwvuZwE1AAXaN4QWfB2p3uSzw5Rjg7v/36I4nW+c
jGkTDTOgVhQE6BQ4KjuGChnhm0418dyvyaSXisFxuy4pqR3G0pdKCHpU6enCWSVaFJJVo4RCaaPC
IUnuTrKIx4gsp5JtdXPyFtieMooAEsmLCWXiJgA5/5m+ba6vNuQsCYC7feHHHBU+6sO5MDFxclJh
mqSsjTMBzAOLnfdfKp+lbDy6HExyY9do2RlyQGyUqoVahgAcSDU4zIAqoHx2lw2cOwpiPvevU7tD
eA9dLz3TBEi72zQ7TiNOtLSxBmbk9DUvc4OySlxOWb+R39jOv1DDPEok272qmx833Q0tM9Cyd6J2
/TfObdIJoctHnnUtLTSb6n5UjkuLaM4uS6bvTdJpbLxRltrnuzTDLx1LgpKdaGh7kIS1YFG6p1jx
YLbuYV6+fX4na+RIjGDNlzYYe+AZfRTpAx4w0WsWT9wyJa8U6j6T8bU4/yvk8zPAI0k4U23NWN0E
hWrLvzXj85lUwodIEzAyz4jSHHCtdghPYn8auqH3gOgQozP2/a20nqHn7ksimJzIXUqDBV+earkq
bC//r/GbLEJnFZ/ZJACVPoznYx1mVfYcpW5v2e3SpicwLq4xqhA1mlW/eSn8dYcgSsmn4BaZIhll
xwiMYg2ZGJUo7SnsalIbU2sY/K2NPQnk47JK4MnB+hn0E9jPnfJ2PrLICXfXD6tXcdoDlxmYNkpl
8xsTDfdXjlZXz1n7vLy2Bw2chn5rahmlxhI307FeYUjWbN5D8qe9QHpWTxD0FXCqJ4TmsFXcr10K
UlpAp9EPjP+Skc680fOHuIJcoayaSbdr1TD686RiAZCHSf5EZnGxCnqZj2uKdKqQtCtL2Mluu4Qa
deQneg+BQ3QM1lbK24t46wOINZgE8lWerBPHlzAmPmgnOgHd42oh/8nc59qALlBnszKgo+d1e5/p
u7PHryAbA1KlUWKa3HMeyFQc9MrI+VCUgDtFCVAtjjRk10Ca52o9ZEB2E8HfxIBvpMF5QZ8qpL1/
CMLCK9dlZoVmYGzukc4xTX9cOyhYLPlNVdPvZbRLl7g3oce4cW0IeFhtmPXDV/BEXhB0U8bUJZqZ
98y8ZVegnqwwXBrqIGyZDEoTLzxxcD8n6qEcXv2i9rU4I4sZ7pE4OxOrvSZ02oeSgeMOREue3c8y
aFS4p/A4mQDRefMcvzY+WGNj7VN/2xi8TOrvo5DURsgHRUxPFge7F3DVrEAUEtBzIMQId5hz2G6S
mBAnC8lOVmaXYQeDs6gbF+GBKgkrFXZd+K3x2FPX7K2iwZHU4U1ZI/nG1APR3n5lg91YwaZDp+FK
gj1YTzt5dmsbcf1PXNtJc6qKBLTqQXI+ktycujXw16VduJN4j0dAHxN/YuijrqsTsWQk2dSqy8Ww
WtKwyBeLQV4SI4V6aVNzCY9ckUQ3fHnf/UyAcpcEHMxv+BVSbvrO2AyyAAEzprX17yoA6TQlrHpG
OTQ+2w/iMZDW+wLvptuSSypQRfPPyqMLqDFEUYyZlxS7kCKldCkZ6sumXj/9/JTEiVpohqITOgWl
HVeTspHF6d3WSujAedp3eJhhuwywroNyYhV6APd60ttATEhstuk6mzm3k1wx5iiBfWyCGmSmDIwT
QOwdG4Ki4kf5T+imAlKpncPmjrlxUKrvl3ngWfvcgtZGscyzJSjeJbdh/GtoM8CtosKroP/oP091
XGAc1IgygSTAkwQghdUG48hzdmfsFKzu0Lg+covUs0en0+NrtnpdgiBW7Tl7+Tl1/SwrxEVtQ84k
ouP9s5yevFFNhyayFV00yY/YgHvLz7DNmiHqpR3i3hIMuj3bYJvhZEP0WgxN+dd/5Q9KnYyd0pGX
N2277T1t9kWuTNYYCzLaC1vU0CDjFs68s5bKqiqBTTQdwXHKUNVCAdr7hDNvl2dDvMF2hnPNn+Fg
h+Q8jqeY666uhXLUSlCXrgBy4t5/U8on0wi7DjROs3dD4OCiT8qa4fUp9Fjp9QHOpn0vP81NnRCM
dhP5qJUTD2F6Ctt4E9sWwU5F1yNYvm9KRddxP1tBzqdJGNgVbbEg9SRk6VJGQmgkvSF8kx8o/zvD
mMI/uQz9ay8Nt30l/fkNxk1O8FzEDb6rhjwZaqlUKYbEakTW9UwVYQmGGixlXVvBR60KZ5DQOzT2
Kpq17pL/WWeqhDQrU2F6gnXvCpm72/CBfqq+QAqd3YGZ4C776Tba4YqZxDFsaEVdM+hwCDj1z/kz
ccJlq5KfzUUC2Z1/USD5eVXuVJ5HUjaFezg6axzr1UHEwyEb63f8o+lJzqbU/LSBA/KEgoX+As/5
EOSHekV+q/BfslONvB60Zaq1ZtVf4mtDpZlKW7nftl0TIzusth3ra31BConSbYmpYMWdnkf/9oXe
BaYwYhhz22I0bZD56wTW+ovxhdXm+g2DeTtwjMnNmSiARDAcnWd7QQM0zKoN0nQzG+f81cDvZz2l
NXM+qpbZA7F4LSG+h34T5jMils28QwgXM9u+o/3mkqPcsxYozFfMq49v5bFDY0RyUhIJtjRznJtJ
Iz55X+QZn9Pn+jhKQYoxxpyTdFX5+Zx540K4okM06m7z0Kc0LCa+fLTBZqbz8OEssk1Yzw8qjLfA
uGLuo0BGqN2rM6EzfEeVBiJy7qphFbBYknESmC8qJqlzyDeVRCrz11BGnxS+llMxm8dqJ+ORLHtQ
ri6qP5iTi/aUZ7Gh7rgQE7D8J4fxlFZnNx+1kbmaVFYlknQTVq2b5hF/CPZGa3rg8g4rIAPlgyov
yQ/hEMJEkhKNAn2x/Th1Bn0HRo/CqQVyzsHoPKaUNDyjfdw3MIhZx6mXlBE5Dfr7x0+NH19p2fF0
RMB5+TukdeEUS6xIjow0fzKdmbnWboSDxWgWmzKv8brdFSaJ9NLsXl898/RoUCa2r7MoOQlSP3V3
f9Kk3kGeWw8j41wFMkja9cB/qo2uxxJFBqjkJqyXi3X/JL5eh055KINeTx5vWnAkqgaoMckQsoTv
hfqmrWqMcjwewuAGPKTEcu3xuZrtiRpRSlJENXSmsBo042Ui32MYXFjCC0gFX/TBQdmAxx0wxw2o
tnc0Gs82yYHgRFEv4kNmMD/28/cupG5UH0JQpeGc2Cyyfr0z94jV4p0BmJZ9Ez0hWba3eoia1lUu
XXFaMLRcXizzy9L7fzyuRfbVd2OqnjNrUIa5YY9e2eqSugPeEJkvuoPDy5mHQiGoNkbr88NHcXJ9
cVlr4Wm8qkUHK9l1+1Mg3KtGFHb7PVPKXTT7Fy32dGhvBQVWxmr/bANblo4ZjSt7T0mOG7yWU6Et
31Gz3IeM6ds4/CV3XQ+VnoOXk74tgv2eB9yd+nOW3uWldl6tdOp8BjJKyHLxqWT5m0I0D2GPNxgP
3bLF//j9zOikXAZskRu/7ubOKrsKGQBXS+Lc186i/HOI0bNLPera9hTI8iD6X8r2Gyb+zLcbxub4
wyYP2Jr12q6jBXaHLjVmYg0cwivdkAUGkjVyWEMHH43VGcP6K2NPa9ty00vOz1sFRJd9ucZzOD2P
5oH0dUHRd7ANAvXjeOWVzhiS51K1tiDlixMuPcGKH4kky62JjneL38g8Bjb33rxCBy82OCIXWNPb
/jwuG8NPa/MmkXCaniZyASeTRMBCQa4ajSfsXIP0iVqlAEQQ3eEp4iJsZGni3xAIhRmpZ5h6YnVF
mLEw9E2QYpQ6/ywCPJhd77ezZHKFhAy3FKsP5pKKIk8KORAGOar5Kt9jBSGRYJSWLMYvdhOvx4pB
XjOAs4umuBnqDwzBhZm3iF/d1djcEElNLN27+oc+t9KvzhghClR1VvMl9PHLC38Y/kqTQZa768eU
l1tVzgrJrR8GLIIzaEZsnkd1W3NKXW1ZNvcUs1g6HWSVSAtTC1OIGd5lx1k3XoZlEIT+HtiDMuKt
zJ2KX16gGXyouzulIyC8wEkLOqu33c6OlX5qlb49CcbBC/KSdZosA9ejbyd/9kJWfC8Bbkvz+xVK
PNaUqy7Vsa/Fbp8+olbpP4QcWM3O/p+O0/fDYKsilPgC+7EV3i7wbdt7MoH+ajJ5P+2gsUNq0eCa
7NphxWhEah0TfolJTyeKuI28BV4gHJPeOzgEz0JMx9f7Xq62GqgiPjo00s+oh3m1GCyIQgk2ar6Z
jvHHlMnY6LkQuEG/CJXgS+Pq+HYH2QXGGTLVJJbVXHk99iAOYS0rkcmeqpW4WWdkCp8Mcqwa7vZb
jC2F6fLrmfiueBElwMNd/AFZTeoHKjUG6HI7hQiXzP11xVghzQh1V9xojXEtAHcI3MnOgI0W0bXh
00jNRG28fXdgnVOhtvwarAEcGU8LJHjunSLdO8VQzmJVO3h7LsGHbRgG+ABZDLsErcrYRrF7D0P5
TTJ6OaZ/gHrtsScZpCyYQLI2ocPrarej6BtwcullW2JHgrQroUbVy++rtOBpIWD6QrnYb1ZNI1tW
8c3Xx7fA7kNSwddV0l/lqESWPhxYeSOg5Au5aE2nqdaUMqMGPB3vQTEDZ7NBQR3k6l2P06z3WxR3
K/cvRU/w25Ovl6HlTuR/lBNelihJC9+zcmCjvgZT3CJqdJy92roJsLMSJuIKMcjmkHKBbMxoQmN2
XGL1etdTvQznSxRPnpBWcSWNNmh7Z1wC6aCbLr50KUmlqbdn7934urKluQ+DoSwSAvdikenZ3o00
nVs3mmo/PQf91BdjqBTEfxGCEiiKqti09joJ+AAnqyY78LhUy4InINw91H3u9Gjmys48Q2UKMvIS
56QaqeX1kjeqxnTJjk/R3BvCwdKyg45CA8Jv8MJWw2XpMhBdFqG0vU6t67a+W11VuIOe6VmReFbz
KAHWyro/L82A7K08j3AJajpiNI5akvuwV0CiVam4cU5mQC77DOEbnQAgqEVjuLChxGrY/6cgYiRR
oEuVY2SPTcvfB47YeOge1IIDoexpdhbIfLUKjbgnRbY7AGHcJYmYN7cwv9DN6uNLANHG6z4EC0/N
CyFVj0JN28Za6tIwGkR8JFChLMlQ4Ef6FUgPRR5+SEndjXXKyq4NP8oD/U4Xna5nW97x3lQDG1qv
RJRCWA6Nl7lyu5wYsx90gCYEyJTKfuGBOGwvcCDUJLfNMFdzMszOR1X9ahXenL74cu8j9iVTr2qQ
BLFZhxJP0qkJ2F7mSQhp/mryQYGjmMnpLqphQhMsU3qWG6gcOneiMGbEgaUMHb2HbVlbVnR6Cz2M
DMv7kOru2wQI2b/io3LkslpRleIetp3XMoXubkLg3IUakMN3RxWjR7eZmlZXyIUW9sZ0GnULlW06
6jA/UxamaIu1Ptk5YxjgBdgAcssLkD1EvBV4UAITjE8YZOtXPyzOcDsLG1fYRT6n4YG7bzRXCg1e
Tb0+5Fd45oOu64Sw6wukNmXnYxSoj6/UuEi8AIUD8Og6mVV3kvVIWtOBJgSIX1g+HDmkRSX9P8mS
PxFE1es1HSXNaPCt3g85+bS6kBi8W/hfA1HqBBUjVKRnN2g2n3sUNgL73lxvVMKbTkjpUNcekc5C
SfaO6C3uu0zmh5m/Qu1LpYbustITDdt9T/Z1LrqOEg5SxHAIrnn6UGxqdbMa0eRuMoHv/KKeT8A6
5tREGQjmPLX3Cfyc9CAV3JA2avJbl25waYEoUrwZz9nV/09FgxjhOKO+doIOMX7/Zxn4aQ/pvWfZ
iy3HpnhEGvY5kvnn1bQzXBMFFfsDfccN2NQCxy06glY5HtxjgINGISUZxGU8af1s+aWq5Jft2UOG
ywoyzoWpjp6y9bviWCk3gn6ONnx0TrriDwIe7F/dPvtQi8qMX+mA8h8zIfvePLEcyL9sTz3KWRco
GTLanA52EFNwgzYvGCrm5ETRtXkoto/j6sEbbFmNMopErzRmrFhzF0413BSbx2MgNPYRVXvzLIiF
tmDv2IEtdvZqWqcubS70F50s7kjxW/RTlx/K59KnZ2Zr1l6aR1dudzImjky7ePvPH9w2+GPo+K3n
jTT22Tdbdufc1EF29SvXm+05NyW6oROFOxekzMNI888iDz0OV13PDVUekUjM/OKOPRTvU86F7N++
LxD/Glm9EgoBMxq8IvfR9zvnQdx9z3WDd4GNse21wF0fpWZDFF6XU/j2JWbgbPbG3kJ4xNf69gh8
Z4bdkujPzYhi7stzHpUshyYMhCO5TJPWEaECuvqvUveeFotNExKcHD7042Du+Wyy2MkK91864BLS
b/LHn1i4FbqJcr2eYwWSdkvwIzyuIhvEmvPWWLF3CslZSTVY3CXdP6mJL6E2X2arFyaA8eClO7in
4TsIQSdfsD/hwODjpwkd4JoAVzzj9cmdUoueHAobvxjyO5hT3XhHaapIAGFasKeck3J7VZyn/jtT
b3BOePoYUx4+plKgikq0Yho/aHECqGSwATzh/jcjxKWGu9DyXn70fYm5ULenaJdNJr5BO86uc766
CC0UILM38V/Ilx9HZ8U/QyATCnVsFT6+H14Z1Pe0MURfLXZB+hF1GeApL5IVYoxLg4Pz3rkbSaVR
6J16nF5aDEqThm3yi1shPFrNFzM+Qg5ukW5f/knsP1Hy8VhqBvWMhr43qpirDIYKBsvl+Z8VS0aX
DNjEnShNVLaPHfPDTwRD1UPJkFDxceR12DC6EnkWJccq/MT+7gDMbgyuqZp4uI2rD7phZwY7q4oc
YMhJ5Y2D0tGqef0g/YG+eOzCM3rwJh77Jb0DQQRvVSof6bZbhgNGT5N3nUP5QAEqeGT0NDVFe6ov
/YYdmnRenFqfxHIJ+i8M2n7bSjl77zg2ONyJaPFNi/yJYLQ/+SuSYBeaY3fzLsRu88TTvvF9A2lI
YdXHqTAV+iIqtx6SDaz4OK2n+pRq2aDnGxjBIJ2tbdT8s71dYtSNNIoMEuUF5AEGd6/qiJCAzrEZ
C3jqoCzmUTsZ1wj5clYayMJvZySZuQAnpZJn4IxjMELiLArT98asDHZb//hcZ/J2PY59TwdBKC5M
rx75L1Ph7qzb8oc4EN6xtI4jz2RFHbxpRQakcji9eixm2xnhde7f3m1orgyhmWMExfp4bIEGV2z+
JhSJV29Px8zOIh+YQ9pvC0HE7xDryWKf7mihHoqE67Ii7o79qVTerhHGVkUJJ8OYxqEMwOtH2Xte
9uKLQVkcJFQkmQat8s/KHW3A0y5AM6ifBT8J+UP5Eap/qTKRFp/hKNm36O/yG8e05P0089ay6HWn
zursM7ocf6cVhn8n8eSNqNDWSKvjYH6f2EV2rYdfZEpEpfq+fP92eCYhdpngW/aXn72NYtwvCSwq
XLCVgffjIYnpDgLyZT8cxPv8WY5Mo0dRR+F+MUutiVTI7MJxbT8cTKBMEu8zjK8UbkETwTotcIWk
Yypw3LJ5qtcaNcJUumFrzaBiVqWmqWbQNNWrVkESxui9LBvcX3kfHr47IUdRuWMAvJUEOiNnUnFp
G0JLsBmCQaqh4LbsbKshDmfbyHPI+qRKMR+pUd5KQ47hzKi/vMJXXPuJug2Hk7sH/a+XIBqxr5qP
iaLEbLMb+WY2j70v6SF59xfj/Pis851YpMOCaDlcJWFJx/z5gnPs1P3uvZc5UOIatruSXcpzl/B5
eeJxpRnckgqucR3vbu79RPkKbXvbNS+dC4gRGtQ5/uyoNYYbyFfHWPRyXW1h1s0rVxp2Yy3/eRv6
VlGO25ewxcildFRaZaooS8PwllPRgejR4ei9Dcw/3RGfsAqjejgbirvvCaSJfbVw22cyTr3u0h6a
pSh9vxRgnzB0tjn7ik0lGfmPGO+J88JAtgZmQYEjZICazNNJGqxnU9BqL6uttPy+5EdyWXopCd1b
rrOnIrQXmXFvNZCrkngWH7Jy5PIc0wWu5SynM1xp5wfpwTuqvjpBhwjk1zOxd0NLcUzKVqvCXpDf
0swG8/zajK8YcsDG98ObhkC6juAWlpBBhzpi+tUozrHAA4bNSIj3X/amQyYFLRYl/PkhNO2zfFCE
PTxKTa1F2qxcsMyHF07j1I37HcLeV95S0hQAniNGP0AWYkLjj0iFOVTcQEDmveUgChbHOlemfyEC
zHWTBqvFtPzlGxXO25Elfhc5FbbaYeXMWHXuErNNzhG9xarjJfjhcTtaM2eMQm8oeAdZeKhU1ZPD
DHIfQXpgujDQ2hV0Z1rfzEzfRDzVDnnVtrnRRQ+Sk7bzOfpp7ktKlEjImcAZF3vfUIadiQ6Or+hN
s4KVNgLRV+F+mmFx9UePXep4Dpiw7YaAzASTfGFimaOzNgCLqX1icMTkEzGbGCLAIh4/DT1xTlhb
FBzjDBUFM9iD/g6FTPLxP2hXJeVeX2uAhCxZj5gpblF+K3mx72ii6On02c7cdzMVqPxg6lnIJ0z0
wlMeihboRMcGd/20OigFL965YN17Wn4x7B/UtF8JXUpoWhDrOJ2t2RlQk/BtkXH4dHjg8O2pvy2Q
he4hfJTL8UlBRR/P+5qjwOmoX/RbRb5tk2EXAoIeAL4x/Cm/zdZ9OFS0vFFHulGaDvKBELmEqv9p
2mkTYiymJXIkZsmySbITOSTBVaOr/p/F3NJb+BD4slTRckKPHqAmfNn4FAczN3vMDb4hzhIDUvaN
C3pyrGe7MlT5SAylcs8A/Vt+JHxE+Pts6D/S1T1pNDV8HtIhHJnlL5l/CHAdWXdgECJRqfbn7B+i
c+44kmEi7zFr9F3Tg88u/S8/hdsFwY6Lw+yWhVWXZ9SNkiZOpmUqhF0z6cOYxtu0OhAPUNXITbIh
CXfeV1YDd1GwxSecJz/AWHljL9KERKq+PRZjUMRkuylNAqw4A9lbI+M7Ix7tBASNWeXeiQ3SmvlF
pEecgCZUPOxyXuGrJkJuu5SsVG4VPlIzuFn56uUqi5WuyvNeW6ptWzqrwo0gyXhTs8he0SXV6tNx
oXkGk79kJJrcDd128Bi1TaKFWeti1zds7CU4Jr8KOvFTbtINauNziAtc1TwCtrxBSFhVXuFBwklz
ShRO6owkAo2J89ZfXtbfHwIwqBVUXBP1FMZKIgpV9SVAZUck9qhqrFMZIWru2pVdKec93m+QQIYu
r6YPbkv+P/pyD53WhJc/xX53LMpEOC1LyrilvdHFniCvDAQuN1LSlDii0M5lNK0mx7VO7N0IEDqv
3xkyYcAoojyT0OlSQFYMCG6Eq/rR6x+O9GLmmqPelzYw2HDvrakDUtl975tOK6hatQzXYk4+GlCs
8pItGjkGz8jcHO50WshiZG9OJxL/yLCeoUEasFVcII6fye30zR3uLZR4akg9aN31pJFnrb106MjK
Fo7z4jvKEcyyloIgqe7444Vsa/YsM+ZO4WnKDhVuqj+nDnTGZNuvcSTDzrHYH84j2g61NoFRrzii
wE46VB8lY+AzvYwPRjjVg3hSkzAwyWEDjGBPgxuXQqRChNmsTBc+7AkHCIErvwKZyRX/xniOZ9ge
ylMQt3dMqgkvaKbb0/RT2N7M84HoWVlL6UkekyfeKM27V45ctlgP4F8cgN5Y2/U0Njcfz+C0CYbD
t/braxBvQD6qq10fa86mNInqlpBV5gznI4Vd8gofK71r2jUJCyyNqgg1K7kbjxZS73cfscCAoLWD
ByEm9QTiU8Okhc5mWpdSQ0KU31OH/Tjgncur0Li+y94Xs51PnOADUQMmKUljJA8BUJyZ4TKfFYML
BQVEfngHQX9/s0Sj1W2NJlzLwyohHfptIBXAzWdnwuXCrFx9yVJfCVE5SD15YU4YZ1NlNoEcZrUy
XiMcRl+792EHazh1W8yIc5djtKYT2sG9OOoRVfSQRMyoQCogQVIMWd0cBcfYp8etQZm72gQA6q4Y
H08U+oEjQ5517JhglUuoTQf8ALZBE8GfO5ZfTM7YTaGKAiYZmYUObcpQYxpwOaN4uEvS5/7neVNK
AlHku3V13TmfzwHawj+Mouu/AWPU8QbOprNqEW7XLQeCPmN2TjbrQ9KTrkcuWqEAzCo9jMPNPKp4
6NqV4/ArLMpPyvTgAJmiCYxjbV2dbscNCo6Gli9ZVRXh4oGHYL1qBPPWHV1I3j6Gqba0IYxudqzY
0nMeNXRo9q1L0B4GJ12Tj/xiEzhn4vAzM71PjiWHgnPA7pEL+KRv2nxmG5Ux9eaKMacpPtpP0uvs
WJ5sh5+u92GbpgeXBlB/t9h83LbGvtK1hfLH+KLZqkvW/b1RbJhsEzuJX3d2nBlGZ7dnUMH3GooT
jsNw7GLCZO68fAJRNrVDga/MM5hmeutVULFbUijSAABHz1N9V2ZYhG6/HzXxGWDfbSP1JJF9XdHe
0T1ZfEbViT88tncz4i9S+wim/1Jk8PDz7KsKOs/Eq0LP6dgsadTL7tXVE1XrHK5Vh/tONt/Ju9Hr
ndlvXXw5sfRoyB7TkRkYy/ktKaO9OrzGhuZ4O7Dklo/d0D1J+Zq0w0E0XYKQkidJGlAZqB3GIKM2
RBKDDGaFeQ1jAVJgqno5WzmBrqJyhrpKcA65Xjwt0ha/WqH1sQZESrOy9ji6gPI1hfZYhQ0Dbpvp
02vjx/poUYuF6Em4lqfgEZYXV9hLp3awytl8DldMT03hKUTMG2NYbAdBNmzZTWERkPkqVTDPBN+u
NBU8R42O1mCrkjA/A6/LFeNiHEjSMj2PmL8OHipGN0Q2xLwYHbr9My3K0k0Y4OHQl9Zrp+NP3sOd
ycR8K4jLTDxhE0tRr+ZJYWhEEXAcbe4/dZ3HEnANPHXChFR+lQV8DiDeC1cJmiE29QEQY4FoJLUW
RzhByUqr+cXEAn0/PQGvIKG6ySVmtsfEO5z1jhNuVY9Z6vmmnCjUAa3w0NNHLZSpvT3OWzzqZVtx
Gtdi0K/Faq/oiefZ1yMRWRK3nvdkQ71CCPvG0kk866OvMrcAv0kYmRoLaq5vWLDFa7G8jw95D5Th
09YthAjJmyg1jGxKrkC+L/gtqjszvyZRjqYjbQoOSekO9uOtg+DMRx/pLxQfAL6/tuDB6P2JrKQg
h1sYjSqNy1cpGE281w2b1vT7LErlbyWKKkGStPcuTlGYaCWU57VGehbtsoCy2XVEHgcQoMf/eKUe
vKGb4ZWokHstg51/ec0WydecduTnnFCq+xpF5sC67z19TBx6oM3tkllvQ7eXdHy9/UeGXLM0Udln
FVKIATjNPlvuBC9ecKLGn0C97PQ4QfHlLxMhZJI6Fh9/OJl1yYYBUMxDcfBYdenzUl/5NUDvpDSm
hcc8HexCMf1GOMJGW5O6LeIoFXZNTRK2nxNs/tc+pFV6w5Eem5QByNCzEpnvEjjbhPGsUUbsquwn
PqyCG8CfLShaTVcitXAZ/AC7+dYii/gdcmfm5jopTZ6CjHEgHyj8djfMPpWY0bIt8USUwPPV1Gok
l7NGrsrySk68bYIisENNxkmzSF358IZCN8LQkb2odIOS2kOhVZjTWrvW8mp63iVCArYJCKnPVbHh
vwGmyGFOz5vWJn3eboqMF845hU+zzI+crVH30uUWYuEQR9gsbWElBnKtbXZ1f4fmqY8y5jJALyaH
WIgjLbEuTtbys3ntUyecV3oGSKQ6bgX/Pv4XXEXVrixgblcs2u2KugcB5qvBIxxdt8yoOxI96rlW
MhxsXS323klK/095s8qF5ezJHxPYqKmw1m1jZYNlv6bowdICo4SYuzyuCc/yqR7WmCs6RMdORdgu
QBmIXKOtquVPfi/FxoYq74NBGkSyK2mu2ZcPdSJXs2shvmRY90f2XBzvoXNOVP/pKgDjkhFTH7TD
B+HMvkw7sH2+0xocAzQ6u3vjIDcjdYlJSzx/VYhqC/CxL58QdifFPo6PFYvbziKkOxIL2BtC7Qdx
Z2KhETTDVeyLKqeHa9Ls+u60sMVdt9pcydej9amzPXI1aXvrREhIseuOkQ294zZ9Ou+wkVoOzapM
Svo4/9BrK0KRDgnT4u/GF9uebSz+PIxlnV9ZUWNssQsgGzk/Jz2pN4zxonzmUxaiymhx0tNVhTlH
koTH6Wn35V70N37XQqdF9TAwQdO9+dXq1waHC2lrXDcwtrnkay82QL/gF/9IZ2vbZO6AoTyR6v6E
TCKF30FKEYJslWdLIo/DGjslturJCyuAFT+QE5RFyaGP9YQgjwPWFw1ICKSCGohZnKgu4fgUCg+G
x1B5/9fmNbDAquHO+LLHHtCj8xMz9zjVtWobEbgj1bxC2inVC1l6w/DkhKpvFK42hLQV2XRLufRb
Fwlzl3XGISsCbKw8U0V14wn43nLGA6K/9QJ4cdNM879JTBmEbAk0o0aMRCgySN+P09cGhkBbSioL
8/m0ok+7IajYpbmTsqGYq5Uat4ZbdnqetGd2Gt8R+JMvnLxneGltVESj4/oyF90lQqgnCwOEFcTL
KyxP89daUsmuZlLQ8gMdtGbQKlWQlylpcUPeqjyq4Tfb9FcRWNK4LQlgenhz9wejgvq/0ujhwRK+
nVIPh6/Urs2fBDyLTBw1NzG70vTC2D5IHCWTdpgAhM5L7q1y8PyT3y2loms2HIKctbK7QAFNOEpu
HuTo0vyD4P0z8TeXGVlku/8c6O6JmUBfZHN5zTe5cMfeGAKEm7IzjXPEoDGaYE4IJETB3UXT77eg
IVu6uRy+ybY3bRtfJ8W4HoIjYSrr0chgZlYA9yhNMSJTmNviHDrGkQKkeVLmei0d5ooq0EH5+sbG
2kdxwt2lS/67SP0p9hV6T/TFQsoKJ4XtTKeUZ3Jl3HsfHy8eG7gwmEUfdge6ZvIKEwH4aypypGcH
zAO1TKmauf/FSMcy4Iqu9jaaVZpu4qFjuGKAu3/sQWD7fC3ySYfW/iVOVIi84XLo8Iqwj0FoF6wI
YmBI3f55tgi5Nof/zsyo6qKkV7izt29l+uaoz23EDs0nLMpJ0GogfmWoAduMWUkzItKCLQtgz8j/
ArW0smODbWMGbPimSzbWP7AKNUGwPB6K85ikMqeaM+fRPflUwuOqJ53RVmYHlDqYX1DsTCjK8w6M
Toe/fEjKbj4NnrMIW7OS+tWdZ/9y2dEHHqbR2xbgdXT4k+Vvz84VCoj59lo9tu/688t1S+hy9CDX
dx89BVRUTMkfnK/M3HGXSlpMF6fF4UywEVzlgHZdlVHH8IvALHc0yodJRUa01r2ytyR+yeUB/ftM
iI4sNfvCeCIP844t/7YnJU7O36LoV5gQ6euy0VYblIVg2uZ7oSLwu9bIRDnl+iaP7Fs6ibLtt38C
Rd+QHL8EGc/qarSthytqwmBClE7woWoWJPK2qW8SHyeyAH2Fw+FntHROEslM5Kx9mSNQXhWDLakf
V/L3ISPUYliFv5/AJ6JyuiPc3egaEl5EguWecx8cWc6n7L/j5Rln075uJegrRZDHuvOGbynmIhmV
JYdJGAaKfMX0uG9qOoi2zFYaK81M+DPcnyAR6dOr/GKH7PW6KM8IpdnzehD1E0QFZfjAFz86jCbi
OqXTzvgNFtAfLZPDq1V/DLK72uZN986aHPVLXlS5cPtNvrUnRdXNKqZ3O6JidG/nm1ysuMemBhtC
bLQlU52bWITd9e2bCRytY3SS7wX/Ch8mxeKAeAz3d2khVjzbBAdF89vw1ElpbFJZkEQlH0mtbxyW
o6hiYBCFZozbACT2ztXV/inE5Ik40TnBSG7RAhphmorzUxufmXcJTgT87TDDoWvSBOkqWJPoyf4v
lKxObiZu8duvZ7kWMA3UFrzLFqayh65kH2gffYbEEF7Xz+ZT+THWeM+80TQSeifiPmV0mEgwfOYG
QKjTQdue6mwWobn/KCJjAItZlR99tdrQENDyPkIaY4o0Ek3LSCWs3iEI0tmpHcqCSnMFazLsNLYy
3RGu857bEUx9JKqn+VSgqdCFMWCeHBypBJ/kGdpasqo7RVyU68mK9o1cjXE7tpeeb612jWMu+UIL
zN+8PFU/Rbr1iexxVmj+TSdO2H9ynXcj5y5dVDeu9Hve2Dbq3sGzifujDs0buV29gaPmjrIz5dhH
ZEA++56mAIHU4/etnymYL2FGaVYtAmO8S5PhN6gC8whj5dE+Awp1zA3D2/9LHC8eGDKXrjQOlKoW
ZdnZXzzC+VJMavKIdy0/AIKQL1NlmMl7fSjKRIt6L8MY8E/fFb83FzFTCxSN1xmXpWpnWud9dEMJ
aA5QxBceTFQghSfOWKWZQh6B2MdTNiDkFPSWXkHQUohwHpUKEF9WJuyvkUMWsN6o5kvT7zXI5na0
dD8LOSvrOBR+SjBNWCI6Qa2IaKhK2WPl7dKxWxO8VKFNJXjMF/7ENPFC+ptGRUtvJCZmoJCpjvND
qqYyfcb8LSkcYV0/7b5fd30Tr0wmvIG4KLKyEi3lL0PtLEJVHYmDGvHRJOGugssmDhoNqoZPwws1
tD4Hto6dlj2L13Fw6+Dbt0kAjOT9C1wUoWFf1fsJbUu++8flWhN7a4l3c9dTjnjHkN+MhqXHpvyk
vKKgTC4eNngIvS8Npvi1rkEOtbfVPjoyLygcV/6JAQ0+6p1uRZ3vdl7MD1YeHAVmqE7KQpdhwiIm
tdLmCVIVpOmeArPeBDI7uIZebsqb82KwHkMrZa4Sa4zJ57o2r7X+XSPwzolZZq6QIdOkUdvfzAQ1
BVx2riL85HTuXzgsolphu0ws31O0k87QSKfFmsjQdp60JUtcB0rQXBun8UyNXuSE0FSbnfVEg3GJ
9lPb1C49YsKp6oD53qoH3ccpNtAMVH1oxbB3OHMfH0ZQbdQx0jOoPno9kzXTwFgR+jkspFyQ0XYH
38MuBmJ3WPwvhkBRiQu9Vf/YEJkDuraNjZTm9c25WC+XGXlfVcl4MhW8icHjpMSdK3Yfy8pt1E8b
RKuQwi9/vA0WrPfsHkJ4ugz322eHj36MCEs8dIkQiv2KNk/z9x/peLENIfKtD04qv3/lM5R/uxxH
CmFyK5k38It1wcCtdT4gFZM5tl1pq+Ag2ah/8yA7VLYxmdojDtUHuabNq7k3RMxXkKNxuUsCGzTi
a2tyHDjSU4qvp666QgVipC8uNk/xkFQw42v2UQ5epvWphxBna/dU2sN1TMDlWsgRHGWB8BxOaKbg
l654DhsArCjRV+a9RhgW4zP982h9+HC4o/PyT6HFG08W+jyhDtxJ4/0Juu0wJMhi/CHh8JZpUYFF
EOcwBk8FdKy8pnlDvk9hiR4HBVceEbrTZNM2l7K97EVCbBRO5zI/p/pNNwyvyIuEfunWviWB5gV1
2TadAEuBajO30OSYutgalomURzAIZGUvus2UYXCBGLjhFJdAhVw/LvM4EeIUvtP3Rpy2F0z32x+S
h4iQl/v/DUwOqF7jPV/ukTFwlTDB8vwqu+TpzoZXDbK4zLuPZ3Pru/5gffvHdE38TvXpaF6Ydjgz
86pTxUjeSnH3x2rHTq7y/KSiW6JJDAWolgE9ZhM5ZPIATxv5AuSipLUIbcTwPeGEa1caPsK5VmlH
1LI5t0aCI9qD9TNPjjKYfeLDiVF5spDYD8Wz+VjAwkjin91jqSGY8XeKsIYkUF2uK7zVyHBESksx
9z7iZk2dlvHsWcsK9O+Kf8zAO+ItOvyTmkNtoYCwIvjvhcfeVQX9fAKoXPM8xJAcmsfgTov9cawG
oevBFN248UzSg+hgVTqqzeAGDO7CN2zFKw8uU2OZsdgHByJUI4Imc2Syn0xQE+CGhG8zgBrxzwxy
RICzbRzKg8L0PpWfxU7tZJQoOO68D9Y6aJeoyUVn1+oAYuekBbwuxOAg2p1lWQJ1Ej0bhjz4EaWB
LKjf25SU69CKqmgUKsHkhP/e8y/N25rct24Hnk6EktYI6cBk50ADTqcfP6bFyAXXJMrE2AYOyEQx
1Wrku/h8Z+2n6tF6hpOFRpuGXX7wcfmYLlthz6n9oVGuobBjWFHJdyghdLVr0mwWCubKXt1uofYQ
cDsHBtFXx5oJHCNcrW078XQkFk7FpTtWi53koqEgd8DqsyJROUXysn7ceKT4FvsbFAo7yckfzTCn
p/TnCFl3qDw5bjhfqH2La1ggagSqGYSvUT4ofoJtfUI259/vgiD85qO7Tv24tD7NlzPiBECllPME
x3+Qpw5TY9efG7EyrDAdj+VdGnVgF9UYUGHBWPRAZIOc5rC5VRWoEfyl3XHFraPMbKW191ihRTPG
rg4VUaQb3jUb4eWZEjW6Vrhl+DLFpvRC5oAym537xOtvN8NnDFVsNlYG1s6PLDx0Q45OzBrtXe0K
fWRczjCwG4cAkon7Kh9UBwZDjYatidyXZMBNK0lWWttf52EvU7K1Y1qbGaSNBNuW28p4VXS8rKh2
P7I24rXyWSn0ZpPUPtgWolAdwwde0VJaxwkEljxPw0xFHpNOLaj50IC06SIAUTJMdUtvvjEFCDmr
D6z0yXGCV4rYzjQl3waOxo6XIxvsZ1aXSAxkABgU6Oqj0AtD7xGZWms24Y0oGTUv0Hr9q5fmU8Mc
gWHOWHv/P4yUADGtxYy5xbPDN1q3n0Ff5aPlSGuBI+YWNqM3+kd6dA9yDDPcKQGUpH4CPGs8Jcun
4yaJyLflw+ToqgHuH25C5kVAAypSVMNOvjw6pSV0Hi9ORswAaiSJW1dVSuB1DKApB8eeij2HsB34
76/kylinB5sD2IHfUu5BSrayJlGsT6/CG0LvHsnbnCAJ0PACUEmkflUwyVWQN0Rrrx7/XeVm46Iu
rxfFpkJhcf7Pm8AVch/xmICM1s5B2pKlZwS7/fqfG5mPN1CflFbqM8SJz8rQrMjCOcuAQ65uCV6N
uynYjK95qSCfvq00GDRFV082RynXsa0hFNfVBMQoruKLX45b/+vckgt45OIXj1ipIVnp0yzFhWWB
82JQuUw4oTqkb6z/tNkxEgX5L7cZTtRV3bTwT2+A6f+TiOHdisi2UynMwPZ10LC4wtjk7oZStjvO
gcLgCpvh9T+Piq9mO83eu4uDumIl9DUiN69/NOcFEbISd63qoSAQOWab7q3EFodFKdphR7wWzAOT
yU1GMfsEE5JMiDcYrZeDzAvZCP8vT0epKRnL33JA68HHCtDNRiZkvIn6COsKmENUqqE/WuLayHOa
SLFgPB+0eXN3p/5KJMaGCKo8UbqJFLaOUoy+oYa1W9OXayKja2/jRFXOLrrl4Ef0kfoolFWXnCzJ
85u0izt/cbeIco208Q3F2YEBpkU9sCruSgM7yTWr++8R/fx36icJY+syw2q4MNq75YvmEnzbsRyq
QPBFYdeEP2I5NWUOBPcPLbPPBMH47YRc3xBzJMIqJOmfmr2pmdEme+Mvnp2gjT4xpXXmmZGCUb+D
IpGyoBI6t7Ac2MGQz/8QbvSmr9e91VzDJjVrRCaTpa9pCxrbaC3UHbybpr8G6lt+sqRokkMMfNoW
W/i5XjnWkifgY4gqWfTowRS39CuWMT9v/a4gdnkNjzsglrAhuzdRngtCqXhyziQfpKlidTLCHauS
Nm5Inv5Ctz93/Do83HQFOU8TQh658AA7QSOMno/vfUVDfzrGvq9eKE+fjdaL3KoWlsm1WwZucq8/
YZUFQIXVMZ5tp88tkA7UMUybFXQh/5D4+xMFOi1G2o9QuZ/W19Ocfojc8lhZJziWGT04+1x0cGSm
Rb3aT+RKsHSrzxqcr+Bz/FU+98FlYwGjcIpPjcX4aZWCpESZ0FW1ITxRo7ahfMqU67RGwnryhwII
kStDfTydOUa8UmR9H8P+iKqONFc6lvUV39eJ+mBOBcaqdy6dm/1ZxW66BgozxzQp1XTP+dErsbRH
73bLg5gP+IRtbUL+yMsrRQsww2P01IoQZQQS1M44E967vwVBAQxHTyBXkPtcUeph/k6rR/wSn/ad
YtS7opSuMvE47HJYhLr0SM4IYslyPzkw+rtBOYt4564dsMKyLT4vuHMNUAxx9d64kGfMnWJfk3OR
5i1Y7u571kafWtaskZQ4NxnyxHnNFW7EsGMgZoEFeV8T6Ltro6moZaL8GQrsQRaHicJsYy8Ppgty
JJyFtmD3g3XgyZ3RcfzTVFwD0mobVYEnM0/ClcGy8egFRSh9i3HFjH6Ybl93/pwMfEBcLHV45Vz2
yJ7bWdqWVQyBw5NMhWc5VwhPLFKzR+xY4BXQBMFfzmjp1gpbwz5Zd1TazaeikCwXC8CUhN6AwdrD
4uXIIZccZVtUtSVCfDC+1fuNH8wPZqkhOeKffMEypm8U6pXYWW5tHwDnn1B6x4wG8fFV4Vj5f4Zo
HlL452/o5zbg0vn6eJ29KpEVcrS+wcfxfoFM0FbcN+SsAggWZHHiAlV5bcFHCuaV4q+k1tqWpF5Z
ELcXbp5NBaBh83u/E5WQ01G46Zy2u3Ec3I9niAIxaSF3nFcYHEFwlvIxwPDGmAiu39gBZWV7VQR0
HbsicY5Fo5iNFvviCTLv9jxcxpWSLlPzMBLmCMn4U/FMXHo6DEt7/SHbQkByfD8Bu0CcsD9l0t8y
rF9mIRsxv7DxHly0DovNQVI2jfJAqJYky90x6xt3AlPr4Tj18wVts8UbHeEzK53gxrgeIH92FZG+
YhvQRxBwzseoGXqjfPdAfgryPrEGjqYLQ/88I8buZF+bZwU3FTpTInlbBKJfY85c17McueHy0sy9
0D+6ToVwaF0macxmuD98QcwjNP2KJ2DuqK3PN1Yu5KGlBAoD+jKvOkEx6Q4s8y+we59iLLme0y5h
R9XP+Qiz3qWPI0byzrGxHxzQ37x0MK/DNmqxLHvQXvJCPIUzAaNqFSd2B+w9Tch7Fh6zhUI/qYFf
BguiBCNQOorntjx1zFu+3/dcGClWW45/Dqse949qPPbyJqQrpYh/LstGJxLAPikTu+cUwnDm8kTV
0TeGiFtiiBFmoTeoNPuCyWBbZNUETlTRTRCaVD6FVyKlthVdXm0usWx+vsM3AwQ+HHZIgfw8UENj
89dkmj9iyEahO3FT6itF9oPcxLjP+XM+fHAIGTSuWSn08UvUArwD23BdFnvYHAhFT5WBHUtS346J
IEorysnmzHCuD9ILnBeXKkWKCP5r3UqJ+sfAwhQ+s7/ZqddzdLHD9JLB0m5BCbw3sa5jF7c8+vL2
Lcid7yVFigd6xfEQigv1slIuKCX8WfxkBOIy1wUdPQAXjfIiePmdjouqVhsLyqd41nyaYy5H+1pz
Bmma9+93jlwQUAx9I95t2993hGZPT5i3MRf55p44uEdRD8qTt77dNdcX4BtlrAxKl0bxZkLJCckl
YtqDLQNLcy6qKjmr1fT2a7O/vJ6jbPvLWkZVl/oe+x678JRItBngic5H9SgmIEwP35w9cyDXaRNY
d3LSyx/b0UfI++q2D8BhFLV6ligvT2poen2pz9IQgIhIH3YxQv/Z95HBIsowhOoZeWZrnHq/mWZ+
Y45Izsck5zmln3XUC8TEkA4DJhDSivQ46g0n3FrpPfVgDlRBlgkB+jmo1e4quCzUNglzXXR3madi
fWxbu88SJ/SVICepcH4RP4NffBht9b4tfvVabXjw45if28uHdbbosPMW94rsC/0lYh6+Inp6/Idn
1PqzrmmNkxpSq6XPxTmh7XDKBcN7zIx3iIODn9BIk//YxZcgpMaXyhvicbnKoB8jYPGspzBEHBCI
d6OtFtmg+mA4dwDzrtV0AoDAJwqOc+fPK93tgf1XP2Zxp3hDVXb2IUlIimAde9zXLWxlZNGHeb2/
0gM2JLfeRTVsGxWGMMj2585aZzVupgL03SC7RemL/1ty7Z/a05oiendLYGIGP4QLebTSQFWphatp
G2bRwe4tqhd8JVWFx3z5xdxDvh5C9ObBX2o+5SJpI665BuReXTPgIjKYkK+VwZPc29GYOI7EUrGP
CCKA5gRZDrk5fdq58zk/00iSMRUXzef7mhcV4FYxfx0Ytc8USiGFdul9tVTToN6VrieW68IpvBFt
RQzkpfoe/x/w4muE91XhDdSWEHNfl3bIc+9gg8rloaxlU1Ad0C6CU72OcAkMQUriy0mZ9rj6+Agm
Ii0MO24I3Ha0q/AMJol/Tf1IGcmpqTnGwvN0upPiLWj64Ilnfqd+WdMPFJo3aN6pVdqoFd9a4QZW
bFp6smV3o61iVVptS8ihWdwEdBSSvmuEDhCGCQ6+6TWZm2ehRgrvO1Fl5niGi2Qs1a0yXR0KgH0P
cwDbJsUj6oqspG58DdwDa/+WyNljpmrZSLJm8u4C7mQQ1BGa0jP6VMqeD52I2fHGE/U2XneMGqp6
OWh82RjgVqXBS7K8fDZUHUkgsz03+JEdCzgY8do0SlOWGdyDIgiMrDsf7kjP9oF/AAyA/mygTPk0
paXtoOz1Q8JJH3eSbVnFQp+lk1jxKxAyjORkEY+sJgQYXh5aSqGN32JFBJJz+vIodKQED9zEzD4R
u6r/OppZyfA7Tjt+zdsCMRHQKEdzVs9O3nYR5hSBg6zZJk+tse9hOAEXuYLocUGmMHoD7QWZjl8Z
yXYw+g75bR8SaNvVHB/GycR34/8cguiog4z+Lj+S8FmD4icCIZ/gbO4zccihPE6h0lI/PLmvRiFy
Dh++0TVi+T/dEkW3Y+0y0sKoymTpAbMz3qSaSw625VDDcx9+HgP/zlcRDL/6JSRbAdtuUPoiw3Mb
5CqbSrXQuuPKZF/FQRiDL5Qth82ucgh50T/plQFjTZXMfLPImm2Wc/J9/Df2YNU/+yV9H01y7lJi
DjW7/dNAfsWtJJCi1euolW7InK28h/e2rWlyXXO4eB6LYT5MJppE7zsQfXXWARcSW2GO5T86bJsB
cUkgDRrurPp9tlBebNkNsZo1QNov8ERj0BkEjQacC1hP9/hb9A1qyW4ov38qJ8BfzcKvgeP9LUgA
T1CWHhuBdoN10UwNhgN7jkgxsRzrW6KYcVmPp7t5n/P06GqhK9fQLOxSEwQtZQrTAZxXdbe+O+i8
Bec9wWivefYm1TVFKRYLZfrj0RXRZNV3Dzs+0Xr1R889OHaSJro17oha/OQb2z7WFwrJJbY7UAft
DN+rZwYHPm7Hb0KDegGk9fUWrvFmeMqWjj6my4AazhnJpOX2qVbT8NjzKSSyJiJlpYyXIhJLt/g+
Q1bcz6Ce0CGSWRWN7CsTsjuvQP5xqYSN7JCoQT/iw8M0RJcMJNGmBukbYg9U2stgDF6ajjZiPH/v
prhX490/dGgwib/au+8qfpoXpCa1asJFHtjfyaOEI5ygVdzo8ixIebC6G6rLSqlA4bYZzN21BVQa
xMzf6zmAiAYz2qGDpsbyF07FygbCfsFouresyuavMhCF6ELxvHB7Zuke5pzKlm1QmWWzSqU9xUY6
D+4MxhydItk5jZ/EWAnz8/w2XPtfZ9jvY+780BSpPmFXzTWzOm4Cu5zZ/+bX69mcH4+XzLo94jHM
ZQDoqYbQJ49x5Gc8X/f0svatLnaJ0WzSo9q5wH9ZS89jMxUioIGVybQeMJfAw2Qi0dl9Z6NPfr0R
UGZbIPiT/wjc4yw9Z5h+ADW6iWVYN2MFOtdZpA96w20ctMGzCmqQJBs/bES9+ZrvJxA7pgdb0TrI
vxwXrqH/SUgnIzB5diexuu1YOkI7BX6j9i6S+rOKs3P8hJYqpead62hQ65HUWxR+4qc4suP31pot
jSX0YRIoIvwOgtlA/Uc6b49xoryxuKDzM7vPP/Cq2A6RIacpnac4N07FAF3OE9rIAPoL23RfrFpR
6NipJYC5Cv0uO1NHRpnaiPLEBkhf+8FEF6Sit/Xa7wAheL9run6QMPnQNKCHQ/q9c6uiwRPr+wii
TmqM9M1J2USU9sAFCMHZ+4Am0EKScIiUHqg4iP1yt/Bza6bM9CWx3QD+/38FCi8iFUSzYQRWU091
QTfTQxsZJy5NovfoEiZDCmpKBv8Ag2M5YPwoUrAgGc9c8UvBXak52ElQRM5YQA21zxYZaHdfvZEV
JRZcRjV9LkkzPLiX9fa06utrNvUVh0q0D0HclxfZFtwFjDDNOtPq0ZbjzhWSNI5HHvds9KccyVra
T/CMRzKADu/vZfCUriJmZOEd83FygDWnEIESDHziz12V3TV/qlA7csFSfmgKL3VK9XMas/ju6PWF
EdlxwkGQ+Fg7upWlGLH/3xKYu/SqsoBeqXqhzdjaubExHNLWlOvpemUR+lt/hX3nedUx2myOvdT4
CVTmVkAexFiQ662a2ps+9FjbjQ9qGyac7aA+VbEX4ox4JOoW7jsjS9aBL4PgNu5rbIcOIEIaGvZk
7K+CkKf3OIooL5tW2c4JfQZ1AQIKXZL+clxUFGSl8SEjAsbG6kH4lGWzoL6fjA0xRm8EoPSiNsyk
XbN03paKZbI1DSGNE1/eNjJulp88vJiY/D+AfP1vYpq9yq4TdWb4a3/MHEOinjdEIsrKPJJqKAUe
s1LyJ0jLcqSF44cRDxwSjqhv0QikiZcU4CRbRfx6LcHWKyJcwK54IwplZ+cF7OpAHn1LdNJ6Lyiz
UyFaCmFXwELbrG8NX4f3ARJUvhCkwKtUk7MZ+AnOQ50Hg84Wqza7LKLChtB0toAB+NPpGsXHiBBj
SkTddbsw1iRWWvmf3KPucUaR1p5CK9VR2G7NH7VzN4haq+vMpAKDWvqv5iBNSTHNNE1BxtjPwBYg
3WzZaampKOZXICZxT3XFiO4q3duCnJY2FmjQMzKV2DddMmUJHKTGWmHMnM/FI1bgWRH8O8qiutpp
pbYa7PBojewrqKD+v1bb4Zmm5yMiG4mE09YQCgV5ZS+LQ9q3mxkh1uw0ypthWXz0mw6E91P/xasm
TC1QKXF7YnvLHazuNyMg/OYj6ufQPZb6QPC5zaHBVOYTTl6bX8qh0AK1roy5hWOGmhIhj+By8IVt
KIVwWA6je5IVEpar4vh62WZBGwSSvQ5SBuRwnbpINwIWCUa4pmgpSsw8DhZHFdFxq5xwf+odCikE
9UbYU5PcKG723y3UTYGxo1yqSwLrhjzJGOO/g42kKaa/frM3p0bUaFAQ6BJTSwIfi/KdQaQl3UoB
CVI1Q6mu28TZMcsAk9/hYdupa9vBhXTaLA2vSuFgry9guyJw64iYq3oAjyQELoTxwOXEHBCMP/04
oKQ+7RCUh+4uTvH0zHu6TMlzUjPQYBy8m0e77AYtx/4oyU3b8iSZPi2ltnIdisAZdEtMmeX/xwlw
qPCn8DwsiphQ1lTYdtHQRMh9ZcwwThM8hMhT3/acSNMHH+IeTb1OvUw4+aTYp+KOLDjh+sFZjv1V
IaEwtW7Pd3ehKhXnOKHCJ+LzvQLzIDeZoDzQT42/pgPe3HIX88ZAaYTMjJBmYQ7fP+xuTx1P672w
MaJSrdXXMphqQ9zTF00o/qKc63cSm52XrPi6DaY80lOYnymfv9MFzs6fq9bWJ2/LgVN0H+e1GReE
IWU8lQOooCHhZEqbgzMC4j6Zs02U52RY+qwS3l6AEw/KElqgxGPRHoRuBMYKY4olX+1k/3It+rqJ
h+MXVEFIqW4kwsG9G1iW1lWGYQeyq4lanw3OYKsPLf27UH0GruDgB7+NisP/V1kCSH0Gpro73v5J
4PVO581cMYKNG2rPkG2ZkkRwWwPzZRqz4f9XZns/cNpzT1c21bJv0JNjNWd+fbgjm4eCVreWihVU
+frl15JxhG77KesGQ+TTS+joGgn8Onh4B+v3tKfG0DihYv3jBINK8HrOHoti+EvsJZxKdcXAGQMm
WPQPmgWab1EszLN+U548xe8o38aL0v4kQRH8ZkxZr87U5BY+8Ek9agiBVew0gwbIhKb7Cn219Ben
1cBX8SL4OT/iNWjWm6wt9bFNYATWpsfhL7fv1P/CBxnlVbGS29ez/SSJqg+1q88lHJYHEMjuuIA0
hwi2Ihh/hppM2cRjfWzretppf7nkoaiM/NfKzi9JffBit+uchnCfTCoPQ0tdY/dcq3kVsqe4JA2q
PkbjNbP5IniFQ43p458ny8EriSUpiSaz8WQydcDSvkIyZhoZF4icua1SsfKRjbelcui6ur8+uqa1
TeAGm4v0GyOEb1KF92cBp6XS65meS6m5v5y991lERJ135ilhRhpfEtuIGcufzo0Xl1T7HMUNjqPH
f8HiEtJ9YKXZdLlLPxH7cG8KTedcpEufrZKeUaBuriiskS533E4i1gx+nzbv67yTsosMvbf1Iq2T
mUnoFS7ERknDEDcMo53qMS27CxCq02ClMdMgcio4iHEU98FMBjQJjekNCo79/1y0n72T/U1AtleT
RYj5/7iDqj+PCn8jJpFEqKAZeTxqheaZ3770X4VA+rvhzPySF4Tskr58tafbtHrTvcje902MjSZ3
jhbGIMLsBaWaYvfRVadAfsbgZZLkQJPvenjXqLua7dotB7CVoUU3Uf9037R1gjQqNp6R6CyS0bW9
TpSsXZGU5lv3JOGA+6hiyqTbpO62yE5RA4bnnyT6uQtp+VcaXVbbgN6K82Nr8/hWJ8ybtkKySzvL
cMZ44lLDRhTjZ5bPie0AKITLj4XYdYjfeGSru3C99Bou3CJ+TNABW3pjb0ycSplzuj/BA9AEAda6
yAYB6TVbYM5HjuPrZRlPIRz7xwaJYxAPKTSkq4g+ndaPP+NZ56rD+R7m/T1UUMPq5OF6qFSMl2j4
teCJE8BrNzFnaf0eFjG0GIHHTEI3bC1vMBz728kQLXSjbW810uQ+vpw2gmrc4WqGbDJoHxJXsco6
c3fZo+sJXn1eum01DvDzwA6zj3sbCaJc3wqbVoSHG1OnL9ew4TosuSWCMMvCqtQIABOOjeKFoc0F
Hozv9icyGlIbT1jx7ZAd9/VJ7CvMBpWDtg4EVb8LxfhZp0U8cBQ/xr2ZJZaRj5RUlWmE9Nc+D9e2
aXN6oKqqVjACtZex3k3kEpFqQxLWtfoygijdBg0btTVgjoKrUUVAUFgwBTcctS+GJp8s73D6ER4O
0HJqCgexmCB8xuFHdXhe7DqkvsGozIEAcM1/RxrAjmy5FGQim4GRM1HrTtDtH3EW4PBqjlNSq55h
PskiNL1yB8MV4Ni/pNbmn/7/fFKNlblif4NA8JxcUFmKhZtpSMZQkOb/eAhSbRF0lefa0HSKizW1
PQ00atV2jU1NRxTJp0D+AmE58zRjRouR5E90J+RqPLlG0n/WvykbDaH69qmU4Q37/h50z1FjBdKE
tPDfS5WOCjdXdM7TUE0BxgYF4OuKFU1pBjCg3z4q15adXwtGTJ3M+syil9cdIaAWUU9I1mSUSQpW
87LVvu4+GIpFXCoE3fXvKpg5/DN0K/pHEa4MxXSdo5V3PP7szAYKW0EiBRpLpLh6i0CaegWG1Um1
CxIWOSJuS/24RNwzVv9WuJoQnjP3EuatlXHuBjziM3uE9QITa/GvZy4RJjYZfqfXiymttL/kQ/wW
pDmIuhmAfWJFkuwRKgtCbIaWTKlMLfKnX2zAfeT+HV/qcA6wv61z9ZZTeNxq7y9I1T1MGnxN2IBz
Fj2+DcgI84k07FSMAVFd2KmNZESXJsXVYnwpDYCwF0ydcEmLEP01dkVM4Bu9K64vSH2Mmmty/1z1
/bZW/SXWTyFgevy0dHEc4BciUDflPe1G9NJBbAfcISJZU/WUMjXJsV/0ti0YtHXeRjIdjPJJmlJh
JqfNcV/5lPfPR8YzRgpsmbUKF9t8WYzczP1/QZ32dZ3Jk5+HJra0qcssNidniyZBQta3gwHhJoaD
uvKSpKvwxGyR2TafFOfk9Qs3X/5lYYFFNc1p5QhBfeUUN92D29U593USo6whh6FVuA67D1k9wibw
Y7x3VU8bE5Q9nb7B3wesn+UBjB7f9YMpvGIYQFMLG+J0goZEsKfFsEcVJMjKfPnyfNql+vxgNx6I
xDL3J3ynT5lolNwDMO7F/iwMTsiid5kcz03uFn+zh3BGbZakEYCD0bxNmF73Aj/W/U4YH/ZmbtDI
rTSZA5gF01IWFcyG8eBDE0stiisj6m5PB7GD9b4tTYGsDPVpcEm3wCpGl3BjXLY35mdxKJEG9AjZ
GCPwK3glOlhDcYh4eSKfUKFfBNiwJxLjCp04vXVzupdHv+dFqHopUjqHp7Td/J/XxIOQAHunboTv
F/EA81f+J4RJBlr0pblOPY+UIgHijDnNBJmLR0+IzjAriSEYa/A2XG1pgzWvet6PnS4FmyW7Pwxn
CspGfLfnQU8dBr3O8nEEF26z5p1CPhsBzIRaukRWfnvN0y2ojiESOwTXzmat08DdKGD/Oh1HYdi2
qeQ2FoVljdGFpzvhRlOK9Zw2noGXPzCsrgLWCCtAI+QjujOFSBL27XtPJMqAeCnSqpTtd/k+LIM0
FTu6/Y9kGHIcFSztO8IETiTidgNMy5LwGBXM6vq6W74KqtX4OBpY5e3fiey2MySmz7SGk0qvagf3
T0E1WKfFP/Yfw8NhQhWr/PnWgiXxsn3nRYGYInExzP6MrEHCekm+Zw+Nczm1JrqxROebJGqYeXCM
O+5V6GsxkgB+WGpa//MzVM9Qi1D3BXxldqHDGeOijZy3+8w2f1o0Xww6WYJh23qi2XoscmYCeS1g
9FtL9Gn/c+eFLFUZ4lvYTsg6IFV98l6GWvRDY52HNgtT91ZEqmsDdNJ3tHbSIf11jFkwniPQc67e
xjeWdqCNRNW8deVupuhi3y2iq27RokUMkL2rRjKm9wbUGsB48Je+1RY4QsEoFvMR5R2+mOzFPLb2
ofYDRRzI9AFVyiiK0qp2znR94bhOB4hxHUwMTyGb43ZJ8QhkBbobnnKY/npH82lfgxoSh+W2htH7
SshtGL0NW70SK2pBtnsccXPQNHVMLabDYLeyAcJ9HQKde5EZ74ifSNZSkruD6pTShLdFTErjwsZP
tp/eonjWcuI8Pme794/z4i3xlhJEqVloMS2rIbCFERO/LcWaAM1h2DUUV0/QGAkH4zknmv1T4HCY
WhmQkQo8af2sW35SlMUp9zlkBugpe+yOuFCfS8o4auekSZsjfKkz/E+ev5+UkmHXm3Ufy//5ytT8
+66sGP6MtjBQKLe15dszxYBQGeb2bxMISbRIB4JbiIgcGufT4/q0rvNr6ZkSdC/oIRAGFLxm7D9O
QNX4wwmDsYIrcdhWu1Mfye9Xn7/wpnlgzS3Xur2iwanxTXhma+m1yJg0xXMNXWjAHNFI4FKbf2fR
XhdvV6jxKxjoE7bndaQYar0/THfYn3lGLA1YDPFT88OrcUOm4xgQqfmMfyLmqLZ9RU7VkZpzsty0
Gzp297lNwaojrFoVJQCC0vYvBc729vWW+5tMPJV16ikPrjQwIKrs+BxhjBjmcwRE8bMHCuVMh97p
xMb2HrnDw2PVQ7IICZgHavvKNT5jWC2ki6jqeKkyPA2wWnVsJXJ6e6BDdeM0c48Ih0K8+xAZN2eN
YiYPCkptX/VOJR8t1zMz3LAQ+XFSaaq6Ra24q9pJc9zes8psFWIAa/yYFk+SjsmEMFKsXodEB+Pl
xY8M9AjzqQrPVDGeoL0XAyHZuBKFPPoTVrnnOOkcz1EBgFsdp4iSUo7jsgeUB94hlStOPST5617e
mlCk1iBnPZ8mIhbVMpLHN23Uh0+UsAtybNvFIsthdcF3vtUQxfnXu3sLB8ALqSZmsH7bjIpxqBSB
O062lyHcHm7GgKImX8WDzQ4tDaTQkeqAm2sZzt+F1YnlLCrC+GHvgK5DjBnqyfTgheZdhCtaRuPK
t+27t3vyAHkmkzLI1alAa3BUxQVzyDHCAXfNo+5mOEEwIkwcFxQaA7mFTZPZBG9ad+4XyeK9lqlI
xZ7tOLEMhWj1HEESN03oRaY0CYM4PHMFHE27VsSR1+WmQL6ldkKaD8EizBuDvTC6L1LSoypPmBpu
X5p7fMU/cQT75TmLlEzrq1AipCss1k6ISpdHr3ZUX/coVKkkoCX7daV5+9CRpEw3T81OPMfOUP9X
YCNEEkxBs85BfWRi5dS9pvT2rD0B3I0LFmj0vAsvlclYZ86+HfyBfngf6y0ESSLPciMaC6fGj91+
qRqJMnGVMcM6EyODgE1Cp5JYKszkbws6gD017hWfpNe1WefbhmzuybHqaCYf8oZ2/rdY+ubdthK7
daPUs4WOHzozlFmhFRVK1J8bNYyVcs1hr7Xz+cpmp6QRxv7s1I+FYuZ5hRPNU9j3/v337rVY1MyJ
kQqyb69x9AGJDoE8Xeh0dJ3Dk7KTBy/BR6ipUuGSd23RItZgaD2GjitFelGNS1QkeD3aXl+R/4bB
FTFbHHMPEms7/FoMVb2qkdbt0Lxk7qc3sPwvEufSp3ldn9157OJav4yl4bE6hMmih3C8CbS9AMCT
uoxX1CNO3rCPmaDsKF3NcWrQQbr7ZJUGUuZ7xm5GksGvnQC0rkdxWTimWXUe2RWaJThgSC9EKHkJ
MczIOVDKoCb6o9BT+kz7wfpHEJmgAhKjT4JKv4tAhn0H4z6O3gRQKwz6dU3zpSGlYEjKWqBxSUxz
1BL2iUidOSFMigj4tpS6CFYUvpYwBR0HMjVkwcHZFuJmeqdgj9bqsHeNCD8x3P1G6jPLqgdLF1un
9xauWc9Xw57lTFGnfqHjOUYMOakc7Scq4PTbvtkjfnNDQkllCvRbiDF/chQpi9DTXns78K6cJ1+w
H3C3A24KJWaS+UZt1qpjVrkUTwA3aE3KWo+RqmUMAgMIA+nxP604kvJ4Ihf9JxEP+Dypl9Xz20pY
fROnm313UC5VKXkX2609bEc6vtIEuTKSgxHq4fHIHaye5bfO3sFnYAGqxtYjaPqSfWRHMgRfbID4
T4Vew5xG9d4bTvSa9rKHifhCnij42EZXD+///QvkIFnKQl/VFdUMdu6MoSnjws/1nGb1tjsKv3C6
IjqoAInWU21TgIZ3V9K4m70diuBmGPWpMStUptTAslM7aFwlvhBwpCDBP2XsGHfeQc+kolNhzgNV
phbPUb+XSpOXhOjcDfRrPGsl8p5qt91e/KZgrAN9RuFU/HhBcxr9BQTjSieoYd+JeV2eyIr+i32O
anQjWYJjvsYx5RZemn2+9EkUKY94Y3s12t+A9Fp2w1fkl2EdRpO4SVHh9xqG0FbtmuHgK2Rhhv50
Vx3MRbK3mZ/XO/NopbmFk8yJBzJfAt6Je0QDc5RXU6wIVF8TTGecuxH+RDEoSt6lyEpiLHSZZUPG
i/EzqX1ZRPI0jZs494lR4KOkx005ul4PwImCpJSz4keVXL445zCCu2vqql0EMGG7Pd3lMRm5Pnpt
wrRmxeImmUDbiJFU62iHFWkWjpP2TeAzy7HGDE1CNnhLvzv5Hwdn2lmQia8434KSlAT6ORMnKPZI
ZrTsT5K2IgIlwUgs/OS7Y5efhfurnNStJDGqGOiGbMbGXgD0um3/SQc6eTr2GLdtkyLoMDSLaFCO
RctF1o0yUtnZkXtZisFpdttzOPITYFjKZhz5eiOa5nRxfBhAUPr7P+iikqJMcw45GH9j6LvJVVK/
oxkmcVOTebZhVy7RnPW8oU23jUT24r1dI0uVUwY2Ter03DADR1tGG2CRNDDs9ImvCESCk58T7AZ2
cO0/feoPFxtN+HODqLQJOBw/VN1RtK7tSAAHzSeNpPXEl362gXDw7JACOt9JuOPzEG72YNxTc+Vq
64zH6wihhUJV70hZJvKmWZJArBLS9MhhL3/iOAt1PQaV+2Lv1+Ke1Z88nHkFwWhhb1QxynEoid5g
IYgUwRF4sAT/C8SGAYIcL0eOhgv07U9QJKIb2ZOq0NXHLvbLVccx+YOmuflNS3lFK15sedniojkz
ek8EyInwm/cO0oYfnfsmS89pTAM0++7bh0pmsQpfgjfT5K+dSKNX5vZ8y8OjgMPq+8G1jclBFXmU
sEdRTkrRDA/kEeQJXHlgn8hMPP7dbszUOSZLDdlcfsC6m6FEWV0y07rVE/lD9uIVfTIkYrn5X+1h
eMODq7WBaf+V/ZVlgReE8vJAcWwZB0Z0ky3as0hOIS6A+qWADHC2LeLepR7V9miqJgoZQcSZHe5v
AdRme5yrN0W75HAd6uduc4botw7luAyvuodySeTPHYoCkn18ZqTS8mNE/ty+3iiiUM1KGKqN8kcs
gc5WT5RK5m9ELx+9Enix+lmkQjE7nQdn9O/HepIc1bMs/JgR5Mp/sm9GrvTzQjKLkWPYN4oGGrgX
jgCAv7mqdeHltUgNycVNO+el1wexQxuGjYxnHnCeFxsGpg1JK1uXjznjpNWUMmL3brX/k93s8gyw
HOhV2DZuCvLv1baAqBGkLnRMbLnqhy4AFK9DFKAyRNyqdBrrMfFVYNL5oGfr0DyAuFH/d1QsHwkJ
42QbfDQ2DpcWLzaljV3WjzAaqgPh89pF0bohEXfsfXx8/KQurEjf+vXQcTsajOgsRm4P5WXff6fg
nOdioVheCx/I7FwZU8g6SmtqybPDsFnh7M87VSTAA0tVmxflKPUK9fXdQgmsPeuzkhNJjirrVIT0
xRqV8BasL0yXL3PSGO9vX0UA2Duw7Pfg8FaLmhVa5y2mO33UdXasVdQA+TPehYDNvpu01WECQFSC
9+2wo+HBq4n09ixkrC4FgsXVO6HRsh5zma1+hvKoJZSopN/ucQleyHBr8ilMsSuX73KSNyVZKMj6
otcB+pmPvp7xPU3NZwSpiUyYKF//uTRyl7R9K7arB0Ex5avP2IuMldftvhnFdnLSIavqHsV3BDVZ
cSUHueuxwXRAq1+bkuMw2zxxsKTFjCAQzlE+ZryAbT//8XbyhAdu4LqOlcwG/MwL7WfqJGqscVtO
pFkS7Ta8w7s/s0uXPI09eNrnnJET+mUKqX/NKfG2JYv3hwu5s8W/+2tWWvQqAFQXh3oXBiOmBO/z
xAbP4eRiC/wQ6UoIxZeOKrZtxWJR8PfcYYvMvLM2CyqgK6mS+PdGNEAsBwx/NGJ8Ewxq5wq+Gul2
nlWLGlN4ixxpscRXim2z67wpDTEIJDDdnxeDjdRqbVmRkU792Z9xb9Mc3YUNJsygiacWlZ+Q4etw
5q0sho4LwrazlWkJSA7WN4wH2dJJQFTsmkf142kxQhHEBgdpEul2LNffp6wccVsoZJEuQ3eGCQzK
+YF0xjTUodYBkZy3hij1eWNj1UpkEmYJnETESA0YwU0Wfzt5oOogHBID0usxQrR0EQVKSDROpiJK
nKfWqNVrI222cKNO/5UB8pLeApXGbX0C1qFdS0EwWfUr5NLBrHg8ls4rqpP+RlDJ/bUAVxU4oTEe
FJWnrpl1CThFsb32SrhU3fC+VwxrJSmJDCu6o8BTw8yEZbUBd2CxyO4V+y5wigurufk8JtFvIaJ2
EJQ/56w5NHf7Ft7EU00Xm3ubVDJlUrW4ur6oyguFgYD29QVXpNSikI5l8Jv1vTng4tbCbM/k/3ps
QIcHKdueJ4hpLxCBvkvRkcMTXY5w6Aj6mS/otwAIoNP/VIH3C5BBnipb0nq9QLGx/XQxYjraCh1V
aX8STHbwgzpZaaWaPCNAUgMoXqghThbeRsqYIfguSXKuyE97JHmRzTlKJpeaHVJA6mDUlMmbNh2u
XP4FTG54HWpVGGlqR0Mw3odn3GzMeDQdryIx9P2UImylUqYQZ93uvX5nHfmxlVNnXczoVZmB3fd+
eHd+luaptVBMCVRFKYx7Q1dILsIEynbgZGlBsVvVY89aovUo/MIEsJ1SbQ1GPRzsSM0Q6KHLFigD
IB55DPSP6p5Z82KEqWEz0w24Iuzh2dkU5yRbYZhU+YebP2oteSx+3cuux7oBOYK2t/FC0Vf3GrmT
cDlBovaiqonTd4yvOM6q1Cu4piKMxYSlm4LvvvsghWCfKN98QBBh+KeBOuVM7RyLIY1Kl+ABlfA8
t/534TlAf1Y0kZTnV2xGKfU/b8vr6QU/JdaKxmhUbja5ZzlEudwo8+ATk1kj3+K/q4Mq2bmHowvs
oOCXfqnmUGC7p2qUg2yAwMu1ApIljL5bfJVYVtss8PxOBpKbTjq95gd/LTobSw5rK6aCqjZgguBm
0axwcxilUftFevVcUu9mTRwTZzAJTNicsnhX58JAq/i7heE22rv3MRGmzkNtHMDSw0z5jrt/dqbY
hPfSpj8ng/webR68VCVCcz7T819JbNqFPSU9KvvUl2/5IMYFYujzsAW1fWPiGU6gvK73TqYYBBsJ
GsdLD1Bv/00EJPQkfcAW4iB8TY5O/OEqdN7TeAsjR4fTqXBkUR1nrKYkCjV9R67tZAtPfowR6ysC
z2oofDfz69di9znBnpyFV9n8SPnqpW+zu8yo1dEfRwDpUHwTbxgQwaYnqUJ3/kEwNVB9z2sSbrp/
6Zv9IaCpGZFZ/Bc8R+3UgMnpoJCXsSAOJps+6nPE56H6t1cHed5I57O5qsIjOYKX7WHrxhaEilxa
48tCm7Ojp0gXaxUAGGXz/yytoKoW7Bbn5LXxmod+2/FXVmJ4GT2ybv3IUhgV+sqPlY7NQNBsmvDQ
W1yjLzDRi8AOLWBbT9AE187bLsKI1bJwPJUyLMaqEKFnigV5mnFnfbuloIIyzYo7LXOiz5wDCQxL
YtRobH4D+EkizzUz4Vyz7CChuF8sGpK7Hy/tEds4SYtm6cDAdkpq03lz7nUsOhoNp9ciDq0ScnsY
1WFckHBwMPwbQXQfkQ4aRD+LEhdXdhZWpSAbTY3CFJOUgnc3Ypg6a5I9xJJIxPJuykoYxDDmTSsl
xZmkDaYNYk54nA/CrjzNU81CLmILK9QXd3x76YPHFa3gTQjHXa/f49lRzbcuC+EEmUYdBwydLbSr
l1dFMP+8dvbSJt7r/ynI2Aw5yHUkwxnmU1r56bCgk8/AO3DBBO2YXnDrIXI9ip/IPDBNyLbuL4Hm
5s+vMXtbG3K6VyAmTLp0ONx0bsmYiCLzihVE9TxccG9cWMg+tkMKVxAoH6AmNY8XJ3k1B3/P7Dm3
9yU6J8er26xkb5lBkISDa1eHeoZmGxeUH7oPTz1UmBq8wCmmVfMIaf6LJkYDdeVIEp0F2XK5KnwM
EITeMqn2In+opVJx+dXfW7UIfZThKAx/eWUFuKvt+Qf9luEK2ssllvrqOavdDvN98YPgfTqSQE/d
ElWwsLBPBiRDWghyorSTxRe+y+VBH/UB0nBB45N+Ar1sdm5FwLDt6lpeIela+PWWnMNLLk7ItU+M
LpPM1uBOx8roRsc3iOAHFbIkwAIVcVQSHANCKRh01/G0YQ7iviQqCOFA2uUi2TOPeSWJhuITTcM3
83j77ZOL1qBU4Wu3NwjwUglQgyxjl0gUzl3s+tNsWeMn0NN3T88/F5yFeqkqm5GMIMmQUuhgLp1K
vwAZyN38sgXnUDiQV/xXH+dFR1iY4CPy6DM3g7Z+5ON9AAoD4JND3drQCVzjGGr0Ty79nZ79JfqV
mA84ZVlb5fWaZvvJDOALptQMbwgKRUun8E+fC372MqoFzPyy6QkolchqU8B+7CuXJAIXLx7p0KrK
HQJEaV/n1Bz1EW5sOrv8xCQhN7mD6aqZf2L0iPlT8T99YbG3crXXuxm+sD+NTgOYc/jor48Ksbi9
8tO3fVBGLAIUVphsWnbDtjmxk8Kc/+AbmaLfH+bEHGuZarynCnJgcivBTRKWA4dMcBw/qu869iCX
TMORqhYqcFTzO6//Y8WWxutqITZ+MbaeCMFjcTEdqX1H7Z3Yc67jFKE+d/7jGEdRosgyIG6WcrXJ
sz8akiMCvfi/lMiHSG5DfmDrl/a6OuY6ssnrHzV9ECdymbPOpkHoByCxTzANOu4MYxbN64jU09jC
3Tdk1IuRwppWXoWiS5psahhpjjBlS1469vIzMHvwQqk1t0l/BvdFfOQkBhhKjS53Hn/obROrJSvh
J+ad5NpZO+7Y2L6EvjANPwqO19O5WxAKosuL6aaNUBUxxjLL1xHNjqPxs4Suj37SpUwm2q6uJsDi
J4glpWZtajRxUYDvkYD8p4Tg1HXvdGZznQClVyWgl1QojkL5g6OxFr6jBW6fF0MFzHLHHlryYcCj
P1iMEHXp/0zIm71+G4bfPyGeQEuFUHfoS7oDFqdTHgWO35ThIe8W643RFUEqBCnpjnvybUuutDO5
n5sAyKlAoYdASqJE7Ryjw/uMyc5Qb3o+RB2D8vqv53BMHRq87cj2IYahsq/vwW+/pE/0gBGXt0hT
0XyTifyIZRheSBQvWBQ5cOthC4Z4byMGwHZ+keEW9OYIlVlEB+sYNXHRJkqhcpYoEp6q8c3AQiIc
oD7k+JL5mGOBxMv9f9g3L/BBQlYfnTmqzWH4e+R0l6UT2txxVey/tDxdWZ48ltM6F4s65mGOUUc6
x21xpJ1lCJxpFAVSGNq+mAk/s1xb1gpnmp4onvM4bbtBKemyn+fJHKXT2bm6+8uvIt+hrgKeyP9E
XBl/rZGBu1/8UY7281bw0RpwBeesrejWxam4MOkq7Z2j0bX3yOAOgzBRQK2clcWSdzpgMxlOX0WB
uxKNaLIqNEvW2KtNSWKbwUTUcRheJ30T9E7MkzHn/tXpCBrDzbPrSXbCzx1dKxUgBJi5v93rzPQo
pAhFax+dNbwBiJrXWVuvp4cRMXm9JsddP4+Dn438kYek6kt3aTW1eFLZ1Ns9uhPuRARt9F+f+8gh
6p6EIKqbLmR/dzj3/a5CaCcAwEYJzK96+sY7CDmGoyQBcMiC8wKC0P1EOZ8ZsUDvMc4m06mYaBlL
b++Zpp3DyvnC15zvIU2hzlz36jsUG5I1LHpYzqVqBvv8w5Sdcy1D2kNso5Xk1kOmBO3Ga9NoN1q3
fUIKSSnVaQQ0On4iH4D/J9/PGi03W0jFHrcS3eS0/7kDO8vpY7cPvLCN/khsn4jKpZohaEa8Yqtl
VWzCzwGQrsxvTtYI82dmbPV2Oob7+XPMcIlCwoIUsi0Psbyq3QfxRWY8v/OSIUmYMVqAeF+EzqlU
LJpmWGkEyKT8yzR/DJ73PzDyqlP2MjkcrbRvsctUyFA791aR4r5MMI/Okm35Z9mG2fCejfKLbakq
7nb6Pe9s4cL7vTfL4KAY9Gycb0ge/iMrDSraKJPdJyr1j+L2PGSVQza8242HqCLeVGIJKo9UvB8T
It3DmAkNvliDpcLNVyIux/5Kkq0CY+dO2v0XGOO2fC2SUb5813Ctzm9oyhbu+0g2+DP7IF1CysVm
M4FfqvHzkrcxgxUMYsr9NY3YPtvYDWoRz3Jtwl4uEutiabK+1khfu0AnCAIg+rq/nPRkgAQSHhjr
1YWyGkU3Vu+6U8vO29JkS+sCcQZYYXnYhsqkxx4SVIvRwgFRkYf/NBsUlpAj5F0X8q0WU7LsjoLq
6P3bUq1DfKDupKK1Pr/ZdEzJqq4tf5V8EZa671EJi/RgIcJnRCgA9uSiwBkfW0PvewmHFRknoiLd
IVRn4w0rfqQQtze4l2CKNb+BI5AdOKXyrMd1MP4BK3Lyy9po/Y+3s119Fk++JLLFisDZXKRJqQOp
OG2gaIMScQ/FVBYhnTcCM2UusmiUXOgcxlM8tjOWs7df75qFBAZahKwMk3rKynTn7dBOo173bvwv
fd/CeA2THlb1UlJ8rVzx4FKrtBIqSIpTnV6TPpzNfzgGdGUAcNZRaq28wIXRCXQ+H7PGHwHfqhu7
OvUBS209Jemk1fdCa2jUrhQXO+3lDv2nKbuvhRpc6RyVRnI9rmAJ9doU28sGNu6IKvkiiM0i6RdP
Rl2djkqCUKrQkBOlrfMd7F2oFwyjN4KU+PuHhbFYO2/vnnDsEIrCIiiuippJfTV+QuiKd2iYLmC2
N/b9qMO/PRYo3t9PzCjpUgGc/Axl8bUjCmPXW7nSr9Scwr+S9GVUYi9AjH1FTk9/DPDZE2pW1MVU
1+fhoERfkvhLaQwNr7oHR6BvG4Ew9oVTLUiYdehualbDBnb0k50IEw/y2eReANIpgz0BlfPax5mD
kMJ/iV3bT3eD4YThbynld381OjZ4dQ+vP8b5fqPmnS/vaXfrHpHQjLUryfm85DKKG1wgnCDiN3hS
gzpQvtAO1deic4zisK0KOUCMJff7fTigqGhj6B6uHS86DTCWi4/V+wLLw0tA8Y+QK1yTsdhpzL0O
oMu1qwOJJP70oigCAkptFPmOSlTfdQreGnP2Vea41jHYQ/GIwxOa8osRsPlY8amevG2Tj5T03Grg
hG79AW8bDVEOvWgevH9MiAv/uNW73wkexXjA7cDUW/isF6z+VYnDdUYPOccIqVXokRzLQkEyFGYA
nuhB/VmEhdKTuQk3z/gp4WWulPE/QT5nUgalhAqPRBoUjGEo9Q4SIN9/3R0M6cGIW63+gy9pvvN7
EcJ3av323riwuiwa+3IWVwLBV8059r1334L2Op1iphx4KIIALD8+sVFRHrOw0BnTf3/MpoKYnDI3
/KJ5dJtLA3Xieba8BS/FHnZHla5iloKw08sBsQeHZHoI7L/k4GbVjz3Uf8NWMYAMq6icL+TBbolL
/IlXWsHryTLD4U5Lq4EF1JR+eOS9g50FC1nowfNItBkOX0rWSq9zC+pjyXY6kmfcInVkdXWAWHtE
+lf+WHtruTWgokccBcvYHvKqXKCsNMtc19U+HfcuuOynVorR8hGJyOAE6R5dXyjmaNQstSxkPYIh
j1PyHuIQK6/q1ehvofw9A5ud37o5f5XDWVU8CHU9U58FWRDs/74429cpnskjME2XpvzAzyCyQW7X
bJk94Dqma6EQFdZ+LLFQ3XxZkHyl6KNxTRNZTuh260P7WPjGXp70UPaAy/R6BvbGrysKjZ+dd2S5
uRcPrjkyVhnZa4RJRV3xu5WOYWx0zP7V54DmGXatL71BbxzUTwURTsNhGaLTa2/zu1GRztceAidl
ADFm1cSBqMTYv+Pj3B84D2NMo7jWCsWpu6WRwRVtreNxnlvmJDvwcGcuqurM01x0MoQ8kfsjVeAJ
ZUzII3fDH7uIu0M3kbfMwx71WyVX0R7OVRp0RIY3V9JDKF9dp41+ULYDEIO1upgFxkKmhYQTmwPV
Rm6MuMrjvw9+HAl24wdmyqEUYTzoSDfD0Y8jtJqSfU4DU+lZ3uhuLYlYo34JGWu8U0+nLyzSEhQ/
v7QFiJ6cl/V8SAIrWfwYIc4kT1K8cz3OfJmYxcSDtR1vgvjHIZDpigfqQRu1vz+OKE+ZGjspSgiL
dhqB+P7h1kXFPglzT7ID3JhfzAJpY+ymHYva/p+pkrlytx8HtP3UauC+AuiQsyqfWMRujwVCKeh6
W4I3cBQg1tsa5GpWa37lJZXwuQJDLHgvrGcecjSsb2C8s5xtFovmuof4CVxTH82VH7IBTdbEKG6/
eoepFWnd/DJO94yJsHJEaUx6C9Qv8QeQ+ii9xs5uK43ykDEwwsvrmHGUH6p1vbPkjAEkwD7Gcdyz
Bu5GTXkLNyMTzlPjo3nmSOZ5OmTCFqiLFdeNXeymR0Z57p2uvS3+ljIRj1V8IZN80xFG/EbEfVgV
h+McsY2iyMn37gU9dTCOpC7f9ofTEw0HaWQ23SqiQuJI+cd+OOZ7udEVx5njviYJ5DQtlAODO/vX
u5mbj3NWtsjFa5JUDrAiZ4ShQWLpT2WSxCJoPrY0Cp4/bzT2jDVglVes6e9He2z1M0LNayf7mxQF
8Cro1EsKXxyTSYJu/xKGol5cwNl6oVOJkJTG6EhpxJ1o4hRCD3mp3EyYE5DGaiBJn+MgywCq8AtE
DFwWdqy2Lq+j+NM9RmMP3Igu0JYMmvdxzMfxqe6fBJRfQyuS2v1zjLl7ftiK83ZkLOuzkbrQWnnO
VYPsnMhwmLmm1TkqtVZ+aDul3i5MxVmVI16eDKZQxCjKLKor7BML3Uk35nMbC/dxRxIiTTeFkI90
zlEI498rv0Nc8OMZF637k2etp/cglWKlyHmyrYdPOdhzP1WzrYL8CZXraXTFmUn8mxl2QUAPXIeg
yHudbAlNDpBb+1SkJF4H/Wwxa0c+TW3+QeQ/v7znOyHf2TZvwZ2iWsIcQur5gGRrkGBM+gACCLMq
Gz2iLK8oDBoq7I/qSicOVzJIA/3IkSxVKBAPO1RlgP/+gkNuWV7zwH4fpre2445UaiJQ/JCYHtfb
wZ9Ef8yfLqNTmc0sbyaFzrzB4iP1iKvQ2PDpoO4MnuR7cti+dg3PKl+VifbQkaZ/5F9GV2kzuDpU
shMxTqZy7Knswzz5ZtgJEeaJX4kMI8TPRkYcVNv/AMpXh3uXHo4lmax0Sxuu6sk/O+bWqsxt1HGl
ie3frswKtnLD2rMNvg/vYKgotbQiYzb3TCNLZ3JSkgZg/85PkvfVi92mq7eEIG/buq3hHwgi9ZoK
kGOKqgEAZGVdH0fRX9/UEXb7FT7bWoBd/fZw4/YuG5Wh0IeZ3ykE+q9LK0EtdFcTQo2WYNC1ufzP
L4tW9CvIJpAXL8w8Te5ESrzmM7G+AVBZnUOg0yfOjQR8R5ykHzgtNdCOVQYp8/OFLUlollU5iCN8
AXTKrc4IibgJ+F6mgeBWHBldgstQlNApWNkEI0RqtmukC3neP+4/b0lniWDTibOxOYBG+x7KiH8X
Vo9N1yHNLBuh26r+adEx/OAQ6xs3eC+0Hfw/lSbjSqCTKLbpzz6isZTkFYF6Drk5HkwFqyv82AtS
gokNQOkNrN0hD7BoHlVY3SjGrJXT/Wn+bZ9M06ecTxEcz5GwSzMvBI9Doy6oKv/78xXhiFlimU+9
yEo17KzyX+QEwi9LkwoFx1UiFM2OwF501SxCK86J+CMptE3sBPf7DHItnZ4mkFnhIKF4SCUYlhY1
XY5NaZvp1TlAW8lYuls5lqF/FjU3ua6JOFMDlyoFepcz1K+qyhIgpFo622pFgW9tsS17mn3GD5xJ
DJSUJtpDCshRVWp/bMniQJXoT5ugyM2pWsoTBBBwJ1qizVW+UvKME+rBMmAi7a+2Z1IZ3bzLlkoW
LBlUjAVYGwyr+3MCILXSsBebS+ryXAP9V/S+5+5UzsDZvcggIf9jneOhlaA4lid6+sAQ0Ae1n42S
BM/9kUQPkt89gAgKi8YACgtOdE0Q4imEvRqCo5AySShJBvvKZ+SJglrkqgBP0QH4zpan8pb1TWuk
TI6GO5tZ6jh2lmnXmb03b+eFGIUsNBXqNspgkK+IO9/m8wDT1K8k+dczOIq//zBYJHBclTgMdbbV
XH8Uc0MJx+M3QacgaL/tqDYAa2lYod/S8spOsCqE35DuXYfuRwKZk2pvFWl6txpL0QVlVCtb7s+C
IqOgfahMRfygWNVhaOT6DwXZnurXNBOkd/4iulbGtuN5BtUsc0ZEJpo1txJN9sihdk6R5/UvPlN7
vbrrbbbND0XbjeZPcoMdyUgUz4aQBmw/vS1rROeUutaz12Db+sXES/xM/h+BU3hAXIFT7POVNyBI
z3aSSAQYAaghIqzKDsbXFR+j7h4vlxxopP5LeEi514tXg1rZdhiaLaaNyu4dxo8Qb5z4B5rAY+y7
JsLJ/Gw4pfBwDz5ozGAGQvjOmWo8pLm7xyG4hBq83ycmKIpXZaQZ0KFNVZMuGlTnqzmgST3dm0JZ
v7INjVF7NOksoJ16i7lZVgoJIsrMGbZ8tI7mpFFqxL5mDVUnhUAwxRZ6PEOqcUWT2KTYQDa4RA3T
iQqNWOtSBCSebTIhXpxbviJreMPwCv2TXrUsKU1FpOvbmM9089OnklnXBRQwU/zaLOqf2/WyDQDy
sr788wVXCaDvVEHqI/M/lzrjIqg3HTJuzywEdz1i2BqkjiR1DeuLuUW/Sc/WIQgchCB/XgYzG0oW
MQDF+c2mgvhRmdpBAZYiVPA37gOHTpzf5RNl4AkZWj+oArc5s8TZj58TJVDToXpW30bJEVGeYU8R
UoRYt9frpyhC4Km5wPjS0Gp+eRTqbkFRygqipIUyl9a0b4LCuhq71/ZhAgSm64/D/Kzzwx1ZtlwZ
SD/FdnczIBFwPMOe8M7/MydH3lUcEcfEsiSIlI15YOI9qHqzHY1FRxwKsnALIqX4O6SnqIe39RX8
eliaDOWkVLombWq7KNPPwvse9nDyQj7KgpYjZFw6DRLBcv8B1kAU1IjA1c64EDXoy7NKVtf6gJno
ALWFTeskcdT8hMEN9xLGe+OtYt6nj9P6o+Eh9jgZ7Ng6rISA0yOoKZqnPn3lvA2nWkzryqEWYyKD
ljTyBIcxUqGKWe7NkK1N++mNvVMjLJWBFW/9SAh9ms7O3B7+SnJO9NYhAxcoRFI5eKwAHuejWg4a
piAJlWh3FTsYijInVmO1hqOOvO1+gCFP+4PqPNr56fAESM2R9oEQ8+zdZlly4pKki5RQ47lYzQ6m
c33GrrFZixKlnKd2a3P6kWVOX5FfDt1UmvS6WppQTcXn2SPtJQqKI6cukyiZZD+xFicoBFwNuE0R
UzXFB36L9AuIAruI3Udr6GcU1wc6VMm6O0WDTEKiYcqCXrYEhGAT1fv4Sygxfaxpx68dHG9o0hEI
2PRxgiFVqbIJ3IB7dtJP8Txo0Q5uIgAls2X99GFlGW/sZKB1Hx3xh47MjWKUsV56G9LIeBR0FBq1
9U9sruFnp8Q+tRR4uzRwo0WVSQmqpc/pvNEPjQy8PBdTJeqKxOqo6AhB2eFD7A+kR4PtvElpZA6a
27mRIkiPDj0na/HHk4kGctpQrh0DqIZ5yD1XgIUa+xyQskiTM4Ti4DGf7NPVFMTQ6cu4EnawL9VT
GJf1yygVySUAmCC252ToHRDu9aVY9X7oAfw2A6FnNQ8VRFfcwAuNWW6qI5J2YXsj0+Qug0JQm7K5
qUQbWDTMC52yh8egukwx1/ZSrS0FdVQtUoydhTCPgZdf40HrREORdgb8MqeRGlC82+VxQYePyOJw
Mc9tzru02mo4oogAEvHVy0yiTzsIjGBgHJ7/has7610SGkBk3YfEpaZ5fYwvJac+tYWdt3vw1rIl
lMWPcJ8ktYKC00LKz8UNOgcZ/rgMEofKocr2CG8vGYQXyruj9EBFRNjX1DpC4vPHlsKD20/K8oDz
RdCm3gDZJep6glavw9SHFMQ6sjUbzPOjxkJPx0lGNrW/KKGWeDkuRQGjhriIPql9tjWCP2QPtcNR
zKUUJVexw91w0WF/t+Q2fvjr5a1kzDAC7Y1eOSWXCNYuS4uXLK+elPZa2YyEFKpMnZTawagmr3W9
bDOxBs4Mlq5Z14GzVU3YqrLY3IlY3U9ansi+tSsEw2YykD1cehEHvxEAq9lQ9wgX0iNEkngtz7r2
IwObMelXfka3Ij7kEUB2qFeVLQY27b5zpgjDymuXd2x4VOh+KNN8AOk3Dgqv01gg315vxJsvVA1s
rdr8VgrlkK6013pptgvX/W/N8jQvvqkd8+7r8wyo+j9t9JMYWTdzdcGN2zNdRDUrydK7QYDeLIqn
do/3FIOI31Bt8x8PVbXWtTGhHUETSWGTtMnSFHywsVg5uHxMHHFln5MjpQO3T13hMJESTNyhmD29
qhDe/Gc2mE47LigvSj4RluPSh8gynq3WoVEZnn2j2fB4/PFPJjssmveYm1s0IBqBOau/n2Z8LGVr
FOz+yrh7CcyXjVpg7MVmTeF0miSVEgAua6gZiJ8+H/Batt8YFLxVBLO6u0RiA3VbBm4WgsGhbq47
W4nrRy/JtXMTqvKGsPRr60H3gy7RNQ7iN0BIh/ixvb6kjACbr+6ZRRjdVmVa8M8tLgMfSYPxCUJy
Jtad7f5wNcO3KJhEdHOUVBZGhn7tYVaTl5YVsF0fS095siKG5r961E2yAkpznfjrsQcZWixWFzLe
rTioOryqPf9toyp59UStf4A+CB4Ki7qk5BfK2CF7su+TtTCIM+4X+T2lQ3ZV0Xo7ixkLMiHBIahi
wEFQOwp/PutyiiAh8EfqZVEa27JXEtc26CLN56InUSixgdXcMesGUW5Oc4QB07vdTfVk59HrlAYt
IAuFvHXQqnZvIyVndIyuMY9GNYt3XlH4rSW3DyqAI1CztHVg1OzIUvx5PkqtqrPq7yCsAkBX39IX
r4ed+AogiNi21pE9L4lgk4g6qhk9ij2jFTzdWyydGDqpQVeUjLBg2XCYMBSu6lH+79HTkl2Esyqq
btPA9mAEJZq7WSPOVU+OrgIXe/fQUHNE6V2ZQJPiLjd0eyCKGLuFIClKOQ8oT+qLcSSdQPBjaIi5
HJAsthE6KydhX5jK6dgdpCzupcVrdR9mE3IQ7GFA4PP1/qnF1bqG2Xjhy24wcv5u4u99CPKTyetP
aUfdvMkAp62Q9tjw1T1a7HMzoOD/RJyryPpFH3XlWOpR4+bKiUBrX28axzRtHM1LSKMAwGsTWaz3
KCgiPmf3tGi+NzJ9b2yRFD6p5zCB1/KVI29HTl3K/5XHTplfSN/eoECvk4y6FKYm3wRh9D2kjfnp
ZhGxj1FcbZWIHWK0zGxqo6zzOw1kDfexQXVCvtcuD+MVNu8iQbJVU3Jm0V7cK1/wH1vq00cmQ3Nl
l1bqjGoA1DGEdzs7fKshZdd0r56krHtsfZAWGJVCkrIENky7NVNxMOF/2uwrZngRYyyFncGbFzxH
d3HPHG4PkyMJJEydW0ZPH6Szv1BALKBdnzk6Py+HVOlNZ4feahh1VauCHi+VI0OkO6aflWfvUENl
faxC+njyQ/EuXFY1yZLYCyagABUbyWDu4uCOx2FrJS4YoqIdkR8Bp8aDcs/WdpcG/1wojzg2KBiJ
wttus6lHIKF3gv2VP8ICCsKG0bN6zAGd5lzCUPNtY1+NpIS/gjbwWhw/raiRRPkIPQhntGqP0WnA
fvtxKzRLJ+fIjiyTMGsdkqj1uacpuoyeDl88msQ3LDtP/p1unfkNlOGqRqXl7S47tYEHMM1jeZgD
ormDsQTrSco7jgliu8lXhkunJndfjDpo2RvpKY620OgTYUXKhgUeNImJBf9/aGCmTPYFSbLTsbL3
JanNQvX93GzJSXM7CoCkT8s15+9niUUzF2vdolps0y6pppGkRhf9MkqnzmpCxgsRyBruwRDBW4Hz
54xu6rTNbDnhqueRcWGD9L9esXkKPo6bE4MIUmZhXliYdWfk5TnYrjGYOt1RHi4XxHBuNcXtdKSq
+A/H45IEfXb+KS5Abccxio+230EPdhBj6ASnRBhPRRBb45Fn0TdAHud3qbYH5c1Ar88KAHa1wT1L
Y2aSkwjEkAhCMLYtJGdGtlm1gNmpdn3fWFSAjWvfW6SqLxo4NXwlO13gmH3OdWSH2monsZyRSjog
Ysa1NBeb/VT/0/47FQaBII6JuQjHArcur43cgdJmbSzrK47bXZiajaWY/gJjUwaKpdtQ2dFxBvZw
paLCoQi7+zcvoppRIBAriu5E+Fkhs3zfBJ2/SqC4NRoANB7UN+lf81pstQjdi/mnhdccyiGqEtSz
A4H0EZLkc0JrmjAd50L0stePAL7aGFW5goDTqSAvui+AgCPUFPQn1vaVLFwLD7Ew4nP7J0XRn0BL
wl/XVe0steyaugTyjByAVtpasFS8paHWirr73c6y0zirMhqeAUDs+aOY5BToYEWQRFIOk2wIuIga
m1S7BRgrOpPcsiuQZzeDlptx+c8capTaNsmNyHSVh1XBIoZHI+nrIezCo2zfPwY3U5gDnCjvXWgk
qz2XAXxR7INgsiI9GiMhgtMUg9B6FzJGKNngOcpU/jqklqdZNvDBzGfXn4y6GzIrLCqpT5Ep8PHe
ghkyNiUVUebG2pwbCZmqBj4kFjQxzZWty0gq4C0C8To4QfRDvEzKrRyzYCLpZNYIc4kbU2RZG8Wo
GTIbvu/yGcLuPGBO7s1rXRXzHyhdQ+TLMzyMV1xeBsL0d1wbE+QjY6RofjXW4CmchPFHIzTwoB+c
302Ogtj+jiXKWpmV2NAkwCR6nyKa0RMf5ynb4nvgK3iNowL5hii630en3II53dx8qu3FvU0Msw0X
3XzGc6r9oaVkAgX9AFLI+1LSWvzsZAruyE1yAUp3Qf8tdaNqHiC87cvrSjJTB/VOgxlwg/JjNkn5
8N0vW57jLuXCVBEIx0KAf45k5R8QAlSYdoJi/XcZoCRUAG7nUh2I1jI92OqXrciggfp5Oghlc/IW
rE0zyzXC0tdUN778Z/v014IqJOJ1U7qySfzm3n7wZzVpOY1vKFB4hrQhxgud93nPeaPzvLT0pA73
wB961NsH25XuugZlxJRjPydNWbtQLKogdUWK33dt+Ph39xGmFrhcTsWdUefSbB/Qt2pK3duz/8gk
s5/Xh31TSWwN+oBScxAihQrLL44jfMdcESIgpna02MY0/QrtUByOljDbTz5F0ibStek3ccuGfuTf
giFhu0HhOD59qapuaQLbyXDdYd5tPbesNsqmGSGZOC01Rq6awIsTbPjDht7poIuly4VUc3BLzkFB
v61KZqmGGcbcCJCtlvIk29L+H7s8s1VMIq6+Y1+gadZw9CyjSoaze6ksIYqJkj60WH+WbqDGvYcF
4AGtGMyBJ4E8kxeb0kbF9xzImFRwqH2tgQA18ZDob+UEjGYyrK3AZizFRBonzq53BA9K4YhxGmeA
cbwbikwJ0hrvTAF+lePu+5IrA0BrtBxz7itEh62MvQC68BbHSFh2GBJrHHYacwJpd5dCMBlEQPcA
xQ4ipppt0ydWl0dV2hcAGO2YxPiuXwMQHxbebGxOE6aCnJXo8JpYc/3e13BuTwc2uMsqiJx0SbxV
lavFxm6J+EBeDQNSSpWzU6E7+QuJQy0EF4drBT+wn+TmoYUFeG3aRZ1Ai5DYcBlmmaqv1kDitsgt
O/rhEYBn3R2YlPjoxlKQbkvO/ZLl0bZiZ0jBQ8dlH/8tZO2IWABA+mHVmI+UezphtBkvoAeTDgs0
qXb5dKXJfdFeBSbV11yMnsO++RoW8sW8LodB3WTWxcwTYuEHoHkWnaWI2WSZCSgyXNN+gZfQmYQY
pu/WY6wN8zICzaCU0RN8i5vgjHk1OvfcPQFSigqXsGlKbw9LoHJhkLPLY6x7nqTN754/gdYuQCaG
zXgnBVa/qxv7kdtgQMx75L3ZdZU7DppmcXRrK0FzYjqZVUDMGEvboX1vOoj1HcesL+rWgSR12yZO
JerNKC/yQYK23DAPdy3GVJqC3cdFm+Pv8nXc6OTz+9tZYKG48WAuhl3hGC4TfknFwjU3NLJM8KF9
Eg70lobgoJJTdfFfo3csm14G+Yh+JkmY1XMedMMwwdTEzJCfvhLat4JwTtuhOcoZBv9O5Z6p9dt9
EsJj4vC5SwWVcfSE3wAiQyH1jm7xXYwkGptTNLIx5o+CTLbuynRPJ4yOVAX42LKvdSKJ9GbH9Yd4
Wgbc+j7hbKKPBCi/BjvV9PFiQmMcJJFUcEQ/euYk+fWfHRnfmD0ZYNOpYVmJa9civzpRuXpaiYCL
goIb3k1vAPpj15gBpT33IVwJcslIz2XwPEX5QfdO9bHy09MX/15XrjQU8BKDkK/XC5x3z5ut4Iz1
da+FHLb1fD9Qc4F9Jds9vsDvVmQc1+bwS9+DvS3TT6WxswVX8xDJ0zDs0VOS36dlXim2WS4EZ7/N
5b6rLbcDBdl0S9LGR4metEvoVbgMr1xKYczLMhDV98xfWPETzvGrGHLVHSz7nfGXAoNGm7PusaNr
UcNOeOtkinzMklHIGXRaE4i0L1biKQhT8OilPdEXoh4XCUmmp3kK71bP9t7JatCuQlCBa+XLWGKH
w7yM2BORG6W2RLymCXjBEcIcj5KqkesgRP0sn4cr/FzrTO/enMnlBVaJ24IvpHp7pjxIcam2cUel
01AHPy6b+lma35W+CDylNTGwIAwRmtfqzCAwlIfDF2pHhTadiAIFukohk4I2hbT6nYXq1XLOQz9W
Of/C/n0n1GUmuGecO0KwgVSyXCX+AXIdgv/YG/vaK/rJ1nOAYLWfoEiEIgnxivH7zKJQlKTWvre0
prL5t0Mi5p8YMyEQ6ArjghXGg8Xr1GaVzKm3ao7I2bUh1/DSeWz1YOdgxGq2ml27zX3Dj2JxROa1
iowAZR8eXqC0yGMRlzVvMN2RD1F6/jXfGNZyor5MnbhLv8AEQcuzxrIid9SxHRq/hmpj2Lv5M0oJ
9qk4bUrCyD5agjQaJkb/s7A0c1pzmUYVlPl5C7YdKOYChk45I5ES9wtA8OSAl7OlPkgIrmhxD5Qw
InJfafMA4KabWDJaY5qdHqAeDORuKFim8FcNT20CyGn5+dLKA0CJwOpu3xinKxxifD/50Z+i2OWv
EP/j3B4B2ULjsbiXBGYqtVjsmoHF7NGt9U6u7cNsargXDq/q93uoV7HpB9JveBuNTNJa0hFei5ij
WjCcWBVV1ekA0EViWOCZLaJ8Gan9IVP2mWiJ/33Ls6GhWFA846GNWdTh0UboeaXljDgazSx0izXM
4dC7p7Mg41dcX1fcqqhQ+gThzlq4XxLBxsi2REeL7zpgWGCBEYooP66ZqTGhBD8121H12Xyy/Swj
hDikCTAEIeSH90JXdGccIczTBl/gcJtRI4xJBGl3dncRK3STW994X/snkqlELBli8kWgDpD3mHs1
+z7LVruRTsh/u3sER29tpAVJvjc4C+QOnGoQ3FKSKxGOiV6r5eF2Wu6kA5Xf8wdaYGDqjlSvnvga
IqZ7WqKN2ZuSC0JrMrhspzztnWweHnYfdeN4ioOSO9DqIDyZOjeBCvDqEZdxiHp34Yq5W1TKeKrM
ioa+NhKk9DZkJsyttpDtpKOZirs+cl+6hfDV7e1/f/6gp7MuAHo+AQmY1KLRMtOgcmHW5w2ktV/J
W17CCOEu+W2hVQ1SnoJrqj/f/d+w6PTctEWJW0Oiy6eNM7qFBG/IrbTlKgOhXwH9PIU3FrF4cC2T
6fo261k8C/C9wCyFU/6rO41xq55m+xUvgXh6yUAbODXBcUGlNYgOs5su/70V3rt8LkRzLJ1ITKy2
aWffUcqBycuwJtvRuHBn3NLRXcGve1vSB1xrq/4sE4lKxvVVj/JWxdrCRwU1K+VOl70JbopKU7Z/
F3Zeu2BLnmwcFuTs2SlruXRKiEo5UJ0/pmRwx2ARDy9Zq0EYkHMtaXsTA0DlV79KKN3p2+2Fwt6P
GptE62Ith3zVpibiLIlKIF1JA5E3bof1iwAaerBH/g0yWJ68QF9FgrSLe8eEmra6aZpC1qRdDnqo
YwXjmTxWHtuMBLCgAIr2zhmUEAUXwUl5njWeq99+bdUmTerW/FW+wOpgyz6ygRPYQC/YAFJUsCHh
Q8ZOkuRWeBdNfF93Fd26Is1VoRL7D4SnRMeFDpBRoEyUyGYcd++fBlYfuYxLsxzManXoW/GXlC6s
K8gcbCIa/uWTnwOH/ug5e02Ld5Ac32xEwOG7cP1NBz0mWsr55kKx8d8CQGQuORAwk67TgfFl0gIw
EKLuulNLp9hTtp/HcDdUkQASf6OOt2MP/RQfMMlvyqJ0rh2Qz8xrDnmWHRJJR6vh5H1hK254/Q98
PfX918Vq1+bS4n2XJinGVZwQ3xec+H8mcoF2zvjmge7C7JnE8OurPGdo5sP5DMqf5DyYww+o1dmy
/w41YX0ZtK2u/ppsSLX+U4a1Ap78veQ9sEvb9DVhZ+gdZXKjYJze2a8KeLNJvVIPAZDSe1k4eImC
jPk/d7U7o7zKQvvzWoA+e4YGv+sfjlOZms4v70FuEookQBgfce6sk5m0S34FJLi5vEEzAB6kibOw
hUxF1kFhTgUFmAZffKe4M+V88vrLj/c+6f/86TP1y+HLz9nZkftJ21Una4A838izEaBXg0iC+6Lq
6exSIG0Vx0V0T21zCjBsHQmgZiS/+TUtWlZSYDNVTK/WIRomwCUtvTwJi0ngKO02jFuDmBgw8N4T
qCK2PMpDPsEkA2NXvzPR7tMwl+oqutH2Rjy0Y9djbD42qY75KViF0OPde95X5I5CwpeYSCEltVm4
d+w7KIdaT+OnMEzq1GfJGZ7jkx5FGQIRNrYmCGftmkXnEzFa2S9WD2yd9fcuxfylY+A+oxztRFQn
NkhxR6q6VYaVum23JWsVVuIyZCPErEj6WNVGKRyBb2LKecOFpQPmc2UAW+Oxkda0NhvGVa/WjfQG
Pg2hy05DeEA2UscFeT38AWpWJDWQeN7amKrJwJoLrKWbT87S98G9MK54O1OXU8XqHxvIr9U+4GJ4
WWEEYY2XgIHpz5Wz4Oqr6A9e42qowYq0VMElTB00pKic4GioHPgMJqVi9cmOXuUvLYLpJ/y9aNsp
5vQWmiEU5X/BrJ/oUPkfCSPgR6uUekjWofCU8IjXIzHi+uIYrxqKDeOfPPdVrJ95brfg/GEWCi9R
m1XqXbLZ0bgG+2O4caRQL+VackKeYeXXQ4R0azKfmXVCJnlfXfB432l2YuGia0ZH2FS055lO4O9j
t6tjOk72n7tPPx+BY7+ZKyAL07qi2IHCpgBLDcsie6w11VGPSifchN0HXq/LTmRv54tN/yzdn3WZ
FlsqKytBAUVtbeeUXPxkqyJsL3AHfzUBxDbVRDaMH+zTOtsPDFI/8XJ+C4iTNkl9/tyqeVvhOkXp
c1XLU0nFQZKyIo0CbbZfmyKgaJ+Wssd/pSMpgNKlgfEVRfeTsWAJT9ol6qvKyScPC2ITA4qTKCUp
yL/BOdL7ORkfeOjzjfUNwIKH6JOaVcscUYwHf4ceClromEtck2ZYf9vckQ9XeyKx1Cp6lhKq3JKv
m7eU8DtDHqNh1ggkNDtQrxjBwNCs9fCd06PqR+6hzenFrgU9HnIk/rXtWMuhI2YpVXCFD8XLMSFg
CcErAnTt8hsuLE2ewnN5mADMRqnchbS7B19ufzWJTpdhORrzhjHsFUK9ijPjOixaiijR4WXZRhC5
17KR4KNwGexejh6Pt2iOfXK8nHsWbH+ZiI7svWcpWKXeJGqOMctMh1F69ndqvMj6kevZkZj5f3pg
aWntjRKeQ4LsdmSWkNppq3o0SlURzIhy5p6VppXwAPyLbFDA1BvM/DJulQXDCUSzo0P6QV+gO0Su
H/F/sz+EACUaS9xAfLea8DWNGoNW7C9PSgjek3zaqfGawEjJtRwUFJA3kMTfaP/pBmWAZ72PDmh3
BxGJBF6X70Xm9jG72pZVzOOQyR70Z+RRuCamB0HC51yFVWWhOu7digpNpcw/xglalKePJR8G+2h3
9RcTSeB9NbspsTTdgeM3/4tDqqtsES7fZbdfZ4k7HnGKqqINVRrZhM+NYhZnE/EvM6KMagdmN6xe
I7b1JJdV/hro1qPwLt6et3ibqHeOBaEU8MgBx/K9s9iRuQfzw6iXke0rSrFr6UQjkihU69/gEe+V
HLkqZA7bUf99pac+GLXc2Lp9NtUB/tcgjM54PGaG058gNSrw2SpipfoOm+ECgi9ltThqQy4dpKnP
QZsHDj6e1wZDB3Jz5z7/wO9Q5LkCeeSM5YinKRfT6qwp41QTN63rXU3c13GjsLj1dqRv4DUw3K4z
x8TSX/GlXheo1H80kea8eqP0maHezA+ufxYB8PhwOHkTn8iD6Qlu6RVr8jU/MEIrNlIZpxVJVG3x
TyLzKMgJrC5EZU9AxqYkRshIKuxq1mtasKIrLzOY7R6auD6aevj/x13xz2DAoZTNtUfEd9vOoGgt
i9nO2Rvu/ilcSwvTohRQT3cMyE6V7zIWYm8jcVJfUFM2n1KLiohl76AMFWq7PJHhLEJC4S+zApci
dgjbc2ZFOZdH3YUc+moUDPqBAQckeoHZtA7lQ9KzK1JITLcKcqblQB2HGcaH1vWao2IHbstIfVym
9IysbNO+yOMU639yNiDOiXNo5qNaUzmc5bL2417TVLu26TPFwaf4a14eqdQVW5/+imH7Me0JR2db
Xvd8vDqzTxHue3xy1T+YY8o3l2wrW0CLi9bJ5Z96c/kaBwYnRfaVdM9H7H3K7AL9qYFfpLS/tlBm
lKlrWH75Pzz3HWBrLVHNF3yb8zniGkQYzrEbQtgcsZVwdCiywM2KtAyjhkEbdrn1nFKCxpfkQ5EW
nYrP6IJuzQEbe08B5otWKanMKAbqTrty30XToxePAH9q3K1fKvgD+bnN1nob4iIwqadrmbm8F+RT
Dc2P8JWaBl96O9vfoZAc7H56LXv7w+VMMxQbumq/O4yx1quO/ju2d8Z+UkvZvCjDt0IhqzAIw/F+
XQrUQhn/cVa/IvxlgZIjePbEY9CyuZhBgxk/SmKZOl2MiP5kBwDEjVPekzGKN+DgXs47mdC2W/5z
NF/i6etdOQ9iDZXfpjwHIW0ACMX2fgDNemYVNHvCTILfwuBOeMhLh9NTlEsuhuhx9YT6yhLtmomu
GkIFEsH+Br3A3d61YYu4LEsXkmqnbWqbV8boXoWYNK7QMps8bQfh9DOJ3Wy9bfqGMz99plv1Okpf
B5b49JdA6x/1aSVCVtK5M5ixB7aN7+UEGDukv94FPPEwb5YsWR7Be/flNA9+JFFddI7nKZcdXI54
zizY9v1FAP5/YNo+7SOMWLD5eioJSSt3ilyaMDqDowlc3k2ePNJsfQeTTYKb+taZUHvz4XvilBI2
yotlrh9SrEEBKqmgA864TN9sH6oqyehY9kscSEB1C+pbO773wNIpTKzN28opb4q9WFOHDrBisAiP
Szy6eKuJrDVwQyRfuU1ntz/eRiG6HNI4P90/tYo4UOnqDHEhFJRZhQBwXGm9eIDOFxhM8W8eHkgn
2TIWm8BMotPeqtS/neZAlqZMIBCZt1PSQEb5Mv6YEjq/hjTd2jBS5F7xuYu5RBjF1WNqVRVdLwPm
+myBUNFrjDi+7Q/e7yrqSqyH9maKHDFAwqeZTID6+mKg34Jzue5DXpJmBU3C3UjFX6GfWA3g7jWR
GtBkLq3edXMX3c8Mqea3Wkdq43AbVcbv8OeB4KIw4Rfv6q0/kowYixYD7p3KQUT1Shas6DAL5rIJ
tOqUhLKcJ+x2K33enZyIu304zxU1it7YRA503Y66nlnzRUKnKi4dCN8zS51dro7/yazvUqehfES+
T86dnJnEwfkuDtCzk8P9el8cT3sGMi8GCpMsZaIrQ9brtDrLh6M3rOWifbIKje/j0/JPa7Fko5Is
/6xb00FYFjwYDhhJXLFwHO2pLuDXk99o/m05gdHBf6AMZBA8lavR4DoFNZbaAjG4A5Xv9YDEqX+m
1XsGcjCtdHHH26wjRLB9PrGXNtunRlYd9wB4mQ26wNNllNAuMzo/TxADYZUVbMyw7EdmuEzkSLyk
Cz69CrcInG+qVv0Myo3EGH+LUz4sDfTbk4J9jHXAuo1as+6CSxEGxN6kA0sjHHiXotLWf7wXQabw
VLzt+pQCCdkamqDVEHFVgZJ3sgkuDLIN8Tt3YyRnFJqpqKpNQBPuqyi2FbiYjtJt3YYTVGMRZmJL
/AJCc/bkLvXHFjv579F3qPzI26OXmyA/OZoXKUtI/tBc1dP02cXoHrOsofCvm/G3xPzZWpPejVP0
GCLdDvDJcvroBTpIB7EXRSSpFjv8z8oHpJMGlafkrqrl/kGZ3OUL0gJo+rnVhqyAU20SL09MlC4G
2wUIk8W51l8ep/jXeWQlmpkSN6A3Nc0ObSHf5hrCLNJIufCoVr0jcHEOCmaJTHdHKcu9oWLvWVse
nHiJ3XN3i8Af+yHAxXRKGYjYaCi8VghUdDmcaREYuGxPbum23D2ZVJzHZiFllwb+rxj//iWPxXT8
tvsEpS79jBNUukrhtfDKkDvFN2F3Vv2JKu8Tl+ALCEGDsbxD/9SFyA2tDCgcHwi1XzzNxfuhjLCG
SE5EAVcZjDXOTNXYEV/UPHToYz0p2VC/rXAIP2XGckil6ncCTJVCMeE10Xo2JJhjno8FqUo/jT1s
IYIfYneYSTQe5x/vjNkCa8AwSX4+LLCUpGymfTPrk3mEqWv8/3e0j8cEIAnMypQonEgv3w0+HM4t
pNVgsno7bZu7+F4Lc8RcXHNmygTYtWMhRVY0Z5YtNiXgARwD1hQMZx6QhV0uVTPmQFIT72mYr07P
cctuwCrsmE1162WLs4tX2yb/Pj/UgxfK3QZsRseeZj0JEDzM+g8tZcOfIiINTX3NZ+aj0boMPj2H
OlnlhR3n2rCWF+gcpple2KjVCgvlboRJnGXl3cwVd+U9iu9vf8LWWA+cskZ/FrFXC/daV/fN+kra
vD0HH/keGwKXL6wKui2O6WralovuXUllYufdr6aypDUp0Z9/MoiAGUNvIUmvwYNP1P+NFuUE4N9S
1JEcPmYbI1ryWvuToOGAzVHx7ZqOwkVYBU5qgLa0dL4ZHTDj3gBi9s0kgkAGBXs+nrw19M8Zg1tj
DoTnY1vuNSTJiwV4L7dTWDGQmiFQ5Of1CR+V+mbBwglNIjMSCkrNIkE55ZAD3WX7nhRJBuTrEzYr
YeqmTNoHKTJUFeX0xp2DSkuZMc6QPucz65gZNteTEF7IJvg/DF03315IhiBlc9nDaHfbBrSjQOis
Wlyao4a5q/9D0giBygbN5RopH07bxJVwPIbBzzTT3YkxxDKBUFo31RXAfmf9vadsiLShQ1YNMRUn
l/GU6DxpJlxz9dw4WbKIPX0tNlcUajuxnqsBf/oUYdlqAUCvQmGRJ9dbRbYMfUl6kgwpwaTdJwVt
O1iIZo0lQZRWTZ6BEhhMQ7UQUP+MyGgYbNDeJYkoYohck1E7NqkTMzbF31mbWst9YbBgKm7WrRBL
TZyXofWnS4b9XDlt9yoA/u2JrFbCXOS59Kc0zhRQa3wwa+xWg/msqPeKgD4ConPtepjtTKOAsZ8j
mWt8toyzETGb1Z4WOD7RUo8YsYPSs/YvLzer6wUOHhIsHbzcyDaQP8qy1iXyuYb/mMhcx5wz/7kx
MQv6wMO8siMvXSOOSuTcuj8+DztsvG5LJGDzK8791o4MjZZo7KuSokwfkjsq1Zg0u0MJY+Up20Cc
+LBiXYDwKE+dWotW7WZJ/36IiWG4gUtXWJpoRzSoRPtgFYqVZpAQmWUGvoIAmcH+in4P7bCq9YMd
cvp8BUKmgRj3XW3xyEOw44Lew7FkneJQXBSaSNHv+OB7qNR2VPf618NPf0ioOoHbDns8Z/mS0DV7
jCkrsIvMR+HmMf7CVW55RB2HUEzxEHv0W+DcENXmB3KIQXi97rWm3ahvWcz1qopeMvi8gDuUrItS
mwyktiauJ3Hf58T8BM8PVyBdecd9COVvDKmQpHDbd8vDukGhkkCplc+/rV4N6CNhcbuJFIVR1U1z
LSQLYM9z8Ypf8qkoxBQiZj516wcmE2T7wDsRe9TNJzsK3pJuOlfqgOxrlRQ3Bp3l12HhjGoL8UZU
sOaRJxgi2zWDvpvKTS4nrJmD+xL57304TubqkkhAEgpZ3/V5Ma15XR9PQ+pUAVSuVKFwCeTsQT3f
s97r57S/e4/zW/y5tYsncIQGIDXGYuFuSL0uJ/r1xPfdEMeZvb9J+5AWdsPThFcY2Zn0Kdm12PJS
xo7T9mrgi+mrbD1f3qjpfAs72nmafW8c7VwCPSKfwDUykdCb82PChhU/qp4x94z8RMRQuq34qBiu
XBBPaio8Qj6mmrP1T/0BE3G1Lg/zK8JxacSbfOVF5AGWerVbuhgHCBZJ57Y+5Su7e6bm7cANi1Aq
8kFinqE8Cxnu4zf55EmbCbsReE6o7SVj0ePBgKVG3wyC58Jbun0urtidTAu6uSpWljIBUMQvNxBr
3wlqsOpZrsoXq+4dMTyJw9sOA0Wsu5P20qMMdwRPNjyQpyf0EVWY7OMmbCfDiv4GZBED/9GH9NMp
zf6jK/ms3Hz1u7yXrPnKg+pTUqj/9M/iBWOxDkZXZDBY1zo56mWBDBqG2dwnsUGL1sOmYtlqz5M3
+xbxZyTyjNyPJGUzm5DDVBHo8GSSRXOFDCkFf/J7MmsHtEy6D1syWXta8rULEta5hww9OodoC9oj
UgOK7rnJFMq8Q1D7PCmx+Bmw8HDVmsPzDWibH2oCWZJR4OmkUBRzaTRSwC4/GiEpZJ62+oIeaisr
g/E4qqS/S+7hj1cAvvect/iNs8EWDsufTNnemXHgKnDuFDCyIcO/wiAFV6T40CHq7jdDullSiAjG
8FUiNyBitZcgTfP9/v739nleNPorasctXOhZyimWnJ3tvjFEnZRs/8S7qUzIKub+8/KnI+QD/Sat
1Q2uWJvWtxc+ccLv+oTG2MbUvV0xgxyH6ERNuHMvUtgLskLyklUHJGoBD6Cf/vQi6of/zBaRIkK/
FH7zGt+3Jx0ymULYRNzIXCUTKfp52rqKOQMUFFIfCaPF11qAgxSzm/WQRfTsOk0zhgU6Nes7IhOQ
sDdURlveF+nEcI8ixHzL57KtifataZAETvwt0e8TezrU/8Jr2OCAOfaKDsIs/KiOK4B9XluOGONN
iJmxjKdglwzYqNpNH5OrsAfyyx5BqyjpUepSdLuLIMVkpE15rDY3pLGXwCqQAHh69qVGcc+iAGJW
s14NFc89Oos5NAvsoWNnoCXQQ7rxma9BB5JeufDOe/dDkCIcui2B5uVC1dInxh0MBsCmugReWkda
lW4ch0EUeTS1s7/BWGRYAWFAgaTjvYUDR8TQJN+SZmSGTwBlgUNjw8V4H/E24pFJ5N5b+XwXR8nY
HBiq9eiMzG4d9dL2hxvIbYA6r9YnY3Qug65bCoLk5XEBYMoxLQeQM1Ryi2Jg9/FVLDZaYJjml4O1
2FNd1tgFTtBH6Xe72ykG9W6uV2r0TVIWBg0EeYcJH3N4ZirMKyjA8AXB3HFv6JT4TH4PgCLDh9vO
tVBqUrZHLFDsdfas9l8Rnp2vYuaRrI3rLjtKXbK+fa7G2HdKWaQEcHdhi3gwwmlkCwAnt4alG/yS
4JswgCoKvfgroVywftvksX/RSGWnSV2mwW8C+Wkl52l28O00c7JFkzkCoNbAfgs0eafDrzTmYfsj
gOQq113jnZVkqdKzWitYJuebwQTA/BT9AAYhqzb31NTCz5MBFk18xoQuZcJLHt+CRp5WIdQ3l5oh
oLz6MzkzC3ynMeotbZsGsPCx3RKEe+6ifQy8p0KrFnko6/OET+rn3YUp5tg8aexv4NZky2SC2wMl
t8EAbqFLuzhp46oI9SRnED/uL/FmM3MyAeN4WzNpWgON01W0E8Ospz1w8tGY1HMuYAhPfKPsFWSO
IYidmSmGSx+NqMUHlSRAM9f1vMN+pRXs3+CSlwqGNgJTd41OCInVc9H9KleWlPOFOlQ7wx2nZ1yc
LlZU3nLBTMu54FuTx7/B44iJ74rGI+yZ9dgBD4jyKrJLOnXV3jR4YtvYhvTz6a0ZXaTnaQDrEmYZ
ZWD2XpPJQtW6TQ9rtXtSeIfp7+nfUpvYSZSAQ7xYl28SGzVPlU8HV7L8j6C1MZ3be51e3bXtuCoc
FlppB74royg14ZKkwH6c6FXX2kEBZPGub9GjxsF4Vz+YHRO5/LCbzUWHoKiHWOulTWxU89hSbLwb
l7rtH3l30LfBwyGL5bqw+LZUv6bJ00HATT5aL6dbikyYqbm6toQGxIbEQmdoRaNFFlxoiH9BwjwI
5AGxbIENPzCk0K2iPda3Wz7U41l1y96BvceD0kcN/kCmjK7mock/vNwY0KQGBQJjwwBcYSAu2juw
07v1bTM3oWBnwph2wnTXPHiRwD6t78ME4MCZ/ZAXqnLjE+4PLkQ2e/a9lOtOjkjZglxj2La8TonJ
/TOhi1ULxII3CH0FQ982Sx7PWNVZcXposy0iEbu1RkPB6PyB7orZxqZY8Y5Nm0ouTvxlHf5JII0y
tKzKb2PyxGqMmRAO44R6KpD/C9jq/7Mw7FLqzGuCohziFU2Djnwy9iqVdowQPxy8WF17P7D0d0Gh
LMP2NpxVWOK+rNHUwf/B49H2EN6+GJbPzmFtAWwFJpGB3SlDHl3Hqu5W1TwLL4PgFrZA6Rxx4xrM
vv7u5A6zkc/NNHSJBtwYMQLysEMm9lsUuEig2R/r01cexafv4xQjc31UMMoVywLMAGHNhB7tBr7Y
pANcsjze/52nuKMhNJft3zlv68hoNMV7GVHhBTPltGX6QL601s3HLpGs/6uGx2mEbugaks1nt8sa
tsPGhTvHgMYV/Ptzju84JecxJfUQUasx3LXXtYFTcSXuXpnyihjfUChB/gC1Diuz41Vicgm+Lo9v
acBdWaJfjr7uP0FCyf0LXV3L23QY9vxSza1IrKpi4mZs1d9lHI5wzNxG06nt3hbXZHPYPpCimTZG
KCb1k/dzin62VDO312YFoeAm14pWEKSrPf6l5REbGZn1U02gmYPBjs9nTzBiIXji/4OhTBOY2urP
/ZKxTlyb1tGnFWd9ME1Iy4tKf2pJ34TukHhs5LPMjai8fOSMLYq8FB058fjY4T8aDJBhG96ZlAdz
wgBpI/7rmyARkTTnFRS4okfRWDMg3o0VAjOtzKj+jnXiGU8b3KLERYsfdQDADXrVaK5sJ17IFhX9
OnrmbPkgIK/HNNrMsFT5O6CwC5eZLndvYPjZoXb0YEawU4ZUCYSlwyjroYRyIXRtcWCM7O3Q+iAD
vAh4qzrUaodxcMc8shyqot2laHbb/7AjHeu4iw168Ic7hb4y/8oxhOTA6s5136Lmso58ooyzwGch
wm5J8dsjtyKQIYzn423bwwEWkV4m8W/Tz7/RmiDAiAKSaMebr4CJkDjJYCod0x0UCHVvQNzR6qUi
aKS7KrIGSR3jNKaZOF78vP44UpgK4y9EdEfMc2JA42xO7dYzOqshsdde9DpUjYHKwXsxxMWa+QnB
zj9aNiIdnS2UmYLTi/MtSZAllRQbH0EcIFEYg+xlm6nxpfwEYlzhbnumsGajeTpLuPQCN/H6/eNM
izKjd31WxBAUzpvg1CNa9NbBG8ttQwF5dXKhwec0imzqpqpxo8UgT3yAylAshoe1oVxeWIii/iwk
YHsl2ssFh98uLijwaaOalCMOixcqtx/niEjl4UaXBQzLr09tGVP3xB2kP32r+/KM+8dMzh7luoH6
XJfIKMGRdAsfVykFjtJs6vaZyKOFjJ6Yk779SMNl/3le1Z13m5Lmawm/SXHy9TDYbXI9vLOka8uo
PT1kS65nHXGfWRNmIBViiN4g7FA3Vi0+2np4+5CQ9vhoZVwQP3MzQ2lZ3wAIhMnN990fJmfqaWav
G9LzEUghKD0RytSwoggFF4zcMxccRcUFT3Q6KnnIe3cPrW7Si12bqlGATFEJ9s1DJRG+roqCOoN4
vLPU0sl+KRB5SOYTXlzRCT03P0jxieRkYN7fG64Ey0hbHsm0HTVaDr1G/ItmzfjZRcm8f+yCukwp
A1vnlLOxkG+R7djX9Nn7U1ty3J7rXL6xzIakP/e8BxeO/QfeyzW8+5I268AXdiy+lPDkxrMIWVdn
2itKQpwKLsurEVbf8loGPvRGnWMbAVbCEym6UHjINfAfuUQyRuMaggDJuk3p5yMvDyNHMOfSwOWi
klXn3I00K7mi6eWz3eIWXo1sXaboD6tfbpCBw5M/RYEk2yH6IMtdK0A0d1VhSZO60yHLgdV26VH0
aiwwiJNZHboySgd5E2ynARuToEhqRsyvYQZySNmYqwCHPon0oWOM9/ezyCbqCnXZIsF9VnXjHzmc
WsMbLeCU5AvacVgZcOEhiJ8x+PPzr3ukKua2B3k2212l9db9l1N6tZ2AtUwkG/z7X8cnOkfegf8M
riz10VIHOaVG67QQHGH6NrZnPONDQkBiSt6AiGvQcwnDQiqN34MhBLzYYLmGEeBr0IyDQ96oDixD
Lwt5dTe4Iq4K19S0o4SE3vyqCt9SbWzaO+Y40DAWJKpV13tAevImCpJ3bLXzQIAH7popXQFYAnU3
1u/W9qmrGWj/xCrVMaQItxaBZkZgBOhufpSTKg6KpYPDKoE1FvUaiZ+oAiNRHGtzyYnySz91UIea
cjuO3qOp7pyW13J826vYMw3kA2sy7ogzlKTJ4zwsb9BtyC4L+oJnHmPReKA7jFPxX8YYBFnIYaig
BRxc2DnWhI1zuRra9eZOi3FmFkbRaIVQfSDmphVB31zoVjb2cAKGQs36jDcn9f4RGmhiiEeuLiT+
GZiSrOESPstzq/kq9gZcbY/Eng+dI/hVn2zjeSxuSNAz9WCenrnIMWRMQDx3MIRCIRyPYjePJ4en
5gGFlAnjrorB1L8r8YwqU2AhgvHPXcZ48BOnWNHEJg0HUhuYLKrveoI00r6f/4kXAwR5/gLafsyN
ymbwM2tgAynqkvJ3EHhLwX5hgwNZ864LSSMYapOkTii1VyIEJjh7ixLd0gr2slh8gljdH1/pVSc6
xzVP1bZrt1MzHkCHngQbIBk55cT+GDQSAoGVgtlol5XmVaXLpWyN2qY1M5rKH4Tz2vKjAGvu4/+9
r73/o3gPH9NCNRD73idkcBpYcmCO+WBmoJsDwijZDir/8BbICdYCJcOBuV+BPN5jpHERgiGEF2lx
nmcvr/Y7pd2THfydSrHoBVSa0d0/GxoCD6tPNPMNXFklO8NSqHoQc+yGVhidHRftNXt3FL3WiVjJ
uPbHbrXjcsZullfc97BY2S6pedIuHXh/utXgWyVPA4zUj0ee3+VnOi8FG+TkEYhBrbnMfFSxm/uN
cU3tyx3gotzcL0lCVCxLjX+WdPHa9FXrA+AJLavTSNMISEgm7K9SbqKmk/uj8FqQosO6AdNgsLYd
WRBS7foocX7U/67XLRW5Lwglo0y8vT24w3uk9vyxon4S9L8MPtm09V1qivOblsLA1X17Fu32gc7+
3Lb9ccl4rkR9XyGzdpBNITDye6dfJtVME69wUK+uZIvshFz0JCIhCAcObvyFdgH/8LbUJFAPKi3H
ajRW2Hp97NsMGX1qbGJotRQuTwm074eFfs7YaLnKXWUO56/lMAofCTaRGSeXWZarxw/xEgiQSORK
0LUASE5YP7W0seYAsKeTZ0iC8QBtjxSGG+usANtOLz9O0KsVu4DPyxtPn+TW9fG9vKjaiBbAKo3T
nOldWZJpnTl1Las0vqsKbzTj0Fr699m5uijzwA0DwVxPVD/t3TSBbGnRg46GZL7ljCxUj5N1jn57
ZM6vZ7UK96c2YvXkCoXbZAGnoXISxMq00e46z3zGSwUTJTD00M1jA7IJVA9zvdt5+hla072xsjdI
5sLyGBO+OIJF1JBF/DmJilTGHDKM2gjkvTSbk8dYDJ60+flbBK/0Z1izjIgkrwR0TIjMGPVsOwUu
rxw/gKIqafjLGto0fEfHBt7JFRbH7mW6CDDYoSjM0KsQrS+qMeqhDRBEksxDotwQ2pSu0gd62duT
cg6OSPi7Uk4IVG/xNPpC6H3vGpa0N4IDg1JboMSjYR3iwySFNh41SU6ew85KAOaZhJqQfTNlrn0v
Jn1myApA5MhsXEyAplo0SxZorwogUXy7GgE3BlL8CKHVaWe+Ar2m+/RPM+xyUwNXwQd9CTVg8WMl
bqiHYXkVWCMMiogiMlesJ2ygYOBddp1DaGl57Ffwc+wkXVeHPCYnIBhaJx0gZVC6JHNUmlHB68RN
9ajQX+ArMe59uK+ZhysVsTn+OJL6WDJV9uxQhxHXFFlxXAjnK62nMRKNcX0tA3+Vw3o4JHb8evNc
Um8fywVLScjSKNlfISfU/0yrSZdwMoitmri8sYKp63VgIQOT7pRJLaNrixv9wp3g8dKLOh4YHCBI
bvmdBDzFfwPGDhSjL9aIm8/LggEey2SrTss+L6dB6vPJgREDVo+Er/N3Hf9aZsnnOpVLM2q80AgB
kAqOXG4PMaKbWfY0bNgcOzBKt6bWkVC9Pcsa0TMFzfdjgoBszWElXMTt8YwSE5ooVetum50dhwEr
7Cli67IpyFoXxPBryXWqC5PonvPqapA892LYVpFv4BsiL6xiFBXdPg7aRP1gf2bh7Lubeb2EId92
DsZB87f+IjUiqIg9W5oP0OdIQRPzfkwICv8u1+IiauvBlADJgOGddCWA0qwBJk5JQLEsbm/+fMM8
KZXeCCP95/4p2WqijSUt7eJ2K021CJ6Zs8F8rtfJktL0tNRzLer0mOI4rOEIDdMmkiFyvUhBTCeX
M/tetwzCfGWTcY2anEYectqKdsLWdb013iefCOO2fRhEBnLtgQCTupPZfIuZujLoIh9WRx2xnbpo
tcYmrmC4BcAaw2984XYkHmvuMGphKLzpsQnrhUp1x//wGmxXEQn9/FhAGXUuDnaFUrbdiL7aSOUc
uI+ZkKHiejDE1ZU7/eWSQNBzhLSpkSq14mPBmlESCM0ELC9MVY4DuIvjz9J78dTA47aTsoPvcYv+
VAIMAojZlEPIdkm6BaGdAIsp3+NdLs6fQ0dYXdfbQn2iKHnfMKbXGBzB2F5Drn+k3mGzqGTQbGHL
7KaDBVIIg6nCLWOC4M2lrmb3z1s9LXpQu6G6LubYROK42d0UMCG1lB+jFh2ZaU4MBXc2t2CHdUoz
D2RRw6uLRtblwQaQypPJCp5Hjn7qfONeG9ZlUKOjNUhOZwEYeX5TyyCOMP/o9B0BW9IIHtXeZ5uD
Vv09nvbUMCET3tP1qpn9KKoaPUa92rUnV+F2xOZYQRCNUvnGClJVr5r680Nn953hdw9QektPmlWh
wPB9P33q8opQ3tNBrZmbGKliCo+OqeFp0m0a9p+hxdKVojHFr9M+nWzHQ+IVTV6tgXkXjfCTm5+m
CLOKaXGQ0e+rF0LoUIlrQJtclZjYLaAjBd6rkNXASqEH4fGaWnfI8g1NSfMEyDFhQ9XT6lGUx9EU
aWsAe/1N0zICyV8oW7O0W1s3llorHQRQlsdasmXV0WbGoDGnlhJgXXjxyT2u3RwxQYB+gh0K9f1v
7r0Ckt2iA7ZVVVURv4jFygi5nB80MQiqMOrMx4bO2jx/oIyM0acdEyEnxi/1il4KDvCeUxpRcjnn
qDO7dJikP0AvDIPvU7hjjS/n10y7GSxzQTje+sa4t9zue5FBv6erDsX/YUGB8m0IASm6Jb3VLJcS
ztKcsHSD/pfg/V5ZlQOrbynrYgux0Ny4m24p3slkuiFdMiddW6+rE06J8ENqjEtBTQtuCm+SOpjA
3kNtoqwtv+DQisnPo/RJBS8YrOlwjZL0t4d9/CXumRwOlcF7ylcv/Cs5sGxZ2P430kRDl3FMhZ2H
5k3JYflTWHANxTfuo7xlOKBe0scQd89bsqDasM/YjHiVBDV2srw9UkvyDeBzxkTkj3Kmrt5BVdzD
YLVPEyQUOCr8Q+MwQpNdQUW6hBWxgoJnAjt/TafKXhGMW+wKUlQSVGpVr0Xz7p0B1BGYPWuCfJc1
omXBRi/7veToFtuue19m0Uy3hPHY8enb4F4njSzxQmz4UPnBhDn+17t1PSmQEq9uk+sXmMzFhQhZ
zaP7Z4wMTECwGSXQVYSBhjgNzUVo8xxlrqZkJsF882EgmxpV8/SKACGN7rllcau23UjLcJzltE85
n8dn1JfXZc7V/lj6rIlATvW5NQTmb1M7B4mLt6qdrNjmBPv0Q1Aj6iPCiAZEIqde4GLsGAGY8THC
X5Ce+ovsQ/vjAsctaiIOYSB0YwlOueV5JulGWmJvdfCbQ2F8d0jISFs72tvDGY5TEqX1788WuDCY
uU+67o1+g8+7jiI704N7vyjK6XKtOQSEtRoFDdyzdX0qSPyQqeuzfXo34VbICsdUXpspRCfQblf8
iy5jfduy6lRoPbORHQUWvQiHrsYiiQIPFWJundvnMUyAT9Opx04pRAflt7b0aYWtNXj2NtVTfZ5P
E2Sp7b8GqGn9AdPrZs9N0BHzwRUjl8mqIKGrNM2Ce0dqYDKfxDLqwkCPQ4UkeD/rUtpq0O0eJ/0k
8RzS8GpcNq38qPDpLoFIrFWMuaxkbZ/tmUT2N78JVWi6F0d78Xhiax3anN0u9XSwBIQ0drQ+Wh18
zVlOUENHABneJZgwT/wvVk1rJ6Ni2g/luGFD1UY99AMfFHdbAX82Y03k1kw+L1R9ijvEVvF/h9wr
spNbAb2gJrS6HNeQ0Cla3QFXdZ0TVWP/0T82XfEG+OW40XPvuleYXx6ssxad8dCkc9zNX/+4sjOb
iV8b7I5L0jAi2nQOiRhoOe2CP+qOSAc+uxsmJg3AhWABG7EDMPSQV8gjjYwtXoQwf971A3Qo+nGL
itg6S6KAzcOZLGNuYeMR88PZCCPJ5bFcFCowaiLDOIdc2vjzksfzZI5yD1GwLmC/LHQ/ALTNfQt/
GE368ZzPB6IRpqjbsPDM1GUfNJ5gRt4L3qqPK3OAba5SquT6wxP2xGLWg5Yx0+vgfoezDC9o+A2N
5NHwj3tPKA9a5xArsIJvCiQAA2cB6ySyS5susaPvxPVUijd65YSPvvARe366wrJeliZ/0BLUhgFV
z3Y+Hz8cH+PMS0/mkDv5OX8U4FhD7qAy/AhHMS2SGQU7+6M8Fa2LMv0em0un6YpRa5/6pWkLMLV7
u8pY24xCx0i6C1WGMHcowwnKQYw4IfaoDh/MdGNa8C9YmSVEt3gOlqEKielrYHTqRoSSuZ7W4ma8
0l7QZuArbmjZboKfgFZsNDLW6CRH3VldC4G56xeMrzuNihQc7FU5iP9XxO0+rotYjEI5i8JnJKtk
LMnCTLYu3wZm+Pxv4aVx8WHxAPI9xZUQGS7UkZ2veN7V6dh143pAGI/F4dFJDvOgeqxcr2VHXPCc
mTUlWc8cyU1wvwR7eWGy+VrRor+T74fpApk6BPLQDeasPbxhCejrsD78GYVimkUDhirBYjiS19H4
tsrayY9HhMGbxc93mWMYUEH2K7RlWjZOj6WpLp73s4q0d/MYAFkjZ3PIDCpI0Tz1U6THfWvskGhc
0YoQptDIwU3IZoiLIXznI0MdCroY1dTd5hTiuUCCW44MZUFUH6nYG15rwnI1QDZf0eQs0KbPKg4u
PlwJp2E8lFaTBP2nxXErixTBezFBcvbeh49/MjGOfZ/GYWsEur/EXw2CQTVohea4w6qFfFH5MH0K
9tX6g2HAeEN2k5elTyEwP+p4yDr1vk5s8/GWlx9ImrtRl/o9/BZ3/3NUFW/AnoQqeo9cXYXjkUph
Tp1GGAdteW7ATaKbiWz+/GylK27oVGTFPOp94YtGFNc0DYJlBANQqByiC00p2B8CTc/aPITdXa/H
ycOTXDicjyx7RMTs4JkbZNrJjBrAU4cPHXbG/+62RE9RyrRU36n6l8y2Cj0+DiPvwtm21GFhRQTD
IQWJ3qOVUzGohSxtn5FIeQAWw7V6XoRWD/6v7hYyUhsESeO1OrBxKK2thmrGrB0XrFECUf319+Vv
4BYiQrjzZiby/1NShQPu4nxZrJInRNmAHjdrkZ1X/CAH9Ua1r1U9e+p8UbTdgHUTRRpCwo9Ib1t+
8XSzFxrkaFHgThN+uUBdS/oMSo+yw4eRkxz/PjxEP6lZYFgRlaswtC4EdqjT8yZbJIoctQJcufab
T2aSKGiXnrztnRIeMHDTzXKAtekKFF2VyPiiCWhZ7hHxjmeWqgOSuH7vxFHA2Qq0VM4qgZQtW4Wo
PK4ySWNScUGHuK89NsB4hsMgvY5M7sPjuiDnXhCofrIeb3ZOt5tnL7eLTGZFRRPWqbNWCoghTIqr
LtPgw4qoGdAfEOm8nW7bdMbjBI+UIT0HcZt5vDI8tucM8dRGFJejf8eQY8Gjn1rdSIJnoFQAY+y7
NeodZ39WJ3c00UvNsWYENolOdO6UDhikyHJvKSbrjAxGyF7LShYZ8a5YtWhFsi1RYJUtsKLQC5Op
DU6wRn1ZsR9p7uCzQsAqB0fPqeqY1vgu83m4y2I3dlf9d285BX9P373M2aCjZT6Klwq+XSri+9NB
FoTDgbB/P1V8kOBU/JT6fXk6IrASyNn9B+KtDyfmFi9lM9gSh3+2FhpAzfJNmLmvhEnEi4tGa20J
S92xJ4XAEyDLoSwfa6BeAiBLhrjfhkqBrF5Ymg7staWmqtPlurKmxUPHs14ote+f/lj5SW8pOU0j
aJO77nLSGsx8G6Jsh3iDPnryhjpn0Cx1hH76au2N7Xoc0Ocpdb1u9WiZT3aQHU7diZlIW6Qp/feN
8iwKJ8rTg/7MGYRHlyB1Lx8t1Q9dyVsC16HEK7hTVwfZSBP7DjUVbLeavfmH3wB/Lv/8T1J6Vj2Y
D7HTpwmIOKE1ASmAtuqGlDGU/LOp8FcwfWWhZ33PxihPom30d1Dd56IEPNIIFljCkh/zoHg/H0Oe
0ZU0TX1GZjIue4rQ98/HP2LGZOpbtJW3sWY39me7fZGonhrOzFmlYq+nVSQZ3/B1y5yQYYoX48mu
uN0BYJnFtklU66rRpE0mSz8Xsif2cix4GTZZ2u1pMPP+Rl8mDGk5KNFiViYIK5Kq0A4LvReqH6Wf
2CWtNCFNdKU7Le8MqMHkXVQHu6e4hH7qCxJW/58olMWG19as54fRkjhiCjJS7LLUFRoDiQkkWauK
k8LOCTjiCPk8hnpNHcuIPGAWvEA80LVh8tCWAWH/pOddV1QbsrP9K3hP7GPHhqbtdcsFWUKTEwBi
es8RT3cp6wUTKZ0a1yMsA+Ox67Ry1cAnfJX6Od3It2BpcFpqqgiH4NMl/WFOcAxRfg5rXvLJPx1q
tpW/UOO9X26s1iep3mirHXeegcQ4nToN7Dv7U7DwdMKoig72HXHIdMCDEfCp0YK+7Z49S1lBXHV+
dh5b/XxfxJ7XivC9mzBz2GESLgxLW0JE44W7p/wd+tpoLBLsrXGqwbOQSuy62KIfffqlNMGB8dxD
WmHfgMo7aA6/8SE8Dj9VjZRBxQHyVR5vba28Qj17wjsIj/4xKVigXE8gK+n9PWwUvMiw5sB9/EEm
8Ul+212GVlBTfgvXsx70rfze0B7CfHfnyaO70GadFlP0lq0/X/HIRaCcwg65rmO+q662Yy4l93/c
HzKXVi+OvhLkjZUdMwcu9jumitA2fI6tVsdC1bAajZPOBesKxB/KIyR2TEZnPcNbu2ObeVTiEryI
ahJil9bUJcTGcJaXH0b7bBbLf7J1UhkZwld8n2yI+qvClDDF78eVtzivHnZd5DgETc/CaC2kg3Ph
SBu6wyXtf1KswRMGdFZgoMaB9jio475dBOQlJzzAcBMueqziwfsqoBBfASr9QwpKXbFmwnMT7rF6
Cy1eIxz9d4IpkEJDFgfqFDsp7q355M4kn5zcQdA7syXfr/WRRfArltmNmCEQyWMSkJ4MpYUUBJRx
DwKyhCPs8vyMySfl7fwJF502xfYZ/gJw4v0VIjUZi9wTpqv20/gf9++QT020AyxLO05huk4lOm/o
rByTmt/sB3/vtBd3d/6oGDsLZYUWpoXWqpNEAHciLEaHxq3RMSZTXC4rvC/0cEcN+bPe+l5F+ttX
4niLKmXhl9vNEYOJel0b2ZgvLpLz4nyQJZQS778ZkfgTaRCGNm8DIi1Hw8J09idXXKenROR/gzRz
SYZqHqkhyo5AJ00kjdmYx3t8XgEW9E/xPrzj9EM77yBK91npYPT65c8ZVboTqL5aw7qudOnaqOCf
DkL0wSXwht1LZR3EEP6GQNd5UWPQpWP2B3+fmGQBeLVP355jDsZhdzT6GlVG+iM2kXNr9FpnDRxV
giAPRl38wwQrwloqzZ58mitj2lYfFEkCkatOhJzKmz26qktOY4udr1RjYGZAZKhZ5uwrEhV/NzMo
KWn9oRHafbeeLIjwmZzOnKbvTteMSBprQeuDBdplIQK6ZYrb8fVNOfv1e1y/ChJroEdZp28RPJh2
mgcGIV8NPHEC5dBO8U+5xLKR5+GdIsRyhZ+2KRf3aONuDleb4bEnAw0wLkWa5Qe/qWaV1p+rPahn
FvkDIiEO6djy3Z2JY9LwFfSs7Q8ULtXsashjldxQh/pYO9ekUXvWjPedeJKxHMmdeVVx8ueblf9b
P4gyC7dNnSNiG7mnYklM+tC/hjngqSuobSMp/rWW2wN2BucTljTpiNZdbyssF8BwdfX4zfUF71XD
s/SHCt53bzvgFa1tZSCLx++658Ebas3kE3IbM22zF8BIjT6978jnndCwSbrsHq9dbVwiEtv618Lp
tw72aMgzaGOKsiuPcsgx5pRq5Rw2fu0V4i4hKDwK88xpSB/DZ1wfOKg70zEHmswiXcajGYCkMNSM
d+po+VGO8kopz2MbbYxjpdp7BnbFJ21CflBZhEKXeJVxAuGPshRD8Rh9yjsdA1ly64hmVgcO7+3o
eoAw/r7eybXG7aZdee2dXjUUtxr9yfJi5C7AV08qoq13IBTMAjE+ToL6aqkrkd+HG7yTADwoYvd7
57/dAAOJjR6s86uM5lk6Lp7xjltpInJy5FBcVaUXtD4eJ8nVGmI4n5uzbx6KODl4JXLF32U2bTsj
FC4a8CXjq26C7gTj9T0p2fr1v0n3sOib6JOQgmQYQ1Q4eouhaJC//a30PNRVjxIZDhEJD818eR7a
UoOjW9nUDBYIOEvjFc+RH+ISRIJc6f+XCrppYz2Qq8pATV3tft2wcqpT3uamIaiPGbBMYjuTk0HU
RcktSDxJ5q2hZb8NQWXidrVRIWE8qMXqQf2t6h5NmXQEHb7UjERCHcG2+QOkMmU0UFdx+DFc4Re3
XEc68cIJXdzxB3JYmEnLNjF7UWLKv25Y4djuKUSP7VnWzmmSWCwQqqHhDalTb5TYCB5+mr8HTBZW
J4UsHg+c5d3V1FA1mNeViwqqBMDvoq4oG8UX79846O1PHnLXY7kIJfy+siW0/L9J3xzGgva9XnVV
2dBBxgFUhLnjPs67g6X3zB8HTw0wk3iIrkhQIlYqBAN5WRPp80+AxhzbeVmJ2uaHcC68usLpw1Sz
VVDw3RXNuUBA/vq+Zh4HAtMievFy45DacfZUdsO0fc/ARXaxiMMxd9W+JyQxVUFVyVNCoIqOu4dc
FMmjgQRXb33MofkwHhO1nFIBab01Fp11rW7J695ilshND273NiUSqxPw9Jl7Zwsb3ItwzHvWp8J8
kk6x2+Zo6XyEeAAP4mfKsod272q2tjkQ0FFVQVc5ZyxI7NPgWn3R9lGlQZhcqEiRc1Fxm+tKQeRh
YCQO2Mu/ei374jq8UlErhJv8o5ZSNmLPeyoEGJNlFB6gBGrpQLPgaU6ptb4gafJrwTDbyCIEqCCo
RSPMGWiUHH0aBP99SH7RIEYUI7twnkB3axs/JCRtJOAYV4EUARnnQDpdcSOiIA4ZkbFj9RC+JRih
hif+JcHnLWAdsZbTpkUdnhvbGbjcjl44V1RZHTOfr5vWmh8bmb4Tq3LysK7jJVdFr9uvZ+uStgTm
meMIe3rDuMmMuslgljhGCAFPW+H2k6AC2SrLixPKF7KUfAEMxTCsHgFAmHtNISK0HCT6yceaizFQ
+6WODvM1OeBt3ol+4H6yWlEOZMjN0j06riJ4kURYusDN5Z9HXz1CcmKus1hKXJWlb5WGVbiFA6Ej
FpfMkpMpD6QAZRqM/5gRX/IQ/e4yvEfOnr9BSWk3+TKSOXaZHwl7xvIGRmtQ+AVuC4H5JpWqm43C
dMKm4uzp4HoRXDzl7tS4TCHD5SsmbmvqLn0DQFF1Pzy32vXe88Y0UPashEaoxvJ/3ufneGyUx5mn
VpiyVy21GtcMoqxti6V6z1T4VtDf1sY1lvEZ0SOPjCL4VfX/B/2O0/by8NBW9jz/7idSecFho56B
WKr2SfbGFY8jtHyDoHq1ulY6oKKMLejJ3GLurNX7jsQDEE03NK5y13p1Gsgqh3yoHcJA6FpMTeTz
UxSjwlDPK+RhOPzwb39P9YoQ4vRSQmS6D6XQ92wSK/zKcWTVi3hCed8JJhIqwy//rPAxfv4TUFd/
0CRMl+e7yW9VpGvrGyZfB9JFX3zRdY+ugiD1OGSQ2kojHGwtfhviaWo73c2m2JZdat3kKrPomK6E
Q9P0dvJgcU5Ow8B0v/zFuLTpRBwXcfW98XNQmxDtIM/Mpy5g+vZjZnAvPiAhPTWJirlzyDFsjtZb
drKUDPj3CRpa3oWXyCMYxkOT1g5a3Ju8+ny7XL0xBQaYdpw2wZvezWqRuhglmY3Mb3FobQswUZvD
Osa4mIu69zyEHIQJETw3Hb2ENxXny5bBiZ8rdP8f56yFegwELxb1Vqp+03/VCxiBpNx6RGs/o3kX
a5SEzuysGETFLwx6XdEb/r4BgVk09LyIOErkTCyRuBOLZJjoKzbzWI9FR8ltBUufsnxbwV2Pm/kF
EQ/SyIiPYU/vGheDrbPF+u3xOS+PjB7Zejel2C93yvIL+27+WV5C4TVOj7sQuwVT/v2D5SggJqFa
nJNqAUODP116DVTT37yWRLtzJJyJ/WlIRTzLaENsXF/t7+s8UJJULAET0lmV66r6m6gBoU7h7mIs
SvM+KYm+/ANUpCyWIbM+CdoMBIxDqI2rCzcMliqWSNsBU/5kpatBKcQrAyasyNmx8Z9RzatJsweY
exYktBCGzv9i/0URfJ3Q2Cyf5OlWEkzkoXDOuSd6YAg6Z68rNPdeGsw5zvcUKgMwMwS00zqcNFNb
rp3s4XMgdWBrx3z4RYXwq1Vi8TPZAgJhDub9j0ieoBQNp2RH1c0KWCK9pRheXUeQwNET6hUbcP0k
RzX4Y5p2JcyVbDFVHNlL3Jw+SEwHs5Txy6XWiO8kQVAPuiMpLA1qcdG4wUgQSCn+N5WOhnVumZPu
Mi193OPQqD2y4FVwvXczX+dwQkyyuZZI9o9C6l5KjHgSWJBo9xor5D1YlwaMd8j/x8n3g4MIg0Bl
2AmPETY6wv1K2rbN/n7lTu78/B6kPNyJv07KkfiQQIlePXCfPCh0DrED73lq+zQRCWFsxlp0/WS9
LVP+hJeKRXkUnuCi0JtPCeIRnx90xxHNXHQMGJL3xa7TAFvx0zGuBjJGbNAZ+DqfR0KZzCn5/hZK
rKLZ+GhXYpXsGFtewcCPPy6WXXrk0oFmXJrVPoP2zXDhnNvvoTZDNKvDJLyLBsow0hNLWQiUoDZD
uYBysLnis9FELbFE01ufrj1w1GPXiHa/WLq0/FP48teMeexaMZQGy1pBFW15gMANmhfH523hJV44
nB8fIu/o6J5Q56Qvff6peBsBfvIZ21F4+bRg5Egux36o/P0HrLARyd5eufVUqM3P6D0kao0nnM9L
s/vOhS3tgJLR0m7kzdn4ba0AeGwMgwMK34A5TuLJ209lxmiZue2t87OAQfx9ef/M25M4b9P+qDgG
zzP0tONCHNwG1qMkof8tMgul4m9z8xE9cD1hpigdgN8BxN0vgki1vZhsD/s4lfdW31LvCx3oSwT5
l+58SSZ48NOIZUjq+E7lIdipocswxhaqppYDEI3mOG8NnAX+riJMuOWbHGiFhFfpgFtFV60IxWrh
FUg+N05y4Ug+AMvjZYyYjJqCeh6mjqJssi3Bm9PrXLf5s98m6+q975anKbRXcEEptCv//AkEb7mr
S5tPJGrLJdVzec5MIJQXk8rE1cD8ekft7bx3DM4CaQXXG0uD/o+Wd5TP8fstNrzdckBgGfdYjkcs
644a9fFMxpeS4fNymhbVGA8ECCWbrYl7YR6Rp2lzMZ8W5G3DwAs/O+B37W1XdrjaYFkQqTi+H/9O
sOa//b7AwK8D1JfLsBN3OhaSFeA1gISqf9WPRI5/CM3g5blTjZ/ZLbiSCD3ZAyhr0gjIKRa+l1Yv
GcLoaTnTYi7v6fp5h02A9oCXLBJMAG1DRfZBbM0yT97W5UbfPrYpRq6yYuRiT3b/PStgUspR4V+b
wjDm8GT3Ar/jlNNWxM4tAuSyGew4DuKAp6TFZwOUWWUs08MAHndsQftGoDEpGuoRva1Y5IXUArx1
PzJEHtWnq1+kFnelOeQaMdgNcW5Gd02fpdjJ1yCOjV2lNU+vRr5mffjXV0Cho9IAT4pnb85ykeCW
SZDYXEeG4vM8YAFgb2/lIpXhJs/xGgAUZvpD4RZR/xxM9qjjbZwSsWhmVklY5Y+hUcDGfbj7JWWw
4ISM+Ws6PGJ78e7x5ZMP9VSha8vC65ZW9xIl/hC3SxzXXiejim61OhL3t0A1Qmfvfiv2DwkB3b2q
/JnPGckAQuC7nl6F61GQU/DJlj94ABVv3XtZrwFpxoqrdPQqE5WTZaDDFSN78prDOUMH7hgDhslU
Esv4YaVDKIyHxHJwnPK5e3+A8OzYVNyHFLPcngio7eN4jHEHjeAzg73iYuBwdJECRjSSCG9KLp3q
ZmZfC5gl7Nj/+bMz7ow2QIOeNyV2igkW4/xByNzyp3pyYuHulzQoZ3lFIiyAShzD2ynB3qa4vYfG
ZWG2i9Y+ZT4HMnL00Abiark08naZuighDBZuRhau84LYrP7IlBd+4He5XYFjDmZqi3xo9YJ4VAG+
7iXTAVL5aFyDNoi2oOdcTvu6WhGdeyfVCxRc3Q3yIk3yMaPDXbwLZDQX/H0muuBgkW8enfLFf9mh
2zJXj7kmSo2nFYZEeNE7R/COKTGWWKv3icSsn9St59fVM1wau4C1QPYrDfKRsqrBwb4JOn33ppw5
aLJ3BsfB7FegRG06UMAZN4tLPDQa/bTpO6ITI5MYhKQeOJG9y306Nc2fY7b6NJ4j7Pr4bcj7S8Iu
MLuv3XxbJmTknBNmLwqgQilkRQO5oOYTtktpnR3beL1U4Uqita37qlmnbqdcsbp/LgSyR66uLQBB
3mXXjkqhWT4xNa4J0t/ytERNuowvk9SnO89lenF4IG4kiqnW5655droVPMaKDr/eZWKAX/FcJQc/
aByT10jygcqg3KX1cZGSKv4GvZ88DAvc2TApeyzqH3RShb5xTAjxwynoxpplWYnNCDhSGXHfeewC
zdcPqOXZOHgyXhWU2OSNWVJJ5fSFDH6iSjTanqaAnkZ/X6TbYqmqkJ92HuFZngovb2b48zinVGuC
pHvxdJSnR15ruEUETiSKb5b8BDnpBzUZb65Tus/3mJauqzrF/O8Qb7h5MmVZ2isOn6FCWFO1WRYJ
CczueKZ9CNezbnvRoIhDKQGAFfwYhdzv7BdyvA3bdjZ1il/l/xtjrLaOOqqeaB6fFEJYK/3BU6qe
n9/d8AHdfP8Shcs8H5fDseoLbH34eYbQhcjpc9SgroYMwCEYIBV0IdfbhVUSKkuKTTli/SMRri30
NC7rl+wgNIG+EodzJr6t4InbOM55n6Kc2b5gRLdnwMTRftKoUFsfUgyLcKR6o4aHHVOFpjZfPA1d
lPS7QX+ZXsAwqjxRC7E1RjplpQfTgYg8DCtLc88sIlwTvDxcuYxLGRO6qENs1MwHylpO/tZHm15/
se1O16kdkE3MjvUgnrileOA2k7hthcnwNBlZf2ioosv0ABGqecaGxc0A/lhDjXGLuVDf/VIqUDFd
+EOrUeGkoD9xWVw/Tq/I4/Wd4EDFMGcR8gtWUxGQGeI7rrb9I08GiaWwMo75U+KAiWfxp5TrD5CV
W5C/hmFYm7o8KhNy3NzgQjbGlKuKH293BWm9em7QBhwfOfNPmtFUimfTEIOxuobjiAXtwhtqFiMc
FdZQEsFJJBI4OFljW/LyeAynN45sgWHy52hW01Ym1XjNKAoLe4obIbKz2a/s+C7Tq7wtByXWVH/Q
gVmVHo4D2MP7iaqvH8212Oo30XfW48kAybHUwIu6Yt854Wxmdj0T6oBOWjLhwrqpw5DtL7ojftoa
s5FqpG5PWDmSJtvl3pvdDdDZxoPfxUishceUA49D648DWW8//pGEqPJT298o4W8CMPIMZ1S+8J0+
7SeJJ7Bwe2jnL9CjKOlU/RE+qfqVgTR5bV8rISDYuNey7gTfO8bcEB6LSXO7vnufosAShAXXaBpw
ofwrYqO27CUf/pGP3uHB5O+m5jJU8iPQ/uy2Pq4Wo3NcXC3ReGSSgsn/X/HzOyP1TEUhdXPrtu2B
eNhfSk4sACwNDmwB2N/FQ6OslyCocBH3yfy/3Yb0rxLajpiXVWdkXyZFTDKMFEkr5sFOG4s2fbU6
tA0Lwma/Lrr7Ci/G3rDw7GtDov58bu72SVYvGEmHxh0BkcDMw6USI9Dg8e8kOczcfHjtpFYLKGl5
+bnlxljvzsp8f1fOwDUEUC8vvlcemcPblEr6qgjjD8/kZR13qn1od3F5HWiWCKQHSmHbvPDt3zCK
IAni0dVECrSS3bfZP0nn+dqtJWSjvmYqPBfbbmpZqIlVAFM9xYwPYNEdKSKUzUDav9PHGcUCcZL0
so9nU1utFfqKBvqPnx1BL/ZGeN+sjpp67Mye/FRymmv2oM15y10EuS+5nHHYxW6/G6w93KhGZ88y
XuTa3qdZld4PsUEA4loHaaH5IzGrDZSXr+HQKTZdJMwx73bWqd4qMV6QM8tbcWY5sZ2O74zotxr8
ca8KPl+iYWJipwnZgvkuSerfy1v7B0bNzIyeZX771B9QQcOmhKQLYLwHGD5pskaqAJhxehHUaYiB
uqDO8RII8NZ4z/zxsMUrIEbxr3wJBBtS9QP3sojao2JTh9tCVTRXTriSFOwadz5UE49yAH7m+AC+
Cjh5TKVHyMymNDDiAOz+50dszG49e2F98tFxF54cCPL35pcM6rmHrnu0gujc+XveDU/s3kFOJKJz
sjhDeeg0rcyTeurAPDkdxLjIgGO5yobIdWWWNLZr7kT/KIEZEoFH3OGhsUQx0/FbUZOVJvreBW4/
nFcwwW4VJYlH+5Q23bdXbish3em5QEY/yPfyyHcUxIgQndtW9F8/flEEOI/qNv9xtU0vhX63xHgf
nXPdZ4HuNrg7zhFb7+wdPse7ONahYuqwj5A1w6dccWluUg5GXW0eUvrWeQh8g4j06ZHwbtqqFmn4
expe2Z4OMqmZe+HJ/xagsGVr8zPH3G/rXRS9lGo6ZokMtPjt+EDWasdM5i4wpOWUdYy/w9PEaZJS
KOork8Z+PaHsYKczvmGJFTaPGtkNSFJocfOPKhTIsIEbyzMLk6Ym3jmw9O7Oi6kYxt067X/quqZs
sC7WX6UlGzCzURFr6YACtzDoEVtOM6fpgDTU/i5edYMwxow9K41aVwXRBao8itSTrekqsxonMCHg
GM42peZdZKrt2Jk5erQR2bG5aEomJBhvWF1i/R0jaTJVVfZQf50cOiUsdSHmgqzh+WYDXc9RzKNs
9NkLsWYn3dN7gjEqzuCGrsm+cfPOExh3nXWJ9t5NnAOp4ej/GJzZuajG2Vfi3RNuE5EE0Pkzwxe+
fTQezHvd/SVPLl9yEqgr4ynvgZUkD6V0M3540U8FHgu0WrC6L6x3p//3ZEuEtvE+CBgpnqLHNBkx
lBwWWE9xTT0yDm8dKvtmi6iB99xXS6pU9drxmEoaJvkFwSkCVwMz9gTL6xQuq8kmmKcGQ20CnFHq
pwZLiBIgi1di7GPMaav5+aFZeReKLyUTveEB93JMIENtHgYr0T5jyhJuJzzU1UIwiVptdH2k3y/A
gCebVpHS+QcATuxLsgpeM+6Wz/kH86E1oz94ahQyH19IA71IFAf+noHCOEC3lcQkOFvSNhmmcAF9
5Uc8hEwhyk8BTGK9cADEKdAheO0z4wvwjxRPTgvmEMxBthOcIdl1fzGeP5yUAoi4zeUMGWQFcLJ4
yxLq90PyUOAnoCOce6gdz6GrPMnKvdggzxNG3Ui4h7Kuo1aMHsVDXcjkqhz204HjfNeigLfA9ZAz
vjryrTQ4hi02GcHWBrN8CQDUwvNDpHq2CuI/Z3xyiu9gwSZ0wnECQuAGQ0VHmoyKXygmjFYdnatB
0hu6VbYMoR/8PtK+AWaY0/2NfekBEIzPIiXUxDeh5csIAfhM6ABJFC9aWNNn1D9/aj43k5YmFjhC
BovuklR8XZCpfGuV+d2vKBTVNT/4g9XjJtXVa43zWrAfueZ2AEJlPw+DOQlw0x2DOaUeUVIkBrxm
p3/R6w9DMK/ctUrhpHm+uq0klkQoqLQMn+H1ymUAdwdZlndqz5Ic5gFsHC2SnvwnnhrHFIJ0S5Em
Thl5XiTiDdBU5yuk+5CIDlZbK7HfhAUDgBPe2Ah84T9dzisITOJmBqWgCGCr9dhVdgqcTNbpcKja
4DqXbEfNQMkkm3HFrXVmZ3Ac1sVh5dFBbbbOzlDrMuocrmY9hQTjNEIXZM2VhGzR5rPKzTVlqGbK
LExNRk5Nq4yJJIK26UquEszBUq9LqD53K41gJD5vZQjWQ30sRQY4DZOcshFSmiXKgVkS7nKvB2hv
VUiBCFunuiPCf1MOMhmq1QRuYF3+9qZQUfy1P3QI2tnCoGk/UTvbMBaMtyxNYi92huVRTRilQ4jN
jYUhduaLSwYFNRPRgj6/wM21PGZxMzu+ILeAmGY0Shsa58qwMmfSf8q6JyVPAzcAtrleVDoBYI4A
gyF3txw9NBDqmkUjd4Ndd0wZjPOOjlixsE7AMFtBWfwJmXCAQhaQ5fCPK3gvQeThXEy/2FeH7uxj
8IYEDjh4MmrTt4KE4oc4NOGoy5gLmA6GG0/bEB+qXFsdoIiNOGERUDEKuBQ7yMJicIe/9rXJWv0g
PDK81frDnXFvChMWYNcKaYqTiOZXJy3coLSFStnr/+ugbvGtHMJw9ewo0IEWHpbtfgHQLsWtZKDd
HpXrC6QRAHSk1RZLczEAUB5/I+T9y/yX7OpfjbhCGWVRDDHar9wPIZ7ztpx59NZX+3OSEw8Bro5e
kB1+QG5gi4xHLMX9m1gWm3qwmSuog8/mj21ROkoPZu/rTT7naLlivveDxrGOlSn19BkAaVTNq6Eb
iiwyhbiai79p8CCcjV13YcqoyGlll6gmEjYKcxqsl+KgWZOFG0eYxExKm7I4fREpY86zRr7tsRmG
TBILTEDLSm3wiMl7vjA888CjcOji2E74j7q1lmeviABKqGfDWK0jmXqVosT6Ad8PA40xHU0j3Zmt
FG+eRnrQfS288lBWuXfcapWDfQA7wunwmnuztXWa8X9OOE8uYL6kR+H6t8mSWMmAMOO3Qsl347Fr
lRL/UEbzdgTGVKj/b3hWHXnr6oP2RSbWZQQ81LABjbt21TVWTXlmZTS9QvsB9m9uH0nBqE95sqDT
1a9LWBT0Swa03IRQCJBVI4iL9EENZyH2R4Ob/GYt1gk/lV9zcDDLzXYMvLeXk5aauZkZMph3pa9g
afhh9IbEDE6b2bmDDoJaDt0m6aRqsk6xxfRSBiJNw5ihg40bPpHSrZ9uOHTKtj+YBs2FfokYnADP
YpDvxIChVHiVrB+CLZurVu6xWgTaOyHDw3ekbRDiiLJckAk95EwqewQ44Fv+BXtS9CgCJNZieQku
NDQSRJCiTG0SmHPOAZkA3Byf+97WGnB7xfVNRr6RrhVCcxskJD9xAfIb7ziQ55dxubgc0qwaYaS7
c+X4poHm0STewkGr3tkCuaig6NwngV7ezEPF/G2nfK7Yn4CCgoJDAiEPtzsP1MrNcIArh6QsZIP1
H8/jc8L5vj8k8BuNtdHy4hv7E2iFOngg2jbR5boF3sSjKRV9Y/mJicILvda9QeYdkzX0B5Oa6AvU
VACqOD+I3U7w9SXYUMCLqP9ElxWSD6OqWQywdo3rZba+h01drmVfYqCA7fTCd7aSoT0EsMIp492/
EJU8M1wItGJ0OS1gd/rLrY+Gjl6dHIF6vU98xYnfA6pNK/tslo6ONxY+iBL3YA4f2p9Zqt7Nz40C
U6ktbqWeCrCmKIA0x6CNNLwd0su1Ka9s7ZToCmIrmk4BoWZcvl9zPHHg7UAXsxzqnyaas6hdpNIz
rT3JovAU+vNlZ4oebPCRayywAVmGyJ6r/+qxi/6M+jRCWDHGieL1LVaHE7MuEhMs3XXEbADjc7sX
99biP5rW+wYitI1XmqV2TyAbDXlINGAPOzAViKX4OOKH+UjmlGFS2n/SEjR4tJXo7Q+COboRHwpT
QhnmFE1cSIbWITZJcZzuKT4WA/F577arVoVRo3g63fIwCThsFjcyydn2U9Sr228fDI93acBLYPVG
0CJDUzwjEKkO3LCMgMUU97wzD3NNkJf8YVztDyM6nzWm/1vj2WSP7L/csyqsiWEoUENOTisQRean
33t2nPXOO7uZKB5yUGSEcc39KQGYNl7E3qImbc+Nhj6b7sukqgDV/csIqfNHm6uODb0ktxZs/JgD
vkcOjPqrWPZXk5Qx5MZe3DDOCTMc4Yp5srQMAjrrKibiG/h0WnxtYdpJNraIwY7Zl7FEP9N8KUwA
a4rX/kvT44TYj1QVBH703/eGF7WK8O3F//OpY3nhG53cjuiKygzbdu4KrVyoXFWA0KXgbZ69lvzo
gr7LC/8feGHae/qGV7VoHpcZsbJLqNGCZtTlQtZpV4Zo8gz/8na0hXCA3cSkm7lCtV2Go+LvJHLl
WfLmBgC40IBF7FEAEMCSVcKTfBwZ3NbQl5R4gD3qwrOtGlx1OwtQuuBC6L6JAV5w/A1NdI1AWi/0
OkvsMqc73s2zg3i+uvPxt7UyxHnBE7p0u9jiAmMeHzVXTXejBdFdZJZNm15KvBps8FlfzpKAab4W
VSKh3h+H1xL/OLHCNI/UNLyptHy25XduJyAV4ujB0iLq+L4Ppv28YzcciYLHqIqNAoZdV+wx3TsF
5jRVX7niKlaxrY/kJ5iQKBMbB0F02nbYS1sDV7Z8NDJffs4IfolXfGAKVKCzflYiguFsRleFX4HX
B1pf2+SKKrR6BjU0jL3nQRrumrH8vmC11gY61gSI+NgTLIpEQriy7Yg5IGv23Hv4+StbRRjzWbbo
Y9XD8XcKxymPeQNllsYTYnhFnJY/za8EV76WNTWd9QZXAjugdM38aJGz1DKgvo+7kgYnv4BdpqID
zlq1ZvDlmW4lkgkjJ3GNwZBCIcmd6rRkOvQNAWRT/J6haaehjK4Q3ylb2OfM7VW3164stgGy7+La
TmU+fm6uw5mVLs1SWKCxjCqBdt20PPe70wrAAGPAqxK94vaas7sQSvAH6cuygZ4rEj+P7MvlXA6+
audEHKi+FlUzBNKqeeCwFLOoNjVfoILVJkmUYOt7qAwZazi32fSqnw0VQDRidYiCfHR1oQxgjhWe
GL4RRIRZ5ZFIv3j6gn/GQEX3JPX7sFV/nNJmJnmMC+mCA4VbMGAA3duBpbFhCwKZRgtIkQB2cj22
P9WyvXtbL68HSzCj1Ajau46/ccMeoB1KKhw0BrMD++YAJKYb3Fd+PWZr0RIikuGgjgagAmPvwnSV
97ECIoBKVKkMFSWgS6+z2sgJAehUHC47tdkVpRXnCemFOsgNkaaKyWd3hCVVc/99C4g2V5k4hBzB
XbkQuVXCNyCxz+yK8WXkcACO/u1gBk8Vy3koVMOJBvD28rct6iWtAnuctBQLj9yZAei3IdDVx+bY
9+1rP6ON5OavaJ+WSoQhKQZiNt5iqwy7B47/DMFMF6FATmLJJCL4sq1/TsGjaP/f3i+7lfWduL+g
b6D/w9BOVkL3VB66HDrNraoVELiKyFA52Tm8fv0UPOihTKrzkEZLWcukxDKn8ZeZuC1rkoeYIeVp
t+dNTYPsy0tXvbG10Gu64hP5JXEbWa8zBCQ3sExPp8bO/olw2bX5lcZAgbKrzQ6sJUaQY79qlLwp
o6WObFJZ5KdbsJ79q2Zrah+diHH/zbYkj5BtOyHYuM0EKcDfnJ0D8KoHv/TrwKr+lSNwhE6U9hS2
hfcf4x3AjOCtigH5OvJ8D2Rfq5Ktk0O9bFZeI5r9fWkyL8XT2Pv4yK4EoX9v/Oivai6Xy3G/ieHm
HckB3xhDtGO9wjqLEMiHwe7yWhRIjJ7Iz9N3nJmNkR1Iqqv74VvJyuhF+HSzIjwDZbbbN44T2KuP
hMstEUfJmDQsbdo/XMyg2R7Tm3savDh9ZLs0Sfc7WjH0gm8PnNVSMvko7WIrqnOiwOjG5C9Tfwf7
sDYcd9cidClZi6hSSv2DAgi1+74GgBYGV+rRUggxFEDvT2g9eqYq1TUVkc7HbJs9imSzrCzoh3WE
LC46s195N2C5VRXUCLkXqe5Wg1X5pyjEkYj2qN/rzqq66HWwXUrm8/JS65Lu7ASZ7PE10VdJfHyb
0GXs+tOlwoKh9mmWux7yRKqNoKuqUjR1Zs+ampXju0QujaFLEzrJNf4lYdAGlnlx0RsGK+vQug5L
xIOVrLLhMHbnz34u2lZ+ZeqdimMj0LOxngl4dy+nvXc3OBwLPtnObSUh7r57Ml4kxTE1YjXQ6Mwn
TtVvjsBerNhYC6141RRZ7PHYUfAZ8z40Vg0TG4l0hRJS3HvXrqHKfz4SPIErYNwAMav4tmgyZfWn
N+bfhOv/DNbtzs6xiKZFraZ0vxxZqF9Dm3p6LQIuL/IrBr71DJlkqUXXG5PTmNiNz11bBGA03BpM
21ukMXuDdvQfLSsowpJURT8T8nASj8CA8xYRXJxGSTxCL3n4MqawZGiGF2bwKmoXlw/2d+CXItzo
ik52+AKVOV0HHQLJIG00+F41lXFL8htLbnK18plB5XBQo2KhmmCrLlJRZILVn+jMrcbQHlT3hXOy
TLLurH/BpDv9R3oN1zgl3B1pTbagNNjcz0sGxp9euiPuclaj7tloAEa8L3zSAPUBci/O3PujQ74U
BtLBhcYolN8W9daOW1qFlsQr1sLrwRC7QEFwgfH/Kqt00xd9qV8zQVSqESz+OQkc8eYdXlUOeQdd
r90J7ZqoxZeiWMVRpdd3EdSgudeYdJ29x67HK1o/TZW3N5rFcUqfA9iy9Z4WTGIdon8WANd7CnBa
Qlc0oHKhMYZRlfs6Shwg7gqL0itxocXLGIMJpjWOVleQZGOpyxIRBp1DPDzK9zyI43v4i+ABNJMF
UEOmQXRLaEuw6CDzJVkFNFeQiWDUQ6sjSiWGU92IREhsQmgdnFaTyM7d9ilUYPBMOVUEwWr/XKfL
DZn87lrv4VIRL+K5W2lpE6D9CnQVVb5AolBNgdv9pqEpfpj/55g0rC6lmf6Nt7B2qnA5G0R9Jt8F
rygL17rMijLMHMoolFsveslmuBQAArqwWdD31jQnwSyEJJ5oDJtmyGHonfCimYJn8drLGD4irRaZ
FcB/1huROrVb+HHyLAQl0O2bVLLyDPavxPPMly/X0H9SdOMX8ZdOcP5cHwoONf6OTtu39wrkcjNJ
XPuJsTHmm93WrO526xa9HcVU8234uGkoFD/vs7qIV/gZ5Ds1yEDygDnKOLuZTvPE6SfriRm6LJWC
B7QERuEYBt/bXEUDkjJdcjH0QS9svbuniBbB2bfpip/l9wu3tKmirLdZej7hzetWJ+keycZ8JgJ2
n51DHQf2nMGA4CNIB/N2ga6+XjrfKkS84PjG+zNqgNgnCQ6jw6u0sprWKk83ykvZw4R2swJlpisT
L14gnjThpOHD0Se9xWJQC1wE257unIJbqQD6jrwr5mwqVhyfLmOQF5hua+6goyh2dBHe2hodVA32
9klmZAHAfeh+4g1I77GMhrhMG+UbVGozi3itz8hhwd+iHtyzP9KjUXLMgeZxrY3RPhdGSV8fD5Fl
80jnH6rKqt2L0CYq5S7M5tnr7Oc0J5WTQR+r+1Y2azvDllZE7NQpzu88FyNcEEfYWpo6BvIaVDoF
OdixSc8BKVnr3dSY9Yn7RqkRiQaF2nMVbdCVkhhUlH2rvHOPxBcxekZ/VpYcuyOKbumi7sc3Mfdk
yPIkCBlWvx8/i5NpIxxc0sd24VD0PY+LdlRjpcv9S9gLz/WgUH/Q2tOUDC0ZThVM7vJkPMkkyPSf
rMXXVr5dMRvp0ie1ve3faTlE3X61OVMKorNqLMzzxvkukZoM+eV2HMeMirORr5YYCaiy8+ku4Z0k
B4OzuXnDmP6Dxl3pCYaSZAHuTYmayqTXwJiOm3FIjDij43wVD0mTzZB19bfSXqqwQC2++EgEdkxg
XG8yCBanMCLzlYFhwXbU5lON82jfHUqtFVOcTAte6fQ2quM/amwWooasgu6htGAjGChcZ8bbIPWk
6co9ub08VsLC37mzdeuGo00EdsX+DKhPxfx1GETRg4zl/WfSk+LWyPI6vgo7D0V6++W+avs6+kAA
WRCrpjP1QeyD5GSqLaEROSkf5ONRpAaBHs6kJuwfJ7lSU5snfVwLIYxb7x+Dlv0gFTn6eskOr8Gi
JontQzbYCNT55qsmqRA7Drb0qqxyE+0/t+yYeNC+nrUzatyU23SuKF8GxkNC6hI/ZNMsuYcqTocY
e/vo+3QU2kKgqJ2x7776dB9tHP6Uk5Yk5mUUYX1SEbscBP+SAyc9glTtybmgkV+gXMZe1FlHiy50
Xc37CuzzPe8KUkFlnZeuPvDkGBZgLrKgeEoNlJ25YWBeevcGSWbsDV/7vNRiZzWO1YQfi93eXXsS
4Dhc0THHq4PxkMe+lXNxBfk2aBQjwm8TWidwDxfER14xkUQIGA6y+gDE+9VXG9xt+7soQ7jkvgSq
ZMouCtWHNM6CZ3vj03ZBg3Ez0sFy/BDzhF3fwzB+ky5G9MCOWvdeYlw5WIZKn0ihIlWYzEm7/P2A
WhhJaFFT9xJjXjUt4F/QWvGmf47SkyUvMS4OPZ6SYMzUc1084yldJQEoDP+TerOR5Llb0VQWGpkm
zyvquAYtl/X5UK0w8aFcwd2rhQhfZAxuewsLouKIsmkC2owgy/3dplPsrgWL9Nn3Uon12Ftw/JbR
tPnmspuGA9jjpXFhdhkTe0zQ6Rt9PuPFZEETKki9OxhWIK7fqsu3EEB+gB6BmmvyuXvYGu3xxLoQ
G3hk0UKmxlMxQJK1LShmvpVAuiw5fzeTMztkH4WbwDMamDDzsKj8XLsTEV96kKaeiOBmncfWl5wh
CQJHt42QgbPLrL7oBUPmEQxESyjPS1R/7khGW9cAwy0RQKedwOB0ckJbSGxOlCxO1/Vq1WytS3Bs
xjOLj1POVK6Y/aDJY6GSH4TSdWcuoBRIt8dRF2WhLh+LcnL0L0uxtA5ynVJ9aup22zIFfUMMY3h9
Z/fC35IbpSCaYGiwfSrOLUpXQnDPyibvPP20+44gu6R+01hJL6A5cVFT5772v1d+UPifKkgDOSax
JQ9uJk3vdh4nMi+eXSHxtskXd+OwaT6+ZozNedNseASLrhvgtRPlwK2tIACUp+vk40sThLnyG29z
x1+aErMT9ozd9APHWz/J2jJJdEKcpbSRdgfZ/a6UqxIuXxPHN5HNLw+9b6pWFcFmrh8snX3J6jwo
u41QdTWeGJpdOr3quAhH3hjOpEdVtoOhw17mPdYk14PLIotI6hPelJCGKqoJ7RPRGV1P1RCcVYZS
Rqxe0pKR/kfHaqRGHW8dt/2Vm3DQ8bd4vtHk7J1F+wpkGSPEPL2Q7SybL1j0rhNMo8OaxipkMsow
kJUgxQrf9GMtxa+BUYLuPJWeNyhGnDKeXHjimycwYiZZxhCt0VF//ceyMDUE5JsrzY9f8x6mJZbz
smJ9oqaM4gPYqhaFjrJ7a62TsbaAAPzqie3RPoMJIvNSdmQ82+Jo+P+Vvi3wjm96Hw1qYEnfnPAm
frC3mYvew9C0VWq96yhl9cOB2wqhH4IvLo8O2HNUcFpitADASC5osAmT0IkYCoQdW+I0nmJPa8kb
NZ7dV3DSmcryl7BgZ9HeUhWGxMLmod08wfxc8Jb0Dkl1qGby6Z0fHw7x2RsJ7Jzadg4P7uri+MSN
MDKOaTKa5xRzdlxNOZ8+zZ34QsttqKeujRetOq841Q1tQN3eKidh3uBpEr/AVQ30K+MsMP8MFMYM
TBjXWocRtv8HKc6rZWa5f17ZysIYXFL7+z8de2WmKfnN94abXpE+0RNoNRIwTyHHAELzTmx0iBtV
IC7r5e65Eg7p8EpzOfSV1/L/yec7WMNj36IpgDxttYlEubdn1YCHeRt5FPgA0X/fmxDRtCgSJc+A
ugsDF1+bsv+kHptSYNQ7ayjGwHqViozcMrTZS7sYo18IY9fUxFQA4G8NTMfz1Gufuj1DlI78byHM
opWMVnad04rL6H+reLnnSwdUoFp/Z2X3zXZe/u+JbhOZg9RHFlry6v4ZAss5yRUjVTTWW5eWJNdf
Vuez8Q1EAnmpx1L3hrk4yj6Z0EYQ+Kp2G5cgP7mRh73Oi4DZKbhVKTcepTejlNJX2I0p18kdNWJV
MJ348Nt01Y4vBKMUKT3CkRFwaRQK7KvjvcFkm1QuSn6+0g9JRaJVbm9J+ERbjVXoh0enQEuRbGr2
NMolkugcJCDFue9Gtm3sM9120r3SdmlAeBl0L4EvUO2tAxZ2/lOUcGA9mGzoTLy65dfbXt9mHARP
USxTlHlRJu5k+sOxI9jSIGa46z81L2/fbn5u5ntlqSExIl7VszsPEbhNWMPcwJISOM+eBl8Qv6mL
Cky8GBZObdBYVbOgHjBbzQ3c4t1pdlLZxJ6P8h9HQN/pnh9FdFIu1DzqtC53EuJPiMj5sE6efPmZ
K9813fJ/xDM39AM7/V4pTdgRepPgQj/oQVbBY3Zhj41DBPVSvB7AipLCN476tX9k7uaOABC4SW9d
ah9/vyrBD9SjmMeXCqfi40jfqb6UoaDbRBUpNRQ6Qexa4uwWBUNZ9n/Q/K16I6011Pe0ui7cDwJp
6uXAEdOgnErFyAs4s6+doNUrbDWKJyvkRHlNnorx72fANV466O6v1oRpA8NKjCjdQ4kdgCe98hAU
ip2Wu9PmIZeNyfSseSNBq8zRRmtgQaQ+hN2+4l7+AF0HLxbCOtPalowdbEcEr2i4ssaBohZPO8j+
tqe5bbjWojdQcNWg6vHmXU7AtAKu9iunEs0C5m+4k+7MaUJ40rVpjSESD6ha+QoGAOle+Gko4808
Jrcat9zApGSCZMDYmvLIgwYYnQaVkbAtQjgIHtTk+rqR/cmHhMq9LWlB6Ijtyyvc7llYpv+naODp
BpgTwKriyJqxdg7lZI/OnVZRgrxYp6vQy/YBYB1yCZ/gmTbtc82jkNB72yTwmW2DYIJd/7wACHaP
/K7lNehX3pu7n6E1qRDyyTz3cqTovsj3wpII9tOqRC1P6CuIEd8My1vwJqyq/pog7Ryx6KKEcc9b
XHFzaFZ0dfKi1IB/HHm1tZ9fYDEcYn9tOQOddx5qaCqljgrzc10QH08WQCzUjnSDxrEQX7ryQ/Nq
T1IORu3BlXDL/pMnJAExuP4Is0Tot8ceQJzUNJwfNULnmgm2NrH9/qEmI7WzULJ/rHzFXboY40JC
fRRC8BRVaUHy1rakvICUZko4+2gpGV3JbTTCO+CoStr83w1/9tClQoZCKoRPAa1KfkgQxNiJaRbQ
kGh03FaTcOl4zNUxVIa9oaZAG+JgXNeXee6UedLxj0C2jJTx9GIQEQ+WMdcQCLMRpHOtBckiCwG8
sGdh/BPyygVgntqNGulCipSo9JKBwG5juH2HrLgJfwCNR2hNIdJspCMM00EpYp2eL8uSxZZmhp04
NG2Q4YAqowRYmFFEqub/RlO6NMvlOf6jau15yVViLV/nqh91wufrBit2Q/a9gShs1zlDc2GcrzDK
NH0TeFkQu1YXsVDa3jWEUnIQgDCl3ZZ6rzEY5SLozitNgK3i1xSuv+H+PUtN79Hy1NtuJrQVYzwr
y8WP7GYwqr3gm/ELaGj6Ur3QnqwxLQXVyTXrdCl+2oWFfqoWRXIyZVSkTobXaldWuHCHP2NAeIw+
YLCG36PtSof6CkmKAnSBoNqsCpeUgwbiD+UjetG/imJLHBCZU2xTRZVqzVYdtuSiB+ZGLUWlKBGa
9RXCpGN054/v7UBMPqA6JiyKIfCJoJC2uoOCVy2e+eZcNeuvYgrGGr1t75XJpzASq8NA4XVlt4R4
pGOxRDN/Izh+kta0JWJ/y+4cmUIbE2qXAxHKQ8mk2iPAVLugEB+npHfEkKyCy9aIWwXhWHUQEs8l
+zjxOsaBFWWnImFNStCrhddIf5j32TrtIYgGsGkRFqrvWarflRnZ2TODkhZ+UKafXm4UkTmTW8PZ
aQvKVbVpayNYWvXjprRXxlsrZLTFZCuOccyXCG7tMex4yqArie88M7Sno3JzGRkyDZdbJVTALkLY
kqq/VIVB9F/Z5evZiLaKQ8+U67gy6i45RZHx6zlPnRp46P+VJLCGoMG9tiHGo4O4qbrJj8hGnW1V
l9rnmvdJSzIYQ5ZVr/14DFdGWowOLkksQ4ghMAc+RcMuGjV9Ic7ZmXaNaXy8xM4gq4Bu3UKIqHYb
hQ5x069S1Q/+X81qlq6zBhcmopJxA88+d7Ml7sX7etzzF6x89JEtITuZo+adtHPNEMkn1Q69piyC
sGTUBLgE6Cu/LSh5sfh3nqt1wPVURWPRALeLT2sG6TN1QT8NR3crhpGFLRJmJHEQL0pdFF9PoHq5
QHfa+KyhKyeKT1c5AIWVT1sDh9z5b9L26ZecRvU5Q7IzXALHyU+V/AOcqUnfIL4YnCIhqE1vKywS
JkOsXrvR1c21J6r7N9KF1f1eOq3C9y4zm/l1SBWV5uFR+7v2SQws96KHcj0eXCFDwE3BeJtHcEJs
Bi/QX7fb1i7IpiR59B/wBHOvzXCJWtyHNYIdfRS+lponSc9B8JU3NgEat6udx07PhqkOWDzwYxv+
d7d4JyeSjTcXy0Qz2xVnKG8/WOQXmm1pXPTREXUDSO9mAtb28PtJz1r6nS83cqZjc+NahKfaRmYW
nSJGmMT5xaUnVFvyj/FDEXWEwBui0Ew3BkI64X9hbHvQKbKKh9C/UgAZDlK0HPbcjO9MdkWyrFBH
w/68NkSDkBF/oKqm8PXDQXvmdbLTLKxnV5VYRBphTCVKts5j83lheLCutkCRyOXaR7JehYL7mxAx
ISWY0Au7QGA1fGdzSQjiozwSLLriKoK010vx+EmKX4G1OuEvo7vEuyB287VEWjBn9CU6VbASR45F
54N/Jd2/+TIsVEo8obJm1cwSjJkjhF8EpZiYS0wV8MM1XyFqxViPU7MEo8aaqh2xEN/VIMp1ava2
ezkLHLxLdLGmiWPX8k2QvWzKSqTS++AZEqjTUMdfdwNH74376EuaWz5JpCDlnXsPtX3zEaJKFm2y
D1UgfT/DhoS04epu0pZgjEQogdNCvykOcbj3+HOaxk81tf3BQMwG/EKnp4ck1IhiyDAggbs9j6EP
mpvI5ffJXJL+DKjIGF3IJseyIu8bauntLNc9rUkZMmEvDZokj+a3qMvzcVvHsplF/LNRLbQz6eCm
+vgy8K8c9vTgQTG+onCLiDWVxTKE+PIJp5/FLRWlWdr71Q8Ff9Q0ZVqPHOsdLtbl1ZT8O+pC5wM7
1U8chwy8zlR6YnM7ERbYBNtjrCgMAqjYDmLlm8xFePd6J+1eyQctIwfc1SeiBOTafWLklSve5OAH
gCWFdN/eTQ46MPFKtJsd/ijigmXyDV/5kMytiW/+TDcPaD8IoSo4HQq6AgbfK2Qtl7T+S4hCAdhr
LlZZb408V8L8/XLFIDq/Jetlwf5dL/RH0pE7DLz8a3buENFo6PanxbYI9uxDa0y91wjAL+AwgxQN
Ms7srTBqCrWraKIMA1UYQoJphbUgpQV6wg83h4ftdaQjea6Pc+rLlsFlxwTDUjd9aFBMTOKHtV1z
eASBcwXYMOXUmW0B4UwNKbOM4Wt/yBftp4cKD95ojEGhBGdoZpqvW+SHFbhAs1wSrTNlvB1E7PxM
9EHMuqUt9va/2Gaxa23lgQ9VLs3Dri+dkHC4dm4Qa1hBdczgx32laIgF2FIo5vf15lMzQ8J5bOHW
VTxTnzxJ4COdLNswRyxHz+5s8rcRfmaBlYwDtAD2ukE74S+l6Ym6jF/awvlTHqaktsWpWC3byh+w
gIXCBLtP9OJnlGTriGnFarbIYI5rAgdrg9DczzBLKlYPPagNHWNftuYq2LbsMSniZfNTFnkF3JiV
om5O3/JsZDLiVnl8qtUsU07iyd9yTujGFZCmXH+MXSQz7xfQyVEVKVmcHnFYoKHynt7pdvw/tn08
rbIjzzE0NiVuwhrcKBLY92i3j+UEYXe+z8NAU66Xg8CGdD5k62hVNLxBKM5/tQqPHoj0GT4D19D7
o/bhavW2Zt+UsN0i26m6RSeX2roOzmW9d+hfS/DQQMP1DrrJNj6vPpeeWb0EspYR8y2fB3BoRMUh
JnkYY1nJ11bBM0zNzDYUeL4sYh+l1mO4GGbU3C86kVnGfu0hkikIVkShUq0ctTd5IpVZWtHW4HP2
4Z8REBund0t5a28aOFIxP0F37T2VoYtcgqgf368/YNhNAqlFv9RCSWoKCL8ddPD5x5vTZZg//6M2
ISvgyOYW1ozCICKtuHOKaYEFP1aDlZdyZYnjSWEaNh7sf2+wvkK3hxSnZqXO8eaRDRxUU09hrQM4
yKCi4vGXt7n64m2C5w6m9KDMXVu60C88i9WubRtGzDCjtNGgPnG5mjylN0CG7g08Z+D5FySjMaMe
mDJlaNd94lY3abddgoDnETpJYT2N52kDejwWFU7CxRMEt8ztIw5JCnNlrUzwfpApigJymroSrcgj
F6F2+T2pHzUEmdKuwvQJuDFxFF5uLLaOqEhVCRMoJzOHqxjXaOnCzVyMVJrEWcJ0Dsi9Jh3kGSSd
kC98INZT3zrQlxiisk8nGKbzuTGzl3HxN79bKyhTDXf9BF4OXXYcrzSkhfniRbARfr3zTb+7kDGC
xdf09hR3/H+GCZiA05K7JEGn7DHvSrxDql9H9qu6g//BorsQipr+JlaQ2JMbmJdPD/3E/VXkvfJx
inAVPagLczRA1cj47NG4j7Hv/GVDIR5nNO6VrzdUYUBmuXpD/nGXfZPE/rO61405NTnHpWskDp6P
5PT2YdKJZSA9dVO04Eu2gZDdi8kkOwBwKBaMwnH84NA4NIr+izxh38fSPyR5yw0NPtm0ucB5eeAY
CsXO1aVQi7qtLupsygvgaHtQHMiBkJvidJC2afMVfMnl/tJrusMuETL/9khOASYdaMsbuxTBjg3v
duN7JhihRCk7qghZ/OJGdbEY4p1tteuC3spNAF/PMBRQgnTO0x0RjEDCXuDBNosnADFmjc16IP0p
JIcLJ/DP132EeyiTRm1nlqVyWTIKdaeX2vA0F03MUWIUSmxn99aSrHLbDLd/kr9GMePpE1+kithK
PRqaxQ19I3evkqaAU+9dts0CI9Lhn04Bpcv0yuX3jyHEcCPFKCAg6PdRPEW46Lh+PhIXitEH5RMj
ulebM73t0ifeBimPceZfoi1z54R+Ng826GeVcvnXJR43QFuaPj3qV93bIR0SWWKAXtARBACu+rb8
9gkSElm/yA3TDFPs/jRxvXInQZYbcUib0YSUb8qLtD74N0iruUtKg7XwF/KbR2O/dyHTtmPP+0tz
34p8Ca+vRa39/OkN3dkAa3tHtvy92Gm9PBtZ5Mo4aiPsgqUAENY/PdHheSRFqDbrKc0rcfNeYFrf
3L7KIR+oUOPnNJutf8zpGZ6qQRqZV2z3g/5U0L9WtmBvtxLwlZTtxFEkdwFaE06nb3udMKqj7wOF
vX7bU+WH2i8iFjEg56I25l0BjEsCFLy+UBWZD+aiOKqrYxzRSFnJroStS7gUXCJi0Td2P48PpLLe
1Pk1bKy0L5EsPuDT0HLIrOCFRYgZhpKDMcIiNIZvQtY/zJW6pHbKHfnuPG2Ky9e6sxDKCiEfLWPV
hlzLwgMBMTZipJLTaA10I6Oit11xju5wGI2nl/jUV0Jdig54HvLbjdhGHt0U66NGjz5lh38dst1N
g3tP0pBcJx6Qd7dFIERO70MY/TxIZhfbFa/+OlFpCU1dk2J6kKne9tKOMrOIJcseb8TOvJkSW5Ha
aYq8pEiwnwIfFXe5VZunCtRWY0uBKXe9gu/YnVLeCPyRR0xI1DYQ8N0oCww45fXtLqp6DI/KhY0e
QaiZE4x/8vsvaY6AY7xLuwmRO6JXVKtxudA8nGlYSutxLPDAIR6QuEIOd+4U5krqG2bI0OkJXZQt
xoVtSOz5Pxhc2VsbBxfpIaF4SvwBQvPyMAHNGJqUdI0pOqQBsnZbQGp43Su+nGD0fGH/MEm2gfE9
O3fGKvzmdjaOIlY5uDWFYpT24gOvYPvAUsnSXporX/TmTSLrJBsMyXnNqKfLIRhHUGngBgG8H/Gg
GebkRg9yDrowf6945OSISaPxKTBdP08pEk2b8xG9gDbOBK7DoQz3u0CB4OispG8TS8Oe7buxvkmz
WM3F40OD6ZpShG48HHujrIp1bKwZOWTmhkwRtV5w4uHcHN3RcaA/xNE9BoX8gTUhBXSCxX8r/+ix
8HGJmi03CqgvAQeeSjrT5+JAdzCmnUb7kYdCANQBESykvKWbGtsDq6/Q2i19+/45QwepHA5hASxp
vHbuZAa9AOT1EBJNPLpY1Xgob3xumFJ4uS8cZ66C8M3vkJcPHa/W6iOO1z5Y98kGIhJK4xWFaHIO
8UKjPpBMm4tGNLUwvwETWL7ONK6GzEgYGTrTCTgJXl6YUr73DVZfE2fks/BebStluOKSFr3Q6V2S
Q3D8dKUzHQQ/pJTf1UmkJFOhrryJLtSMaR82U6mh21R7+efZf/fZIeAPV00pt/jwGC+vQQvgJBem
EyERGJGnqchAxfRS+9MoDe00Wc/t5ZolhvESAcNaB51H+bvF3kwAx71cqPDNrhObfKvboz/d7lpB
Cl03JXEbWODdWIL+lYC1CA/Lmtqucfxq59bgxmCwsAGrmsNlLF+0HwXOb6duw7we+sEuUDNyu5rm
new4AedU+9BOFQKs8EI1vgijZOr4YYTjb7lrhSSvmFuXImEinHeqDn0k4w1gX3sjBDzhcVcjlSAb
oBmlt9YNIwsdAZ2t2ZrrxFf7lNXPCBVFI5+ci63XsrB8SGvs9QLzlZUWJAOBKSBbFJILJKTMp6RG
eg8JJPkbmZd/UcpPovaGL406QKevXSf0CAwbqdMTiZv6A4Hlg1T8AgPnE7YkjL/bVuBF6cLx/iZB
3SK72TKaEu5J/3s0p4+xU88tNkLACH717ViNP7r8cP/9GTxq7sffIe+E4BmPnaRdo7JWX33PS133
IJXdlBMhMi/DmJOoMw8NykNSJrXwEY/EDn5ILF/VKu+AO7OTJMTIPwHjSsyjzX/9M0pf2wgH0nOY
89kAFS0APn4IrJnVb9exjUfpcCG2QJKQ/Zkd3zWZ8RgYYC9epkpBWrluJTTxuMUKsaUhQOse9eCZ
/mnd47dJyteHDFQXxpUiQRowlgkDCDBKpTZzu+nkGYERZ6xt7ZjUXcW8ZReVkkLs8o61CNp7Jql6
q1B0vaM+WUQh0g3aFah8UQ0r08DfvNgzr57nwvYXexL8ws5RNbaYDnu4AiM56ibPOLuPCSAyJ5eX
KSHQNy6/QHJ4NqGKqCC6LtIVQ3Ae9XI1E0i2T+iFgM8b81TgQZuF5LNBnbGauzCCydt/taGpknHI
cc7g9R8x/YxLjVjOgA4ERHO+ZuuDymiTBvla+Z8mpyySEmiGQZIjb8x8mQPfE+2eQ5WEbmWv4GqU
PHY2EfAam5p5ujLFdShAuGgMi4kIRgI0b60wBF3QkBWQ/7tuptlabve3mO/UAfAcrFlxqnWAPnXL
a7bGgea8wNjMlTj9Mg2qx2wW4gEuHqAzkwqIkSYdvSDI1uH5fVTn3NgnyqjEC5Ix/nOPQFyhWP1v
n7CC5JwZFSfsP62DiwhGqFGNY53j7L1fi8FBkbs82QD17EJ2LeVCUT6OEERt/0FHQZX8m4V+xILM
3qigYamAIzo9VoTbi4kuGeRSyMIJXIly6CuCV/h/95VmFcVfjOBMrmY05z4BVTUd46N8xZH7RZF7
aysH41+jRrgXCjg1VTbPdcioMI7FE/5+Ju0Qa9SbZl95CXGQAeUqAQvZjQDCW7P0Il+O+3LevET4
wGSS4IPWoGADccAs23GF/Qtq2DTis3Z3/YsP6PCsbJm2BgrmWRLVURQUmVYCt7YY8U761URXOX4U
vxfk0IhAS8RWLd2em1eBDnuYXhZWkrXjAIbzUOXdY7XGUL/kpzNGhjw28N6bO+xkeGhZAETyNY2U
MMavEimKQ+OWY5lXqH7ApsyKi8z2CTPG5Td7UQUjYZN2ZfyHetDK7bU+X02QmzJkBsn3NWW1+Wyu
oJA9q+J02aaI6MKvRnPYnyFUld4y5HORSVXvqiQv0eoNxsc/LT3+LyokVQJoUhSHuNi6HjA67lVc
zjxpLDuc//jgMsdzflkTj0Q+i8UVETo7lXo4MsNqlQdJu/1gGhTEXWZyROjzAkvM2cFjhgv1t4Xi
/7mFqhS+O9u0pIQnmo0shrojItoq7bbW9zTUqnCOw0QwhPuG81pIHcHy0Eofu/YfTwe+HnMefmIM
vUX+M9oZXAHd1eBkfKJ4C9p3NdXiHzJ0W8FemXzFAa+FOz8VTggnLAtFxTtbhZ5a+ivGAC5rK9op
CNzquuWvYmld1JpOef+vVT6cYsR6VsNjHfDR48v+ZyBqd00BfxBgBpgxiYSv/UTOiMsJYargMFa0
TL6bFxzGrNWVcZr44wb9iZ2rCLDm+IQZZcf33LraA5quHH+8cavOhfDLjPGyh9O6+ZtKHt9tEUvr
C/p88SxNYQe4Qio2jc0tGkRS0/MVIvmR+eCIEhSh5/OFp+LNix+ctINV0E9er0H4R/tcDpm0GfHT
bPGKv4xabOgea73O+cmzmi9OAeXcbbr1chLK7YKEzYveT8jXLG0CTbnpCzo54bqwFiWFRaDPae+o
uNtL/+Ipnv+M0i+Q8i8ikJmdQz8+PGhSFJphZ6Vc42ekObAwKBZmKe5CnaiipgQn5E8fylO3dRa5
XvBPz1YY9GACvGs7obeqhSthbkIoyIeFtvIk2A/1R2wFuRube8mMTzi+iAb04Swzathfzv0cpQ63
L7Gp3BEt/dXuctxVgPks34N8Vpz+JOSxtgXrAdJvQpkcwxhC1ZdR2emBX8mNDgeVWHx+rAvxo9v1
GK9o2m5KxvGl6xX+3ShSC/ChHmSTRwVvjoC3cIivoXX74jL3ierxrUF9UDqxEEl1xrp5ga8o+okp
ZW7Flo8hl2F4on7kl3AOixoOqdBBtTcwy22LEf1ysivhDSf3HLtp8AViM29HZu4ssUvKuYG9QA6t
oBBUl+/w2NP/plTyaEXDoV2LAY9LIaHAP7M5Iy5ytBZEQBi5N2m2yOSIUhaVWIqf5JyW1ryLXtGF
djL846CmdDB5m0Rz6P3YoyuqdlRBTfIiiM0HPjat1AguhSETJcNk9MxNdELUhOBKZJcOn8P8xE5U
wQFgbGvCnFN2rZosbqN9+taVOviVeDfdpOXClUBE8aGBib2jO5GpTaVmMd07MqupapTRrziNg7Oj
XDmiOiRPjZrJIKQ31RaByKrWxlDU02+GL3WWBgIKqYoVQ048DAyT07f7SEC+umUtcikLJUwGfGLE
X3Q7xaJrZPYWh1PdXUmfV9R+KKaCiQAtQwrma1HjPfKnVlk4nFVm+6PfZy4kQjkm1hBd6Ij6uv0w
5OhU4PvC4SwMz4F5KEBHSgDgXe5UYmTceHCjewMlaAU9NC8S0jUOdaF34JN3SqthfUE9VgZBWtKk
5MC7E4ee/cd5/AktK4mtj2BI1e+Aq0wpCzQtceiP2u2j5MH/2JpQHsdW1SNZjH8foZibfIBMCO7V
dmEYAkkfS9Om2fCAEooc39d/Psn9JY2nl725UtUa/Co8YriOoThAEbeO8tg6WVflx/muS30uhRk5
3ELPzmTWbXAprWeJVoLLoBcdJ4sJcxchUc1lYwTu5S5M04QBOh3QpWvk5URUeKGpzpxVqtIDzI9g
pWojl4A3n/cm/6XYHrDz/Eqh6DWK0CDz6J78Cn8VNdmH7XTjbnDLghK4ooo71zOYkL1du7+w5S90
hmsdgXWElfFD/fA5kfIn+sbkvaS/po0A0lcl0RAF/XJrAZtYq+5fe6crRbazHBRpNSXtIPs30cFr
guwtJD0yczh7DCD2Ajl0N4L6YeChEKyy9VDh+mWJ/oSV5R8yfrX9x4n1+bVtErgyXBZZxclO9gaR
B/kayrap4cZ0EvIf80vBBwCc37m+sml1B9/5o98Wp82HSKC8IrNB5ijbamAyxPLwBnG7sbxI6c36
8VvJHy+zvYoe0JVMeIuqRMLTFEHuj1H3iq4yBuAAv2e5GpzuviH68ZPi5bcvOZiKRb7QsVB7Ql1Y
BQN5ZdjhXaMPvqrWxp/6om7cQUINaTR51eBa0g42LvE3HBLEbC4vdEr6hvWeP+yYh6YtYLCL2OjZ
19oI/LBB021Qns8OYmevgWLKo7V7IWpw88h2HA934SYLvWLYxkEPLP2wA9qPL3H2s3lJ9bKjLxAP
ph+aWOPzyZCaiVpZtpoR9pu3wcTyE713HLABAcBKvU+Lf8Ho9LLr/LXLjOWCtbO7au29FP8XmeGH
npVoRaqDKGSrJIh62BFseZv+XhCZrXtifAytnzrMkN6rtwniwPh9SEEyPcZTNQHejM39/PtfwjKO
C1IT9avNg3vcZzXSuQ7MIZv9rSjzPbfEYMjtoq+nhirw7x+zuQBYdmsCdqgYwGlEYO2+VJ8zNJTw
0jQ8k0u1IrDfiC5FRAJYxxCsCZbmDUnm6b8/bwZcFPfCt1msjRhGRKuVfKYrgX44+LnPOMZfYsNk
thFw7fBC5z2KtnsGMhqQiXo4NVwZ4PX0BYKh6kd4ciww8cbOudtBqZkf/QojbVAF/tTZogoL/fo9
NS0/eOS/PwJhvEOlNCR5WyYAKgalJm1ZYSYNv+6kWDK8nZW+P2Qb3pCVAGYxRyVNHiT0DLUBNfu9
TrsdOplNTqTnias9KqL13abqrvlDf+/0K0gGpO/5YHnLosM0d2zKgtrgSq2RYVCvwlglGrq/ycLH
O8eb3KgKTMOLk8f0as5n4JsMW5gmqmpHdXHZRosuzE5xWO3iYnvrwRocuvYTC0Wpp0sw+jGwYQGE
0wmQKA87scv0yhGd3Vy51Xo7MDgzgJLvrykvj3AFqkbFqNiClEdPn5iMjXFoJ4rnE5uth4LYkMbx
8yaoS6GgZ60vL4oJPXTN45eE2vdLLOYNz0HcSRUNTd5hSrxO0ORK2nzmRykeeqF+Q6kb3RF3x3nW
H6BqlPP1pXc8ImPechFTMfaAAtWNgXcEp99mBhbPThYyBoG7hRS/YyePP5oAckXElWHZvXUYZLuV
Joc8DzEvLP3wifnc36N/nVTg/X81nfpBSVNwb75LLTkxa4LU3Bp4yF8Y/tyVPJwiyOpxEXCmUXuI
Pnwqbq6Re7BbLinAGVmX+OPNdcTc9rnXMkomLT/YEi+lERJczWyrJKv/cnvnV2x+UjEURS6OaNt4
eAx8vvbeRQ6pwjA+94WWn/scYkVPfNZM6DOwSWCrsa2nAmN78Kl12tzJsxN4AEdfDEh/k3yTepek
OVf+HGbZnt+kKGNemZ4QZGz9jxLyY7ui+1kaKxWtfiW8ZvSMymBcPxgHrerAopou9KxvPTxcmhus
p2G/w0bDXRD/f1d7GjuGhaegFrY1JA6yZS2rZHL+cYcVNaVgzAWfWfft31QdoJssKa+xI8SxuAcV
9JFVMGro56e7Ho98dpCg3gJCKBnpb0LF4PoWrskUNcpjrj9Hql1jrAk+SAHxR15ugRsfKd+mDc6p
wHMPqgJy6wo8qUQnEgab3Hs+mVnb6u+cgAR1W3PTGQP/uT1/g2cx8UNVnACf2210CkFGOxEOsYOP
IHmk+GryvQpWnV3qkBthMDmQVHrVjn7OB59Ya1Sc8AUHWkg5kjS6H/eX7wWXFrvn92tNpBbPBKiM
vlD3wPhJl19/0Mol4SaINo7W2ON4Vb08nL8YbfUHJuQVhJE/SNc+imHXKzr57nfvV+Qm2mn5VvkW
BnwtT6+a0Ej+nES8NGkk8izHUj21V5oXBacBWErSn2Wdp8mEAxwjcz8yYSshJ9pAwJ5jeiuE1D2H
ICqqGwvbn83fZRk2urlDoDHIDX3z8taNrs4Xdu4Z90f1UlbjPl4ePJhfl8aydJTHSOZyebG7wS5v
aY31mCHC0Zs/nr5dpTXNE6rpfkVIspgzX9GJ7yZoY8TNHFCdoH5eR/Se2xigjFKELIaw4jXCXxDP
JoqRaYGDyk/UpNkiKgDuVDjMGM+P/XgBFgYfmhm+8kfJhKNXTXSo/F8RlvMF7VyZRMcUT7N6O8yA
rUGKXlTrUfbN6Sq6NjmMRSdIy7Xy78n4BxdUcCpwEc+4NgDWefhu2tbKHoeckiMNtQHqTMcA5N+f
Wy1ozjg2mN5BFnDQSoj9uI/k61vW09ctx992LWUEOC91eve0DUtYiADlw9kXdnXXw4fcG2bDPsIG
XlnBzRwgp0b5eqaxqqQxE1gpilUtleeAzxKbPp56qAjGtUzQ2sASodjr2qEytfKL29T0Czr35P7i
ibFqN4MES6Ed2+BbIHY8VjhI9afH1AIJdj2TPY3aQaHXLtSMhHxnf6lf+gNbPe+6A5j9B6+jj2Xh
lyxKjRJpAjxdXUUHU7EZkS/dH7Sfz/7l8sxDkkgjvS+Topcgz27ViTY/iojhbGYsMWYNtPHiOWTa
X4gt7e74ERmaJHia52APsA9Nr/W069GrM8rqHiBVsNXmubgE/axs68NEtr4tIEM08VJleOkEbpgu
MEv+XbC3VOcDYla9KoWW1G1WrPY0pAuEhuvZToV15rGmi0jl25oFl7xfjzy875v1bp4WjSR/WdL5
trBRtVXSlG35TWKAE+gy0JA1Uo6zkpgvt6vvtwDKm51/D6Cah8/1PT4GMB07nQ66DcA3L3gh6zmv
+XDC/bL4NXf22o8qmuAU6gvHX7DRtTFZkr4gF7FurgQtkZgtgNNIvGqkT+J2qV1KzRnZ0abg011R
ckGZlkKKaXFZ4docoqJPji7LsGDpLb2Y7+ISapHPIjH/BpZKrgg7mDOLOUENg78ZCr1f3TqRgQxL
adDUzHNj1Ku43GDTkj+JO+l4LCTxsBQNoRiDMgRZ90LT5Xu8yjZJGcsAXC+Y9PpsN3SFXqckmazR
JixYkOknu58THW4qCEz2F0s309Bs8+pEMxE0QiAbDi9E9iv53pTtZC7/w6WascTRwYma/4da1ySX
5LWjR4MDZ7PjpsjKKTecNRqLX0xV+rg5NwavIhSF+LiC8f7SFcxNsVQi7ERZ0J4EgMUdr/VjvdPP
U6yvUAx/SNsupoysPu3E9uNmeHr09fzGqhoo05vFd27vvdIO+3U1t7J7CjUbxNPT66pZw/4fGV4v
FxdtY0fbNIU11k26uEwXn1+CceuRnr0QX2a2EpPrxxv9mkA6z71piJpZK+MKADJnRaTh/jQ2FoT1
OCyjbOQQYJW8G8Jd+JNgPAS6/8v+0EtZOICHNJV64HSqY26zoZaEc8h8MYNX7MRkN7H1yijSWkGV
lHRFDkChTCmdzmIO0YhDhINEpdcGXjhgpaTYyl/pFM6gCSMFHs5MjawlD+jmxCwLZI5AKT+H5joU
ZTA199YoySSt6McNz2bAafHpL60wDXLyuGG9lALI0jumzP6rZeThRqXEXsiHdTdCeAZsOcLXbrdf
brf/lr9/mGqhcLMQUPxvpMkesYKFk6ScBPhl35X0XtLcK8OnRPcXIDF3e0cVKhe1K3aVmPNsnvGe
g+0G3QO4FINpBY9Z+O6eVo8GfaXm0kvEnUnd0EoNI2yPJuYc6SaHNzeGRycOGXu9jFK2yIczwrqH
Wwy7bMnF2edSCYd/UtqxX1Ta9dVCd9DV2YQaktPd28+CA5liISrFpoCjNCSRSy7AMF29xIYYYb+j
fYa2nvZqHH8U6dzZZdIZFVvOlpGZv/Wj3cEYxSRVEuwldfkK1Ppv0jWAXNkkr8pkeKb4RuuVvtlI
lTnHfX/zKEdn3jj1y3hFpun6O6d28zFOaj0GXiJx9YFns/OCkSHQHXdldplcjrRJCvfVjJyCuozm
YSgWycF3lSakzV473bgIhgPHGA1LMNImK3hY1c636eCc+Z+00yaIyD+Qnb9PzFNgH5iw1FJQefsD
g7nZe9rKSrUZwWKBSTS33B/nomHWzAGf6Hmj9DL4KYhgdpqZ+6SyuxMR3fRTDoYsbOVshDpSJSKt
jVaj4q0mn7adNjHFE8dRrfKaf09o9c/1owc/dLgv0W9TLJ1L32cikO9HxQIP90yXDhBOOG0rCCYg
eX4B273bEozqZRz8rMxxNofhptJCXjLGuUkutcEsfZWH6MAoOhc7hDjOL+m7qK4u3lxOKARwOSFU
Bv/GfY34kCASItTHReL23oAm+GHJ/5hWbWdpRIzbh6MX+bzpKTV2+C3ys6UjxQTUkc77gzLq4SQV
kDKQYIRAK0RFc1ZPHWRFZ7P26p4JB6Ri1/KYo6/pGIfPUfGo/Qas68dbjr+POlQwLEyp4hvG2uRs
0LNHKIAeFy0sy0aCa/oDXFIjExCqBQrdasdW8QjlXk9Or5xjb7ixKHDB42Slr0KRjBL/qmZzlkLQ
dxwC/wWK4U5PVrG3t1JmCR2pMYXqge0Q0P15C0B5jDr6c+u/B5e1wCjCku9hxAq017MBl3ha2EQr
0CdXs7sXARxfu/cwsElB/i31oVpYLGjZq2i5Ws0TABomgdm6iVQbRWDkvpahKtxOeVdVJxxD4H4A
VhiwlzG3/3oy6/ibhTrhFgmyMhdexpbtE/0vf5gmTshOB4C2HyDA18n/BSPYGPxrcmsdW4PX4ALb
ArDfD+P+SV1690saJum/roYvVHmS8BuGUNkLBOGM4MGGXbYI4rCGK6SCVp4rWBq4NOeK+mZEts8c
lSLz67f5Ye2HM7GPZn0ZPcMJrngEf2dh32q720g7vSGJz8rXx8/Zi5KskJnPOBzuhnzGtPG7PhGh
LLKPC6lPrcaTQwufSkm0Aag2RAgM68Qn3pMIQ0/usFCc4q0ZEBLy9d7R/dhQ77FRtCUm2hqBotSk
6XS9OhyuKEjGa8xnnnBjuxZ+gxI3EJNdbUU1UCA5zbmxwPxqfbIEXyo0oyfS65twuptX8DeCjJIr
5kPxZe9g6jH7XirSWh8lG93UBAKUIXdzXjhu1Q0TXJtskQQ7UMi4G/jYLkaQ+X9wjHxv1fCBkwou
xJj4IkpRfdBJG6A345R5RnPV3pAoETTJVfluOQxZ9GPgljaQpZ1LZ1oyqbZobiyDcj6oH4QMtE3D
TGy5IN9lsooYgCDnM9SNhlpolZmn+5gj9IcuthzRnuOBUtW2sZHia+33lT6lJsJHPqNx7ldN4zH/
1nLPWzfGc+1FUPIvx4DPfhKDjl1IfFgJUlhRfwmPdpHdEEDrSiLpghVEE7AsT65liiHeVJCVu6y7
Hi90zuDPTSeZGSxgvOEoDib4LTDkxvJDPuIZU+DZY+/9n7kj+o7HDZ6cWfLiBrS90Zi1mg44SvW8
+abrbzIQZSVqUpAhaEbiZwaB/u0jaoIyVitLOzBNllFlOzmYEQPaTvKh4pd6TflZ8nsudi34KMe8
eTQmKZi24nIn/7xg3g6kWigBPecQ1Xhigja4+ylaieXMRbouUnuMNfp4B1eyuIChS4U6bA6Bce+k
atDv9pNYrNmIha9LMBr+TEG8LkzSRV1QfqstU0+RhK4NygVZ7/l8oEwUjyEd7iUjPdx3JeTr4Pdj
XdAcIXPhlUAGRb48PgrK2huzJH63Lb2BFo3RkxBq21V1cNJ7Rz+G2Kn4Ar+zEgsBhEb/svKhCdTB
uOPV5BqM+fUyjDtIbaw1hbnIuK3bZNEYTaqXmDwjhFtHx+YNToE+7xzfDPAuhSHr66xSEoXzMaRA
yo12U8Q+llc6t3RXfrl08DFimD67T3iFyMdjOdbsjhMH/nYOktzrT+pD57sJ6v26z+AQxKpPHsnc
XVbpIXthhA5zD7xyMFJ9I6mt1qCaZYNHzHKQMUIna13PByOuxtc2u9v2zhypyILctvDj6Kf0G1nG
6lc5hHe4tBidnMoQ42qpgAiZatsNZv1GXl88KK3vSofU/W1oRYImJIEudaB9j+jEPvS7hbAUm97M
vmdYJckDGRhXJw6tDt2G0CJxVG0LoFl7mWhdP7ZnmZMuVrniF7+1xHZmP0jrrGo1Ntf8jJ7+m4EN
7B9nlSqHl9PihmvJvalB8zMfZXv7DqafdecYWNFOW7Atm8xpF4/lSo+7B+wjA1gmxqME71GBT+ek
hD6DEZLUQIlLV38LiupYRcMpRBX/RAsGtLaebF88YwgP0/pVt8os7SJw37Sv7aY5yIfZaR1zpOeL
L4OvzYoTA6kzTPQgkz+7f+l5FZepnC6w0IplCRGYLH3xW/k8ymF4WBH8LA6r5Z44QxHUoJyZEjhl
2/GnwXPZ/0NEtOdyVptD0WokVBi4Me8/dhG4n/UOGBMz5s14ST8frlr/KoMiUT18B5B0N3j8fqSL
CJfxvFUvzpQofc6NeZ0Yv5/vGTTCe1jny8KoscZF6uvGVg8H5frILWQChqCMiFIk7KhGOk4rs7ZL
3hW437+dGpi0nQfLfbskzowQj7Q5v5IXXNIUQPPXwf4O6czmHfZn7/S9gOKwJ2yrCd1KwbcCYE+p
FlbonlzCvaoeB0LNlUQLhwNBKlCNqoi7aaXHinAzs8H/CHLd9SwZBpNJFjYrlybw+Hlx95RYKk1+
jcxPl/5fzScJ75VYpEiix3gMJbt0rVPRu1n3dmIfdFFSiBLBqzFT+eK6crTUO04jkSte2KUn7u6o
M3KYdlegjZCVK42jbDlzq5q+ykxSu7FP+KYS6epSLNlVmeguehESeZHWeYfgWoX/yCnMgM9ZrGt4
9c87LRKgBVgIWbhKHYcXiZVcAIdnrDtaQ4rkzLjhVk8c7EKLfA1Vw5THjwyp2oPWVBAILNuspP2L
92HhWBrGiIXYpeEAjGduphHcNCx7280zOa+BQXVXyjC8IRyoYGYWdw4ILc4XmOCS6+8Ias2lpWu0
PFHguUaiYA34+NurJRmygWXQF3a9XQgd/U7P4Pm06+oyHXljI6r94M/etE0dG7rFETUViN4XAkJY
GN2YyHVGX/VWNHZE/eFCbjAdXoCkaFsS/FKohQfFbMPNyQmjmVDFAMIeyEk+YqcxikbDrDTbfrWF
Loxi0rx+j7zPkJRnFf0uCM2KsxhVp6Ay5h6ZqJAfH8QP1pcMCQmZTqVLRxx76yx2VOE28/T8vzVV
sPwaKgPmNGEV4t4Vu+SGUSGXrdxd5zcTAoyiPJygOTysD0v6Qtko2C3MRNbd9iiRb9upZGF4JDNp
LLDgdDZ01g9SpLPYsZWZUiWl64bV9uuZuFW633mxnERKLlkVSHxyn20hUz0o1TuyrF+Jok+86Hrp
FhU87uZ1Irno1Jaz4R9feeBWxOFR8aRRUYK8O5wVmkZgcV41dLHTsMQz2ej3v38NR3x4cVaErKGy
bJlRKJsd7bxtweASAo2KSCg6An3YWBWPFNuE2rpVr8wUakNSwvtTS9dZWavuSCBp0Rd9D4thv+BA
KUsv3kw1e3YrIMGwDWv2XpSKl+pMGw+eKENtWD1GLnUHLQWbvz0rtGT4KLMOWyLpftmtumOA6TTF
rm7jHuWiUQiXIvZ16FVCEP5J5Z6/FEK6aFY10aft9VGarGi67UNPz6I/5RqkZABm3sGij2a6kybS
XSWsPF4JvaNEAh6tEs+Ov2YKdLk1XRv/THyVu9OQ63lgT1AzJZl20fJ+V9ME+USqr9bqTvPbovax
sOct3u+miEfqXEQAdbYvaPzCoN+GLSdsio1eJc0YNK97hombLme9/d91S7DN/Aud8TubbDTCh3IB
+JjrLx5yTVzLPjBQEuc1wtTvoU8l4qfn3TgiJWYR+jBwfKJgV/QTu8VI5XJ8sDBwt8HATQ+86uWL
1HsGuCLyvze1Owo1W+Au6eXzKbRPk+Bd/Bad6OijFWtgTGGgjmFfpR6xKnhLa48UvvbsO0oH1f6K
JixEh1VaMIVIDj4QdGEcI22WrLNNFxJhFp5SpDM4BRy8R2p9aWmOIAyTafRfOnewSfwPK6rUgaIf
8IrgDBQtdbvIj/nyB3RZXydaneeoa9Y6X4uUxgZU4rfUWcCJEEJ1zTU2geSlEz1XLx+xVK+H1UkI
XYwXqmckiaP7R1KV+VCLgfcVpVa9c1oFhakOJN9PzTCWSO878Jc8V3SzIF3EYs5Ot9pSCuMoWlWF
QtPenK3QeSSRIV1MuVpq2QTZtxKbfZAPorHIvu5PmWvGezjdk3tGf4j+Pn+1XFFuWl60VblRdYNU
2BG1OGYvuujzwHYfXbNWToOEgfj74K2fNVoqexOM3KtQ55NXwAhctXMjOUSS7SqtqBBW0IGNeCkG
RhzbLn3gkAozQSx6DiGJAVok7JtB2jNYAA433ZsZplGzbGjd+DJz+lYOU2z40XRV79WThA448j98
a5T+OI2wlwWSaoLjbQjz5l0HrGrMh0dg/5J5zU+WNX8Ib6eiErMQTdIm3DeKIcUVbYRfApphXpT0
5oNOYqUmzgLyH/OYjjFdSFdnWKC6mMjvXLZn5GQITn/aH8EaeSZM1fVZGuo6ZtrdImCC7Vffk2b5
xy6xnj7v25BLaLFfd5G8Xj+JLsVYexvVUAZt2aOj27sUtJKpgYjsyX613JT2qFtgmwHmb/drHxnd
0WstFGQB+wZdxOCOjHoCvyYltlF5QhEl/yxXKrYgPwFi4CH2+Qzv1cr88lib03RnOdCEJIjdxzwi
D89WIg0xSojpctpirlQP6rY0uO4M8773FweZmgknifbWvjGQnQUGumEkYiebuRwYQSp3O8aoXz54
drZiPBQnlkIk5UQQImry6D3HGB6OOMEbXldSI/81o3olH/qkj+5q7SOA137GU4oN/ZjyD+9B1rf8
4komdh7IlWtyl72Wpss64V7xcW85ijpA8g06S+B4EXW6qmaIfI/vszXP3qMWt8NGghWriMJM+dxp
1XRbKOVdi7e90SxQk04k2GtlV148Vr9gpCtMZHuZU3mzlNkxmUPIYfeYB2m6eT53sgNNDWiSBueH
0j48yfumOj6VEGyomg05EJyFSTRLMjgN+KY5xGs53TYUK4lu0FxOQ8jUy/iESzkdOI0lAUk97Kbv
A3XsEPPDdwf1MPeD/qOU1o+dUd4kqdSKJkw3QXQqzIeW9xaGggYX8aL8qw1lWVJtEUAJuBdTKSAo
j/H77FjlqS2pELRqbMJD0GJEpdtYB479Ohl/4a3lvIudW6XxPevPH7XtBxmfboz7nXSqqWWOZW5n
OEC/NIH6f7ysDbjTjrGWxTnDY8UWa3BotTD28OvH0tlGLX3ohRM/uyOsxgmHovmOtjxI1L3vv0Uw
4FBWaq6azWW/jxG2mrwWTicSPH6BFSNw8uDWSvJFl4A0jUJFwXK7tvNmzjiqs+1a9E1CZ/xNI8A+
TCzpeAjqj/T+cWZYgU0qWL/z9wBGraqR8EGkdnrbgr3q/zXXySK96OQ0BP+rgWFocSH84sYveRF+
OYoowAdOmYlM2WMUoNSHi8wkMsXuRA1tXoumpNfzxlQwcwo+w32XyBMUcAEacHHvy5jQoGLmPFC2
jRn50cUnv6zlT8XDt+OcUQlO8BGb/fOGHtDHVFSgetgGr3joqaZxaGiJ0ist59grc7BjkbI992MP
74a9Ucb3dtePUbAqwtR9Y38S56yiiWIvrKRtA5a0eSSLOKrIo30fw83WFTSSmJj4My3vSliDWCXJ
TGt5OowryJyNH5A/h6LmkOnyPyJnrx5TBGIKaIdR30F8poOBMJ/0MJ/CG08UWL//fUK/yWuXEcLP
i7NmeEsIQ/i8OHUBQfWnMtIaixMadOTn56Kg0M8zbsawEsOZvYpU+Yj1fBKw7N7/gV6GJ1fQYvq7
Dyt1V5U4unHFIZWTLiIhAC2GX1vu4xxl7i2/s779oiZkunWE9mtvVR97GUjUIBhzgQfhzrU68B5E
lclZwhxKdIiogmMk2QiDrdrMFOz9NhhrSZfSEXxg4ShC6CbuAiF6bOCtqmSKT5lthAbkdrB2pzB9
e3fKytKxdJTVhvrOY3HpGcWuZl+u3X9MNQmgoFaFYwIfMyffj5+mqxrrDxHykk+/2oyztf2IiALd
deOlNEuQpjJ/rEZJ73ewWlp9fdmO4l/jJGxSHBI7OeL3wYgOpdVcnu3gGoR8z6hhtosx18XB82d4
ZO54R/epHgGNDeDLX/UemqCcKJT1M1TcXFsg4P9zEonaoJottqzPaEMDqrfSDb9H+iEfcmtd/drn
TvbHgvt3GZch16K1K7I38FHwKsPnqn0C7b47JmaCXdTkbyOrkZHAB/C+W4/UCgPwr9HzfAQAnSZR
d1+SR154zyEVn7nnXaz3XCyboyHSinBazDa/EJM8TKXXltvNOP8Uyj1+zQywhX1GJg4gx4yeHpg8
0EEIqaBg/SchwLe2qREr1oBD0AMGOJgLJi/jTBroBH2jFs2t6gRYuAL7IEEAkCO5zNKd5ycJpXgf
rYd1Xa6nl1PGQ+rD4zaxp6UxO1e6FfbnmLOvd74s3Vy8ciom2nM2ButFarjEHHPmdQmdN2grrE5n
pFpkpAJSAlzdY0E2IwoKfORp8snbpmYc6YEqn9OFVwjoO1WpS/K6Jls9PTgu8P9aOwPnfCiBQMCq
caMLmGt3qsErR0dUV472RWS4xUbqdnfiAOcDZRM0QQW0lPcvp+K6sKnHnuWjd8pPE85TNQZ5Vl8A
xRUKbwD2xHK8j7ffTGqDmStKeAkxcZLTk7qS2PeGkLjMttSDfIDG3juwEItqEzpYCEvChpYjSaFd
2YcdrBGrgav4cg00YjcyA+cxifgeGroEH8uEXsaNN1jxOeCd+b5ivNBbOKKLb4YKQxR3zP8X75GV
jqMuJi49vXwYtcKgCXBdWu43ZDSJvnTf/TGqTjzc0G3RgOacxknv4NB7zG5cNM/OXIWbVOsCQnvE
vSlMOi0Qj0hw2ljmNQU2ozae0PrD/Z9CYiM2zjmi2LCh+zKZTGOh8Q+gqtCQz2hPrvTe7CPwj3aA
bPRn3TqIGS2oYATIwE4H8hPmp+6DQKrQyIVrR24nEoxuYHt3oEaSQIKx+Ted2+rQ3BunFaiTReMC
T4cyHiQZ2aPh9i9qlTmKIWQsxeIQEPZB8seBf7UqF5nlc9FLkHAfEuwayNHS7RyY9ZZRAC8wiJZI
CihJK8D8dGOaddDezk/o2SNwmegx3BM1vqMx8lZaihDApjVq92bYTv/wl6f0Crh3Fs0qkBBOpjM+
8bWT2M13pnCvDwMeRcSedIGyDMd9GYoulvxLWwkozX6xXFkMkMoVLlqidwxSDX6FYQdjvCCFFGN2
mtk+2kTA1w6e4Qpn/w40QdnZPVi6m5805iOV6r+uHMNJJf6pGTqsVfy8UhNZwnwbb9+1XsiFrKiI
rSDyP9NSK0KRT0P7cqo4hmj7NhfHX2RIcidHZl44+StDidnADVLmkXhADCYxOmfFpwYtYl36xSbt
3Zkc7ZPRe8NDCCX2rd9ZlWlig0a342vjDQ/ummo11xrGQ2CMXebHaQJuLVA8LoEmdVbbWsbVrX19
ryroVqW54r/x10KLK4B2u2SzLxHhoby6cvFiN18a1kmOIQfUD9QFjIFSX8avQ461byeh9e3T4bja
PqcVnuc0GWKOqO2yTZFkAtbn1wv6DKF2m7++EjyxZv/Y+cYgWpluxZKrXIvXE6oN3ZH+vdlTR9cA
LHC9FWkRl6N/gbQ+N4Jhp9aFeOvAMaHVZcGexfrwwh9jKy/dYQb3jsGwEl9GM1jsk7Ab11RV5J9Q
LZEtd8jcrJhUnOI7smUdgE2PpwLVPWvBRAsRuZvzQlKtJJynwQv3kj7ucz0iQFGoj5RsvuSdY9xD
+xtR97suPhOKA1uYoiMRomMDeEDtubJh3JCeO4dIyzU83JJrDRpSFZDxKmGpXQNoFU2aiLySpd7y
vC4pmn/xUgQ+wGO/Q42elFFk1RBTKcEha/bYC1hMRpVWh8aaHWchFltQFoegrEporDq/VimlFJgA
tMRHMUPoryzo4nugJz6hodMUfO+gLJSAQLz2eTV5QcqP8fjF3bgikvFXOI/gOzhxDIJUGsjIq4uw
M7+igQv0HUWHzEMc1anFmpI0EHE8thhZD5EWWUZMKT8kyMXPp13g5Nsi1uBibzNSk7w+D6gq2u33
MdTHzGaNcob1VBdpZdFvGYN5lCIddcaFpWSbTtfIQSm0O0hvQknA8hyoXcYX50OVdSgmfsMW22We
5e+tboaaCiODVGtlFaHTcjrh0N5h/W41QXxYdoGAP/RF29i+RG4J893NoP1c1VMh6HjqF9pmEJBP
/a2BzVG8yJ59jv5rIihbOs2oXZuPF/4ea91aGKcKuokYimN5Ta+kNIPuT9BgGHDDIgRN40SsaUbu
2u+lVZsnzNppBC4IyauXnK0ij8X1SvPFiQbCp8UsXWuKvS4yM5nDnVQMyKxedEjPxUMOHEZCd9qe
7rBFYog6lxhRceund8eVQfi4x2CxodHAY78s5clbwSWwV+lYRP9p+t9BpKzxWUkpLR7Xo4Fxa+ut
1vGYxM5IL0Wz3q7WYJgTYowUngeW6wglw1ceCPKN4TmZAjf/jX1CSy9zOTAJtRZgSejBnVm6k4KK
bc5A1F5zF8cD/MfykmqoWRbc6302SbtAW3SeEuRHjN+AVv5l7rxoK4gkH0ak+4FLEw77i/xipJOL
qtUh/ZYVgiQTzmMPdagZK1kDpSkc0N68MkBpdDdOgV+iMgx0IJCNxHyt1o1GoRNGctJXFtDN5vQl
ce3wHglV02f2tV7ADvZB0VN1sAAQtHXGkuqiB2P49tBW69wFUppymGOCMOqOPtNfv37kfv/eTChB
qnSZxerqji/BIIuykp81KMqy0z6vJ3YtCGIsX9AjLqwfsmMM71rFqndI118G4Gqc2Ft8xAPPj4bM
BzENgjWb6hqvQQ2b/lwGQjAN1bFxyKhann0mAdIjB/Khm/UG/psrlqpJ1QM3ClL1Pz8WYpUMhmNO
GWeJKM0nzIlxC+bnmwCtSuhepURu0feyzUzD361oEbWj/HL1HPgHpVSWqYWI/SA9MdwQnF5OLwdd
f/Lr8f6GMXq/H5h1eI4DOyp3GnV3WOWTfGnwFKcv34kZysVvN4Y91Y96NmTBw8FpGmcf28tbvjLm
SwwZmSHdBLAVYqvjs5oeMXo3AoxAqlzEPWlBsFXoeNzebQxAHBz5KOK9rEWdtAMKhXvJv5LG8LG5
x3H2LLPC29gzrZuCnKogtDFLzsH74eyAOUNa0lJrTridC7LCh2nKX5wSCXYPqQLJzAx1CEz9dn4G
xZukbwL0TY5tzYPsl0WkqucheivNxte3HB6dJu5slQOCYHXhQELgUtVzZYNSBFTAwcW1M8zyHsns
QN0CJBhgTt46MrEivBZ1O5+5LErZ/IMtSh1iHUSCxOgVOkQYQC6zPDXciZL55hH+jMkKTcHmRccf
nqD+57UujpaDURrdM+QWNL7EunvCTxPBCAmHWhyjVeD7RrPUrbrPx3LhgvsAIqS1pqJQ8T1JL7Os
jdVD77Gs5p2icFIkrtEL9THO5XE2z73O7rFkK21S1zoVHvCau0HCpNA+iLjnPFxiy66qGFq1wtEV
as1pIYbswGitBWkc9evCSgxNVtsc5D3tNscLQ8kFaoLWg4nHTmHAHMsGsJUgUeYd6gjLdT+KNgd3
zE5ugS37AOzsYuSsG/ErOag1BMRJSp3UfG107rAc9Sbd3EPANGqSmZpr7pyaXgcXSKFiKOw3zooe
ExREYMsOurdkyp3sQQAYuan7ztCYtDrxgMBAdnhuDHzbVrmBcYIhapxEbQEe2jgpyXCxBdMiUhQu
qsB9A83HRwp9Gl/IPD2r69EtKadkpDcPYYaxG8ro/yzPhuE0axTRe6iMU+zzHFXzbvMwEhMo0OuO
jPJmRcWN7YPaDt875+7Mo1MHztrV6DDRC5J9YUhqa4ibdsjpSNXU947IA5iud1KRlnsBmMY2pxNZ
+M1ZylsFsBA9gTuJ/Hu8Ur5E0WbpNQIfmWYQ58SEbhcrQkyQC1dBnQKegJTB3jtOAtEphJQvsxbz
eJ+6kv+s3fMLwGdkA7IqXZtSuobwMI6MCdGGFTHnrnd2aXTSbt6lWu6UWNO5t8puvSgLNELkDwkS
0Q4sQZv9RTIOEmrpBo74Sedf4LUD/stNPOHHfw1hT/Fou4dlpOW/qsD2Eqorh1R8JDr5SXqxt0x3
83AO70lmqaQxHK+Sltg4wTIZ8AUIhf3mv3KSE6Be5NBi3l8Br9VGZ12MfqVKpFdCBpsNtp+qGlGc
V1TY2/1YfG6qNPoGv5x9f75jxxLh+FQ9Cnlk7CKwWYOaIqD6RXh3Dokv3v1JPDWczZjdami5AaVq
8tA+slpLq+35mYvA8+O8AtQhaCsKqgmlUvfWI2icr7Wej5POff9RP53l6mvK14bsitowAMohTbCO
N364N8wn/53br6Ktut3+vkpPi8qQ4JhFrkwG2GBUgpw8z6IaUt2TubDWWNe7aVt3R5YrVCCrykxm
ViN3VZtlksSU0TE6nVdA+4R0uqCRnb4b6bsKAvhH2qupJ8koDPC5InYN1Iz4JXSQgTwRno4dyRQs
RJdlisPIokSZbRdOOH/sFdizMlIdSgcNjN59r6HLFRGzqKZDVgioZNMvuIC/2LVcmdOQ6lm60Drm
8+YBE+naGUijX5sKrm4K1IDzJ8MKBaFyH+Onuop4hiXEZqT4YZyUokcu0GQTcmI4D8GEN74K1fL5
G7CE7SX96kmtg6HyXdRiIOGwwkFdzctuJ8g6wMnCaElnDCjbyODtN4NwHdTbLSHUPO0vO754Cm1g
BUSF9YBn0KD2AcdAVQqPgR/Gx4mQlUF8lkq7zZ9DYLxhEZdn4EQq71d1ETuIppxB1yISNxR+Wty7
VAwbpkipDGYesyiT21T8hOsuTNIStS1pd1w9BcYk25alfEIS+0pHVhrq5pZnSIgWfKnbxDrnsJeI
KZPbqfOvXHzhE/SZf5z8OtA3+PNwP61XmlSedswqgE9Xesp4sYxswPibnPgnslMkHUBbLq8jTkeX
/1A58lUp/EarBW5F8DbVHGcJyT8zplrMM+Pg5vsoJV9j0d61rTyFzkmt4ZBUBSm7Nc5l2/jnFbtP
7nf46qUA9GIB1zjkKE2LyCERwfwWE5c615JS2h5dx+KlvyVJKq6fBtpjE7QrYsfGQnQsnfehhNTb
sKLx08xfv1m3zt6nmz2g+xQ4zxa3TWrFFFUw55gFxX++Sqcw5hlgZ+ISv987/VbkN4Lc1BbBhKMZ
Ng5xXDFy/iJGQkntCvGL3AAcQXTpgrRRCCQ9sRGbZuRmfgQLd3evv30SZYmSyMoQ+dw89HT1FbU2
q1OJKJNOpC+3O91M/HieKjA8o0Fms3GSmVxDm12D4U7XFDUlDtDKZbPRjUOyYJp+Oh/pXHPDhirw
eRI2sD+WgoDx50vuZDTfn87AJdIZviFaiPS6k14hwGnISUvViDUGzym4E4xhTIP16eEEGfleLCVx
cQ0NGLqi8hG6iXyCtWhoUzuakU1N2pqG4SMxE6lhnETS3hWLDUxycie7mDPd2fclSP2j+7ovGJC2
jywL3kVIVkoW3WayXcahdWvoFUW4aDTf+t32xwH6NRAqq087o2/cA7E5UJZNUnVitGLZ6dJC/so/
AQ52uHs4WU5LPbIqSAOl6T1fxXVK9QrPgujDFup+2r65ih/f7jBUv3zZC6gdVWMrmxyp2J0O7wB8
13T3MG3gGG6WyPWItLJgR7bjMd/tOx+N3rMdUOH6KoqLm78rwgp/eaYAhDsqcjjku0BjvLtDC5ja
Lq0mvZWY5TG+Wq9ondgwv+b6P9I9bTRTBbx6pqgsL3SPTX77THFOmhVbnN4NGUw82ec+Y5VIJIUS
6kbNQ++DUmKP4oFC2uviZLRBga59EKKXkAOEOeehuqb6igSyClKnUpP1X9L6EhyJ0hj50pi4s4Tz
Xx06Gc1JESxm8g58i8VjNV8XkHYPu9AuGTlvNL3BJ8Vr6J9xoOVIm0Tv1TnUv7TpH/+fCvTVszeo
SoFmC70H6giS/0+/oadd1qiRLfVkV+La7kwkR/gJQm/HMW1V8g1aiq0U7rFMFIGJnUntWBWNfZz0
d2EGEjuwiVnvYeWNS9RWGpkEQnIosn5mr2w5vzF2BAv2Ss0KMq671RUPRtqxUP31UPSzLD5V0sOA
wSzaE1JV6qlJUOkYrKUYQx7kpt5xAAZ/czIYw7qVp9OgJ0jrQXJ/voTal3r6VxACyT8m+hKOcqwh
5fuBl4fyqsFR/om+KUo6ujlWXPh24if2kH15hUEnCEayTUJHpPE7IYrAFt43izBZ9HU43a+ZKagm
QohjwdYovgv+TytjHV2hOIOqU4uF+tgPiFRjNRUHZ7ph7lE5RmKckv+WL3+r/D3MaELduYtwxsR7
HAiwgbRsi5enPKCCsXkKrp2KFy4PRCg/AUA/nuxvrX1UJOkgYFTjk3T4qVNECQT1AIUKs4MqVj+O
yU292XazFVr3fa0+pGs2IVvMQeYnWHH90kPJJjIHs5jTeBpjGrIQyDlArIE24HkYk0H6Jm+OQVvP
7VryA8im76yAhIj6ZcQEoGhqLoV5k8Zbhr1PdiZjVoIj1bYvcaAB/bzHcbfUxuzpdhAr4Cb2R8MG
/fn2F95ez7N19xNCNCVqqQOlCLPBzmx65Ws3i3ni4p/zFyd5Bkwbo2FjdRTZUFDOUoDqNMXn/C2y
p30gjqkZYk62x4NBjpt3LXt1psUctyZ2+cXOnvdFeueGiEPsYrqTcRFvCQoCNymIbLyz6uL5SVPu
JbghwBRyT2tD5HLRrq6LKZ3Gz51wv3BWErufVpN9pct7+NMiLOgbWVV03eh2/KUWq4OrwOGlF6FG
JWNDlbWYJR+qha9jYpK08g8GREcqMlGwdXKyrhaaMUzma2I3yDgzBALuCP6euHO8Qfb7ZgZF55lE
qft3u5EROxCpD7DAD6uvFODpDCTkYeYiJIGSE/U+C9l/EshaKx0MXwwTMCO8zqW2gLwwmvZi8M2Q
W5aIO33Wr0pJyM5O38uce7Szrg0JeTKULIur+c8uYWn0awRjOO8e+ExZwdJ8WZdWjjAwNXL4GGC7
0l99tenAYJJyMLdnN4LzLAdFRqgA3eR+lw7nH+3woZ6Q4tncwme0MtsrRKO8FIRoT1HUurMOd/x3
dDzr5Tv4LAwbvDlmOIBqQIi9GI2kZagsKK2FvsEsQPEtnhehKcjWTGAE/M8KBQgYuLO58hiBc91x
472ZKmt5a+YFqsn8YBrTcp0yalxqc3yyR8RSlQqAkuFpvRPuKwRdS8YJOY5FTYkQFeJ7vOeR/Tvo
Y9g8707r2qcKO+RI7rsOLEJjeonjzwXsVA8Qovyk2ii1yoa8hC5NbbLROI7oVMCIn6vU+mYl5Ba+
8UGplONZqLQJjkxG8vB/uOxCqCn8DnDQk1161t7C/ZXdsM320R6ukyy7ZrARBZzD1aYYoAzfnv66
TReN+HquNj5440XWBNWmb718wXSzJDBceUfR9Zke22+li4kSBWp1hqCwBQHGn9qmb8I/WDaPDfVV
RME7KjOxNvHSVEgR30BHR9w6dfrFmaTJvSAoWVAccoZZFOIEmdKBK/brp+Mu7P4SaqJz6Ep/b35x
zOWEqaZPajRSJ0e+vG/zQsb2Y3tTu8vWVIGsLa2H4oFb09Dw/Dxjrt2eNWeaXF4fI6sdQI349vvg
zxi2ZCaQkj/+nVV2OFHC55kj84l5rCSiuZxewYygO0h6SNfud/V+Fwt18h8yHSbOXPrHzJNFZrI9
awR2p6Z1tphNP0/PG1xgeXzDXRukY/umErmu/aBNTJg+h+xt2LivReOIRr7YtP0JWTN8xXzLkWJq
tPSJV+yFWQ8wHi314JzuCe1eJdEeCPRfDqDH2MlM9U5+mKCsnvjbuOHOqS4ShgSkUANjDoj01VVY
yWZxjVcRCp/KdDZiv1RzGO5+MFOlfx7LBNNPaSK0g06sHU20O0Ri7AJijCqehzHAPS4bKgRucaWP
++UrQJ7Wahjh8iuc7haQn6s2s47JHEyUGmKzP9RjW/VpSAClDV2twE9AtzykDh4wOT+FTX2d/8vK
Q6RBmpeSe6h/a2/kGj9DZUGWWfz0jNkN4BNyxEC60HRcCsa4U+kW24oHejEgS+47/3Fb5trimhrR
WVdoM0MdzOZsj+pcJS9i++xcaInCjkS3/YIIu7tuZ3jFRIzE9ej5MclwedQ72m9CtkrWdehrK//6
nz6QOhf9QXIcaID/+B6DGo9MUBIzJ9hvOlFpEBTk4hTuwSWYKgwuDxBTrx9PYaGksiKs9NC7nuYs
qBaLJDn/f5Y9ajl1SOs5V7RL33mqc9XrbfLlomD2fcGoFDStshLxBz1KqIEib5zVrBPT07/tTPhT
s89uzRZHfp2RDf8u7dLwmPacpZPsrJIKaja1phKS9p1iBmNhx1tyHvs6J90WMjhJqqhKa54BQKiC
ACsJiugOuFvfTnecEoOwUOEbpUqtlFzqBrwBKzcxMb1SBDLh7zMA1dukeDladFg83Wc0aJWY72pY
dhSK90osUqtpPwMvo7Tphu9kB0sDA2TIp5/Ry9c3y2BWPOr9pGuJ8aYR8wddlVrH/jI+qWGrorT/
5mIjY/MBDyJP8JpvdE2Z6pcls84PrNwpYbx0XLReyWKkwsGEvj0aL+IwH3OI5+fkCzbp6bMvLG4L
6rkeNACLrLYA/f8ZKcuKK/jEYD3wc4yqUGvGzFNFKHCR2x6fTBLOJRJrDnq9oZhhmcljdhqk/a3k
TxzI3oMC3IdC5iG04NxWIPMOHDh6s5Z+euxH5C03dYSUN01Ba4ec1N47sNqqphQq4yL61SD08Jqe
ropXORv50HMgQafdG07KCWV6gMIqsfx+TrxY3QGxSGtbYO+Ab7LFhCiMakwIy+urRADuhptiGveb
6iFdtQVNry6QEjsurrRgNPDX5KOtnU9qyG34uDjemgy9STj5MdaxGUqo78zSQw1ydWY4PfCkQy7v
a9omIsAXkG/Ccv7BtIE0rGcivh+RGyLtVscKJ+heREhvzZF5G5QWkxNBEZXlmfx0riG+d5ewhORe
9WajsPlGTgYAD3rwWdIH6iCycFcisQodGjOGhBvgV5vslqVATkys32iKUHNyd6bidDxb87kIdJo0
IRVevAfG64KOWBQIhTD+2pSqFtaXgA+0pQFlmi7kbccYNHQNODHNnZu92LUgVpJHgAia9sAjiX9a
VK/GQ3kNPl7QdwUCZGekWvC8eU7LFn/7YTpO4/wsaCB4HxCOv4+Ia5G9kyyf5IB/nV6JyYFCR9js
EMlrvAWD9O6XV3JbG1cFoIz6DskGBZioaE/kxeu0apu9jmVZXZ5AJ5Wax4kTRZQSawymDAFo0X3Q
Vo43xy8wRzX3eX8BigZfcRBh+qD73dVwA1vW5WqFsQW3eBQ04ddPApWi0Sl08JWkFNabZQfRexCO
M6YIuzutzB1tmp8NGcVmlkdoakIbsdAFbJZIUkujmoD8hli1CItkLLdlbK3kQUOu7AUn+5/ddvN7
9awgLwC1dJHWZfKoIcQMhLJW4DIRFtcdZM9GgluLhbybdSyJ/mEiHS/g6MuBZKHNCJ6YAvrH++7E
+FNzjt4T9P7oPRY47DpkHtBvisEcQZSB7UkgUV2MwNDwLGCPeVC+kTOe2nAVl5Pn7tlBf16D8ksb
kwz1jN/nB2rUzax6xee2ttH+cu8fYML8NITrQGH7YcbHwVcxWX0TBInGiDwKFyrbYi8JM6FPhKpo
xySSuYKw2isLoTt6kmUJiIMp+vfJETtp0XA2eBijaxc33LBebM9i93dKXXYznLu5rsn+eXtFd2/T
4I6W0fvsoSR+dgju25VjAwQ9HceFu2j8tjCmjhOKW7KxeBC5/DRVkloIXQndrTnvlxGROE1iGj9U
+SrOE0fg7ZfXVujKrSub/Y5YrJG0YB1ezB+U5o2Ppr4+2VDxrUmTL6sPHlQyz2KL5Mezvk4kNAe5
ry8cHv5EMK5XpVsXKjvMVlc85ST35oRwKjqEgMCVjIvyCKd2/4Cz2COMM5Y3zIkfrwzgCLk+pjke
sR9Qz4LdXb8ZN80uV2vWgrvTIfJWNeB+LWJVtO7cYNCsDiuiFQhmbIfe7gVtqPblFTYX6pX+109l
d5pqzoeRYf+8sGNJsAR4jgqcEhz+qIq5AjHjq1RSbFg/N8qso77SpADMS29MQLuyUyKjwzZvwsf9
0tqP+aVXzsFBfhgEuFDzvkSWXyYXNAkq98vl70TU8zae/QXA4JUFFKmyo0qMTAEFHyDDw6g3j0Pd
p7ubdRWbasrIYbk1dA6EvnyQ13GUT3qWAIQUqyad1byco6e0J83/WZ33vGM2+DkHp7LSNYLUMt2T
hdswgCSgqgY/du1HxaZAWOnueofKnFiZwtIveSu0ROlV40O3AvkxpEb7OLHW8VNdEM0o5EGIrfFG
eSD70/L+SotVkiKO5V1p5bZVDzelnRiBrgK8QLTKzZY+iWUZ/EQPTV+ewTBHkPllLNkaWgDJ84V+
vZ1Kpvkh07AneL9c2r+7JYh8YwwtyC7/vgsiXMsctGoOFz2X6fIkZpF21gam8Ziv13mwyCib5BYT
jGQRu9hNCHUwfswgDVQ2di+ae822PPWV1SIwSq39V8A5aH5D7WOtEODfq8PxmuFc+7KhgVndEOUp
GWv+RAheOk/9CzWg//+koEqe4rh3eaSPQJpIeevz/hw4Hl4cwlQWyr7CvcSpBtWfT35YrqyKpMG1
4PphtlMgwqj8UqcQxdLUftWubsx/tgpGbHpcINen2ORoVgwX7XH8PbfsirCv3HsZqPBiW28Ov2/8
IZdCZOC1k8uSsYOzxNmigDxUm5bP6YJQxGByTWP2uCm+nX+ExJpcmm475/pkqSqv0A63wZ/NlSOt
taDBDXXT0TpIHGgIEdUhV8h1qM8IfIY+73zDSTrLuI/2WXQdBLCFvOIaBMgC33p0r7ZzgZH2fghL
13ygFrj2KT0EvfU8EUICSzCHMlrVfTbaTrAqXcjYej7IjBOaD7RT+axctRrM5d2EMrnUCesHHQPD
h+5Lu9v/hEqREM2KMFbtJ4nKTN3gHB10KAeN8+0IZo/GXxgPlePt4EqFyeqlTzsOliFUggmPklMn
+JhP6PG/4bHr6Pp5jZiomZZX1JwwcBYjfwslesbefwreg2qM3+i5lnTKvVLQ5pF9gWs4srPgk+bP
ETcUGQ2alQ39Sr0KA20mbrzaMkIbYDJlbhyts7mMVkQEj4aQUGm+IW+yFW+4Y0CNz+j2AkSJdSre
ZXaE10vPJPy8l4ISf+XvY5JUWA/F4MXb9dJfIR/a6D17UJ49OPCrYBpQ0enQoPrrVYFNp2EoXOMT
2ZfcwwyPv+oPDrouNRacyeUxGGvBrrHiurDPM34VoRl/4BPRalC4Ck3/PvaVawueQxyYRKf+Zw2r
YUiyeZn8rPfLLmNLqTVB9kev5KCbtW9nmobUBHWMGB5QafgvAO5fViwrUHBDRyG7FbBJYO3QMQwQ
74pcE/PV2AB+V+FqMoV+s1DRhkSpEyn+DeRIcJGXtljfxN5+8yRzWtxWwuuq2zg/KDGstXsAOYOO
EhOiwlWBPgF+ZnrUU0Wsy6VYm7XlHAa0n0KrcqvfnlMEs037iuAY0H1yo4rCnsFmNTfjAYEXfrMk
vGQWGA/dozF4LXgubvVk1/7loTR5J4AL58GQTba4Dgls/FGL1msqfXfGUuuBIBdxDbzlB1a1Q3ae
rBkDKQszkbRis4fatF8suNQhWlR7i1reGGPlJ2IBguPbjfisz6mwAk/00lzj52wCt8EA1sSsEtdt
jiw6Ob5qVqwJlu0PJNgul9CGrm3oW4FvsTzVgW+K45Z4l7eQhsXYdgzZ5QBPXvMRA7ld9Z6ZMNkh
vEFfFkctadCgYduRiQQCySjMQk2iCNEtKeY5iHMyQbbB87fh/xT3jpsnIaEmAKJMxJhT9Fv+c/jE
/4Xgkz7dJCzedPbWb4ekeBz2IjDg0V5voSMiow99A0eLIDTMwaYhoPJ9qGgvp0tvRBaCHD47Sttc
+PFsef/bFKq8N8olL7YJ+ylzhq9B/08oA32PWRVPpfWO1P+iPDhW0FXpEVT9uY7AHPQr3+la17YO
lPUxBgOMIDZ0UP/vaUyPa/JMe+RapvINMGU5xeOBoh5bv2Z89hb36DOG5jtmcK3oPIJfOdnK54jV
RRnOb/Jkz2RLHS6T3lOBzBtmPapvp3PCXO1VJdXExRFyu0k65k2+FxDxwpsfQq+wdixKb6WrsGRm
FL5rAT9vFvh/42HardtOi1dP/UmcT8vsR+XI6uMZP17aSC4Y77IqMohOfu9jVjoP/ALHFHn4f00x
020vniS1ppbSam7OR5s1ftgA/CM3XxnTIodi7Hza30d0FlwciDPoRpAEXqdYdzIracZ/UsHEgjH9
wpfw9Go/HB4z3cYvUPV2ZkcVvu4jwssA8fo9k6sI02LEdlSxr8ri82bRCzgMFOFFrxVGKHh5iU/0
3jBSEN+wS5Ee3Oi1fk2JsUc26AlFEOGfMIYS06ah3oPLvSUf1f0oZZbChfTFylVzhFCeNI4lr3Mt
uQNd1EFWeOttNG6kY+BRVf2GP5Ngur3ZeVUPc8kmjjtPnKL3v3qbn+boWWQyxMkY17OGpS6/8c0a
hy4g2pc1Wj186l/NYpK2hl5baZEEcn68SKmp7D1drKrFvS3VSn0B6Vp3cZEqCaf+QqCD8r/hpZqi
LhEYpJdQEPzzqkhcmNV5ZISYCSdy22U3J2K9AhqQIddF1VeHxDBBw/xKQg8bAzb9EW7V/rmfDRGC
ZoLfLyJQkk+TsVPT7FZol4WR20ZGUQVxZq0JVHnk9vNyvjjEBoRswlvH7+TPbisvZ+26PVnxXSh/
5RieDJRlP/LPAWFata5CBLiyvh7csRJPBVwWgfgJ0SUBvEo8vUuriOWbUmhE8sorAif1pvkCEKfk
y44z7Hbl8HDPuPknlFmZOtulPA9QiwykPBMu7l+ya/sLTUMwuqv4gdWsoJKCYTLiBC32xhtXPllN
ruX6fq8hTMwLPRBHr82QDCK1JQJuKxKsPcgU5SN4wm4c6pizUQ61mO2LvIsx/HB8VXNeziYrel59
+0mCqzwGcTmk0A6N3E2ckp93uwMqEQ1W3kpOHQlkba6gLlrGYZsfqowOvzonFC/h8VRlCSAf6vhx
1zy8ubWagT2zm13riidY0PWpbyZb+Mp56OEQOUy8bIm406C0PfTvq8cwrlnnAkygHffeTPv94aGh
o3EHVskZiBAkCUZUiY+iyKxv4RII9dmneG3BikCbO3ypv7fjxSraLqpvOUwi/Doi6TGrTBGuGavl
J0jGmRMCimOOG8wv5iIiOyZJkcKei8uq4Ldr/ME6qTgneN85YwnpcW6O8aH8adxVK858/afHuITT
N7hJwPMyS4hv+i4aFwZFLIAIusoO9lbj5iI+R9bpy3GzMR4USZMXyWDiVtJOikDizCHiDvry0CJh
rX7Xv519nxPkjwS8fDyiAte7NRJeZYu5MdhpoxwaN13a34uQJXeDe5loQFpGydnEwzGXRDTEfrkv
MA4qL8Nx9dBNvTypEyxxZRUGueduVv/iViBKvdp6EHGMqyqBp/8E1na+LgHapLmgWUf3aaXmVlM8
v/s/KPX2tviRK19afCq8KuMPKlmoWZCz5hJtKeOESgsHhwL04cenZbwdKIabht9One05+ZpzJHsD
HNevdxnoayVtUXXbHhCOYxUstJ1yPKTeFO0NkWx8BiU68ifq0XFmv9u1cCzZp8uw4NhbJurA6UVX
xsygsFUkl27rOjpKcjdzXHyIDLglqRfZQYEDcjdMlhbZ5Wcd+VA7zFDUdEwmrwaV/HbCAO7z52eB
GDIbB7lQbA35mNqpievdgNFB9zp4mjyVEEB1yJF6BoE/ZztdMFtv8ZZguDVHIOsYKm6tofnQvDx/
3OaoFjH26+RNbxw9TcFhwlV9kKl7CkLS1ofkW5iqiWAcnsIO+ILv84W4BBv4oDqkQ9aYG7fYLbvA
4Dd0Btz5PNO4ycxwwzfCsDOIe/PYtcLfAivfO1SQTSwlwM5qXiPdD1N4GGmPxm1A/8qVvMEL6QyY
jfhf6mf7HKajRfGWuAlypO7H2OiMx1ea+EXvZJqojdbS2dhyaUKUy78SXaKf0VLrUFZ2jDybsesM
gFMFIMkFUGX5htotquEaZDyQjG3eo3J6NoPsGKu9X1luG174agbf/DHgFcGw3qG3HxV7poti+D2z
tT4dcS45s0Ttdk9q1/Mnlf4/sETbfkvqDYkKKA62w57mjA1jV1lOyOBH8G2kfieMS+/r0DAC+MO3
zqg8mlTrjz5rXQmrghn2VJDqphstUAYNVieW0zR3ctOoGlasMDD1hOMAMCTmCTvxz2OEXWCGJxEm
vnYShwrJ5ndOvbpxkcG0cgY+SFbRaGxsmDROR4W240Gv9p5qpFgZjPSZszBVzHEW/Y7ozputg8mS
p2RRCVcu7lZl4EoDaxxV8EXcFWJVcezR/vrMB6FEHEsk6DR/lRnd5UMO8BeaNL4W+vUGfPuYXVfi
P2NV2qB+AKsQxoMiF9tXzaLrLQwS5NphZbptb/sSngMfE3fm4wgg0UyWCnag/wx7w5NKQr+SAqKv
rOMW6h8I/QP5zwHookdtSYPQaJ1t8OWwTcTo5TTx6bEY9Dpe93y4moC8meCsA1qex9Nz17nTzaE/
UwlPKBdlyWeKUfhxDlAYPbZmig/xmVZlqGOz0o35sP3du84hnqtugNlvTXHp3yJ6sAUKHK19ebKU
zj6Szardolo6QZpr7RnQwCDCDVLI5Vu4UeCJ8MwIvJfaN6RVDSQbnmokoIP7ncWhTkTU4f3YUJVJ
ibOXDQ8xtpaObPMsbOhyYXiWFGbrSIfGHL+HqQsyzL4Da6MF6cvYSIQQsEwqeqcDl0qfVZWXLT21
dzUIIyyehLTTL5JtKoSMWmFqWvP4mb7veQybfxZ+mE2s9Jflmg/AtzExaums985htbpsT0PnPGS4
tR35vGxrFoPsIdwdsSkS7gf52MZ+vyNzlUjNgD6i0i+GugWDdkVTLkVAaPcdQ3KEkHIGpOIffLO0
/Zz3Y77wYCdHlZYQg8WIMKdiQ0e2w3A5wXqRLcoYvwxpOWN49X0iVzRVOKaUqe22yd1jWW29edf2
y+BEYXg/2AxLmd+kOy1HEHLFmhIErjgkq3OC7sHJ9C0JNonNzJmdJKEKzMqMvTmHEycsgUcnb0cv
E1xaR/SAwZiSM0kKJqZ+yUaiZlgJGO8IOX3wgECsxTj7+7SChtJhxLphnmh1272dInCdzbds/Unw
eypxI9jTURXl+Tz/iZ9RI+0PP04aElNxol/k309fQJN+QdxRAJAXR1FA/t/9ehltYOdHn1E22fkx
1VWyMGdmE4QCMFVi1UXdm/KIBdwdc4cvUz1tjVgRxXbfeA8kHrVLqq8HAdHL7RcazjNjMKA7RYzB
x2TGy340+Omhvovm4b9iBdl7NqJh8gWEI5KTCVqQXDKqcGJr8QWCqx3Xhgr3IGyXV0F3X2pXd7ZF
H8pj6vSLacgjFd+DLBrKLfCZGpgKifD4jslVbxmGdyiyq2r1U77PL203yper0qPYdD/jh9zFKEzF
N34or2PtcteR+pS1FtaBCmQr71nqM4S4b1PofsQ/XGrmuYZKja1nfcHM9G6NXxmwiOtLMGLnabMF
YVAEhL0e9oJxJMc7ZvO9qRFHTqVGELCGHdJAbVod2Jk9uh4TM0nygCFDFYCbsAs3kLf+5IMu+Lti
0Xb1UCvkJMmc5TRHI7JH26mE/W72S2itDojlL0ZDoMlhErNL//s9fjGCU4Ae7wpZs1rbBWeYu/Gg
P/st3IeO+PheMRMkVULGO7z+uhcfwGtmgM5B3gim58Y3zzWdcc9u46IWyKc0RV1c/J43qAIwnQSk
GwuaqcesP4faYa6mJBevprjFqJMj5DeUHPElf4z3UssQ999ssmIIVYYH+FXRq5YvBTu8ofd2TUH7
TNgkbhAUDURGcI/sejCue4xg97NEUs7Olh6cJ+5Flm2eXV4NWbNB4svGIxrWfo6bnympOnMR8TMY
0NqGARqO4oLjRQ8jJS699PvGHppi1u0xaI/ayhqJEKBqWrLRhRiPV1JQq/qtMV8yMYYm/BqLLhHu
gI0aFBTHKGWO/hrgivDTt3jBCQQ+xzmxTsCzm+iabpwlOTKevhzePY7FqUAq151uOd2o3u7rTdbV
2C79mWqHRBV0O6w+WwwPVwTVoeDz1lsUVGvxX2EDK9affFPnm0lLy62QWOcbkLLKaSfo7uFrHlfw
HBssDiF5Z1hvFpKtZx3sBKHOWW42UFc1SP3P9z5FjjJnXknmU4exjcgLfuoSfwuYN1+8wjGULgJt
jyRRkl9aZdWKuZtRVFg3Y7hocxqVZ8Td4yqsF/n45Pyy0/XnJtdRszek0bQZUzaN5nV1fC52GSuT
PMKLcDwy4v4Fk4rZSxMrJ+uMJ3v8KjSLBvi3yboSMjw5x88Rfi/JdlIm/8SNgl221sWa93cglEoZ
Cl5DO/MWWTGx/2kf3rYPh/LKaTt6KSZMxcKzvqM9cML55gEKjusHfv8SYJz6whG8DWdaWM3aOx/9
mYtEFnMVJ38EIAgB17BeGicJ5O+mE9oWtwJbd3LfFdAerXDdOJbrVN68sgHmVdx3IIBp21QyxN0m
1OzYbjchrcUjEM74kQ+A97N77aXPv7blq4W3MOpeBCvYSJu2YBp8/GuEZHu2rjRwsdEAp0SlUEj4
P5RB7P0utZO9aBsAS/Ut6njbYFeJT5B74HwSk3ukZ8X0L9xkmFMZpUOkL/geZxZpKrB9Sp1N+IDm
1GlJKqH9WsNaPOy2faxAA8LlasPgh2ED9V+HJvaHeC2jv1TtT8snHgwBtC/DOIiit4sfIs5pGgQj
OKgrlCQ45Ie8a/CRXTpRYAOshFUlCdshCB69REhGB1M4dqyxv2pa/TW2up1iRfQpirMDF3OlkRmp
bK1xmDk1LJR21gdutLHApbwrNe+wKgP4xJIpFke2uieoagyH4S2RLsMWQmSSFfuVA1sdVCMAOpKs
1H9WX45cD04SxbcbYH1B8YSMPO7sbxIhr6D++Q0HC5+OJnSzAlb1Zc38na1iV8rTbdk1tiakPuMQ
D1pF4yKmM6nAfe5wvtnGA24/8kiq1hgKmUnLQKPU0Uv0mMhbzSvVNnRLghXiGrJg6VZ2SFjUAn5k
m8m52LY6RN59vrNi6XsuUvzd7b6wGSB1Fhj9jHjHGfndkjkVcx5Xx81b8ZGZlBTaBE94JRJw8lfN
EJ1mLDQUQqWWs4H4GsFJ0wMV6PSIsuB7CdKmBd0dpkrqKCTdBmausFa5L82RO/iefcFx+rUKrnEP
pXWClibE2mi2yN2juR0mV0WxZsdL7i35NhnpHiA5p9XXUZmAdelFBSRGjGQBVRDSNLVlGnFwkG0o
fAOVjY9KuFjXrDhWLRvLuwWgb3O8W1RHxLp2/k3LJeeKe3vydzJsXSg3A5170HVRIft8Tn1fknXf
V15lFaQVm8sCN7yXpq/kYs7Q5IUUbcq76Kq3S8zc7/FMKIIqMCo43EY6z0fEs7Y1zeMbcp46Ua8J
6Qmx2yLUBWOViNCCwZ3dvZKfuuf6IHDaFijeET6ik04qjREKLcBjx+gEg6LaBLj24LJS+tDK9VUm
wxTlA+xWxLJQOAVrZwRMNgCOFCj7v21fk49Fxk5EWVLwVH6o4Bq5QinZzIdc6y4ogZ4l6pHt5aK2
bY+sKSvehJIcw0ePyc/5NgLVSnJ+SslH54QN/SBmTz6H0fUxJ0S21PeIC2DfIaLOfuF4ZHIC5O1L
j4EJSqy44Om+ET+G0Gww+pkKfRB91z9dJX6QgjQEzQDvvCcV+5blFeNjEgd9020oilfhjEBmhym4
5oN25rmODcIKgCK933GyfPvXlrC3hYBuX2Sjx3Suha0n+jN/WI0DxS1dev0kbLm6bDqIaCB6DRU4
uqq84pz9HMhYlf0uvVDKsNJ/lg0Xok2qvOudBW4JI6N4tAYU7tN7DzKj68jq1ESgBvh+x5mcrarA
4BP1HH0Dq7RLAGf5Ttrva+O6DFOP8AFWr486smzOQdqzDysLNuM9sOHJpnL5m54XOBXy71CHWA2U
U9s42WSSkpEsb0FdZKQUs8MDViZ9fD/8n2Kh6C7jo5L0Zflmh6xg17DMgzPodD0rcCnsZbkg7IDg
/xEkrBO/YoNU0S/iYJNj7VGuxUV+eqQR6p8L6uGmuyjtGgT4/qzIRBadXq6tbwhICyTfWC/ShbcC
QIPG8d3zzVCdgfbXDomQW/kmj5NPQYOUn1I7B3rrAZaPHvgWY2gNZTgtpA0EoYZaT16vv4Fss7+U
Qr6JGpt8R3IF7mwXacyfOtDGGwAizmdNcqaBYfVV+vLhKtY2I9sy71WjdVVG9A9oNCY0VYTPQDhC
ahCx5hE3nJ5xwwjwAAPfsP8R/lA94ZJniCPJz2//vZM5y7r85xa31y5j5kD4v8zR7MDpI+19NXKE
6yqc7qJukal2NPpi2op0voOXLqpL8CBu2lTEj4xfeHoVy5HPWVA7n+9raaHmP9CGKN0vE4iKb5Ix
Rt6XSoVRLNHAeAaqYPA5WGEQNx43nMyjV205e48DZlvEjDBUBmZB3fafpRAIvZegno0eluCNSNtv
wvvY772dUoMYbkJM7mruCdfJ0O0I+DvGp54aVJ7r5PVYKaNIVQrch3fTCoLf3EMN6tKNO/TQDR+x
EJzJ6LL7Vd6LmUpVKnPGB3XIlPCHUxMKchmZKcR1OjEdfLrLsZC+16XnSrbVxV7ET2MiOn2n548E
rXq8ky+kdg1oVlNnm6P8qP5hU8BZhV7dIb3V7rcwu6PjOe9rYxX6Ry0LhOcrhqpwA0jiLzPXjvEM
9SxhHCZjKIHCVJNAkWPPoHWniYWWKG8iqosZ5r9As760GqtA/gRaidjEC6MCrWGpYzUIa1Pl8FW7
4vPmU8SxdwqkZFHuUCFWuJCrE7yBT7ejBs34Q5XG83Q6wt3BJgQ/i0IYqZ2tmTjrwPCQaK4KrwoT
BfMPbgMZE6BYcjEvCfPZGNTAAdZFgdTY5PIaKSceFHxzMyE2wiZXntYZjp44yri/38KSGnXWEn96
Hc4vLjdyU8IriO5YVJlu1k1soPu5J767cKjH3FAUc5Vyk34wwLZAaQgdSqIFvKyg5qc/Tg/f43ye
h/5ZuY+mWTirvIKIIpLzocXg+0nWEk9JT63go6y6jBiREN0W4yf0Xb16aoSiUyG07/1w6/NWWjCC
nhk/IApP/kIqRZ8sY1FMjWDxn60jxooxO8Ods8tLl5F2EcP+q1OMJdX4O+8cnUTI31F0B+R2EL20
JI2uBsadv6WriYfg1PSIwomyFv/ygMU+AMbSErloU/Rv2+1v+jbggtzwY8e974AMLvcjkGR3UUF0
O1Xc7SGpUuMOi7gWv9p3jwhjwYsRYN/9mWonk0Xv7zb31JnJBaEFnnFgg9tfIalqdRr2T5gIysmv
sNPKz/s1VfS8GDg6kmoJts4e1i8hwINyRyhGOMAyVhQUOxIIYekfzhvMmKLRuC5ioB2fnBmXhosW
bS4G5lWQQO0gOULRBvvKUOVT03xCJDj4MrbqQHoAKhxdoHrvjn2M2PoNBTSdlD/m+exz2Sn9lRty
osDCTRiUGQtlcHDxec79GVKHvCPkfwUjY1h/tbyKB7l4B8/Xc5d0YjkwdQCUaOE2eyYqHQy66tik
/5V/O0XEjLIpn6O3xQG7Mfpv+fcXIoDLPFMYL8tdOtvRZfJ9pC6mOa7oJyk1s+Hzq/BwBCA8XLaq
msnmdxyrrxN1hvw6l5XbKLdlLI9m8+TaMqhRpG1TGZu5zUtI07HIrTh4bmO0jlOlKndlChifVeyY
9Kkx7aMLYLEXx2rUaaY9kz/IU6XsWflmO/tArdtedeXuTQ3wktMSBIQpu+CECDRtiRHlkvVVwl6l
h9agJwviWc/6JOjdKRxoT2DOl0SDJsda5TKcE7En3ZPgNUAfXRtuBII2hGjAoxztCXM//m4SBWXJ
prvppRs5TK7PnipuN+hGG/9XkX72MDjpSO4xwjEoLnpDuWZkmAvdOMc6hiF8xk0HxLTtHvawj8ji
7YWN/2CE6rbZnTgZoTqpqso/AexriMT5Bj+rEwyBONgE/rzJzR5XNzjM9Rg1ZM3DFAMdioDxpUyt
mIWgcGCGAYsWdxERcWTKOgauAqIrj4jjdPtvEt84k0QBaU/7T3rHl9sZROMf93zIYTqr465+hgPz
MA688li8LRyRdXlpbJBnf5PgrP3lWMxApa5i8A8LKclc6HxFSvCzkCwKa263Mf9MtI2YI9Sa/McX
5hbCjVL/+SL3pul9KP3AdE0jaOB89fGb16T7sqtJKACZl6/3JiDlKzG3n8DCCJqzmD8Jk22dxkID
LCb4PlBHg0PsiQymfTaFShUJR15Ale0hTjygxd8qsGf+5cjJQ7sRwftQRZWhoyv5in4wwxolxFb9
k4SySf7bvCTzC8D2tOipgHoHSqnlGKMlSUTtm65RzLTEd6MoYB4iktO1FYf+i+leOMGZjeYfzQmB
6DN4HLDOSkka5MaaVvghBnAXS1KdET1PZXNVkM/KeILRkl/ZYicC1nM/FLiix++nEdtmTK4Rn/Eq
68prZE3Eq/fKneSElSNKf2gck3gZCpvzP+MMleDNQfAgsImk61VinEd/S3nwohC4RRwkiKgClgUX
Ej5Y+UlJF8bqlNEL8j2QZ4WfUc7t7sLWDAW1+mm1hUulQsadYq9gT9087U6G5mAaSinDPfhxLsWu
fq8r0+8T4JNbiRxXOgpG5abT28p/NRn4Gie+1eWtMBBA2W5Cc4gO2tecWS+fT6+qG6j3cb6iZeoq
Ft7IIsdlm/DNtuL6DAlkiI4r9aPDMwW65Hi5s7nehz8ppZ/LSNilnrParz2tZ5LfZ30wILbM0ryQ
sOtgbk6awWFKegdeZpI4DgYZST9ZunM0gYcaHdEBiz3dh5K2r4x3W30iRy9SZj/xGVGUjzN4twya
bjbHxbm8P/SXIig5Sna03bDgvz2gnZ87lk3mQwLZ3pJOTskD57t0CEtFN1oWSV/0krA2LMOTOsIk
H84Q/Y/zdJoDaHE1PmbodeZims5HmBEFQIRtqU3YfdTXdf00Wwmzb7C2CnSw2mvx5kp531B72/4L
F6Gy0Cyxd+Y40n3BVxjVY+U5EJNCQsj5G0Tdbirx/XSd0bO+E/RDbMHaS4BwsyLVjlyV0sNVbqqQ
v6qqDidFiC27Mx2YyxPz5fgVFdAhOJzxh9TchnuBWyft0q/qufL8MRFi1S9E0HEKMKxY6zS5QBOG
YXPPS1UrFyQbcWGNnA5UT98Z9xsGanZO9lKuWA3+583OsbfGWF7irN2ITJwQF4Zl1GjoGhuHlFKe
Y6cTnho7zYYOFjDCgkO8PN3tuSS+TprAFqFw6gxnYI3b5PJnoRqcRpRBiEA5fFVNkWo4Dz7o3fCV
FkH7FOkMVHjFweMMn2S+VHXaq3T9T6X2/Xe0cPNr58euTsJQs+WGGI1UXkkV6oGeubk+o/sriOhf
oZEEf1RWdrkwF/mfFWGlOmJLS6mxtV+H1rfqcdpF+1WkZpUfArelE6q1/mGO7tBvBm/2zgrLVaRc
GRm6oHFLmccIdDTy6eRgwrPPzCCAjpVKFwuA6WsjA2y9P3t73BSfIvIwHi8lhofySdzaALcnuU9F
TlCm1tfizPte0Lp6ufA7YoUdJz6ZBo5grq73a91kis0S8+DDpZYJcYuzsbUJBS35NRlvxh78PsRt
kn4/D/54bbZ6ImeSocUbCbUTtCnNNYiSZ8zPb1lxiiPmvybZCXPWy1vX8QjqnQJBngSGAcBZVAxP
yJorkX44k5dzjHX82k/DOVxRikDi4E74hedYqMI++kjf80KAeVzpdomsAvCQlJ4VD8bDDQgHpmYk
ztRyQrD5WIfBx+zlpipFJiXYf/Vj1+GQH14kNHOqyprCHMVpKdvgEHQweIPvVoxOkNh/Lcbr9pBA
M+pB+ARpzOI5irANRc8dyTzj30JPEal7qjWsV0BfWzHKfzlckCzFPiBoXmY2+DwCLmCicJsYMrrt
/7SoD7E4EqUVAcW1l99nXO2FGuFB/3R2WimxFdz0D3FeIeoSzWeIKXgVNUdUVqLgaTxZbyzaUwKI
mGLs/olJXXDeN1VdcLUJ6v5yQP1ECYfdPbVStLhcwJIvXsYRMSO34fH1q+sCA9ZKC3M7btueNJ5E
KaNOF9yKUzAQhPMzDZWDCJBIYG79NchcANPUSXAu7jKDCumkn2CWF+B4NQzPXCFaVKv9hHvhQ9ij
0IQLrm+HL7xJog7ajuhag9EVE6yacRQrKq59qJmsMh0gjBRCY3T1PaaYnADEp1OzDsIqRmZt0xrD
VPsapDNx9o5mf1nAIBXEeyj/c04s7hmnZ+FyhGvr+dvs2MFWkY0BZVId6QSG5OI8XzZn62zURDN6
5Fzs7pGHjCtxsS+GedCCKli2cnFCXAxpmcRr8nWnakkV5hBLAuQDzva+VyqU5dun0NBnRMd2qhAM
a9CpacA1G4Wh1swXMnNUKLaxZ2WCMQYwEVITZVfXYA+xPXLhosvTdI0+2DPuFORLb3ZOptZN0M72
KTIoyHAKRUQsPPMqf6hPWU98v2rP3ZW1OQzr6UrrNWhyQuBBPBBATBkIajnnIyKlFPVkfv1Q6pOT
Bjx8Tu0jGWIfFh5iCcCy28CvIPZHL1PPYrY1VPuPovIdAh0+hvyGMNVS3xPjhCXXSobwpPRYhh+x
CBEuKLyi523XwP4nPAObE3+o9NE7wudaaPJ7V1fwlvapu1gwnfg9ckv0Z+n6tci/J6+TtfC6HNO7
rhoZAyCG8P4UPRysk8osa7lvOlF1D8yJi0d5M2nEvyendDAKtzetfEaNvDU/RLLB4M0uQNqz5ftC
aj1dg5/QD8ftZD85Ie3pUmFCELIytEpo3da7/pwVserAfyzVgzPgXBplTmirGoHn1ZhSu6v1lBmo
yNPI+EMusFiJpsybK+NkzHsZGwTI7T8fKcWh7TlePtrxmYuhuhgj0wpFbsnBHt9T7+Yw4oI+vn3O
XmLQwpmQ8lNr4zvJSEI1S5Y0HM6UquTyKAUG0VqbIDweE/B1RV0mZbKqhpYXoCkbkUwAlUL1T/kG
SEXmVVSO/scYmewcp2O+sr9thvPfj2YW8d0P7KXycraTlaq4//EFvg7ye+u+5h9fx5BThl5yHn5I
yjdZnR1kchpRTdq8xqSrBvrE81jMS3yuOv9wOb38fq1ZaA+xzaXhaxkq8lVfNRFxYuXKbKAZ2Dsd
fDHUIIu1qWunHRFq5JJN8Lir29pL9FoEho6+ETSBdLuYS2CLf3MdVppAZoogFdM1SBDqrAi3lp/M
tvuayR3rs9P7SofWPkMs5VeQFkSXILn5TVBsvJtpQ/hipMyEiHthyS4r6bEYfF1s9GUt15qqzvoJ
YtB5X6JA6uu6NoL+5jS+MXS2SjbAUw7gmzacm5LPLPJjRZzKhOZ+wu0dJH/+l/o6kOBjdJGJmrBC
rQzjbLPgxwr9T4wHKa+yjfg4IkCOxb9eGUROlW79u845+sSRfiA22ksKl9oDem3zF8JuwH8d6aJd
WeA6zRVqmww7hSOjS0ioXcBvSTbDAxBM2FRbZO8EinpGjG9LKKLiXZDVPajGKZhf9PoplEn2GIKZ
pJ83TU2H36EH3LL3Dd3ADi9boodO9vyc8rR23qq8hiQiahEerIauegBqpuxfiz44zHXGO9ayr0Iz
2pPWMy9UWkkzdUk2tLF4eykB6kfUFf7EcmTRUWMalm+YOVSGLjY89WkzFNJ3NxVMGPt5lz3ornr8
63qtAtDTxWN0+T71yGUGuQKTlLr4IZ2acLF8vW/mMhQ34YrmLUDWcZ8cTjxwR+0davIwihQLsuRP
fMY4f8aiBGZov9/yCaxEGcwwOF9HeXX3S8RQKoSeJwG0RkjwgXEH8fWWshjJYEhwalnABGqMHR04
dSeGDOs0o09AC4HA6+9l+xmt0HLwQ1sUpPjXOcmP5awna9lG2qz8HDT/8YmaPYxmW+nd7fRKUj0b
KduvXezc7hgdLjEKaJdlRz6He0i3eNJ/Fr4SRn9PuPzZxhlYpwHzKjSyKyicPxTNKA8Q6+KD1vcw
ZiakZBTUJSzEgwyxKyLOV/tp2MbG8s4wooFgYhWB1xQOyVhsoLZ9CyNlcJZNF13QbdGWBtP7cxAr
ZaWrevZv4gfJ4T4HKaTKYUctcyi6FYPwktcWWEt/A1EYeLGrM89zhIO1hhnJC113Fn1yf5M7IhD8
LZ1M/hVj5poP2wc9PJJJGaEXfiAA6ZNy3yFpNNIqc0Sov9dgWtnMZn6ABpngt9SUAivWDs6XbDs7
NlCLy8f1wXzzmzKvCWV2MlfKBq7oSl+PgvRLaDGzUG3yoHr1YEx9BJ2h5DMtdinbyc0diy5Uvl7W
GJS98Jd2poWhd3H2HNdtlsNhioGooWIkE/mbsUTzDlGlnQOluZ2qcVW5ooq6u7u3dmhXEoSw/8Ly
fXSFh5T2rsNP4JJZBzJoEC1gki7IBUiMIYtjwAjBlC7d8xVdGDCSX8qEnllx7ndaO+lUBjxlCcf7
d0zEbdhveJ7JV3emkHkRcoIGYprePql1KCB3cfK2cZLVLlTJHWPL3Ho5wOC1gPEhMHRpWe8Vj+Qq
NL46hhPaYITT/QSglD7XcXkW8WinCTlSreBJDIEcDoZdDj9bJ05wPsniWSdn1JzWp+M8w2tnlEd3
f7KBalYLLI7OlFgJE993IVJVlYQOBcxjE6b/+6Um+C6LoNcqZ0qGIm17MyyQuvQfN6A+PH8E+VBi
V4iaT/uExMp0SrgbTD7oEeY774ifDtSX1/18IrtIsP6kqu7aecWXcKOSKaBiheq1J6Hfjxb8YAKM
8M3ZiZ4VAfdKvo+rYcYEPuoDwoTumuwkCk+Uxd85663cBKS4mUpspgWXoEW3uVJ+nPfrPEcNx78a
sH7RkBCc2wn33xaS0nnPzRNhtJkZ2iOWoIVuBHsi7bfkzHz7OQWa6LwT4rb7KTI57u8IyLG5dQiy
KfD6f1OKVOBQ1K3/1Qby5gBXoNbEsFukoMsBHulT5rraoE2kgFU7tIy5Wmz83G66CARd13kZXFJV
Po9SS4h0e06Ssm51kYNO32+awJ+hfWxWE5DS7vwC3QAt7Hx7JnN/l9hcCiKN1AzrOD1BLC/7gPSE
403zP7Q1ApsDchtmoandCEd1mvGcnRmbC0EvcnDhhwMhkek3Nisjn/I/yULnrQzYdTPgYTjJf6pf
odS/gAQR0WYkjDlqskvWEq5XO9E7tQ5lSzgW2Ar8UmFFUAhWEfP/w/IJSOlUGxp5clH2reO9NlnK
1iepPp+novcepgi8QnLd8Z9TrJsQPDdgZIoN1848uWaDMBpySqz/qj5y3hGVlIJbX+UCe8ekO0tx
ralrMy7uU0KcolniyDVEiYbXjYRpUhmkPXiSV4oVm9MVUjV6Do6/JVZnGzUrHOtviT3VFb35BILj
gUugrJ7OH40mg8iLI+g8vejLd7YgPl8Z86cPHiTTlGTDTph0tpKUiaWdKYLLK3FxwFiudQozewGM
Kq0DBJUxl/+Epjgw+O5sQA85MYl2+J6B2NMZQtJhFqBOf/bVmrH4iKQ39iSN5d4fw8f3yCKuPXVd
Po27qeupqHjTkKECPQgX19QzFTwOhHWUjjeCv+4j/f2PHx/KUTGuwAFGrl40C6xK+NmbEI+n9HkC
rIkl7rCZIPLCStvaX1SpIDamfzhHQF9Ox0MEN/lqH249xNa7bkSv8ukWQDIQQswIIXVhRNtH7hTw
LLYVtXMjO6IAMxKIJaMUbFTiImvHItjVDFZoktx7kQg0tQS0Kjr71EH5KZBbVgeO8IFYRq86eHwl
f2TIe/txFBVhYmVQ9ukIerEVK1nJfKjo4Ijw9MtlLixXdtmJYnrr8dF4ZuH0sPkYLOMgCSHwk4EZ
aGvK7dfz4v89/7dVXyTNx7DTRQ/nBDChNUrxYvyGKnnwk2K9M9LNBcDR0Q9xmlsaHpmVYwLhiVw3
viYNWppEQeJIEHSzf9uCunh5YZEmoQaNC8BbnaVK8q2tMaD+34LwSUop6yKwFb9DQyGKjPptWvR9
Wn8B68fgEFW9ZULh2QyRmEtSyYxZo0SDFfIBk5RLbaBtZSUmQnkcPjd0GCBPq+y6EpO5DDW8OKcQ
QT/vZ2g2m+JYPTdQFBbAML/7K6PD/Cz9op6RDNp5HIZMTpI+xStEATqq0LOm069HBaCu3zuc/wIr
2indaOOeU9j0MJ3Fcvo4haccWy4tFFwXqt0cfmTxlWEx95p/LqqPX8Cd4FzDL3o4+91rCwTwdM6x
aPdom1A6U99/fk/xMmDVQgZEnt+xX1MpB/pSpahig4DNdWCSdtKou7YnlQ5N3b0Wjfl3pD8TUclT
fI8tcYowB8dLiV4Srr5Lu7I5AmAhssWzFreWorhf00NoDor3S7v+PBWH3m26sfGjS/7j76Q+0Kdz
/3C3c2//+IiV78Et4BddJBmNFebpUp+Qxgqox6HVjUjSFv33mR9pUzDvZAKjPdZHCUr4Jcx8wVUq
X+2hY+lGJVULA/THPXPORQm9ffEQb9DngnkGntdtoMfnnR5GN6Dut3gznpApNPAOv0VJ/yvqJRGl
INFuNNIZCYJkosm0F72GucGc+qUIFvVedGch3403dDyU+fvudfwKMFj0gQKCtcCiWCD/SbZeHlNm
FxKf67KsU+e0T6iW2Bk7/McRb0KkfQgzR1EQicfOa+e8QLL7BPwNLiUjfmqeDGrlP0SB7n1r8tWx
ulreIncBy506yL4zZr0vNFU4cRtujTu+HSjqm7n4WDWKwdp7zaamxtoq6ohnhUsFjXVb2eF8zqT0
zimDBbto/fytyYMSUeTIb6Yne+gsXaoXL0NPeTqE+COw5d1LXkcwuX2nIi6eSsdP9p/FbvKwXpBW
8Ct/femfYvOLVBFj4YYpuZLnYiLbQUWz+2d6CNm+X/tyID381HJq+c7Df1GFWMSpgOQZ9T1Xx3z6
6cWVTZzDRYSGn766TdRsFZ2MU/m2/p2jFhcRf+8hunVIkYc6koFb1I6eZ1x7pv9oiGHre04HIDkb
ghwA325htwYns9A5m/83wt2wi3JKbiq4XUTtsPMJGvRP3Qhrp3Hc5Z8LAPy6Sedg8PYhjQFsNC3Y
gx/8kqSyQRZuaz4UMTQ/3fMyuexZevpk4mQth+amv3ZOMOMkbM6udh0MjAoJwrfOoXgDtw5JeCQ1
YN3NmNfzlKOdyYOunzLG3Sq+uZtrsqtDXbhAO5ajIHvgb+LZjkhhDxzhnlO9GvssSx+JQ7TPMxCw
rOT3ZMmtsQP6QkHxmn1RV2BmBT3MDjKG+364ex0SfRgJri/1fV+lUdFVAgRdMw90D3r3KdWDQ8Cy
QjTPi/GGsxslT380SHw979UoLpalLN0PjfZdE3SbkXxhG0hkO7JvEJ8BW7v/Ig95C1BGHm7YLRXR
FVpHviaEBlW1q8dJWfao9rHxPDDoOapP1Yng45WneJp3eaQZPECRXICKsirCMN5aLE69TW4aDx5V
xT3t3I0Pw89ATeNeqyINxKYy4SJgjWbf7TN4VEX0IqY5oyBZ3pUieTmfAQkhqw0Mid56ICXsR1Pq
g+91b9wPCMC7r/8QJvdjGbIZ5dy+sNPGj89iO/PhA4G8AFokAAmadz2Nf1NUFvfP8myYbUObaLiE
QosuF5s/+4HLTB9JFFgIe/eAPHYKiGsKZpDtkCeyUIZVz2mkvBd8VgbbSPQeZUEYvYKjaVEYGzKZ
lQso2U7ddH/jOSBXE0jJCr9SSTFPscKw1vjF4MhLuEPKCOuac1h97btADAfStP8pzPPVT60Cy6iE
fGmC0j5UcKhxPA2UhNySR5PS8uYIjrgyTR3UgJvq3D4EfFyvC24i/3oEmjfY0Lur3IfR3uFMd0MA
ODxi/e2fBlvvzQF78AfUYO7plO7/+VT2cX28rGphf2WKzw+CrIsBEIFBZ/Fbhcg3XcG8BDb0gyqK
i8zA/hg7uSFKt0rgTQphLv5MIdsNjfwpGkOofop5sI6l4JbmMRaI2fNPV2TV6VPxv2NsWVGBvLVv
CAokKdy5RekAPdHJBBOjoMrg9TCb+qL7Fv/A0wJ8Uj/Qr+hMNSOBHbAzaWfrE7Sdle0mko7FB2Rg
7/13PHvmIrtpCRZRRU7/bj+042PVgABKTs3kD9pJuTQIwZvY+KrYkwVg5KGGPhL5Mxy2zmLz2xCh
2w5GZVqdZRm2REv9N1TfOor9ciFEPJED2VyRNEHozaAhciCVytrkA2XRAZVTdQfx1YaUkxDvT4Yp
hv5HJDX7MEmQVxWMLsoBoBP2PoU68+S24o7lrUOLtSn2HOnX3oGlsmYfOkGhMl7qSMYKFMUafrYK
QdXPvJKchnl4UD2ANs/1LR4oJNPzHopbWu1YR5k0HaE8mBdJYvC8b/yVdkCvM/QFaTG+nctr1qwR
GMXkNrhoyM8xi83Sl8eUY/Ze4Y72z7RzWcRatNL18YL7kqcAPtUKrrkUymWs0MfGlJapObr9/kFa
xAtO8q2cL+NwhegnSWYa3h927WIw+vt+QbvD2tBPRZKIU9BlEmvKeIyd+eap7GlDX3WM+iMgYh7x
Cu44clo9ErtHvgHORart0dbho/jz9PYUMIOuqB0fd3OeroUmFNSqn4AF3DxjsU3RtFIzjMSIKs6n
OucvyHVGd916oSs3JoxGCkSPskPKD83ysLyCLoCAqHFgPCG8trUl3iQkaatOqtFd1jCvk6oUPb7B
jUu84AtxKgeMFCgqBOnYbnxmdF7LXVzRlDpwv00D2J+GAA3BHamH780tBtQlhjXLb1CxHPg0sY3Z
n0/wuf8RO/8I9NpZ0vRYO1k5j6NC0uIrHnOvW1LaS6s/i3YHckJKbAe5uNtUUtqxINFE8gg3COBJ
ZmTssril9OucMqBfwJadR88/AuU+WOwMVv80bP7Ny1E1Zt2h4iAOpqc9VB/PqHSWtAs057LxstSs
bqPlsihKLCQFS6tfNS/9sEgFRXPjVv0PgwCnG0wwvFPsfJgtGPxQHgQV3c5tBDg8NtYOfvyAPEmm
iNHjqX/quzk9Rf5eEFii9bLz7bYc2A5YNnqWw10g5RlvaN/RlLETrZkF51P5iMGOKHaSkmREhTK0
K9UHCxYn+sGoZ8JyzPSmUk8Sln/bmDcBKUC6EHTAl4mtU9QmrtStfLmkLaJzr8KlyPOyxL4Q8vS3
rL1mU1UUMZrGNN/Tt4Rq9nZ4gdGvJQIwDc8+PmBbPegKokLZoXfjRkoTTvMJscy06t2HdfpuNoGp
ZBby9glgfCyvTA7wjCSSNlxCtZLTm6UorZRaFq9uG3tTyWhB68Ndxix5LI5SrK87Wzwv+Rc6zK7O
gSdVY0Gdf31IH4pRoVH1bkUXrUHoAwfCegB2CstdoATAk2FR82URAdHivq2JdOJLZ/h98IgH+Lt8
ptt4bAg1pMONwtAAm2CoOyzdeWuCDf56E7PG37aRwB1jmrCWZCL+2OzuBbxk0OPakdPiQFCBzDA0
y7XIwNsrGZs5lkVpfjshOjtiweolkitCw0IN+YGYDgjS+1nIxdan01GoUbijt37rZOMCppPulBSH
UnMzkEZfcPKwU86pcbW4t8ZNmLBYXyaU+5Am/gs8QV5Y5pasufAItS2s1yzI2rbxMpRhJ5O2Lu08
p3bo2eJDasffgBMT135vdLhj9GzxgKqypSMwlT/8LCGnRI48jWCRoIN1vmJyv+fbwiDm7PB2KglQ
ykms5Bki88dEj9EHCen++wvHvfIBQLPWYyVJE5pZDDQrhR0AD57uaSLNVRfMFqpBuw/vfr0HhDg0
5HnXAhKBoNEg+x0bO1yq/yTz0+h7G9bJQ0K6Oz0Loj7ywywNeRfmD8IjV1s5p3TncRuNhlxJ+QAc
NNybbRHpDWLcjYsyvU157sYpBbRT6/WFglsPhDdVlkx2Gio6xxlk10WBYujVl2LxfOnM2u7Gl7G+
rDEr3btpevBx7SN46D/I4fGbZihYtQCZIMco/unI09P6gAZLE6loVVZ1N29nX2pQ1bFeBUOo2Wwc
DjlA5D3V5tKuMiF9M5g96BZ82DYC5WsNd7lonnODLorqoXRR56BtRa61CUt8fr3wq4TCelRzb7Mz
HENwHHFSyR0hii5ChMxAASm9uno6nWZkkPWhvJDGVs1NBC7K1qszwsmFvueJ5Efh4EsK8oBJCCzn
XRAfAtwFODRlPrxxnLZL0JyCH0GmPBtovnFZQfkUMZ0Lx4rJ1RFBVbLtyj3ZfsMdjiYwTzbSjAvf
A0GXF67ANuSXUY5khJlxTH5A8I2AG1z8NlABIHQmpEmV6KNdpnTbl84GCZYHCnYS3fjuSkUNZ4Bu
pVL1KrUtn7h8Y7203/2n3LmIzi0asKwveKtvXPyCGBv7XdvIzeJlPNMX8V5qTu6YKfpQ3VGEH8Aq
uHKeuO+ASlkKxnLWw8vXgdgNRaS763la7Ue8Xw4Pop3RjGE4NWMWqyfou4H1naZKuz5zD9k2qMT/
rnjt5eudLocHucfkLo5T2nVtIF6OCgXPJIBLLTj3G66qxJJ9oMrTE9Mj8+Tmf+Yyz5GHivEu8gPC
Q3HNI5NU0u6OslX2ifrk4havewM4vnjiirwljSTIkwFU88pkvGSZMPmGd6w6+ThL7mck+tNoVlL6
J/AgDewGmgbpF7tEEZaGDKTOnh6IeTszsIeCjfJvxMrTruc0Kk1yeRZPuF0Epmn0J27HPMRc95tk
mf2r5/kESqokmU1R5RJJVLjFFDUdoYmsu6+lOzqlnMQ67FhxR2dDyHlyGLcvQfL2V+7YsccKWSBa
NHZ6oKgLsbWN6SRl/ALuey4yePzUIFt3rNnQBaSvCDpabzM9xIAtK8d4DBnmODTJ5COqs/qiDwfk
JJFK3T/Mc/Jkv9AHxQxyuubEdwb24T8HN0Xhf9q+hxSRIGHOJHQh/0AHF3NWnOJtSxN6aAkmLaHR
j+kEfHj8qBVOEG8aU5HxKOXzN5ckSPu5V2MUcc9l3/Nfe8Vm8yiH1I4HP3I8PZxdoeU1uRvSrzS1
/5LVEH/cNEA9hsotQChMvk/QJqGT7onUCxyM7zg6r0fnFzvHNwfNR8hJV0lpdENh5eUPRuJ2gdFW
+0GJg9Jv1fJ6aVNNvyqK+arOHcuImmMExxY8HKf7I38fzbmbExW3vefW681Z6doreFgallSVhE6t
Xuon//gk8v5mFt78pRnDxeTtdIRPDYPADvGVA8ZWLG+mS/ObWOX2xEnCv+pVxa7eXYfwhu4ByFym
63UaOFisO0BBsfnBPL01YE74kuKwKgWLSgIoGrTDhbgTpFUFB16UKnshAvi8N313+N7rutCB3reX
Zi6DeQgOjRq7QzGMX12X0oAj0fk3PS1JZGruJaxSO7r45wSvXS4PcFQ3ITyrQh+Sm5QOHzj/3n6f
WoJawG4Pm1diQLogV/5Itc2iWNtRAWZ6BQEYIfoYrGLI7asqD9mtcMM7TNRpllfDIfUR/X6wnliH
Op7iIzo3mJcKI/FtufEiFIqDibqvYqnDVwquF6hw8fzY1EZBKSaH26JG2X8KIkZcIYVGiS2Mz7qd
50nHbNfrV1tTqcOMe+DgKOZJmMnRcVNfoql2pRBI4NjNmHrtyBl61hEIVmXeH5YwqR87TUPgNtGi
dAaAWsDIp9SzijVgaUQFGotGlYTj4BjY/xfugwwbuQFZDWvqYB46gooC/sDW2UhbjQToIXctvieo
z6YqutUteGMbgYxNYHysDCgZ/RCCJv2w64vNS2pXq7ZdkGIykEIM5wr1NOjzWcPbkgXJFNG7oC0i
tWXyOoSuMwmxXJnVoQgF0gV600355LDr99njkp2792HCPDegoWcgKhO2Jm0mRtlIJPVmzYCQqEdv
AFqtVlbhtDxJwlgeo/T1JumB1tB1/g7LDaBYISIZnoEMaxgxETKrMfL6nq0JFD1LX+t81dW70JVv
/K36vCcAZu88TGjgBJcVCOPGFrC0jv20NWH6Gffzs4gAC+sYqujNwqy1uJeHp315ohXUumYvmzP9
P8dq/VCIbSBaiXJ7qB5YDsggg6P/bJVAspSF587tnV134rfcxLxR26amYivDX9UUIjkSar50eceN
jitIE2EAH1r6u/RWIbm8eeQJHTy+Y/FuFgzvFBk42lA+Bf+Sfz9uCYK4twZrg7KJJrNf/qHlOnwi
lmeC22c+GcxsRTOdHsbOhuJ8/FDl/sWylzZxS0HKQHMJJMHLLCsRxP7emHC0pcSXSNHERv1YuNU3
o1xZIBe53b3SaIzoRdJNfVXFvuOieIOC7RZYHJf/rt3QyxznGNjFURZktRJE5/ax+7kyfMtZ3HNu
uVWjGzIpl/wU3oD7yx7R5PXHYPfPlcikvxzBmw28G/PuHe64mMzYU6CoAsq2osLfgiNxDWNHKgF5
hfhTlTyxaYB7sGOe6TC6MI0GKHH4On6GmmwUp2fduYWKjojWZJB3C/PdNpRi2SnJ/wPGjEu8ezOG
NJm/gv6vkzz2nF9NFKxViZtp2S0PZHLNsjmpgLd0a7+kJ72hJ/j8PfU0AgUi6AI0enCdhU6V1z33
IfgxaGOUMFwohkGM/rtxU02YVUdBoS0YJ9251aBsp5vS0E1xO+W4emjt4sL9fPSh/DAIPRRP7rD8
ViZrGGYgi5oTCOtB2n+q/pdgswzOkHKUmCDyonmGJGI8D12OwLostARz1Qw/yRpQktizxOBy79wZ
FxvBXzaNsA/lwlUsnlKuDGj3Sv9UgY+FkygFuMBSO6uAbmIRR/g4bK2OPogAqdxum6jIdvn2KZ0x
9upZJWJvSNDpH8Bnu2NptiIH8oPE6ZQOmNNtupZZfuuUw57OQ5rqReX0Cv+WfLkQc3p+aL3X8jf0
LOHGJ4nIVs+BbDqPOW9bpsPk7D5eh9QlhTeDlwDRRwX1qrnAZ42+OrjmzinHfG8SyIWoKFKQ1XvZ
+d7iUG529ocnZ9tQjNC5nYLQH5ZWEx44gO2wZz08G36B9ohk7UzDYXgvvSu/0GMpquKihBv/bs02
3Ae8zJLaEctAMtlZOa6wtRNsAMoNvuImjfUbTaTMD7/s9OHWH02Dy+/rWdEQYReNhpFRPDEpHMgn
6/ukqCaTqyeiYQ0YJT35gGCIRMwVZeglpaHcHvFkSMVR+fWzKFsTiuzFxI2vXbQgO/6g7mCOT0y/
KfWhRSd85GUsQm7wgJxThlzrJWqlrhtIassjkLvFsRE8iGkS5GY7VKy7Ks1QAjB2m/aKOsZQk3jY
XgmsHyTHFQKHH0EemgK4/Jk1/oaZ4mQMfEEvCE+S4QUUdA1hXl1k1PDs9K8ryF+dhEGoo8vfb+Us
aOywyYclVI0rmel5R2rFwtR9kLkvY31w1MkQOUDZ4LrTJlmi11hA/WpM7tFdueVPiVZf90FZyBnP
JEblfZGyRz9tZTKJ/Sj7/ZmyxFtAVV5vdhzKfqRqwi3yEUQ6UXI5Y1ytV4N6mBkS4PJjmUMKNJ3p
ZI+qk/opSICv8kxQ8W+fq9JyCL/5Ew7dqmb2ZeOhWB2D5jMgCaGpJ2ixGbk9oRoXOJ/te0Yz4pON
/2v81Vl+94NGde8jYo9pZm6XGc2c61xs/410chlA4Z1QB/NvBEfXjcGycsPtPTOH0YrXTtqXV41L
Tpl4vPGCIRhdbCntR8T66+x7vOO+stE6ULeMkWF/n/SlbJIAZ3hzv6SDJZY5cVFEWahisT2ajdCP
pT9V+5dYeqLQ1LnrUgglkVABqUmCaoPs4W4Fk1hWgN5bYkMmAQxMKxF3B6u4KrmZQY7EO79R3j+s
3ckNC/Sq6fChdOhm1WZ7AIv2tHecVPbiWJP0P1z00r6DFXemVaOwWO80LNoC/xxiyPKNFArS25RQ
G9SCwz1awX3yzVPmVBA73IJJ9F6Lk+inNLo2sSwvDBYIoCLjn0gLElSfv0hnap7Hw75dKRowIAkT
/2oU6tDxgX5AE9Xpitiv+fMWo6dG2ilebssRPk6OnYeE/oReGjCTaVNbc+NVBaO0e/LolEvunHIF
F4EukJ7GDYPF46GhTgIg+8kstioKc4D6eWxttujBrWr+3QEdRmutul9ZKnvmRAPdygKrR8Se4V5+
tfpfv4MF1ghJ2SAvOtg/izBpjRMbU8HX/vPEVMeINPEiMsILmQrWUZtVvyzwXsNbOvr4ob8Wa4tJ
LHMRsW1AXD2ps4mYnApXkMqZaIM1vvYUk0SV7fGtj0KEHlP31wy0SDhE2x92ZTkQKcC/IbCjatc7
Qk0Zpri97sx1HHtYFjpRqWJ5MLPhQQqUJO+JUFULonT02SdJ4R19GNrDdHwAVX/TH0mieX6Qorlk
noz/KvoZ823GvewXTIF0AnL6UkWc5dma/eVyrKAzhjUA5Fo7gAPZVzurCz73OirtpUChk8oZXfgW
uTot/rSKEokzFoEwAvj7Gx6W7wdwxv7Z5H40l5hNul+s0tDycLmFiija1kLz2wwq5trPRlWwGUc2
SPOwFVdG35rEC0Kot/Q97JYC3/6KKMZvxdxSDyrYkVX1yHJgbHkwhc1A3GarUBGuFdn11ffVGERH
8FVnMN/e2Z0KHo3DGrD+poWXHwUl3Gj6wmhqLBgGcfCJ9++iUS75jnkYPXyr47GFz3DM6ZCDzGeg
rWZ5d7RS7jOMERacOoWQupt8hwuhQKW04KjQuzgYQ2Xd6gig87YblOxYXdcXVsloxte9i8Qf+8/m
mFqe7ld34OTD9EnCTR2mBdGlCh0EP1XtuILiJI4svbf0AohaMEZhRS7US6SnygbIbxSlTlGnCWIK
885/JPLLjQnHxBp+V5k6sZVvFY4ZGu5Sd7rsU16hgG2YAXsMtUQD6+kmUnX2jHir+l6sGS6Y3xKA
Fhdnswd41BYgvk8llpktzRfIUDzqZ7iuxV15WD9DPV8f0mWZyrJARDCIOTCGOn0Ewtf/jHgZuno9
miBtkPCZqqxymXw66ogjTrbeViikknMj9FYrJS4NNNZY15rP88OeD8ycXvRyw6FwL1vExrDICDls
Yw4ziljq4ZshzcFjnQY2LaKIStVw+hWqFVfoIhvurvmtajvlPl2yAE3fObX57YD8C3a4VK2w4s4e
bZJbqOdG+hz3quptMmaIuLqWwbfdGgcxEbupOPPWxl2U1M6gLxwWyOox2WWuhFQTOeoqnYRidurC
Bu3srejYZNoT4U3xsiiqsKffRVEJtNVAz6kq/04pjoXmVQU7tQnv+DgPAn5RdhvCQcLBzH1LHEa2
PZ2QaO6rCy31pdbeKPBocZWMIrHvHJsRtn9k7vdtxJLUY9FJCHeHAhtVxcMtoUoF7NlKvZDIzW9s
LIah5cacEcBUdUAAjOEjMEQr64IWQpXw0/rbNYBOaIKzFtAKQ8H//LLz7GKcH+uzuwrprOYXKONX
mQ/VQotfGZL6c4vcLVGkUKYb7PwhLg/lJfJvgfzthbD8UqBSsswqlHdtr22vg6+bYqrCkg3dtoAg
XHO/kvxGb55oMsOVBUqQpRVc5bd68QAogXak6uMblyRZkFihV3lAV/3+i7yk8bqQUos5ZgkeM8ak
YOz0dTLZxgDpnH0ded8a1jT/oRmkWUmn8EzrdWbqnRpkogm4kxscWjo+1MGi8Tsn8pb/l74yJDPx
/0MkdquduKZX1h9wFL3XaesXkjKifsoRZo5VUAo1MY/4WmGuICs8hxb8YcKlXie+ZvVrLf4yPdIt
gGaSaRC++25FfiYTGFMbvy+7wlhOb+xoZkgiR8rScuusu6D0n9FdchjgaSa0wU0Rw6Lwdj0S7dSq
yf5dqcP9zg5OAimUM62OJPbtGqARrOc1QCWRHdA1pxXMJ+ZQakhrDDFvFvIwSLHKVYcnkuzfsDX3
KF4dD+5Vs/QrIefT83ceQjMuxVsrasGhNQeoELMcFkVzZqev3CvDH3orHzSV+/+N967pnYw607K+
ASNGUxHG4lrYXEZdgfpF2OW0gaBqtBs0+xfxxJ6Xf/OktV4y6xShfHjwe5J4RHDknKrLqUjo/a/v
nAIwILzAol7eCgY8NpuXuDyxYxbrSQXEwgqZvXq1Ni/YgdQL+FvviwUyTK687GCBiKQbjsbUNDy1
Tk6IGwjtxnm1QiUM8Y18papeaTsk3HYoMJPbUAH4HZXXNlGupwNapOCwHBKaihO/fLspRqg59rKD
e3hiyze6/NO3fMdvD0mWfPxpP75a2AwqnbCaQPmnEPUZWf7L3jeqc4qLekC8VijpafHOAbmnY2Cw
NZaYgZwooWk8bi2hguJeRrnP/Alijit3sNepbaWQKT66mtoX7uY3QHlWII6ejrx2hGK/Ifgc9NTZ
JuedaCu1JaXYdH0uKKwKWHDsib0IooNu+IoPWxkZNWzCNWvLYh37jJfmqAzOJvBgTbPW/z+K9UvS
IW+u/9IXYYvhL9XSggyzfwzmeW8LdHHYoTp90dAYB0E1pQ9868PO7gJFX3kpDWU/bdGzT8nt3l7N
wGsWc+Kzfm6DCr6hEUotdTLtni3015lDTB2bVR4fQwa9v0DSQO1WuT0qwyo2rW/nZqjtkZYgvLnq
FaBTCKTl4ArwKeHBGLwy+1yzR2BiqUBzXP2LKtrBESHNUOtP2awG49u9WN0dJv0Yo5HZlMgSDKjF
6SJ/aLyDnF0FQJBdogdmXeNpYZ8py9o+dfF8FqQ0k66E748vfzgZG/T1piWZbVvJW3JkIShUkRZ+
wZfRcu+LDUiD3M+bLr8ArjpH3XYzlyk1EdYdD2vUoOmIM0DLHzfWB4PyOvEHoyO2mjozm/+nUtt6
875FPnfmmzoV/zc9pmyczdcTE5TQ0pviXvunaiiDOORtlD5Qgiow+DEGKmNaBrDTdnpX5JnHiEWG
5mArPfoyGMynTgAH8MyfVcJALQSUAqzlgBtsWtqnWBxufqemrVarxrtKM2xta4LmXiRyvlhEzZA7
9EC4sY2+055sOl33IB53hvqC40wrYX14/Op9Fn3BbQqErCJ7CJaw1CVlZ8V1taF+Mg75OF3MuREY
5IP+FhxR5L4TCn190kA88C+zc0ynMvi8Fu3tuY6wJbzo/vSohvnYM91mpBlRNHjOuk2jwepD80WS
qJmaMl+ThWhr3HHWS0rqF/o2gxIW7Xe39E4I3UujKwqAzLS88LVZP3oNEnYKeRcWZ2rgXbjRbWUZ
ZF5tFMQn1Aetq/D840iNZ5mBKnAO0DBhz0/yEGydhLkSVGPUw229oCscDR5VQgzL8DRuls5EiDoP
dTHk2A5ui5nlYpYuGaknBrW6zpiAipmL00eVrWjn4zlUlNX2pOvpREEvFVV9uHuFuUBvZTDEGiWt
O7YTY+kgf6uu9bc8mlm6h6/cDweNy2FOhiHsymRim2/3E1eBPZByQvHVW0jXgtEdK3OIbyRULWOT
5Qb7CZZQkdMLDChp0WbeFY0dezyn8YWWbShkh+v9IdNe5IkefDQFMpAQnaNimv8od+QBlbr/UE0j
arp2x1eeIUQzBCVBcbbmifSgvhpJqYumuSeBUKVbvFM2KvGlQ1UEsEUuJxinK3o3wYZVG5dB4+FN
u2cZIkLf/GOo/iWm1+/c/TI2TNvZ1h1RdNxjPROY1bc8CEh5USqwIIqb+vMeqQfMCHEMuPT2Vgo/
JFrj8oD4kH0BCqet6WXFeY1nncsRoX1MQdopELR/ARTLH/DHuGHvZdVogyXVp/hFjyG9FBnxlqFg
aX1ECjXRy92cHPh8fo9uFT53ooLX9vIvcSVqXmh4bVKfFgqpgZn20iQE63lsmHZgjxRJgSo3Or/E
O3pUDEmY5grsJrN5duMIQmy+8udCZ6be+7xpzzLU3iCkoEZHFPtW61hHsgKDtguSAg7XTqjNRyG9
I4ufPLIYVEuxnJ9/CACg4UV1CORJre45/ug710XeUurU68o3VLC9AifzjtT5tSx348uxioD71rWt
eXqlSSEGTal8wWY9htjpqYOr8PLCcUk/HPllaqXs+hTMkbY0y/zgZfztERJx2++fHG84BEuJh67v
2tbWFOwmwLb9YiSm4K9e68UsvCWTCb+4g8wMsfKBNE74+2Gcyxb5z82azxVcGoBW1s0/CwcV2B32
u5WuhKyY+uB2rYsmDbo5GPw60JNrq6rSkw/KEpsGWkjgrktCEhBu8TRSX9f2EweSvU2cR3ONCjGX
fuduajm3l7fk9ntNBWMZcCKxSfM7fXTTN//3Ar+L7cIOIg608GP/3pTHfu+VuCeu2if35lNCVQIz
dgQiVn04ldswesHAJbrtnRiy1WALvfm+JBBEz4xLUJar1Eub+Hyqbc5mUkLd4SmAOSBdfMPIPvNk
jnp0CcRQN6IzRJ593Fsw7adTYcTivks26CHgxM0wXWp3PwfX1vaCxDOU5scYcTWsSeCbjYadefk9
uvJgnqET5ZnZSE4p5C3fxm0z45QK3m4izx8o9+ojsk75Wffas+RcSSDWS2v77x/8laKjIx1jjjHT
koGHM7n513W5tPgKVlt84L9t4j1caHpLWJGvVymZ8W+zdfg9sBUniq1eJR41gBlvHH9auBDS3T2U
D+0VwT06zkAzoeqrgaMLlKXsVPXM47/pc1GguBHfalmhMjOmmmovLTHLumnfjfiKlzmYqdsRGiMI
jhGsus0xbSfBOZ6eKBojYOYafJj4WmED6RRUKkF87rVGkoyJ0sRBkN3euIabwqCOJSr8PelFrVO+
ueufCfSPF0XzrVoOCDNQCAFUJPCKbkedqNrQJmVCIEMBPvAV+X4FFF9KTkKSE7QJDFGFstPqqCeA
Luwzd/kdr50BMfONsiU2F9h+3n//D2AaVoyDW5ojEAoSmDtVfr+XXoeDagm83JsGXzhZbhjUzs76
51d59QsLfnufPSzhOwILP2lB0XXnxzXC6oQyJ4Kze5oHEedorYkXjiJr9zsPlv11UJJ/t4g5ca5/
4avqAmmYU4zTcwQFrdPzJySEY9hg0N9rShyHdgrRirLAbhoHXyoKdxrtRuZjIT5HfFqBu8blxdcI
gZ3Q0q5i0UAgDtjySQn+Q4lCbFplx0MdOo4bkGNN9yEwGBXjrePhLU0UkU7Laf1297nO8qeQyEJy
Y9y1np1NHhruecpuMfEmxBKC5kZuzEjyjkre7G+tnFM1ziNH4VNA3S7xYLwZdIL4JgfitL/x9VNx
EQE23+M/Sw3kVHjoiRlAHGuYHR+hQIIAPaG+UDRCSM9XnnhCG17sqpc4PUOa3HVvxiQOQip0pZCA
9F1OswW5IsUvahV3WvTgilDTZB9Q6RC29Xcg2EEFzTYOWiOjSWv3hMF2oQb8RjFYY7hIMB2qjCpg
UxMyj58x87CTLCVEwNs4awFzvr59ESF0lmyYoFfUWaC49Obg/ct29d315NVOe3apusOg+Da/DY+l
B0NkSbB5gLu8UvwK8ZtC3LwuUjWRdmXhdjgzeNnB2zCBpUCyx4zCVy1PVKhcCPONt5xK0WvpA59w
g1/64ks6qQ60ynygsBeKRz4iq88zfhasaUHr6Nl277NxsEZBQevjh+CzOjp50o9wusLjbIsO8rdy
3TrGbrhr0IQXhbBe3a9ysfh1ehbsW8PgCinrqR/tzBGJnGzbnnbloSrP+FYNEceuZUNBV4V2yrk8
u1dC8jL+SkkoC3GuGyTvcna3OpklaQVapgK2E3po1ZGCkpUVHst/9t0rJhd1+jqouk/5lLeZrA1t
TBLKkNX5vCAb+qzaiXzjVE4dUnycDAjD3OwRGhT7CCXjgnNQgyWZNLhiadtz6uAMWI76tsflP55A
BP4CABMWytkOnQ0FjNjc0fUl7CtfZf1C3cuhBykJ1DfK8cga+K7ZawbcyjPO1PUS0H4bTfp2RMCs
tVuCbwA7fIOkIyFlWMX566Qo3ykdTa87S/7yVO9jVDe0ydEQN6Z/BTWE8W0VID4fpSS16b23+U1U
ICARNAdiiYW25q7VC4Ral7dTGwAclvnXEQNdeFiUjNG1yp0lPFPTpHjDpE1PDQhD0SAbrQQDs71a
+P5Abm7q3BKRk/FsZ4leAQXbJOeUdE5mfomY7PxyI2VWMug7w1ARPse2rKCjL9w3ffNbM9ztt/NY
tJ8fU9PFiQkZWDGeCQD4W647VC2GzzESK9+v1jrl9PKpgLEBtDnsapyVTHy25LbMLKjug4NooiI9
mORlyEArl7GP+XsBTEfFIcJ6NEYbi6fZGe+TKV/Ggj567ug1GBbtFPLdvwk9cih2TDqEi7b5KH7R
0789723GgdTnvtV+pzJIHoyk1IZzndTNhviKY9BSwK9kE9eCPnPsGN+33SZygFSNARapql8qylJ3
IAgp2/gDwPmctM/iPo7kimeuiSFGWkV+JWU6EGSHRBZxKaQGpLwcnXej8av8Z6Er/ARhD91Ozs+7
A8H51NL/gGHb1qHmjPGpP+BK8Dl7zVFmLqx22anz8TXYGvmQ8Lb8osWbXlv52FXNjIkpjfhx0QSX
KLjYwhGQNxJdPx5gk4PTDEq1fjwbVy717qK48pfHF1uP+D8smGWI8Dt/AHJnUB8Ku5MyV95b8aro
3jsvIOSjHmyQKJgnqvhcrjxce1O15s+fC5PheCFPhbtkzIv8D+sT5DbTmob1CHnRX5wAb9oBstyn
n38Rt772KVb5bOInJ0bc2aAGLHoLymO6V//FqKKcn6nmM61aWsuFhVh7XgpJjiJZT2E7m9293+dW
ylFyNTOnojV0T/NkV6E+4uAxszV2VBDXmDFeIbTzWXqYiWubOSEoA6AaD4SIcwSikqgkI5AnFf7l
CtkFiWpN8OayKpnLlkkTTHjiJEc0h5p6sVX2RsDRvTN+ttYuwOLhzlMIUYxn81CJxsjKDJ9ZLyFd
AHBI4zJh+/MkKsGrsvHx/vWo25W4DZXPl8De7ZfTp7wyBjVmm+D6QyHrD57lFvu+Azy6+Pdw4M6H
osWdgXPGUU1wynrgvvUSbixpbFJxJwVBsu58zyfO8UjHf2jtVfgJG4hAL8W3Aq7M/neoOaYiyTnd
cOYXVgFNcZkVNDnSbmqQVyj+gUgCu3CZPZhhMtdGL7z3PjaL0LGy6An4SnKdJfmT4c1pONdrkShv
K0lISil6Hmc02tL4eAR/0y4QLQ0GJKJyhS+ujxeWkKmRoYY0l5AdR/pNu1Heixpphr7HY3zYLA97
CTjNq2Tpfejl+VMjV/MDMPAZA+IUYqXznzA/5b0vKBsRko5KJUkgst/QhpCt3txgZHYYjQ1FUzly
785fLNSiEdyV527GMxvdZSZYgblHFdos7SAPCZSJPknKBprCJa0A0Nhr7CVjJXqBzahofRVmE9wc
ZAgBfYzbJEEiqq0sQ/VerMvslkMdoK0JRadF2BPD+CHpQehzWz/QkIw6wLsIfOGQ1jmza0Paznrz
0feumkfDqQaXi/7Wacr/xG5VuDxFLgyg5kby74XN7m4K+OzwyUDQBmqTfFgxPSbVw+ZyhzNoTcgn
ukmVcwZVcOhHD4VYo+nWozn4reAkaI9f5CT+XnJfaqhdhz97CzRK2h2E8Wue2fEqsB42xinXeflX
qBbqRy5aDRRJhm5MDpIMZPk8GBSA4dS6S9qbOY5EaJVroW2vigJNyEMSxhMVS2JtNzuyBaE+7vSE
j2+cjKu1G9+UY2SvjjHssH4NFJOqYsYPrxPaXwRzEWqqJvdAdXxIrQL+bPMu9DfwttGNfgB5yHsA
kr7tt38aBRKsakKhTdx5jfe350e+wOz4TXEiefLffugOfC73GV56Ps3yncgw3cj/gJEDnWNmUHPx
a561oy/J76yXBYABO34EdwExVKcaLDW24OgyLS7IKuO5ff85jf5EY+ytQr2knKesTWldU8Ku2Sbx
MHEuCQ6SD0eqsymowSwa74BR0Wv68H9wvsa4e6VvL1kBq4PbZ0xJ/yJ/lY6RELNaQY4IojJxFVgQ
rQhsDzWxdpiwl54FgLHloDqOz8ctq9KXeR1fvMa6MpRclR2aXc4qleaUBNbzdr56FEogxZz0PCeP
LaVvI84fIybhRzfoRcqy2uiS4eMW+Vstzq3OOe0YGVaKJ5qRdCOABEI0BdRdQGd3eB9xgDnFj7mv
kFd5QalUjOohgzXI4tC+WbOVfuDRfwxmqj3CSpanIQ+oHuYPPV2n2cesuhFwuVLKF/nxlYtpN0Fp
c+rus4/OgUVwF46p85fdUvPjNAxssRGcwjLq4E08jO/3+io5PnEQvlUN/A0ywQ8hOPMvQXHO1RSc
DMdEmtdHe4s2BuVV/A9rxqFhHjG3+qUuyVfw+rdUM2d9VjQP4jh9tW0KY/iLsNhWx4bZwirZ6FQ8
V18y0Z4/ZBwaSFDwq9FqNa2yCMAKLf3x1vC+OlJYyH+l/I4qKTRPufIDYEwOPZf0DDbu33R/LEXL
pCPu++xongaui4Oi5QwUSKf65k4/7+5xCjh+miCFc7QK2rhBdsowec+ytLmV6GLQiHaJBMSrxgj+
RvlRa5EgtMuCmJGYPBW2repIh6oD8ZEkB+7lTgVw9bS2fTozI8XdJ6MRxGQr/ztAEFKMDGH6C2hf
hPVvNmYxxxwJpvj26RXbgC3cV3ayNarGPQCt8LlKUt/Rz8zdFFqGnzCZuUqADuFgIm1TQor6e0mE
j8sm7NiT5dfz/d/JJ7wPQCvXUXAUnoGM6v5PYUb/PP5wjylAj6QsXptffczaJ46PUbI6C6TrtawN
idxUaWj7+FBVjzfuJ0I/KPDsB2SV57FZ4pQ3AJCHT1eJ1HUa32De7E3WhbebLXZRrf62k5BXZcDL
sdKENtYXl3Z3NMehFccpCwQs5nx03SAqDPeRJCvUXAefLJARfG/ZIZRw9Mzj2aVLPzvD5kZ0AQHs
C3hMtSD2WmbM5TzC/HNf4bZV+3u2My4pBmyb4HYYWjgjWhF0L+BMKKhTtc4CGrVtoHRk0xJv3/DJ
l6KR31KogHNonMV7kV1NENfHcaoFUsLQOR4uE2lMX5pBd8gZot6RKfn/DjI4IjzkC9VAM3DMVtR6
FCUhOnOFnqGPwhyslcnBsY7n+uEoaqF0TIZV5plWUCU+QDjPuidu6erBkZlLlUgpjPZXLkCKnr35
pwM49oUbFVyi6GeGx07d+VkzkC9DmE3bfpcahrqHFrdZ13uIU61x0s05d3lEPqkod+IE+yRBK7WL
G6Cx8gadoPnCLyD+PZ1gC2pFa4Tp6z/MDT4x8nfpBas2PREqZVwwtzAlMPXyazFfYOBkNARASLOT
HJRbZRqD7whqp76Hq4JgRN1b8TTaBr6082UYAEmuN9wTqjgz443qtzzaK0gSZpeoZ4XHl2htLdui
h4W7W085+DYbXFLVIuBUAo0oOTmtrZu4T8/MKXcToz0351QHGrMtAJFIJFzrbpkag8m3+MMrDcpm
nvPp+fkTNXp8GOEEFqp7rEG7l02SFXgMPq8obJPlehlLfqjRpBTMfHENWOjpLKfhXGtqMKMntm7t
lLHsWNKqnick2JErQj7BrsUlAs4Qe5AJoiORqbQLVF/cPdL8ofV8V4dvOIIWY4FnVtMG1St822kz
8cu089Amfa3JYB7SgYwGS+N8izMpbPRiBO9My3caFHr/f9egta+ko05wptaHOtG77CUrd8rBXEkJ
58GH8uLy9/cxIn+eimXdWD1/sZ5JUxoZ6lHpzG7nmx34u6CFNrh0ctof5J7RmwqMUFZPOs3ISIPL
GdQICOMMAYfcnyhk64wgGxEHC1SADUp1AQ9JP8yUPa9VW3T6TLkHZihV+Gm+MzlcvmEjX39cT+qm
uLh+nruOo8UrXgRgsGE/4/etxKdyXvkKedFb3N66HcVpRJ97isEXbBzfnpAT6ryOStQ43FTHgDr6
ETaugG0C9BcJnFh7jtHLGRWagHwF7UOdg7SZQfyIvEre+y/RzKkCzBo1UJ0OH2gEWdmL5nIj209b
FvJ4pErC12Wa7LWndmanCPTqtVBAGwy77vJziuYIqGjiopB1RGs8hqYhOVAMyj6FtJq7t9xDbk13
NtwqN0q4w8mvprVjBNq0hpD2ib7/xm1iDetsKW5xV9WSDHwYRnEllj8RN5d98YAxIZ7W6KrsfxKh
AVQvIumURemCJ7ZdNWrNiFQPbyvanhzF42mVkXCaPz1oTBwXCu+E9AyG/gvkUcViNf/WN1aYAsLp
2p6QmA8m7Q7jrxYwNRVJKGvzKSMUpDm+KWzQVjJhHFb160OjyU/U/JNzDrUmxeTPKHsdOJTu1Hdz
+S209MVo4kKMj8eLLeI1jZ5Wy6yoxjv+ZhwxxaSWSULDBzZtH4jkVXCrWagiWmeJEFpA7axgUaHq
cOFCrCJGpt6byysU5CDFQzqlglI0g0FY6sp58Uew3g77RUMA9opkZSNFi+pq1+ymga6VvhUTejIF
8o73ldOSYIxTPhxxIFn/7akMwDX12ofvLgielhRPIU1C93Jbwf10RrSphHjxWxNeT3eX7sYQS01B
4PPInncs27wdTfm159fJ0un+7EQmPklMKKGyDtCqZhC5f4hEaBKHUmVr+kdiimnpKFJTXQo8ZyoK
ctUPEnen0kuh/P6umtOJSuNMaPqUbjPiyUVxXPd+BICfvwOQEGejKtuKv9Nh8P8g9+syOskYQLar
ZbWLxLSpW2LBF1Z88FNBtxziMpCN/rkZ6ZQ5DlKQST1mOFU+b5t23R6Vnq4vQ43x19n5HrgzJiVD
cBnh6APoRrgGf8SofTU9rkSLdTwfbV58aAGARe/ZmOVIgLNTy6zvkHPXyfhCe+jCT2Y1CaR9jjv8
uPHbsq1eRGGEhh3QfqoWJ3l0yYQUTsAehVnIV3u3jpZYeO7tL9HSrOQQKiWMqhXdCXLuPE19XHwk
bzF5kxJufiiVy6bIhKZwuoEsMZDUDXoPK4VEPVd/C6fz1tQvVDE7PWHqeCYW/ld/h+iicHom2fko
Fp6mlXD83qCdR5WT7jCms1z/h6wfFc2xMI/Svj3MuGzl23foRJDQAcYxPgSIfGK0LL8Y/R2B8CDC
x/sUHE1ADHJeASyzjWUuMVARZ1pDiS49ZYg4Xf6Hw4dZ+EXOy7h7CUcnV5btRtvsuRMOKD9IDQK4
8vII2rpCqTK7XgqYtsu/Kdvb41MrsrZrRNuTXOJs/KxjiiSk469NZxa0q208kWv7uUorfnpFRdO7
0yrs8jNaJxxSZWrYG7/OJFEL/G8Vxex7J5rEZD1yUa2XcuRLbnSHruKftHA7MvH0eaLDHGJpp2le
E6+byA7KHHwbs358bUGZ0Uvs331+OlkwBLslAluBBr4lUuhcPtBKtNXT4HwnC2+krgspHtMPj9Zj
N9MS2BuFKfiSp11xYy3rbwranpT8Yl/pjNF45fz7tawTAHR7ElsdmnPHCYsrEu3EM8zgYvoU7Afe
DQdklH7479/m4DqX+ZYQIgMRLo+pGTEKmr79bOszlp+B2vc8Q28mEcg4oUB6BTTtcN/kLcBstUs0
nwAz2E4yB5EzD64LoUQYrOXDd8cjNsjFdOBetiRJxon2k5U9PNLIoOPEN+MgyUNl2bre4z95goKv
5WPSJyXwveOlqmfCZjbwL/1K98DfKao+C4Ib0n33e3zRHKpBsvrUNNrDSwNcn2uz52n6Ko2MPa8l
W1XfVugTC5vrgXFOkmMl2+19VEjSNG7bJV87MP7Hcp1SYHrcjdxay8W30Cc+aZ5bwcEruk7pRWAc
+DcKny+VCwzWiGWBzlT+EWfc5K4ovFG83sNdp3mP7XalWJjXlo+yBv/r8rQNNG13VHlwKxCX9WpV
e1uOMY66EwdQoBV0PCWGQrtrrUQUtFhEBfZxU8b4j/hoo10c/7J/nOnrWBfR81ZmSVBGMMr/R99a
HKyB1PQnX0nmU463fGoKmivFdR7jEt3kcBVOzEuOGJYPiOBUX54IVuRe7tW2pepLXHW1spH6wuoL
gD6/AY552WsrKOJlkPivdrK+oklRFP1YZ1F/TOjN5BLpu3Dk6gt8vfsdq1BwmkpYglK0DtCiry7x
SYZ1vuSJC1A3Wie3qQtBxucaUNewkZ4wdfLZnQL6MCAX6lirQ0U8LOtomKFE+nUh5pgCOaa6kWrx
7iS81CdOj7ojkv516r9yC1lP63L3GTWcob0bh7QvpCg0Ju/2+2mp/YJAhxy7jj0KdmHO52A1sVN6
uGU6dTWrxtk1rIhuo51ITVT0J8VDtawA3CI6Qcjm5gSHPTzBbYxbNUC6zryAyVfuZ3oC8KrW7nC1
NxxTJWX4M1Q6kLx1Ub+SXVD7uyMhJfB2h+73gJLA24M/pl/AtlScbhQ8z9QX6qOiL89hn8wGx4wY
NAokwp7vbSf+vG1XzjpjF3ySHtxmWJ4cW+R27+eeyVsJoIFAbi46Q9joKd8YP4w+/jqQoMOZc+wt
mFhgkf6WdHsgSQTQazhncn4tdWnEYhnyxghQKKn60umRF4pcrz+RD9mzfSnrZupYwfRoOR9BstSR
ch2PgjZ8Gc4bozXqPkskC9DUSLeLL7xUU3rDDCqPkP2PeygpU4rwdRYmcKF3yBfcW4IbVDYtiuOW
IDuYspACc65MBiFz5tXUv7cz99rY/8UHDO4vsIaGZi/IFQblWC3nwyduK9gHX9H2v2NQZ72wAX7P
gAwBgIMZ2Qm+OwIYQNpa1j5xrQFPrAqrOvVkNeCRv4ct8ek+3KDbwGp1ToITkeRyCuP+2yLk9oft
8YsJ9IZ2hW/elKwRPULYIIZqCuNzy9rxac5Fshox9ynsC/PvdttTL8fDzrFVF9oJ8EXdk1xpD8jn
0/iahrTw/Yxc+4TCswbBD30Sthef9SNegNgrfaaoQALskHDGs3DF8ZRcKiTY6+C08j0kRDSa6jP6
kh438UasU0PEeDi1tijiD6zzBe4qiho7DUpQCl26Ie/PZNM5x/GgGuqmlGobCo5vWExc0vyDntIZ
j8muPN/dH7fI5JPEyoSCxFTzNsHFE3K1Zve4mdPUSXQfQz8eBObNH3I7Pk/b6S+MOgCbldZRjORY
b0JZt4usfOmAL9zLr9j/0w9o+RaHy7oqQ6WVMzTAYH46KMtFlqAhTgdltOB6rGBVbIjFGwFOIbNm
cCPzdDNITtHi1p9dEtSrYTNJFB8tlGp7We4nr9osR856F/ujPgqZSYfg6scey3L3+amae9pCIAPQ
ImK1HqW07ZyosSnvyrW5dW/Ctq5MY9natRklAzm6MXIWu/zCHUuJtwy4LzMOALjhdCCejrAJFkke
0bdYAv7bbxycDbqqh/1QwnHzSK4NcAy2rWLABN5V3KRAlksDwsvqk7JRk5ahKLUKsrOvlwjfHqYC
k2qIWRFTrS7gb5o5erUQ5KPOP6+kqC5sd6VyBCsr6Lsazn9eh+BolV2gt7rg/xw/hOr6ag1NrnEE
bnsCho7ywe6wEgmeEvyQjb5tZ+UyuMEhG9bgWfyR8qOMbMiWYuFeM/uYb3S9t4Giq7PCVeTf4ied
BoQG+7sw0op1KlRs3pex5CQoLrYgcS7CpTvOS8N3an5FTTSS1gaYA3iStXPGThLeT5+OfP8IdeFX
n0Xu3fVIDV4lvYC8EjrR5X/OFIoXXzN8nRpJD3dLpg3H1jYEfJ+oqFXgSvZfiyiz4UEIxfCEmJ6z
hLeax89q0WqKh6Bj+OcFRfoR+ZFK3rVr+ppQNq/7U7agru0hNBZLhr52WrWP5HnV7rWCeiaVk7mS
0Q1Wgd9dmU9oBUwzz7Tqv+TNINDuoIHwKQPZld0TPjkognyuS4bx8IOIoIXKZp2DB03aXMQ7zD+1
4sHpHOoR+7a0XaYJVEf9of8a0qExeRzqcfZ08CjtMPaTx4vBfLik8jzpb3q4eY/bEFbq1E9IxEB8
RioiiJDHc/YSYHGEAPA4tNiYsSR3Wb4MqHqUCVlCasqf2QLKKyA3LXRmzh1xw7gG2mBBqj/VLaZh
7XO1FICDR8+f5DnqHUp95h1D7hDGSQufN/JMEBBG8dHjMpSkUWMPsw+B7763t9RHsJdkxruzvG+i
V0qFqVt6DC0AHP+ZzY2eHXcTu59FD5BJiogC8tPCpfLpSgA/156qke6ZYRsNTcUhPsf3F8RKjLCp
eRI38z5Os+kESgbBM4ssJtQXaRvY3opKJKcnuzR9pR4fvXtVcVNNnIs0AUPaQl/g0UuDQSYvp0mr
Rq57ika2i6DVrel1WxQAXt67dEvNHcqRCkG+QU7M6TAPRW890VzBrzi8wtzhW9ZC4x+hc5QbmCpY
l8GLLssSTi4+UC1a95Xux4xhiQqpC68o0ImPbe7L9v3832lxcLTcKARvzzkTPQgGmczLeD8VUtJL
dYZq+Ruxy0aloe13pl4cjwYXBjBteUZrU1VJc+hZSYBE4xC6jCxwW6AMn2DMCiMaaqPQIYM06YrI
smS3uHXrgV+NCBtR2qC+0aXIw3Y3PNWLg+LI532H1glcdoCGgYelA2KqZQk10FWzdFSHMf7Exjld
x2DwtQMMqsLh9BPtJk11131h8M7aCMpmCB/KxPSZaTGyxcBa571D9AslpAZX1/qFu6A6vI4KFOFD
0XUbz71KXo80yfejExVTU5dDtjKd42OSaCPJ3/b+NdpIAA1WFSTvIc9svbA87gmk6YUCY+aWCPH7
5JmrmVW+9LSfvdDIgHWaxdwzISHgwWs94VMS8BQoGsjLJdiwykQHitmiXiW2x47HNgZcDiGwGcSB
H8Zb68qe1Bj1zIASDPJKZKsG5nJocaIYlk925I/4vB5/oKTpfcNHMgg8irWtKIsCN3JDtiWi8H31
Ir3tevqYTPXuAVSBGe6Zvb9MJFyXqsuhnN6frFlsa+mMlmAQ5bqpnPzc20N+0IOhra0rZWVNlbEP
7alWB1kZfkR3Ukia1g2XNVgxqVMKEMhzNBkzj5fhDJ8a+vpztV+VrKKxI3rEWkL8uLAu2UvG/XYP
EGL+aY8yDUqk+3G1HVCKbS0Qrg+Ox9wbp8EJzeudpescNrCsyYu+/KJcxx2LpiZqV1Mkpc5iaegO
4y3m8OGVNiJCu9LMRbiocOS73CQs1A2+LCqeCbsPa319xLVI5pKdm37wYE7Jet/p2E4G7xs110nE
fxKmfWFZAuq4Pd56nS1EhyYY4S15Tz5Lf/aT6iAhmuL73FrDHd2tmgb2HyU+oxWua4lbUgG05phS
H47kumy9M6OJtaofNfO3a6I5zCR7aOZIlCPksgb+sczhGcelJfjuYocHbk2Fyi2gJT3grEQPYYrG
D/Cr0pGyCtrBEfUOGv5jWqO5hzK1VdlPWuUkWwdmWnFC9oYgY7vj0vOFI1EykqcGG/ayRnskyWFX
e7uxFuX2d4iSLFUQ/qttoeJd+KyYsDi8dV5kYGwT98olke0mGQBkOhEVtc+ruyJkBy6+OHwyT+PC
iKN3JHN4cVksIra/zbduK71vam2k7FMAlT4KfMX8ACE9HceyNXZ8hVRA5H/lP+6cHgL/47tDH8ZM
+fC1x00tduCSqV2YtkTusrYgOdgFYPzS8ogyxIN+vO+2gFOoTkkWL7hiuDg5OwtEvYio3FuPmtWF
O5rt2ZF4ULw9vZ4QnUy6TPL5Yj/ykUmB40Do37OQllU2mQ8BvYL09IP1L+R9kc/reJKI6XcSV9Ns
12iXFOokXXdbWjI5Ewl8IhdNaXDj3v4iKLMlHTLfC/Cz1OShkXCcAVBfvqm7eKeWnIKzi/vk+ToG
IgxsDGhjIpNtKKKmcf0cQHfJOELAcUVNcgQw7KxKCiyYWENC+qJiN/CMmQvtqB9jk3e1yZRnM1th
aUiqSuk10zblaiocHfaN4ViRkjBQm0iWmSQD1I2/7MwjB22OoYTeMt64OFHzDpH3ZgyzDuOa5uQA
Jfs0UgK9UyCVKkjQvQxsiYpev3pi7KjftTFdd+9Yr/L/4V4nYLcXcZt46yjKH9UhQjZI+1RwFkJQ
kIMMA//Mz4egTijrmTK1wSfapBpJbXA2TihLUEXjbGs5F4soxI9WXLseHU99XUzExZyiyE///FCC
HIGcTJ8dpiHculxycobqPZ2jNxG3IzbXohTzxR5L8GEJShnZaUirvCXQMc/6Fcsy0EDU6W41ykkr
w1LmClkGT7bie+UO7ELGC4zYgqqkpXEue4uivDjS+H15+BWUodOT9wR9d2x00WAnCbq+8kOmBEp/
UfArrRwzE7dSyrIf1BHPQLw4sg0+hi/xQNtzrjLiPTXbPGFVCt5S1Qy/lgdn8qJTHNw/pCiAPzHa
bb3aFGG2OU04DdupDQJyVwihT81TfsBF/6w1ZVhkGwxIwgNfo6gMSfKhS+mzOMdtvXvHygGt2crZ
yv603JU+Oa6I5JdB72xUSNORKTawLR1GB95pJlZHdD9SztFIgX7JP2zEzvc1Ps66md0+2RwvcYr6
kMc0MphlVrHQDBktO5l4ug94IWzAhcoJkOECnRfsDyOz796/DjRak7u1D+MvrdiRT59xhoUFktx/
Xhbp8UFU9YZPwbu8gyXQyCXD7c8O0bepZD8OZ0kE9KPUGfUwdn4tm93dTEbpYKZDmTbclFLuHlSS
97ZPoGJ16DtueIg/sT7aen7eCr8Z1Wg/qEfqlOwtSU7W5gry9hHi7hRTYkYaZkT2xqYCMv2WTqg2
k+8YHA2Isd91uYNgU5Ls35GgMhTljHRxyPGIatg45MjvNzyq2t202Xhm27/gGQxUyHQxLFx+ANcF
vcTHszVIv6mlmHvqYki9/tQxwnK0zLLXFssAQMRt3XrAHztRcNE84tl702wdO00GANfpYV3Zlgdg
9y75euZQ7bp4HLHcDiSBMKIifiDOjCblZ27ZUABpuxVmu87XzQf/cjY2T1hjprtI+3Ku5PCjDHdq
p9F/uPCu9MgSlNNMBTZWrue/oeq4w/gnFjtdOAtz5QrnJVWLDRmKHAu5pjMU/jcuj8d4+6Cjx7j4
r9ES0Xhz8Y3CeZHBwKR3TXQoYftkOD8bIDAzfvGvXUJX/oQD4uOCTHdacZpSHMfTMvrJEMnauZV+
X2JBTBz0xvvRAsytQdtYFJ0dBgr7IXYOOk4j6zqWpd1R4+gATvY0j086/w1WaB1ladGvSCExNcSn
FWskt0Gzq47c7j2zgyAxv+zPwO7jl0B32rBpVpAWSGjuHWe3gIPNV1FUpBAinXIudu/R6fcLFuZa
1i1j/FHmCUWwDtRj4JzSxQVsGW3nU7m7FC7mIZDI2wdYO6pr1XCeE6PlzR6/WfXztC0RWCIpuIt/
BCcRhnALXXbfL217HP+mMMh6BF7MvI+qeD67hwBDFKmYkDaex/G1c82w1TSC3i+TPhwPyp6tOGjV
trWJkRoo5eVCZWDHigAnr4GHtkerqxgiIgiqLjF1W5KlkCD0aI1WEqi8JLK9LtFOV7SHRIZz/Y0X
uvB5KxJe5sQKwgatDDIMm3ojuFSOoAQo4l3xK5G4FwxjfWx2rEukvaK4YlQXfUw+EOjwwfsRWRF5
cKU1XPf8lNuzM/opQgvon6gYIwNdmPi+F/J0TaMs2WWr0INCeJf2IUWde4Byk4mVK8aYkpFNeDyZ
alkJTCzdilrNJ1JdtvKMHdie4F/xbiKGpwNIawGpJdg2zfVLAdMWrwkFDHA0ASYY/qAAEGUwDk4O
PV3uPbA/5oautSNiiZL1+qK7WW5X4Srknh1/tNRPBmKqvSNXCtnP1dXUjoHDaG+wE6Ca3JmHJSRa
hQ45XtsOjKUiOcllZSJtSGMwIPjKNPScDXYkxWdLM8g64PFem4D2XlPjePyKg0dHJRpmrKkbQdgN
8sK+AELl9P9uYHN4jlbjj5M+2XjHPlgxDxZZyqFgi8m+nf2vvGAxvn4uMldpNpHIBijRYemouIA7
p29i8qG8VAXtdvIB82Y2rk1gnStyOtud0lQrF+udBXST7u/Tx19pwZYiLxwP/z7U3owF5kV99IvX
4rnO45VsDJUQpMRdqLwV4X2NflL/iFR6dyIPZexWqONYgjyCvT+tZFctNYoGjlzj7lpFjm2ufl17
ptj5GNz0r8qiICuo1WkTCcHZyzrRwK79PyRgVa1R9NIzFgEwgJery1RkYG3K4uX0hujdY7kSrFPQ
W6ZPksF9L5JymJHNPSefLRRiB1A7NLl5txZu3BlWADwP7RB9y05U4gsJq79m86ZnXBdomXNgVHFb
FeCrz3COvq3J1IhPT4zIwZtxUcGzXOGFmuLrcszav1KE3Nt+Z/iP1Px4/lvWWGG0+/663dL0M6Dh
Kzl76Eh765rZXzNUxUYxqcGKCorPsNCZz0PPZdbiCoqWzfMJPcT0MUMVHIaD7iXyY7weJLFb2634
paSJMFoUl3BSTda3fKtpdVmj7J9hjfw66cRM8El/VUGJzDHP/4+FWFDZMsdNEjhGiJOWqXFjjCXE
CpCwSBF87xOCEylXQQNQYi/g+AhWx78LjV7X3i2hbt74aaUQEMcZFNu5NyknH9NSa1KDAPadITJ2
sGhd3VqOYcvjVzDUdl/atyJwhWrPD6FRvyA0/A3dCgVHgfLDYBgMvUKakcK9BB/hBs5ho10MZw9x
6xtf6jcS/xOyx9vGkSCAjJZYPpxczGgHwWfClbNG4SfNRqcU62QNbvEvqJbZPjgoN2xWW+UlRowp
oSzmpmxzk1q03ad2THZOEq81SHvbJccUNDdGMA2OrZ2A77tx27Dc2ptnEhjPNrmhx+J+BUA6I4ip
kK07cJrbSPdBp1vCc2ZsFQ0iPZq4dFlK7e7RKl78eNuktlYF7M5sWQZTDYBF4MYXl9YHEfYo0Vn0
kPnjQ3MVkBjBY3FlBgDUmH2LGFCK8Xp3w3CjYa9w0EMn8pnqCgASG0wCscV57ULItwQCzWgS64Xp
yQvIgXYe5N0pfFH4DAaPsyEDVhtiJ3GNSjemZfMmT/xv3QlwDdmFXIzmCGWyvJ5ywMOYNJWw2DiH
OzEpRcFXD6dCigBaYgzjj3SV2NNeKl88TtqJ7tKxJTaAxzHKSMEoJOdbLbqZs5+/omyrEsB+YvPL
DBlTofbaXNeWYIukeQ+ynVKbx0whCghnMWwxQNEj7jalJiEeeACbnKUeWFPx9ojbUCUm0Fo1/QEc
rvRPqB6Qj5DxbIqdMWVJshPU/08XIedWrfzcYe57e/aP/yXwXaEwkzPZloZDJuUPdZBTQhtM7J3N
4o5oSBkDZwPF4XlCCuaxA2bViy4FjoQtXp0efNLjzJU0tC+7t1x5eLWzOtwW/wcbdMtP4bXT0WWB
kNPQBM+dqFOCsQln84oY7jEIBX4kyh0cpfyVvuNl6kaWGvbOR4GJmxepVN0lwKsHBgOvyCKzUYYD
LVuLDKPmLyqnw1a3vc+2kO40S83SitYEpegAjduESIlDfLcntJRQ4TuKiKfZZe8AN12dPLm4U12P
JfwEOfNQHD/ynbEtAVVK5qTQQOTp2mgzwW9FhtLxsVj1Iynhhwt20INfdvJ4rzs7hZtpvLrjR2ux
coUFqiX+M+AwETnR885+cNohfY5CDMgDAqbMDYHKfN5ANBnVFFYQlY9lR0bY7VYqgW2DoQBUTYtI
iAaDa4G6Gyd+AYdn9tcxhUy4gSXW9615h4tWvFl31WvPEv39Bhd1dDu8LXSvVWpaicdCnjn4b04E
jGF+RV5GVIipGJVanOwNyr6EBJ2YMBpkAtTDGy0fsp5fHlr1XWbDVkARt/7IctHSboyb8njaXfW/
zmqIOc8HIK8wC4cV0hOV8How4WNI6gmSqyLKHQfwYIz5nC9NAZIW9wmkkCi7z1IjOW9dgLX7yAOw
LgrjAPH34H5kys1wdOPZF+5wlFC2XRVLayhJ4N3JMlJQS/Ew6hvUOtFFefij0ZEMftGH3EgJfT78
LTh1GljFs3fooOMEeQCB7GXVADLAyn9aSkm1D0c9KOgocCDPW4wxIFsId7PAEMerpS6c3+7ElZ27
7mb6Gxw9veDtVWYt3XWukgYkSUbcrtDaq7pu2MDtoXy67E6bIRvBzjd5pN+5kAO6TXfx2sOY+Ai3
nMoZAXmJ92Yj7248nHh2Ex59oreT6nMpHiohZ5aFl7mrISFLqOBKqUnvMZCbaNtwVCtKwI2pZP4L
L2eXl71GkMEnhqhvdnqlEhfnHRt+CEH9+CIkJHlmv5/lv3W5aZUR3E/LrI/hUM651uAx53bcFDWp
awhzb5dB1XX9iUpd744Zt/Dp3HzjKNprwf5UVQeV8QGV/WHlYdzbm5hgYs1Gz88pmtjOgAmR/AF8
ac5uWKPe327gRgP2InisgxGErbvfkbjdUaAe6ZRIZ0cbGfGurviJHwHmqYJDHSpRz4NkWfrqkNGy
Z/a/d5HOq3loDhJLqcohcKQRL0a3R9YVT5pYw1XDZMKjhTFcTepvKUlqoOTQ7v+0FuuPO5Fg5I77
FOLaoeEs4lVOGnrClPbo3/t2jYq76z8uUvkt5Wttea8UL+uZXhUm/FZd8EOOqZE0OG8gaY1gInzE
WPOfoDOdY+EG2S6cY3No0bVsOM4C2wqcn3BUnFFPFK+FtC0ByBW2jLV1RWMyzRdjMD5r7k7qyoXa
IQbNAUpWRmyv02bB3ZxnGxylHClae1CYE0CopdO6ZtpclACNMc88PpCmVTRJVaRBRfz2uRH8vHYj
EaJF2OLJI0Q2dckWY/VkkzLY2pLc0PVQxj+8ohRLVVqJE81Dd3h5PRcnw1iHBXt7v/FwY+3aDMeW
YqiKt9maG94v41jJtywkkVn8Cg9OM0BLtaMsVFh0nD6Xm3gVJX/3JMUuJa4+ZM8gIQG9Rk2CAXdd
FKhhKmKbRjwzN4cXOPP54xRW98b6nWbElYKcV4FZgsWSf/fP9Ln2SuqnSOxLkyQMRIyIUABGyxLQ
lyrcRSIX8mccgZ+GwaAsetHLoUi4VlqBAMwspQ5FJb6j9cnYguA2yl/0Q7DuCbFR8vxzShU5mrg4
FQGzVeAF7SRqNHE6s+XfasK5nbAMgkaMvEy2yP2eG3S4EI5Eh5W5KGfXm69GWzWSWDWdOMA+YJML
YahHEfKCk/FtdYhxAXG+kmMHl89cGLTZKAqGD6kZiHsbKLeHParUg+CuPeanuafYKq39ELuZKwpi
MCWQ6tJfAw0jJ+5BBk92U9xFaG2H1agivvHnFX6Al61S9FlSpuMqzk90oDGFJhxhKbZvn93DYsyX
5qd4VfnjeLA6lcjPbh1mjn7lEUO8QZIZzYJIX47ghG33BNoaCZnV+/+ChSLBBqT1kPgpQ84IT5Fr
huCwaHzFmAcjNABm5Debc1ELrMoeOXGqMrndrqLZ0Tx1l9pt2l0EUt0d0I0CHaIz4ZL+UuUYOQVO
PCIzgPp2z3hgDvj8sfMMzn9S7koythwv3TU/lqZ9XY82uEq8pzVZBtUDrZmk+JtfM6Zicsxami0N
fXSyToMQBB2bzUp+lJ/usC+d1iRlo4k6xMraH84FiaTYnr6/hFwNVtgxpJVNLA3D3fki7HHRS+9p
DQvAEAV2VzpQOIEEUXh6cC9IQ5rodSIWjEhshExpOHNkRKYQPnFLQ7q+ATGFuBqwN6sencCXkVFV
GK7FSKzQuyShxAsR6GC6LxoZ/i1JNi//nV3AONo3d2dYKDMqipZACYbr6P+4dQZJxHU5u5Ts0Hvs
4A6GdZDCQUp9pt7KsxCKqFQTGPCJTgFabSE8qmgJcbMWisw/nascrdbuTrXzbcTmSbUDDEzOr77E
apqAEbpqFetYE9SA4jF1x+TvPex4tfqn8j6hp+m5qo8DGa60fxRMHYFTrt11f5Ub3Or47jtdKxR0
FVqy/m6aRE/IowppHv/JNmFa4dRDsUz6wT+lDrK/01CuebDfs8qvhfJ9LE0vcCXgDElXlR1EVNYr
9B9MD2oEJg7qBQBmyuD7rxqx4pID5qGcXUVX2XX8BSDEFG/jm3losheQU+YHOghC4jpAjNI2tzf8
xUeuE0ydx9d7q0YlZq5maF/YmIKRwym/K6xfIbP+xjsKtGaJZlsjbPhZVV2583cafYwL+LblLIbb
lYsNeBEeRfzy3WvNeGrAUHQDJAFsWJ1++I+1gwHX+Lj3ZcPDeQQS9uHZ7Eec0wn5oUozThGas+bJ
iU/Ou/d0SG3T0ICM0juoEZ7CrtE+5UuzwKyF9KgLN30SgGn1QbHdCEEtRlPFOrp00g44m8bA1P6U
OGU8LHnWwxUTcg08kzP4vI8eHHqmYMZug9PFZhCCY7P7TZQtka+lSGKF/sYiSlaAky2OSYYyifJi
fJULN56+XYB9VNQh3h/1wRqSJVBnOVjx0t5N4fZif3VT0kYrRJdkcftZYkXtJYFp0zCK0lz/tvSg
B27/x7t3LxkszhAv5bDySPOzyHcI+cyqhtSuMh3eAkNR3gmAbXVvu4UiKSvMqFgLLwVmuLdfqlmr
JLgDFsJw9Od86W1S6c9DtexoRKX0wMj/2KAipFSYMSgmVZbSckDm2KW3RAz+jiGmodZRROyNV2n4
ZSZqPmBUf8NCbSjwVrdaHOZMYtxGxJMk6hA3j9H/4th5deb4Kd+Pcgl2TmdkjKtTByhSHI6hlEbG
QI1ephIteBLvmNDFnKsJ2hwwUsTOvwhnWuOQKcMeD+mFJHbF3C6CMPwxORdGUZllR1bhtgEBr0Nn
7MxsohXn98AJeGbDSzjgKBlfADMDCcxSL3N1lMpqz0vu6JswV4krUuXswifPvC21IkkhdMZH5KBF
Qts/mlfamAoke0BuN29QJNFxUYjeyoWab0aZ7RMginXuOuCaW/XUjLpbvcXVtJ6Qc7sDfTWOLkdO
vzzRwzJUuS8mXnEsmxTJj3uMyu1skeRTiVxq4WW4Rw++46XDfSPMPmjJ3SjHksrwVax71zH1CMSa
Tz/J3pwn5QzDb4wGsx5cxed0g19TcsDDjT5UOJtPCIXV4XssAMGxzGTZ7HOgQ/DtAXba/L7wNtJp
r/0ykIs0psAa4GNVdlqCkG+9jyNnLTbEiKhlAvPsgj/5/S9ok0isbKQoYooIJAMvDhXjHcvawBqO
8tJiScbEhGW3MX0I+Q1hyeAclgTsBott5laDLbbZOKh7Kf0UUxzmyID1m2tOflHl4CZOw/Y+Xio8
7oDDkrCyZbknhKDJ6FuqMJ8GXFjnd9lgNj2XF+YhBCEgJ2lDmdscHXpAeeKbSr5sngBITH/5Vy/O
4frIrsgb4cHHDxCsEBWDc+GVfqqEBZVN66+T0zS2YsJOZWHcJOkpRybmH2KBT9NaI9Eg0s4AXIgA
JHnvPx2s4FCEqBJyA904/xc95DxrZ+x9kUhPR0yH6k+Z78uqf23YGQqZGKvKSJemh8lZy5j48cPf
IubNCRScyQHnUoui/0YuCjNhCXHvOi2C5+xn/tKTBrQK7Gn4WdAbcppkp42Q2vTFGscc1XuQ8bQ0
fUmKp2s5uHsJ3tyN6xMN/S2v3MRU64TIw/Tj1e/d0S27XxmjHZrwhQln0zDkfS46+wxO/1mVzh4k
jRdIifqQv0jxUfQY4wxL2MnxJiDgMppJWVvl5Tegc7FGWMoyFpNP0ANQq5IvWwbsjIzcPubHpU72
l07TyGT8N4ynW/1apHTVd3jdCkrJ5SRRAR0gdrgDcbiOeAg/eawp1eQDNnCvGMf+SM/Z7yJMrXKm
L17pVIvpgvCYTSF3f4Y6CVpW9n2aJQemgpPmtkUErW8I2xj67yjvgHfD/Iqr+4V+vYF+gupzL/An
wAiDJ7XZlO5Qi1pCUm4kByESQ1+Lb/c53luExA5esXJVaZMkb7REKcxfAZksZA0704h4JcKXDjj6
0RdBE1rAI3nqMCKQSH40eT/jbA7wUImJEvwbAFiakpI82JKZ+a+YROYWax/iQ0OI0FYbj+4asVOW
NjVRIFzhaZMzQRl9X5rYdzyxI3PskGkD5u776thXWa1pyYjzp0fZZaV81kDri1s3CciByQs9O9Qp
ZX0QEzSH4jvLvXwTOoVfXbeOmt7GYCnaGXDUFwITSvrLjlOLr6bG6wD7mTEFC1gQtWMoUI74io4t
SmUbSPZIrdqBT+jpfXENjYd5oFX60XgPc+K7FRi1n2+6YSzb4M0Dsy+U5qp9N+LSXWShtnkMBapd
sTBrujv0vQdxeZMGEzew6KbppoL/NcvOToYlmJ0ZJTCY1WazYPydGUhB6FlSdGIhawOl4HJAXlvX
Gh1/trHq7CyDlUOPbWQtK5MpZzc7dKd4wOquTsfV9O5fXc6Q0toI7E+JuNU+E+h88eo5T9c5KRJW
WMThcQwmYyuDEYRVJCuNDnh4h4dlQMxwVzkEzkOCEox75aGwrBB9fjgHuuzdtNWIfhz9X+upq6VD
gxDJq2yHvxl30CWgIbYeuOmgTnVTyvauQ64hf1GhR/bNJUVGjCDGBI75AGqrIu4Ay9ik3QXrAZG1
1RqYKefzlaASUxxoEsLGzxC2YRM8U5IBJ1StdjMB43H47B00pi8o7trn+WZeCxGSh5/YoB8xVT3p
8MOxWjkq/hZh314iGte2Gsn6SZ7K1lLOa5rNm2chp3gmSU6oXstjgGx+NBwUY6gFvVn7GvfJGTs+
ZbVxZBFfeAsmzqiVEKFK9mynMQt3F3aTY5iaKN4Bcd68TMLImcG6zqehipdHMeKGzrXFZqldeZDK
oL+SuQdh5EJDxWUK1Vd/KRq1ZWRD0PtIaV6+Qmmelu4t00NfCBw6gY5wHCS7F0yWF9iA3FRPa5dF
PtZZSnkGEhgF5DEqkAxc99jPMgxH1e3Ad9kvmeykmRVCO5yRRU/OLFl7K2ON0hg+i2r/F+EAKTZU
rert2+17pVTLgXNEdEnSN0NkV9CLOKqfxTMaZXVJBiksdDOPqNY9i8I64z1LSL0m1lrSwi35oKrs
1Fb1lmDvXJhJyxkYdlGwQZquo90IvfMSRmzv9c9O+/rY32Rt5PGhggArKphBJvLgXCMICVOjnFn0
zZcDbrp0O8NjI0ux9TDp0YbH2YUg2YEqEJ6Xn0nFxOnijzJXJnmaw96vS6Jhk65uW/No1nwWtlzn
M257klJOZzmS4NbvIjUvz+dnLuyBNgyR4FA5tgYcuDNfjGYxGvd9Zb9o4fVlLQi0ZCpBDbbuU5gh
oCqMdMzrZiELZ17EenYpSKLcF8rHxoxLuu8x7rBUFJ8/SaN3lM+RaVfO0eKjFZQcUllvCUhM9ome
XNZ8sg4gbvpin9UEzAZuCB6nH8KdDT/OVO1hnGWRrgGXXQlo2Tl57xZOGwK+PNxetwLM1L8ZjbWA
+C2OiH2U9I9GmexelN089iW33i3kcNItmzm9NOowv5zp3WSEmJCHLG2R9x/l+NTxO2w0UUobFrbs
5KEpW1Ig7PQ9NnnvJAiUQHI+0wGmP1qFzyO26z7ite8T173E0x01+lXrxHZ5hM2VsjiDeyfI0KTN
HeV50uHFYQhvzU8AFeGtgz1B5ORsAF5aHoqQj5xLiARvCpgRlYm0bpF5RFVUOlrMB8kuitikgZV+
uY/78dd0XZRrZlmdM0SsN5Gl6r6u1getsB7NILYi5y5ZbMbYFLmELtsgG3yi87Z05u6pPBSxe2Ha
D+dooFa71fUiro5i3mTzCnNMO6/Ha6CSF3uqVqU88SIxY/FvV7Hti2tqOuoLsIvbOepis5wo720c
MizM8cp73k9nBrZpas0qafoC6WwDkaLEfYhuXiSzR4XsJIyH7VbGWGcFWx87Zbtih3985l2NRMU8
RJ66RqZGsEL/25cFhQr/lAGJq7Zos3N6Q3QiFEDTWu744SCbY6BtO3xQ3/BahQuzpP036RGGIKVC
E8M8ZEcbBriTXkng20hXoZ2U128OClpoADSBi+udDYIG9HtsMRmL3YVzyS0k6YyGWoWMf6Ogo/Fh
BP2V3Wx13HG029IsniDxGforwCH+dJBFVuEFWQ6o6Dgb/IRedwyIpueIA/7L2hVWcvi2FMFM7kBO
hVCxZu7etQ2J2V3e5ILceSqZFcOueVItB533/6eEgC9eKYKxqSV5uFd0unvBqdHw0BUz6stvPDLg
cZY5z4Dmn6xGgyRVBPy49H/TcopIUGzWzVe/X2D6fyok3STGm9rT19wnwTpzmlHJdaEP4b9EeWmd
i+N5/0XhglCgxQlYko8MpYfA0OoEnyPJ/0wt961t9gJuDGxY3c3YpRw1jJT8/FzIZ+RGp3f5V54e
RfRhnUzFN2pqyrlwJQNgFbt2i1IE5CdRd2LR/mozkW8nyutnzAR7bqCppppWVIOz7ZO8zDY6hFg4
aknW9A7RMdApmjVj/dPTfhabjrQIFy1uPy6gBNjtdd13KqgvTqvOoZ7/+MbcgY+cuzKgYDTl+BHe
5NGle4jp/JuupYCQrdL324GNzs/eFQTbP6JoeLKKaZCJ7zEfy30ZrOPBfEyOVJszNGa41FZ7FqJy
qLyvxKULqweQ+DZOICj+VnU2ZYk+P77/Vopwc3FA6Sjd3nm9erpL5zoBMnXHntIM0n2Ft1Y85m6R
a1n3d2BW5JdqPCR7IJH4MHlCiRHkhMAHljGGo86w0ABOu9P6KwGR0JpzKKvJw9BE3fOJtWciw1VZ
KaC5IbL9mBvAiSpMZKGM3eaWVY/F/OprREUgl5TkYDE43jiA5t+mtyg+mcO2sGDkBBxyRQ4kZcTx
B3p/BWcn4cGE/TNxyYsSe2v3aCgWLrpQDoJp3tzpdvTLE8da1Lcfy4d9YgRZ18ldNhrQ8WD/AHhD
oNPtXLw+3H4r2sPup5ikgjKOOxVzJE/tMeurQ+bAiuFFp8VjshmtvIYzQAwHJiMcyWirU8ypMfYZ
NxOu4+XUncXGdMLbQI/rCnersysGmHx5E2MF1vGUiQLqBuJcRXZERKKv/YuPZfppNNM0wykpZP0W
2W/HclXhWTrbjV+JIMVAL2egQIDH+tE4pn+v54rsqRyhaGslBGpcKmfxyPrzMYZot04krrFxTmFy
BdfbYspolvzXzHtOdak3bC2PnHESD0onlqAfsGWvyu4DUGYbTAKPNu8W54a6OsU5JL0+7SeUNY2b
FGSZdq74tRdbW4V78YtnkgSEofaI+5W9ak4zuMd/OGAMy4gTmWgtIvEXYXZtQc3ctQf50wTQr2jX
xV229cqV9FGtzVM/IcZ4RB32NpjI37KDbJRJAIMuQSvdNkCIOHzM9Xsh6MLx/ayXn/ZjLndRrGKT
+foDXtNQXyWGXo5JK/V7Wbb4sZcR0lXIBRnn8PU1tBXC63XU1BjXfQorOzYriXxEplU0oy9n3B9b
1HNe5HGgMfkDF8hro1nZacjoYoLFFIsHf/Z8OvqZKVVlhwCAkJpKXOgjujhycV+IviaRykZaW+Sx
uqomz257KQeJZAoSPW8FFsL/aIWSwbGf2eWCD8GJp9rTA9Nhal96Lcogz614ECq5cPlMFkv1ohWN
73AOuP/2IbkeGI3F0wke+U3KLKIXqckAFKd5c/Tp5wPOW0lijhNrvnQYpmYjhQv71lrSuU7VuqaC
LsPuSMuPc7A4VsLvw6/EocrDTXh2ZwakKwHefOneGYiI3CDl9EF7Kptt3ivYKqUni/yAYxdhbv0q
7DsmjQ21OH9J5fKVTeQ6GFQcmFTuosZBs/cz8f/JL7F2mxsMmd3EB9bgrVKcOoevRporEiC+34KS
KoBYuv6r1IaCa9kp4rAA3DmFkI26We7qDtKcZ5d6Lmr2sdGN+Z94RmWWJmxq5FfLbtpm5ZDxZ917
uYuL2Kdu5muk9SY625T/A/m0kaKqy5dWuJBKpkG906t2nI10oH3eRsueLRLF8Hd4HO/mha6/V4mN
a4NRw8HG5SdHMOAa3uIY54q/03yksW7tzAmueEDF7gjl76dcElL0HtQiQfljsCiJ+rR+mKjLHyj3
MdNcSpcyh/Lu1cp5bW0grxCNppRKnC4A4e/N31rljbCCPSoU9UoijRazBMLwLQMTFCF6XC5MU+3X
kvuKXgYV+maPtms+EWVkOIAbeGapkciTF78KxutyQ1KeZ4TbwQf+U+lYN1OPoKmP4RWkIYFZdDPS
pV1+wDXZ50zxQs2Gy1ZY82eSA4cnPhN7nOwYSHRJ5hFP1vo8wsN61Z3YIcp5/JtMnPWVTAOdgDjn
K66KWu8/ZJy9oJigLoUGoH4lyM+l9KYbemu9ovFYuAnyvGUnWRDEubUvMCFbYZhu8vyXd3ZWxjZK
+EOyyQ6rnDaSTksn/fh9sxy2ZoDLHA8Eqp/VI29muE57li4Zg2vrdUP/gbe4NKyAfWjc8qABMy+e
rJJZ5WvdZqwQv90qohbcctP+zeIYJM3c+0Mf6mR3rJgI4b7jc72T8lq7+NTy+VCpF+G7udn47Gh4
G8lJw4nde8iNynO9gvTTJvz1mmEMhdFEdCJkV8ac0CtxMA2G75JWqwp0kp5rOGwPk6i4+39kBm3u
keMpD2z8VB/M8xfgmOb9gdQEYX9bTWCLsJVfrY0/4QPy3l9GXyEl6tbjDvBtwTiUAJNGuxf+ItHx
DiD9ToC2uVGkSbCno2BhkOfbSoVbi+JwA3P/kjNsR+onauZQijEUonpf0qToS/VQ528RCxdUpH5f
WtgjsizyFjItHIveWbHGyCC2nAEcEEyiIr05sQWnqCPMQ/gzM3KntUgwCjopcmgWUDsPxodpEI2U
plONc7WDt+NK6TKOtluLGsOBCER5l78w34ZdaVYdCQbKrWiEuD/zpgExK8ZexQEdP9c/5J6YTCYO
C52g8GxQC03MnY5VXXv/ofHdrQkfHXfayXqfq4Y2HbZKRDkwwfBzTfal+ZbpgLUeiRcKw29Q/F3a
1BIeGYJOU0KRcChrcGOlStyolgG6t6REczKg3lsNLh3YMfqsvs+bQJwq9vw4lPLBKgKLlhDXcXbF
TUnReD9Tmu/x0RqY80mIANx8uHHV8zCXJN30GcexBagnTXFf3edcz6gDOYiKUESoy3KMvLy4Sivu
KSRVdv78DUu8MhENa7QRHqFgb/2jRvNo6T9Z9tg9uDLXThW0jLpsY56tH+QxKxaRLgT75NnbsLxo
WcgC3F0510uinNqkr9sEObub0LwlDNjysSwYTq7MaSEYZCzT+1mCBswsq8AX52R8ej4d/ljzcL1q
XF5eznK4+oUbdUAcC7hwjAJhQd0xCUCqxrxAMadad1m2slG7whsa9uGG/6CUZs6jirP2eTXANH/P
6cbEty0o12/oxIT/jiggH2k/joREg6XEKlKsD6bwDTn2h71yNVmWrnfaqlILAsXqi8vOep3fYsGg
mfrZN8Q10a40KuJdP2d/CWikJ5sLwoy4Rcs0rwOYL23sdR8iJN74I3+JstZ1VB0tb2KV8K0lyJps
EAxFYvDPHdo5hVxv3SNHlRIaYbjjeLxRTXb36B7haFrkSrQSMW9PsGfNgc3eNxbpiVOgkMjaFmaK
img8rn2cbRCDEcrB37ViV+yqigyduJpnXl8uO7CXwzckWRgkJiPDwo9+IF0dWLNYhXKfbmWc9RuE
Urfhx2bGqRDgqWC/gnmCuVSJnnUyfRhKotk2ugC0vfPuBBE8MJsFatuin1KkySdzm8pqdpgdP8vA
k8zDReQMFiGzpn8qU+qOx4QPkH8FDHZoCwiWnmZ7PSgqU9D0/ASQsFJGWEN6RNAdyozLPj56diUN
/vIjpfEkE5fanAqIRNJiD+xCEFggPyZAWOhYj64yL6AO3uGjnfXpotw+idrqvR/tHcZawX8yVjQK
XvuxEz2+W7z4dn7QihK72lMWdtsBPPEtMmAa4n/fw/rmeu55XYaprJJ4vx7KuHdXU7fVeQHg8R2v
na51I1gV2CxNzYMoDQWy3rmB56fKnK58fSs4QRKinguVEta8V5v733lxJ3GqGpmva2mDnpepZ8t6
I3/W/McivDZILAenll2DaobiR9JQSl6r4ySQHWWMkwThkfc1P4cxDvxbzMMz7Exme6WqLp+nsNvg
Qr+UHwNJAqPe6P+oPpjN3m5J3sWk2w9Dm+OFJlvJ2/Zaz0ZGbeAo5GQfzU9GdRNoSpBo82EeE+WR
BsPSq/7u3YFtYi8HQ2zFMam3bu4oOFMNaLfTUGtdtPT4GcY/lBAJ4wRUBG4kTyfSh7Jofpq8wDeN
o3rCnvWr712Plv90yL/OQ2MUt/JcsDkVc3LlMmI6ZntzXbVZpKfcXV8e9YxLLFld0sb3ZHFD4FSX
DdAtCPACW7StL36556cnMeJfIRUBXw4MK6Bt/uYhL7s2lb1HeZ+bi8MFqy48t2q7kB5S1OduJ2vO
jDQTq7chr/l4BaSnD4Owi/9n1h+nb9SMMy64gE2VJDeVOv5M63MifnUMDSiP3cK8oXw1Xul6546A
NEHF89utOW+kR9V0T5LgOvT7oReqQB4lvTP5trNd0/icUAi1rH+aEviwncq+SQyhH61Q7tjG3eTE
9MbmAnnd1qWtMztpesp/+vWn28QYxGE6vUklJV0SfRO/3RqVpo1hMk+30Ymd7Raa7M266x5hTtSG
1Utty2GsRSU++nJ5CXUV/wRXD2BDYv1afa3DAxAp99GfxcTHbaDLG9HlFrp6I5lb0APKSY7zYNFa
svHqIaigwEMMNjdvg0WBCk9vNok0/mEtpi/aWPZTQ0iLj/Xij+LvwgFBeMNmDs9dPO8HyoxtJMSF
qR7DCsxZGtWHIXvi3jOajqfVA9AoxJSQb7Dngq6y0R4ksq9U/6v0ManQXT6mOHh5ztShfqV7DRtE
Z+M4nxIoyGsP0qHwkTm5mxfapA27f+RUMCXJppKlI00dRki3MLu2X1vO5GrJx4x23Gv2R++PtNyN
JqcMPAkWWqmfFLB4J7V1dUa4GLWYAY+EANzMK5Oc7PrVNsyjLT0KLBvhIoCWliASPyFljwKfucP1
+DmhuVyEbfXhRY7iliMnnHJQCoDO0+kkKhrVy+Diy6NXb2XZWKrpPmqX+TxnknNXEIVbAJkyjb5F
+CWWuaCii6eZewyKK8hcJZpI5lTY8UqKtv3iXIAT7i4NlaETDFGOpFS21oWFp1sTQLu3ncAS/ig4
VDtpRMC2bGrRA8Dtmbf0OlLTQyoG8wCa07/CV+LWe24ga7Hu7DDY4TbPPbIVOMqjVkmBokVmdneK
Xy6xhRTaEovhHP9Ov5FXz3EVIcc5mrWrCR9Sr05zcDp3rvb/Y7hksWRaLIYzwF26bOgO6/3zIa82
zgLNax4Qd202H4R5j6aDbe2f+6ezR1jjffP4B/wrKClc4025Fwml3ahdHSuWixdIbW1Qfj463eUS
fQ0ycbR9PXncjGONzZ2qHqRDX0bcQLMU+ndLFi1a2jzIH47Bprtr7c+dRqYGkeQBl7GriWhN6IxH
EMrG5OpMopHVwZFMA11uWtVYo3yFISBMijtKh5nm24/aK52oRn6/vmhwoRZHTQW7+AjsU7KdnpwF
6xcqPkiwLmcDCRfBYpduEvEiNnakXpysNQaOcFknhwc6x62e3j9DLmVIym53t9uLsB0mF5g0EsSl
pqjoa066BAZD4F/pn3ixhBp8qZV9mwiwpYm5NlI+oWioGePQ1KZVNO1SFPkWRgOlnzgdP7mO1vS+
PMyXKivR1eketlta+AJ3Bc/aytkoT/BaGj4CM8Q0cWY7+EO5WdvJEupKqy92LBKFDxsEGT3haBpi
wd8oFHURYbFN6mHuapPJs2PEA7bU1+vbA/X2tpKFKKBcTora5/LE/MKzky4R8nzZP4/jvuRMfiCc
hrOrl7EgWelJmbV4tKrJo1VTHLtx0ZDh/HnjdNCkFnWkrzwhxNwYoAmxfLfkNplRza6fxNA+0gVe
l1THHdQevGJsDs7C/fqkH2fNsBYnqHEEhQ98ekXBxidsSD26C95+OpGEKHay02GixhUI4wJfO6Tf
K9bxnUxAByUd4S/Tpkw65wfZtaVBTvala95EmE4SeAmhh4kIaGp+n3f3JHX1csxDbxhKk5kyFF1k
La4SWNprcc17WQ9lsQG0sPLnrD1pHS39EIQzb2WJMSTjYzaiFAIbg/YWB9K8kNY+z9WEQ+JFLPhD
DCgpuToAgkOTiCdO1xFGsK6ExWeurNZH4egy4XiZWpYcwVSYeUD8pSIV7F6RsqwUfvOAbCVTxr6K
k0CbSdW1EFqLch0NjmberLVIzQG2yq6HNS8g/Suh3fU0knrhFC6I8i6huw/qZmLip3rN/YpaOeTu
1CVMZthe2CrvrpfFlz0rlq6B0msVVcmcSX8HqgddVmyeHUAb5eoPBdgXzHiWw/iHQzDCQhf+8HQD
bj/c6JvKmyIjaNKYKsJBPIcQnTDaq+LqhNQdcokd/0ktorrjXQLX7ENAHOQ/nmIGJpMnz3aff7ij
O+hgjgd/Iy2/pTPm99KJfQidpiYznzCt7+ecp7QuMCHF+cf3EkbpKmBLvu/vOpCYR6Wx3K+/BIYV
r/iSTQduZ53QNQIRSFgRrETGZwStrXEfbsDOg5Rf1+/VD3wHxskelJoy7pAMtP+1qOs+N1FaPhP3
ftSx18xlMF42W4cFWSeEZnYez1ncoHMFjrK++CP4hie9WomfDCHtcH77oawcxht8jna84/knZGaX
47WCCt5VVl3Pt3/2Dwh1q7v/Xsg/i/0UaV8h+KOQG5yDGOBfpWNipGt07+jHYGNPWxIvyZpQS+T3
uUwAaVwTBgDz6zeoVsIEcokOISvGsfw+fPHKqffcDKUiDbVSdpn/RH6UXbK9gFeUU0tOkVHseSr2
w1we5fwSJZhJA2pSy8fW7p7RIx6p0eTq4r5MOdy4CDn7l58qXvPfknMuTGQFtzedc5hQPUn55TrB
C0/n3ynjnrnO0Y+Fpz1h6G0xUC9Nh2P1neUwxfjmhxtQalSP/KiwTxvmU8CJjKzKPiLQQw93Ye+W
EyfS2AY9hBpMFoD9AAJqStD4petf09KijCwCrKBJQKqG8zU6ij/ZjpwVY68fcjuWyKgluhpd3G7f
DRz/dWOjBEJ20dQtTaTfEoRlM5BEGKRNGoQuFvuhK/PoNUiKNmwgt2xVWK8n8zfqFYOosS93VXwu
PN2h4gKFg8Z7KsX/jm2XYaifD4QESE6HIi20BDHu0tRs1vNSLgayKe8yHG8uDO2Jcw7JHqOSt0Bd
qReKvbJXLk4aN8Wi/gVx5GdvC5MKDrOHJntwaM340SgZ+aR3AbbtQKcsxMzy5e16k0wbtWMGBxJf
+1RMKbjCHhKZj958lC6ITS9gBLowyj+gyHMirdLI3kfIEi4QWB0LM370PuWFre30QaL6e8asUm9U
b1ZC0GdpSBoKjhHsMuO0SAt7mseRK0TzkAAUprJaax6EEIrUdHM/TtD0G2HurZMlLaHruVa8VKHL
jMxREBpt6g6erf2iVftKqoPrL3TCTBAy32iMAaYi37UmMsreO5wj7Jjf42PeN35DvZN4bkOveOQm
T6NdvTf0uSqkC5ljzCY8f3pJabZrxU4ucrxBJYApcLHx0dflnpw3nwjrM02znc1+2PZErIofzk6n
vUU0TjNicwVnw3weqFYjerda5+bs5ziE6uEJsmlrvXEqxP/kHR1WxfP4HKFYHcSUFzCEFHeAjPvC
F8ydR0VtDW8gOqve1KM38MDkzss7kITW92MYWFRalcuIcHduMQVE9qj2/4LOKiHWuFi20IpjXr32
wevRg3MKcWuOjjxtN1Ef8vrZcQH+avafdDkSCd9JRJN7hQim+uRbBhBPHhLm1p8WHaBuomJETZbU
1LLnn0LJZnd2+LnWEJEIZNrZt4nr7xEJFKAKCl0WNttDdJPAd9LJBQs64LRnjh4Fx2mEb9bob6q5
tB65DV5X1LBIB8PohnIW6ThVEOsg3jRte3ZMZGocgYeqKQbATz7oHkgpmP6IyvIXrkCqfoWOLt1T
Vd30PXR8s6ZRgFuIDjA8peydHVRPDYHRKFWm+xTVFsmFUikyWR8Kqs5mXKcrsCSAlZgb9BcASV4r
lNZEnDqk5kSqaEXNP7qQDoh8uJ1SWy5INxG+CzhnZ/M2ljJIIe9SAQ4WACPVfglzZeTCbF/DlfiK
Tdo8F57mQleouZVGP4U6VQUePOfeYdVdeqWy7kaQiom6xAsLcIpxH/WdDtaixywlKdYg6oM4iuPh
7v7/hKBFiKXMdxyT4Cux2xRYDFSq4CA6J2Kyf+TDntjzEMvIpYaXP5yBiXcTn5jIFTXJ0VvIx5fC
5m1SBJQZ1DRKL/VvPcrTVKG3EqtxEZBaK9sUmMMml4Fz9HXbYJgwnEJzthzbvtHbesCr0+9bjtX4
vHNjsApSwY7wc6voWgPmHSI+ootra+wrwIs7mdil9Dq3WZHvO0UyzKiM45JbpQXVrc5+krVwMwbc
TZrFcfXj9VbQJLHCY8fUB+L0cczcCgKqCu76l0jxd2JMYgO23/ZYdcpJniDWQ3r1DE/qbp+k2AlI
+DoBVVy5Xr20vCzZ4j6+LrAvZB/AxLIggeOwENNXROo7XhArX1F4ZiEX9AO077405GU+MS6/M96R
nbbEl6vVxYtDm1G8ugbnGVnbOW0BecPH6ajvaZ2bzy2+dqGUi5WExM/qfNHlMvtaElSS7dkQVtwq
gA00UrivfNb24J+zGDzeVP2OCB2tFIgDnl1aGVil+Lg+5hVhzTEfsCgH0XrTTrSlw6FXi0DuwrxO
atGX6OqTL/gJKZTJ/knX9bL2QeImoj/bCRZxBNeRu88I+is5h3YeoHdaX+pdmwWNy2icqGgyfz+o
+4AB0Gg0PqW8I14C9sLSkXCM6rvisA5Iq5bHEZE16K2YS9apE5COrFRYpiTusQ858h1NoLd65/E2
MzN8BkEgmAMujqYrNS2cYgVXMOOmiv5Oxp9zoLeBUt/PxyXlMqF7N/LT52N8Ljp7h2zurYTaqDqU
CrtXKTMdEndh3l/7f+jmwpRbMkdChpoHW6HHMsDE543hfr9QAZ+LMeFlIEv54TN6azGEhyYtCzIu
gSV2pcXKFpKF9as7QDx0qF3JT7JglZz4zSU5YpB/v4X3xngiKUXc+uDiNg99dGrjN337nVAB2oBr
GHWOEl8suZ5TDT9IfQu2Knq1ROaQSZMM9b8w0dZNhapqwRPwU4Qaf25jjQBDdlg+YYxHVATwd+Lj
QJnS2wBS/V27AUWs1PhItvXECMyzNUf2K6JBIxceC/9c7ZE/2M6vSjz742ez6RpOaOCS84b8hDLE
8Z8k29P3jyD6K77wk3ul9yAMzV3LI7kmxnuXzigrkyA9A+bWku5ywArg2m7aAjph8mPw+zXQx530
+OJNVIawYm3AT/fRMM1qyAwDzH90aqyRKDJkTGgNJqRtXISBuBAJFJU3aYpBo9bwjL5NDDT8zs6T
bpICak1XD9rZLkzVhBvqreRC32/SWoYAF1k0ooyWUxWbAuW021kY4XnojnobFWYq4AMnyhRlRgSD
qOleVDrYf0cuXpzsPGda6X05ehVLwNde88ehAHKocQcISJUd9l6LCsm5xeWvWtw9iqak7oAvcknl
WCj+KhDgElMfTCEuArKptTS6aCsqEBSO2PKrT81tkL7O898yMCaI0+YVhZlaAsjqpoYwIVloXjNF
iN65aSOk123x1kjg9YIoWU45HbAHh5InDz+T9UQeWSUgVXuTyDJPZ0Lcbw0PtWDRJ5fGlVUH0D2+
ojWKbC59zrbKNCoB2FV4iWkDWAg17m7lq76FuE+fZGexC1flC9uGx3ZgdTRQu/utvMG2J0sNeECA
HbJPPy23kH1RMaPw1UYUHvgQoxFHG9apdvUcqO8lPegJbxImTUyLsrlfSENtx/wCS5rsRNDCHuSg
RaRhzRuNncYj2AwKUo5/IdfPxI6cliw62j07rMGnKSX5ZKCXBoGv8bhehNDrVwfCFzUAD2+sKQKR
P43wvyA6NVuOM9Smr6ViNK3quRReYYxahcqDTnxn563CIZpCIqq5GOLJov/D3I2M3Wy6PWguVvtI
MFacN0PvTMIJgGUp32W+qpg6wOKDyec6Ca7mE46eoJKpCzGZ39pPk3NxSW9pNEF6zt7iPOFp+P92
6Z6IY/RR5sF/Fli4YrZ0u+jTj9YgjQf9zDAqokxxKJRBltXs3PHNDwyLrXUYGkDi/tJ12k+2DnS/
lIOoTkuL413j+O/h7TAchO3c4SjAyBajMAvoqHPi0kk65K1PKZDrYGkN2Q+q5VWlg1BtGEufQNn3
5MIYr4Woyeikw0qHne7lb2VmypnAxnyiPQycFR/EEyuacK5KhqLoUl19bSby4/TFZKrZCbRj8uQW
dw2QUc+eSxaWQ3+KIDMryx8hRxFUa40E4N8f2YFiLFZWimdhGszufQi25SsM76UFqRUinhYNXXSJ
0LJ5iZIKa+XmWhhcJRZaRWgHmnGPmTiY1rLIHwVRG59kSMd8vi8JVzxpK6aNZmIanj1FhXIFhJ/2
w+ZfqpQslemkBIXof2ki66Ls/LAGo2fFJYw+x4MXVSvzFMML6/DycObcfJCKpBL5owIs764gFtYd
zmLWZO6ifo/Ay7eVEY8vWLHwwR3wJXBRb8AQ3axrQpI5LxGxYd9WyE9PKRf/L/GhEZpPfSx7GleI
XI86nmJFigk+LxhW2FK2nQnT6BHg6iv5iDyXc0ny1B6hSCJaJqM2hkSJXr5oPu0MTiW85BGVG/ZL
HgSy0mXZtTHxlXn7vt3bty71IxNicTYNoIoU1mNMDatylrQzRl+atSjifgf8J0PhLHB1HC/o2Akh
h91dentHdfV9PuWBt7jqHOytN0B0bNHKnWEQR6mUtHajitNAQyNWAgPk23Y3bJ7YzG0LYFG+SSPk
1Khogi9ZhbHyYzxr+ME+wQ+/Rw0Tqn3QE02ikIsS/beQ9HO8OCS+rzNo2Dod6BNqQZO0PKEfKBQi
QXIwDWVZ+ny37vfRM/8aDDuAFgwqWabs+O+/BT9rbGz1hNOH/dYx+uOhTbmFnDpKHrLRoG8UP9xn
0t7ewOgmEr6ilXzSvPqydYON6p3lZrJsh35fEG9fcZwFvfTCRKJPuyWE9tQv78ObMKQbe1afOJkj
y8vKlZTr8nYJhogH5owveh24tZVXEs6fIQFT93GTjoNG8Pfx6sH9jPnaLtZrS6EyVY1skCDuGNSb
W7W0FrV9N9ewhh7SCSMebHB8i7xHOCCEzKE0arfMv40QEzwMPfljdeDgiWNwkOfNMVc8CFmSxYMB
DK0FOIkNFCo9zW7UlfIBvLpY8N/5IvSyoz8QlsuTcviqp8m31rTfTs8rtvfa5WmDN4juhfQ4Kf6d
IuH+k6n++Mv9zugaaqwKEndDlPagcm7saOp+KE9OxT4uVOSoPwpWOdNNtzfO4AftHzWUvcMJpMPj
YtYGv4yCQKf81o6g8WdULiRgR5kCr4E5jv/zGszo9hC0oNZmBAbcOXTlw5bZMPUaihI8PWlkxlGH
o7bFM8a6u3l1L/kJiJgkNxRepehDtG9l3W45PU5NwNeR0751UeLZ4KzJ+FpeEFlj5xQYhm7DVFC/
FE+OXQfDVYTilwmw8SaYnfLLvLbtkJZfoQcwWBwIfRjZMHK1TNO8T0/TcCbCO4kgApHLGagb8xBP
H44EtTjbOTh3iuPb3j74ohjKPgbAyyH4p9HrJ950Qc0klCqvgtxcL0Ps5jZ87qobKl19fqLiibkk
65HkZTzNibiCaxOda5YDBQP+ZVyc4YTjBStJDHL4IpyRdwD+xByreLD1MTHfnUcxN3Lb6YSguWpt
lBXqUcrqDMqhLciSGE1v+gGRXQ6/zT71M0nelIdixe1L2qRcqnDRfo+SdIVwlM0cJ0mmzHnTYkh+
30azwEWb1KHVqOVzj84v5ibN1lDMKJcOROl5AQ+4Qy629XQRBjRmiB5eRw8n7s7M4SOH2gR8sW2S
bim6NHY6sqtu5DTExpUVLT+i8KCv40Ok4+owEP4R/NmTDirdup24X7fwwISSzAtLD0vFIYuIWdHO
pb2JKQVNd1rSdxIP6k92jCWghVunfaNa9ROH0eUjBpYDCZi4fRFlNQbIJVlkEOnReIgt4nWPQqHD
48tDwKpSmv5wQfVVcboGhXZ4VP/0yqk1z/roJqLBG7zIn2wA7YKVFfz2NrhWCg9PseBLOZkE7PzV
p6SEKT4esE28RQfpVAaeVOop7wkznuQHFV5aRWYxUAKiNWH2zEdYVBLx79gtYaEQgXItx8dkwq43
vstSFf47pHtG14IZIjjKdhbubqKhhTNGHDyY9zyWYoP4qX/in8d7VXh3T45dzo+8ihJjyVYfigzJ
YxZM5rwdCss+Lbw8x33iWDVIqPgQWPrNriSX6+gQswMx1VzS6XFeYyKaNJ/zKBIhAfelZGa6r+YY
njj6wkiPJ39uZS87VVNfTNSJO7S1cGbpIn0MB3Y9skdCJxyXr8YPu+nYSHHHqw7xugs/OKPTTXTO
q5V143xJ0728GX0m98qr8vF8vQQ019q3fmKigEkJxaqPPCoIb+gIHjroxx3VK4MwJZ6WPsNw3uyw
06nC/bFv7LnrV8SG/o8Jbcnah7cYtrOxPghuIhAwaXq5N5EYWP25oWNu0SC+KQLgC2wfiM1MCOa0
HC8443uujhMCtDZKnULoRytahnQ/+NWfyOwzQ3NfI5KOjYif49EhS1BHDg/xuT3xWCUcxouEX4Uq
0rjecj174OMp4xWT72/tfaM2Q9ZBtUiOaRb4mECrzaVNe0OfOgkKnRR01rMgsWtrt/o/cy0nd87N
iXfluwi/g/UuCpwoObYjfeEkwRrZnwW065hJDPd0flbg0ySRCfbmftvQjQurHM5y3d0NjhMrbT9W
rdenKDtYDw0KeaMOpVD5y88Zep2LfCHLzHMyhhaujVHmtDMX4OBYeRUhBCPLkJb3bn19xP7fRhY2
GHpp124HNaQzEYukms9xDikwMgfKvKYbx2ctxZb9VqV+gffwOtJGHgCicEMH7gIHRDJ7yBHSP9sw
zSEnWHenMNwJUCfHObrZjW7r5NCOPuMdI88wHBO9Upq6U6dRf3++kaKXpEeoGy7Ky+L6lAtkAHj5
D4xW6h+ZQ71fIN04F13e+Ixa1S7ZnZwct1JfkUEggbpSEZLSVYVa8fl/wAVcIKsAfXDrgGXfbEQc
LePQcZewq65XA7sd0RAlEIvIGjzcfycfxGMNl56clI2mLcVX9TVkhsJHUFs19jiEg1DLivGlxVzU
uH5TUL01NnfLaHP9YV/FXwbfv7NkwuEzca8Qx01BL2h9BE05hIKlipzWPYWUUwgFKKWB3zzzCXjh
JXJUukq9zJnEBxifmP3FtjZCLLSoPypa15gM4bTc9JLWDx1xX4X883iWFkkQvXLy+yoWAA0K+UqO
9IwMrBR98UguYptqe9RIb6/iTa7qvvlcuM43E37GaUH5NgnYKZyEttfrH1Ni4hHV2eASN7KOiof6
8PSJ6KREXxBmMtr8qDp2ph0oQObNLCF9IhmUqVRBoc7nxGtMxKN4xQTTlhMV4g4LmxWTAeU1ylId
jIWU7sn45sXSYHCT6Ih6CFzSln3LQELhv8kTkeGq8BnxAb5ELTHIZzcVfBIn2U9BMlZrz8EvBkqu
Chf9/Xo9S8e3Yu4s7OXchzw7lNgmX3we5AoQVA+wM+KME1YcIMSHUP2F1n7lsehaW7He3ZSUWC8o
HnKIiRSA4fNwLytD5JrJDBJdCHq4xAst9FB3I3gFjXfEvpU+juMQFhUkZdZkt5xA/Bwo2q0StV5y
Clu7xhzDgx7/zsgdANHZuybt1Zz+cJJI1s2KE4O7/DAQTuV1NMpDLt2PHsMmIEb6VjUf3xn4xzFB
Qy35+jno6gqaQujocENqbtFoL4MakL/QPbrF1CQP7DHzXKpNQ5vZngVa5H/xn1z/4vAjlkBe4JTr
or8fvXKLOWFSBpuJvqKLm8xxUk63yYhbfoJ6PNsjFHPy87NodTodR9+D7tZ30PvJdkEICmDSnhe/
bs3FIny7+JYIxvDr/Zc9OUVToXQthpfHmEBf6/7WUhgV+uYp+ZeT3Y1IPATMYHCgMfoB9hBlHH2s
qJR7qemBi5vHSTr5IPJL1yp/TvbawMu5CyafkaEbNqRcxVbDxPATdYima43ObZSApMbOicR6loXY
tBh/tQ/VbPAtMgDppT6BTusIjfULTAAz0ExLLHk7DB7Pa9i27OOn3EhOQ0LkRC9bLSWhDXN7aSdH
aXSIEQ02sZXNfG0PTjVmeC+KyYjukZz/MlC6YCCybMcMQAjc5a2MQgQmyvUohFGWwGAlXqSLBhYE
rFGO1Ggx6Xk/+q9LQ+i+HOnF93Sba7xcpSr78bbWX1dsTeK0+6eRv6mOdPiuoxMwe6rLOESbQ6qY
zyRJzdKeFkCSZclKpx7Fstv33nhpntPGILN6rYxkF3Q0OXv9uoo6mO+kQqOPhginYE32ilZgt8L6
mCdzmbJloovLosrg3PEDapSEidMImewtV51SeFNN3iUlEYJXNyMlWtgX5a4O24WUcSRu/eMy1nWN
DckI77C/lVShiGlq0u7Pe0w/jxwdlYEGGQXCvMZWyBKWbfq6s2VoyKgGrkN7yHDqXN02AEBX4r4+
OmfieUCx3clP7ktPRCY2SGob2lon3zSNGLSTCP8bNntjhMikyeSr//r6KteJhXIq3JERWxBULToQ
bLzNbDzUALzRqBvBBbx5+P5wOIX1pZo0JR9SsMQH+dUid/6znOpY2TmYbCiqjMc5jzIOql7MI8bP
UQG39iu4+FZAQAbtNGFLa0SJJ+Nyyp4AP1M5YnGzSURVRkHleRCAFAZwP2xH6nkmqKqCClj8S8QG
4JelOMsBHZv7jdcJaUFkMVNF2UexfpiBxCvcycHPV90mHD1OueQs6uyoStAzg7U5BoxlSMPzjSDL
v6ofHu97dR5rEVAuX8e3TYhvvUw11n+jQEatAL0MbX6h3xznU2pHGz/gHtTkEUydtdjCd34N9r9B
vzaeMLaBgM76ROseDF6nucovfzENYzFQYA6+Q7hvYdVSY6fAsNJTccw0ayzmDyjqFo9b51TZ6Jfw
sAqvJ04FiZht8tE0v48kZWRNcbTRTPlyukvZr/b5gVB3ZGNr/bzhqOAek6DlCRYVmW64gh/YoSXB
iCAuLLTyW3VEYVDEjm6W6DbsQY7sIPRhm1qsrE8QJXpFpjC53fOayNu/etFQgNasR57CxldwScMZ
wRBXSk1r45I8XBeEkqsjiiCVXF6BHjLgItVD5x4FmSzoBlbs9VJV+zKuz4MIz32oTi/JIG+fArIX
pkMVteV4znrB/zvCZ/DI/dBgLtUYUG25zStjDsECJbzb6vqu+IlzuTotDtl8fnWbZ4Gew8lU/ndB
RNdCd+0IcLG7AdY4FpwFdfFb85/K/V4uZcZLXxkSLgEj/wvPQQpBv6qJf8Ko10Ozbcsbk971lHEP
D31f2j4j/vSa+dBHRrzjjuq/DGQNjFGGk/Vr80dZ0pQKjDKKeF4YdItcw3cY+Fm7hDUiu9gH67Wu
9pzgoa6Q2I6uHJahjcFVWZH2kUEXkhnnwvPP7cFfkZkD7KGzLaZM3o9C4ZGcxyfanR25lfyePeew
7XYPv5WNe4PXF4fyNlphZgcs7olRtFOcWFZc4DvRfIo0Sc7v4p/UXMuVstELNwquQRbbuz60+4Vk
PzRQqB8MwHUZa9V/C63yQHZO/QIGIJXlNpChqTgkjXzAh5IaVoBQNokYQm05+ckncd92kRiq5XyZ
VNNe+UNZAOorXLxYU9iJN3ufYpKbcty0TfaZSGSOrSW8oeWL7Nu6wG+vv84ghPlp3RQ2KDGijmF1
IE+Ng+SdvFbjiglYT9ZzNiPBJ5Q9GaPS35e8LYM/blpx2eG5kCI4bONtqJ9tYa2LyWucjTL4u01O
Eqj7Jk2RpXyiBPY0kp84yZ46pHxyYBE+hP3KmYAd/JVTyfNMU60RbQ975/oGaA3z3ktwWA5HI0Yp
9/6SKT0wbF1p59m1Vvx/JFKkmfRxqOX5/pt30PjcilP0idC4xIBYAqnNh6lYpg+yyUqi41E8cnXh
OsD9y34B9HzhNladpjL8NetyPRgoso8H5NYklXjYkBms6AQ0tLEUkzGqlf4rmQOOFhhrpKrPYWyg
AVSJc+i7HHPIyDWfj2oKUqL6t5FRlDMDPMhz0dI+vgMU5SuYxG09DH+jTIHcb3xCxY9BvdagSvRQ
H9jCTKVrytrA6yaoaoiyct608oACrLsVrEK8FcFFCDweQlAjNB1KJTCLc+HDg80KZZh37cozrCAO
tDUF+pH364vZoDEleu0TZdiV1DthKBTbkObxxhRECh+mnSymjYe0EBfDSJMqq1gIYkodoEZqhqF/
JPVCnVmU31FwobirS4yYCSK8zPJpjJMiFNrH2YOl+rL3W4euz6qziLMgWrK6E2BWxZ32dpjAGQ2I
B3o4fUdJqMg6sH82foTGReXgmXQqTcQ1M9/2/5VHYOAieWfseS7yJINNWkegYUtRRr3avi7PF27n
xE3wjVZMEJHXlXhaiDhuv5igAYCy4+gD4Y+eZV6d3zd2voAxDB/vtbSKEDVPBC4gWvIDuLPRpZzc
ciB0m7O+yy5EYg7aa8i0K33Zv62+qJA10DMmceA2DQOqt5rqBVEIeKeVpqzSv+CC0UoZ/83nDdij
pm7QWD4+nfBl+LNQ61hAl+nH8Yo6Askf7qD+DMdFMNY4R4/jcsydJ7wOGsZ5B/P1N6cgJgkvjt6v
PmiZT+9OO/YB9/PXFKCf5yIWQddNw6vCRGiJwNcSSJb5U9oyie20T6yQzvSrlnI8Cbk+cWVD8dt7
onCWtZgnmqu39Ep9vo8NyB1KLEqM1xpW/Em8BH9Xn38MBVBKMe5rbOFt9ndCRuP3Gofob4D0DfzL
DtmQB3Vjm79sui28sGjM8skS7ic8tmkOs/7MEsUQWEFpWgdKp7od/ivxErw3AviOkQtrmFQDEbEk
ebaORbEMmWDoTZ3oE3n78t1skcqIXjrq7Fzs6+YuFDOV+0Lh36NhWWJ86x5b1mrtPOqi7LzM6tAb
jSwknIKP9v8J+xJ5KPjqkOQQw1WH637gwISIT5nd9E3P/cXLfe1v9bjhXhIfjrSJX2u4ULODCoSE
pmMPV7vpq2rFThFiDoc/WrHzS++zCLxU/kV+oMr2zrRqQ/llL0//eIuYUWhZyXX4Hufr+sbitZFG
tTW2DfLElkzQBqjrPsOvca7A0UjUok48vZuTmx5YQNcQfulblayy5FPyCWjVmpf4BmaJ64keOopM
GjBmhrqgHdYaqhZf63VbUTkzbKbsiD0JEgQxzbKHnZFthW51h3WQ2hwOXXN4iIlrH9+oI724hQ2L
fOqBCGenq5qhNN89FHvRRf0KFjhha0pQ9D4z3PEUhkYW4kYFZkygoEGQVS0c5ulLJnV5oSWHwFVq
KlcLM2n6l/Iy8OdDLaptmXxCvi+O9YLl8sXZU9npasZLhKaFqt720EaAiu0UX4pmlVUPSL3QVyO5
IfSLOmKEbw5KaL0flC811uIVt5ZgmSWn4fZr1dRnQrtt0riAFeysfr5HPAp9twrStPkKNuGiSJ5R
fHckJejJLlC46nKc4J7Y+wOXtoY8lwDMXxtYHZo6ADInA/EoJWqm8Q+5p0pwcMM1ymcCTdgo1UY6
ctmwWlv3Wch9Kbm8HgQ7s2dRBrx8RunPgzkKpqWskjUNjgABmislql2Cw7XODMVdw0H2ru5wuFl5
niPEj7cSjaXkntwWYiQ9ozuzNymdJthksAl0mc575Oa95BcjWnIy49UHtEjsFTWrCWf9z1plF0k2
19KVLeME6A65kAfr/ZKhDhISw0p1QsaBDMk3yX+yXky4gUYRsTgKtF4I1LRbuI2o1OrK0PLYBuGv
lunojpaVY7joWaZUSHjO1IFkeFHoEbz41gOMnvRks/oN+kPRKtsRYrLM7SX4/4tk9Qao5C+oCkhk
BX9L7gYjAdqczBCaQ+NtVQxXbAgrdvmpMW8yOeoOnLp4zITTTF4MWXV72c5RDX2qrL7/nmz4OPSt
Is4bs6Amxw0ENAtP7rMLlZVi6gRDTarAAQh/FG5bRF/PdBkNiY0Xzx22ka6DLspCgu6DM+8DOIt/
KqhIh7e7gId2Ff2r+OgdCQxG4X1+iPOwnPajYl+b7msqvZ+9xtYt4W7+c22sxu/KdEsA+IMy7r2u
E4B2N7H93I6Vh07jnTVD4apAmtWMoUbYCm6OOcVjLq+GJW1Kvip86dUP0mwJ/1JFhlGGMrmLc0d2
OstjdxiPIbIuD0KCRPPgWktwwOqcqsGH0MIE0LyolviDSCc3O2gcGPXG63SsUs7anKF/2kjWts18
oiM5qMmJduKzZ1i4oJXfQ6HEKngOqSg9HSXulcJkTGGNyKM6k7Uf6lgQ4PQU10oyu9q0sXG38HO1
vToC/SkUJ94OZV0u+t7d1YhqBrADEFxJg25c8Xsn0Mdl7pzEgE6XxWEZzMoCNEFffIIvSYfRE5k8
NbAWSw84ZiuLyvROpjMqJsznX7qmevtki15jZeULS8xYXQAvvi80eqJLtIo0D9sRHcCI7wz9Gp5S
lnn4JMoM3AnQO4d3URhC7G4SERirceoOI6l94R7vT5XudfaDsdh/bx4Zskfog4U0ev3SuzOcuHSF
dYMmfAuWpHLLfNVWT/RP5+5McWMcl2baK7Gwf2hExJk+4vcG3ROX+8ZmnlCyal5tIliNDAZcqnp+
AENqXxpAY/Fv+jNFUdz43/5ZiagJ68H9mjLdCRV30XkljPsiRjt3gnIoq8hlNUCs6Y76qv5zmQKa
Em8JZDJmtXDMO9qRRQNsvi5Eql9b6bzDasi2HFBS/Y4NbyIMDNHX9Y8ZjBLWjeihiIMhBQr0gPrU
0SPoHPUJ8PBicj5BKJFzSnT6WQWohpg8movNuxtbfPM+C45EBKOVV9al8CpADJAzM31MZtciWCR4
21OVyRX2GmRMuYGyYz4p78CBmfkKlY1p2zOxF0c6pyPXn84Y1VD5IpkUHAj7lCUrVq4ENXonTxMz
JlBatktkVa2iBm8WkTbi7CuVltuGKQIzPiNT3n44ZG1BndtdCTmeleT6aeSspnGUWLNRvnfRisg0
dHJLZ5LCrVb1BPobwy7n169SliZ0J48gAAzUajriPtS0Gs2IjBzopeNwa8ltOzD4XuTjqsQeVBlA
+WrV2nPzKd16UtHnxcGvAbCQtlf4r43/YjJfvaU1OxM7an4eX4h/SO0GyCfUGkVxsbATiwvim7ib
tX5Q6y3RP5qSyidwV4NMlXq56pMCqcAaKWUMQkeS65CPHBSrsFtYwa+NO9Eg9NH4qrHpB+QpLYuS
kbloOrDxjBiBC99RrZh6H1ofa6eWCIVeVdG8XzTpwXeptBcwGKcGIWc8c8GrgbV2cbFI7SwgGK2g
GrhGqoGvwbROggvrPQrM/Re7KPpYzzncafOvbuwqeVYCKr9hdGEwMFpRTn2ZeQrfqcefNoRXSZhP
TCM9iWiuA6ziCoyaGmr9t+BY/H3hQkmjF2THIufc+cDo1t++Vl+RbFzrM/Z3U2dpMurauRxHifaO
dhREztFn7mgBVrpJjp9/3tRrAcpqZ1Y1mFq1AE/PyMR/B+anqndXyDGp7lwuAC9B6bB5LKB0HcHC
PunsDJZ/NqBEKw83e2mbEpxmjXQlNb7bie9pAzv40ojhwfxHyQRa3bdRWzjVrt9QFcaOltptc3i0
vV292niDLCaeemq8w+yt+tdRc7iMRmk/kHsuLUILLAUL5armn0h79iwytm8/oAnY9ePZihzD5wX2
kO+y6Usl0SF2oHb/jDIvXOWxIuBZ0IVO2ZX/UKSr0BI+wFnRO+mjdGKAtvBsos9iYzA2OwT1A1CB
Y88IzaLv2c3n5nOXHqV3D11jjEXIaEkD6V+5egQpfPEr+4mcKLUHjOkndoI3xebQi24h/PVlzSkq
YCMn8HIepLFu0wGYP1keYlag7D8RP0oZ7bfiQ6C1d7i8ZwuIuVuT4JQtDNBM6jbP9LHVhVbBdYgW
DRjaASAX+YvPMPaSxNE9P7mQpNKdWRJElrCGKqDpZ9d2oiXhDgpU3cJ4N1zrJsnVVLHpzQYZwBDB
7iyVM1pjSxiAK8RhUn8kJmi6L7dp//F+TOP4y/yreOj76hM0PkeLR0Kz5rV5zFvcgWYWZq5ELPAO
ml5ZVE7jsKhM/0KXOaqKdNP//W2yUjGLwwvv0hkyZ1f9ruXjk4LZrPKq5P875yyhy88+KBczErj8
kY+raskwQeUcFE1PKoBKG9DVLQBQpU8qeyRygVASQklowGzrm/fkJgQCsAkCxIjir9Yt35c9iUyr
jmgSdYmFcIujYKS/Ze7lBuU/65MkwFJ+g+yRt5s5buw9G3+0eXaQWCTv2VQhIVqvMjgtFHOmO1vS
97UMyk5y/cmSDKuoGG0c4IgYA310hjKTPFqNqlshSnXIlSRu+i3zfiNwGpXUbQmANLccBGJ0nS6u
2DbDShQoN9kXdIYCe2YTruATJMUqm+bzeSmkqFddAIeLcYymlTXDDpn/adenHYOxwW3M2868kVw5
yH6VrMvYE0j5yPH/v21VhpzHtpFv9l3tyjk2VA0Dslye4EVtuMURtU4HzoZYZHhmjk7V4ZUL0sH8
/mBOSuHR/Gb7yEt+3jWohm3xUyaahCh9U3Nobd+Zry4mkx7LtZ9jsOUs90ZuNGImrb7ALeQcnSAJ
5fO0orF9oQpx2a0L4ikNXS6gppg+AZAKwXlHdj1gdCX386rMFRr7vQ7kjXbR5wAuOc2fqAtPTZzV
ZTcH7amocJpSoSHeDzD2rN17XOm2lQZ3DmuGj3UxRnM09pQE611Z0Z3qNx3E2WSA2eJIyIQXOWIJ
sR8wagiVwW7FfFsaeTaJUt08YtHMEXeVgKfpLVO4QD4dYboded1kA3z7Avtn1ZDR8KbzoIwMcDrb
KydcRtWyPd4U0jIdfoMSQBRY2ORNwOA1/sKr5KreHRXUrhIyfO/L8UyeCizEnNU21CforlEqiITE
7G80kAKqt+SKMwNI9lhPJH3AVsq1XJaXZGeevEtB7EXOiyCzl0VhaiKC/96uPWflYzDAP23DxjeL
qQldWqRzhOgmOttxCeCVgI8S1uXdU3qVeQJ3ndBHDo12SmwiriT1Wxv6K4fslJWYX9sa2kOVroYS
ZBL1Nk0qV6rglvc6hhBV8SvOdw9ipheSiiVQlLYgNpVhrS2Uy3mDDNIa/M4wcjUyo3VInbo+26SQ
BnHfqrbP680snDRViAgAl1EKDV6mWAShEGgGLl2lVgBC/H3xpqBQ5rwH0PSiCyOonSuIaAoD6xkM
dqM8xXIkadEqMmZb1+qhsTGLw18pw+gB4R6v3JgIdTq+4Sq19eM6phXKMDvwWywqt4DCpRAsMnPh
lFyz6A9ExG5XaLh2PxWfeWA552ZhfjRoNJZ4/0zcMjD8XJz2hxscNGpKBEClGDK11EHKvaF0zXSH
mR3I6XKJidKn2bjq1FmMOHLbrt5Toc6CBfUaOEcEmFb6aOWc/A1OLbG/3/WeoLhCq+ZNDrQTA+9j
KGODhjbKNKdNwmzvMul68p7uCZE9BWuegFb3sMNFFGrEH8n+4GWsBC4KBw/ChYaKKXcNo+Ur94zj
kE/+geLU0q96wQ59S4wWDy8zQg0a+Z9OOVi8+6Cid1WoOlVYoanBTCcWX8ZjbFqNEXUvVNWsVBbJ
rOpeuoeNyiAJV3Wh5h8e3mRnJ0K8bBfz1PO62KMd3CeKz0pZLJ97b7RGTQTTFZ9JXainUO6wPvSq
C9+KHQVdswr3NYTHf3yL6fp9tKlrobq+zOZLz8nGbA50o35ZnDfCyldpvjBcXvBLqN88HuN+SXvT
9qXxgBUeLHd2aCMZttJ8E9u121NlKFCer7pKcbntXZhCh/FjA0OCB1JB0+1ntxQBv14mzXmdjzXR
Z18tViDz/UO9w2SB4jSuf6WdsYhHoLJBvttBLWmJQpwacsKtS/7nuy6VuOfOtFXQWK09TNFReuh3
HnHmkf3Hox/yriIEn3JGaCW668E1AHVQy7yFrT9r29vNFH3VTX8e1HoY5K/QC9NbhHW22D0BbttM
g/YtXCuqZLLb56lxzFQoF6o9NRgbMMRyzc0ZvKXJz3jcY7PxpzL6I4ZGyXtgHjX723FirhYsSAhK
p4yaHtP8ST/lUAei/UomCOtwuMDfpXPIrvucm1qMEDBD0EhgsgsGe/n3n+1WiFKFeifxCpeLbCYy
rsHX4L4BwkJB7N4dl398TucgQ4yozIJxeLFsbHOjCF9JB3PwxN1bTt7qvEj3KmZq143k2IffYqJF
y/zOGJfQgwjZJkZtD1zQMbRiL9RKyB1gzzxT8Z+lquju/89gcDeXmkFVoaZ7YpshXeKcWqPY39Ov
vOuhLQuIoW7k5ltGB711aHaKOnvQf04l3hnMrCLYloNdw0w1hq6DzHIBgAqTpXT8NB2BVBFNqFjT
ehubTW+RwZeVkCAcVhZ2q5tISHvJJqQ5otUxLF3c2fv3BVtV3OuT9TX4oUI9ye8VdrtHduv/G/9v
xgob4TbEAyTEtHrIIJhQsxb1kiKmnSFR5LU7Dx/D/4AwS6UpqHpXADUC82V6xdlZYoNOaoLyVxce
AZEdHJIUbRHR4SKDhKt0C8fcY/SOr9OBMcgkjioFc24RjFMfxK916fgJgT7TgicyGW9oaOQghSOQ
yEIJuAe6amhOn3sI2xVs+z2Fna4ZwZPoBEwUsYiOjzdNuzOiasV1Qs9tzsXRAWwpkmWNRLIszIlq
zCCalKEHJLcwrNAURceBP9itk/U1ysx8ho8rqVwqqN2L6ikq4q8Q/9ViV4XsQwpjV0MtZb3qImGh
2iuiY2EnuT3zVcZN8ArjlswEgs3Lqj1Q42MiN3kukXcjXoPm+VLxsaS34hpVU5OXieuuDqpXTGkE
u2FK/GPRgez5XaaMqooUEZTRJxZPB3Ux0g1ma1K0+f5AszfyAIqKZuuVazMMY7j8bKaS7JdzWhPh
zJgCsrrLovT6Pr8vY6ij21jg58VztS3IDJirL0LrcmYdScLsuOuMbK65JM2AYxbfu56RvngOJPpp
Wy8h4FjdpC2bxtxcpBZK7OQmxE0LANngStr9pPDOJZKzLxNf7q39E6YK1psrwIP+tj1aOi2Duy6s
4Hwz8ncy632yQ9hQtAnQafNfHEb/IaMe/N47YoKLemBitwfaiENElq4EqvCho3qitF+l1KEFywcK
tuX2Gg9OsOn0pF1ikeBnv7rM7H0jOmAAImEzJqgDKrGGaicvdlQZqWrbgQ0Mutd2VSOtaxnimPYq
vlPgkCJrJTtQ06rR7J7/uHYyxd+jBSmmSz8/5zBtKyXUGKhzWh5Ov/pfCSpv+/d6L9/Tnc2Y3qpP
BVuBOWyjzvPg8GFFjU0eW7NHBBS8JymwYwVC/WkghXWEFWDlEozadirZKTdiRD90NCnErXC/RgQu
xMZFwFYnIRVlCD4Lt/8Yb7RHhYJS8jNuViSt4PbN0IenDPqPi6G2JUnz+ll9qfZVNV1q5fbx94ex
XI6eusgZVNqXLXCWdKjVY64PNMIA4St6CKxuKafUjKlpiElmuzAxRATfHijCkpbfdVJWjyImxli8
IAQnzeuftjVVhTRl3jyKj8umB0x4onzeJhf60PVtxBWAuHRetKCjv3pv861qmc60M9l42epJb78q
caTrA4BhTTolF30EBeEmGgNQUeVd54e+Jw4YGkgV71oNKW2wNaK5B/ciV5RYwB5Z0NQxw+jIk+Ws
cuQu3AHu852lry1MsjSEqZceL2qMlGuF1oz0GDiwoi5+vbs5/H42zQdsa38fwPHEjdk7GOgV+pBs
PPcJuwgW0J8Z/wfcGeIkOiOmFQjHlndB/Pr75TmUEksReM1RkQ+4OncO4oddWs3iwCkQqIe0XB2R
aLJd8JPr2ETS3xI34ePIfTqMWYocFRT2Frpt4H4tE4v6+ZYULQ6UKOiqQbOTSnvtCp8jh36BfGh+
PrFSMMKwWk93k2/lHCbjc8BFWG9NjzMPR9IeEJF82RrSNQgqF2T+NttlOOD3WXzWcBWKxrJbHkVp
N6tpBt2dGR5sm6cyuoRBmmwo3QHH5DD02mDQRrzDG3PC1omI64tHr1EJb28HiIIHJyeFdVCnbsCF
JHYnsm64vjPaZWSIgS+MVkN2sIdkemG+0hRvCOJZoBsMW2k+2nXvK6HFAkmMukXG9pCnHbV02PUw
XzL+G6h6fWjuvXht1squhXqPGYhfVJBNglmccSm7S5dEJk/Y0LhXRYdk0metZcfqmYDE5xLFwAQF
7s6MPAN61+j5eVQE4FWH/JJfehlhT9F88BMysbyQ+MiWtas5v+78O0XIXHT1UXNzHCbiDVzW06ih
FcOjeR2xAN6siaDYJsjX6Q5G/1wDYOuf5p8kp/dHLwy629LmPMPQ9YxMwdst8GIxoQvIvpUBT1wD
C1wXikdkpD92mntJuzBGFO2MNgd113ZA380jdK/3+B0nXKPBt6HCpQR3AGyHy1XQyQiH9odmZJQI
y/jCCxCgL10sTS/H1nbL3SHUB3j0Ew3I1zpWg0LHAXr1df+TaZxsOc/Q2rjrWbklH2L3qjfHkFGV
kHxXtTst4+KKeRA1bIquk8tzOKV2ZoH8upnGulYMvKNAntaG2BMzl1XYP/48GR3hea7X6PoaA+mW
h4UhmaSyHiM79vlCr78nf+Xl2LjktgvWNLOEQj4xTfA+fZLfWjER6KOSb6KZrX6YCgkNFWUkgaCl
bpInY3H3e3BC9r8xQ7jYGHPF8MSB1epSsg8B1ZkKKPjRNej2zSEFkEzaIABxZ6BGv18QlsWDUFzY
nCIHUX/QPIstfKOPqiSrHf0Qw03a5yTZRKUG/stbflNiSw66N4XMObaa0kJNcUQ8VCKZmwn+m/fD
e3gDwx41mV4BZfK75QUKrlld3y8cxpRE5coQZyVQGUjVx4uXUjliDAiOPDxWwiq2rrGCQq03jok9
fzA8Bnp287F4+7ukwwFt3AwmNKGxAgGRIaxpXs1wdblxCm85VTvKPVm2Eemw5bfNZyasg7HTd8/l
O/6B1P3aYTEVOvn0n8iSHE3d4TK6lAbgARGQMIEvw4VsvSwt30RvE9AZY2Ywy1qEyMsmm/fdyXIo
ZQjQqEJUfdiATil45sw2kPl20qee+aBXEwopppCHSpGCfkMqeDLGhUsYEr4HIWZiObTYovaOs6+G
Je8TEXt630rTEvGW8SaQhYHnCmajT239OwTnf+2lWkBv++/AcDJAy4AQNZM+DvLJtuqAr5vXyiz7
DYzV6cfas5sZ4vBfCDMIepmWorVnTAzI47/keiZ8LfITHhXP+uSEokVCYCMpewTZAFOnlxfYz1Xu
S6RgeLAvXXgKf7MmuLN4nPfm5qNHFEUwuNvywElFxpQX+lWvifRK+TqSVOFSZUT03ifuiPgvaemd
ES8s62a9D91staE7F8EfsiPPYBQHFpQA45scKJ4EYy4Mmn11M2z46d9hGHLwavIHjqpP4xUysHMf
VYOkWxrqX6YWsEFO86hfAg2WP5lPKI3jmLWN3G9JPbGabXL7xUfFKGurD/jOgX1osw9MujvMifWw
gYRY1xtthgdPDdyxszb4rBvcZH2crF525bPzvhP6Abm/G943Zy+BLm2KE6ch3N+5zzdUtbQFI8AC
fjfVDSiYkNoNr1/ajSf7l1/VSu6KwQfNf6t7OoW4uJmnCU/JiV6Z49/ZkFLAXV86YlO+IQvotxdE
p8iwZ6qpsivuyWUVwB1+lF7o6eqEQC6ACEBBcC3soKs+VcYQiINVXk/Kg+0wMfQGELLL51d/twHx
Cn3D3eo1Go78Ft+EJ5bck3+9i65O1RktbZ7hD398ubcB8lRv08W8WEAxufGuG38p/T7MGqXa7/N8
DED6o5OZW2AsRa9PVqfSRFyppV8KmNxmG3m+ENIBIa3G8mIb8rwBEADLsE9qcA6IbJoZhLMnrQYq
juEf82ifBnpggFm3KtUUxPqG732Vlr/xcb/z1EjbhE1bcvK4WLORybmwYoASwyCRBNq7RA8rJlCB
7N2GsgMi5ZJGEZu3abBMYa273TJNuCIyAtDopQnfJ4e3TikBT1KXEvZCpqn5Ri/GFlfA1HdGjhmH
Hnvl5U7Pstg4QklzMR0YWB6vQxvg5joN5TOXNDK1PC0iTH6R27Njswogh2NxdMtMDq8I9rhgkY5O
Ahr+XOoS7GsQrMGdqq3jxBT5IomAeSctEUF6qBKircaxZkRbKx1AJaF3UQPJz6gJ8XAaYTsVILLn
HexvpyUMQNKu+d2a6TgoHyY2rFC0V2FRhRp7rRhQj88l+0rvev23NfMU9v9Q1kucOhvTnfxoep12
WDD0jjXkN6mDCts9LyTWGh2oH7C9LHMMXdngCUNAn0r6U/8xs0vSM3fHgSOInRfoKD8edTHRTrRA
AmpXYtgKmGnMN3Mylp5ggV79BSO8PlP0xO2U3HTYnskbWBbPKpuuVGmbqCw91X1HZCirEH3pJfQF
EaSiJiEUI+i3LLPkWvjc/fZoPEOkCTopS/kvtRTb9N8sVS5xWQDbLuj236jkePqHbscUlHTNkwKc
mRlAMd/RByPHoHaT0D2iPd9gIwPvSV5JCW+yfHIQWhiaiIMZ0GZ4+k1kDzvIcsswmwcSnvCeE7Cj
6Ba8IcL2C28sEvuVohKmQgd9AmROFHADbFIwbNBdzKm/8WXXejWSQsQ6HUEaUeCgdbVZ14ii0Xsk
0umHqFuk+gZ5cuSgapmUZ6gKFgxzcI994svVqzqZqmpVM6/353Qswg3yMo1PMlWSp5Doe7hN5a2u
abNwoBNlrEN2DD8i2TAdkSMQWLMWEIl2yzP77OU/Llat2AimaZKn4VOSRsiggz3VccrhqQ/GEk76
thjJgcdPoJBbMsOu7/naTaYGz2tt0FRPaV3i1UWgADXhxQoTUQt8EMiZLiRXxrNn9xccxAK7eKns
37HvN2YCVH8Qwsm6WH5f8CW3zXdeHA9UbAHnFXL97TXOYFhszZ5pRBXc8cr3O8Kf3UfhhfCAHmI+
nYmeb7CCi6OaD7cY7loFXjyjS3dLBgtzfuOmAQMsrH5GhzYIQV5oo/y6yPbJvFMj9IXDTUgp4Ik7
UUrOggZmHXDJqwQol9nUxJCIggVretyb8q60km3S2CA+Rutf49aHsGezyk3rte3vBiJiOZ3W8uHm
QvR34N4zEp+ZfJN+yEnKImMdrOhyAdxLwWEIGASduJrSjFTdhLuz1MzNnD3O+M5MjD2gOU4V1Fzn
3GvAX+ADcV+VKyeH6nOz2dBcl9oPGearQ4J5BxwAsgOFLOfo7rNXRqcg3H5FovQmo1oVz72/DNE2
5gGnTwVREOzd5js0FtQAi4T/fQnPA108dtFi3swSXhtGUURYPeUOuRDaPrnzOBnoURtCGMIwkJTb
j57J5zSSdXRpgodsKAdIn+CgcTaXED6D+irlGBUKRyGFUwLQRBED+hQta3zS4SOTQExV6HKLMyT0
6cJ423+ok469otIU+Qsa3I9FuiIAuFFkpXsM+/OeqsnXMkD39UgAQ5m4pb0iyuFrKPW4oMfXqlTZ
6Q9eqLPcZSedBPVh/z5RQJl/g0vAJAt9yagCh3JTxdCeskIOAUywAlQQOM/lIcpIp5iHsg8jplST
k5TuiKHQfST2hJS8XHnt24RZ/Mim1xJt7nry/Mr22Gc6gXdinf8646FepBADa1AQ13ID3JKYVVQZ
rHOVtxgcsl5GxJXHsPSxRQvud+VVVfGkyggPXgtrC0RmT8+QIOEeOzcEXiscZFMsgP2HCQ43dD1y
0f1TzXdR/cATGcrD+EpkuzFcHXKJWhLQFl1I+qeeVIWGo48cgyn34n+GX1DTWiuoMq9764rBCTR9
uQvpVTbto4dAxqQXqhkWDdO9PP73g1i2hwrsUzdOkOa3mdqN8GvCtcb59zMoVdxL9rUH2iO5xULn
9fnSP+/KfVRKPrc2+Y9wm/icjXcTU1Iox0qDWVNeGuSxbkRPmuoSubUzxIhfMAyIWLH+wwSvaEzJ
E3oWKYrGtUTMYRvEWojAGXpEStCSazt7bITFwKAc7p89z7eGwk9tHZzwc8dpX59FLL+y+9MWt6mC
U3yRRYbZEfqNZuYGyoE2QOjUxTjopWiUNR8Ndgz08QTWldWN8l6EIksp/2CVNQ9DDAfYFjevVA66
COzwcV0TcLzbDyq5mygWr9mApu+gXvby5Y3JakMsub+dABo/uloRbjacAJTjZg69SrMcTv3geXU5
M2N6K1birakURpx8cp+fFmxHimuTlSwFIG4QeVPW4VhNBvE6d9wnNWOY4cKL2Ad0JxzsJXXgnsnm
3K0AmzsvF73gid6RD5O/qM+0Qc2rTZe4zkUO+i1VCxm/QApQTxLdDRTuzPxcEadFgURjDHN4kars
6prdRJA9SdxBIWof4qfVaEhPJrQ/xl2/xQYFRAosgyXgpBp/139FEQv6gQWb26NGlbRwzDdPbRMT
fgevn40ZlsJhJOS/oG6w+jGuWguy0pqpveidfUkUGhzSYhCHkEHayDcrkYe2HkllYTrSnDIDf9p8
TNKyQz1ZiZ9TUkkbQpN7cKC4chIxiCEotZ8pskbxIVahifQvytBGsdFVHFP73QcCz273zRssKni1
suP7NYAok/x2J6LbKCinpB0KfzjsJ89vsi4uLySY/dYkq/alRjb/fuEQAU5NF9btD1cjo6JG7I7S
gdsSeN35/b6JEmFGRzqej2JOjJb6I4qjJvZoOiQFBwp87fO2tgmorchzcU05reRPbAI0Tha/1DYQ
jKBoKgf+qshMoM5FAW3DHu0mjkwqLyIR5jHSnTKHRYlaz0YChbgF/l1gnDButERJCBy1jCIm4CYH
Gs8CJnqYnoFJypt1HWDccgEsr3S3NygjKjOyzTjJ1nv1izGpkfUnqXe39cM+WvL7wWhg0iwJsnwc
2kFanyGYcVgIKS1nFZo/sfeOdAFosWjjv1BU5DlLHj0eTlHoz3czjt6tPjJXQ2PDLT7qYCTkKj/e
jq4x0B5J4ARX93tfdCGNkd7sFTyTfm3Jx+V+4MtuUy6ULJkyEa1Oe+K9TMsVIXnwbuMiw9mClHpS
xiL7tfpDb/FiZfgsCo4XcsgIhdd8wijRbJhSikAzcYgjJPP3anqNL64RdODgFZOiz7yU7xnNDKrl
YS5KUIWWQsIxpvRqYUYujzlQrtc/mHFW+zD1mRsRHdlZ9Q9O9gk2S+P3fidG+hre0tlJ27PTN1dA
LZCOomPBOu4eXMbhEudwqihaw2E8IpNgCFlEWEDLpJHObXQ5TZZnLFzb95yBRA2b63d31mX21/ex
tfrtNsSgzkFtvBdoR4SBwNYSgT3GavZyOmT9XXIfu/q7mqU3TFQNbMGEQxcDJD1FaUnr2LUGY3pl
IFkD2K/NAK2vLfXmrXsmLSxI0Q71GPQHqaJ5GYWnKVwv99BTWRii/a7tL2h1+gGlKTCZeqc57kv+
UINs5JTPM+Z8Jit8r71oeM92vJEKrRy9sqO1zZmz1fzbOKW0mPn8W10OwnLXc7GRrgYW6RoghXzC
8hxTfvmWdTLNgaohiQIVmtrWyVCaxMHnmssIf/K3EiCpzC2REzJzbUWSlS2K+QittDqrW57VUdEn
btC4kwTc+O5IDpMz8mxiD6FTqgTaqEFzHpIHvcrbmgYwD1spdWdIoHWVqh52cbKz0EesPpzlLAXK
GtnWZCgJ+WO95kVsu4aUD43WzgIOq5iS2zbqvgsbwpTo3owv7ABPpEu7+4pv5spxvRj67aXchGl+
Jv1g2fqV2Fvm+aOdiKEluwj2TZIFWcAZtCgHW+90EtLjC/gfbLMjfq98PjcRfzLESa0/iozuGeKB
/dbV1GyQyew7uJGmEegyGMZBH5x2HjnLv+7Uhm/FD32jDzBojZNaBA1QlvCFDi24yEuLnSpliJWF
wJa723wwWlQoV/w5DDM+VCgy9KH7bcrPWC/rRSvhAMbSFcmqFVfWnQshCqLZFdpx9O1DFURSn/vf
IICrYKKRivJqF+/Iguld8jh3Dz1+TbGYyz94tVUm6+ecYV6/628SGP9sMUWnb47a9U1BMrOKfx+w
7//yR1V0Wgn1fWIRPVDL0kj8YVxXZIxrBSzqYlpVeCYcMKsgCx1ftT4FEJVJi4oacznt+wgbNBmU
dGViRSvAN8UZGRhw5JXsQ7LyVFFDyI6fknSoSjSCFjNQh8nVceBuuWSuFGDHU2XBr0ETJLlEXUIJ
1Gf5bpMJa5LPcSJoEliWSDx0GH37x4aNeUMTS+eNY9MsmKQb9jS4Jxu/dSod97PIrzjYqTy6RPeY
Ul25s1HKB2U4K2+Y6DUXmaNdfrXcQjVVx9o5TZWwuefBlSY/rDm1cce1+I6rUGgVarEik9rNCopg
64LG8nL+gUjmUzU2P1B7sDw+PIBF/j28sMD3TDnrWHMapbFytKfYh36x0NzFkKaS+zlLQZARSyHA
U0BpbxWYcaSJoFMHAVOUnN8TM19a7FEgfwekvbsMvV+g4BpSyw6HonhWM8ZfiHnsv/dN8iW+NleG
Cp2eIJPvlkXAUYTdx+XrmJLw8OqZeAIxrGYpHLk5uGm+bhNWnKvKw/QNyddjU2qDLeu5SZ7djCI+
lH8H3j9doTh0dH1i/0edoJ1wgCVzs4qL4k445kHyTAONIlkgfuFxHibJ4iIwQ3CM7XeRNecP/r/1
Zs42Fg0F3S/1ODZbAU1300cqfPYjLdxML2tHduK4DoB74VMDH7GMMocwAMl+MHrTMDpG6uvA287f
Mb0AIoNAqgLxMzqiEX7loQCTpv1vXb47bxE7S6HKzWm7g9lwOQv9VwFvkLULlZon4ixsjer9s1lM
WtRKDCXBIeXcipBCObsqzPQmoMVYHJuxMEvgq7Dk5V0uXztjNp5cS4TbjCudPNnVpPq1AMck7Vy1
GfTPGGrAynzuOlKWwrXBbCc4wAuTUu2pDzJOmy8biVb0q8Q8G0NBPNa0lzKF0SXCuAparL/FoYXZ
uYrtvWsZvBkrMeRx8cN5n82YDv9TBQ8eHt19klY6iYpGPQ6rzBAcbMIFzXdOqoy3AJXByKC/vZvy
ywhpZOHiWnERf2iwKg2z1UzTnJF0yjZH0Fn6pzEbTAr4znpxLO3bWkX2BNm4e4bLCzSvvjuGYk7X
svxF9W1I80ofwb2rymzZwzV/hCTfdrdtVPUqW1jRc40bfYI4KipAlGHftMwy6dl8ozH8n9mlL63H
InSZ4/LsQK6d4BxgAI/3s1jnac09IUUcjONkob7tEYUwXBfgxsSTYjYl6YKsVpwrrD+L3tU8tfuM
BAbnymriSztg2CQg6gNA4mvbUH8DXe+ZUivK/S0ZguL/lEGeEajCHqtuXOMOi4r+Mfxc+EF5vVxc
Fdg+sKdoaU7DxyxXJwDck3z2JHbkUTQgFXyu34/Q6A7eBY9xsWSoFnpWrcfTBf1UHFdoopKxZGuN
v+k4FZ30X5WWEC4nZ24MVeoZzZcRSdxin1BGBeTIX8cGc3K6IKhx+jcYpdsJmULq291KOnljho+7
gN68GV7h/uwdxahEErAKfTEkc/WlBCoaTVnlGh/jAqo2mkvy9tjHa/aF7lm2NNn3J6CjeYF3yYWx
93BefS5DwpC2dvqBCoeCMmQvEHV394gYLZBRD/f1ZkdDzY6nlEPUYiiNolyAB/8MHJ2qfG55Hilt
ok63A1UgihJmnvhABvBAuyYSDxemheCWHC2dJYXYUWucKC3Qe3bK6cDtaOYkhqSwweR1FpqavsHO
TjhmkxNEf/GwdaAXZFmHxxwB6pY0NfnCKMDpIFGUhRF2Vb1bDveMRXG4gvfy23llKF1UtOvaXU4k
dNRaGj0Q3RSbW64swmox1FFOMJtwF7WB3VfILldfoh/vEKGN537F2XIHiOee8vTGlfiGCYEfm70x
nX7DXNWNND1c8eP7r/sxuHUpthR4bUAvomLDJspprgKLRmTICbqaRKe9Fby/n54Q8ZyOZzxLsDwm
+Lzk1juthVrUep/8AMhlfvcWWbr/5MtdQ9EsBfozfd7FzqUHWijRSiJQgS/5BF71pW8kcjj/YQCO
5UJpDqQxHOFDs2U23r4pjQYfb5f/WHWmqa8GXEh4YluUAD9uhJg0w5tkdRFliPUVyXm9Gc/bh/by
oaSTVrqBmpot5hgtY1v/8/MiJWI1/tZhhRJFSrc3BSvMG/+YO/Bmh0huXk2l6rvwEnXheHu4Vi5T
LOo3hk8zMX1lpzVABXDqGJPuNrRwIZ/LiGtTiij7mwkLHEr2Qe2+G937OEruvFwT8LNcpZ26ecnb
Fco24NI2IIdQYXnwU8ZxX1ROkq/V8t4nL57LkOP4kKWLu89wlFkaIMPtttSb5GkxAgIpajk4lJN4
JnXKE/AXQbp4Gxl2eJkGOygMq9I5zIZRy2LYg57XN5Ic6d8DTOPZJk0QXDbQaHtSMec4IDpYpbim
zZQ+pD7jALMUKx8mu3QNE4DSDvCIDMxxyZFothT+DXsdJvRInGmNyINa5D9R9JyfaO0mbqs5fUlF
H2/NF52aDWljUAkPvv13a0vEmbAEZbHGhQHLTTHVdP565fyRsfXqjNxpfsx1EjzsuAeuT1KJme1W
oSVD0J1AVjNlsnSjWWC+q5qxIuIIEB6l/bVd427ce79tN/EAlIq14T1jZ5bV4akdK/nSQZv5qG8B
rpGGbs0hhuGmqir8xNCaD8X8E/ytmyNFFAzwGJ+P1UGrhM20AW12VO8q9CmXVJPnuarmbhVIGXTS
Xgp/LxfcRX9mQI2zeqPb9+KWiVraqFb8erBXN3na4jOg0iiHdPOknNNJ/e5oM34OMXOfvzmMoY2M
YeixiSaanwGfpFn3qVB/76oY/VAYxkzsT4GHJxRSjwrC0e2//H5eBkFVC35vHxGanKnvhVIVVQ8Z
RQufejE0TR0CXeBL9E7ID4BRcXPBTweeTB8AS5CVjt5pL+irUhwWgXZvbCHTrV/inPbLhaxUiCYO
20afHl+hMAeh+m3kJFUOqsh7bW6ad0NKj5TlJ+Ca2yoL8KWUHQh6VvFxNtvLSVjEq9s+etkI8+0H
b7gKOMJBE+KEaVqwOVSYHghUw5oPuX5kvG3Lchz5Z0BB6izuj7k1DpExtG77o0PByqc+VNJ/5PFI
Xgp2YaoINLzSsVOmY8cNHyMOuBUJttFZM576jJ0hZ6Q1OXq0CfLIsgMwzFyGnLiVAcwkZS596pb3
WklNw3FplqZUokT8GiwkhK2Y5cYJEPr7qnyUwXEnfPJ/gToKhgabv5+yeKQqjQjXjTrdVEiY5U5e
x5ZOMmq6opEyWn/sKsaeS8vy2Ue60FTIhpPW1R2EcPNnblz1gE9tEjRg+BEH7hjB4JX3hBtTqiEW
5FLisC9BLDMnShCt2qdy6Aal2Xwp2Wte8xfqqBM4mw06kw+YzZEqg6XepqjX2/KF6T96MjIjkSIV
+m2PTc+F4AoRZXjmYQapmVxJEAZvjOUO/6MPmbXKCHNyMNsEM91XtLKPosrvaKAXW0BRMXxhH88K
Ik/TJlA1Xjtegr3oYLs5k07VUYoVsLxR0mhA9aS9HM7tCVAsmhVUvOB2itHMTbowDdjp+wafUZW9
eodf8FoZIPiKp7nRDIeVWotr1g7x9sgrqEfHezbcs09l7tweHEhO8YCR7q4puKEzm/TESxTWR+hB
OmJ1duTgMzqxCG4lqDbp6u6auas7BAZF/t1s3F/tJhP6dk2aqCv1rJWuFpRTilydDVTiEwOZtotK
3dz1mlVlSIQyj/lXuM2Ln9Gs+PN46wWsTGjNEvHifLcEdNhPK2+mPHkDvAayaTlyPanGxfpB0J0x
74iJ233c5fOe1W03py/MO9UhRXDEOUZdLsT2f0H66RM+256E2wJTruANIXCLYy4QfcgQsgEf6rCk
O7NDsCJd5Gnho987rHkMPiUWc6oNVfFFsk4+kDfNRp7Tu+xqUQS1eAj2j10Xbdlro/ARUVYagbiu
z72Q1fo01V562nmwyHQJQ4Bg7RMnXNTse3sgDKuXjWgayCX3GJfFdehr8T1ICQoxL5TgbV+VFVCP
+VjXkbdaXrDwv5leeYIHy/qq1a4MaCnMgCvyWJEkFfBXR92gOCVlV0EPy3M/CmS/1+hEFPQYOrVy
XSvBonc+z+dION+w0m/4NjQYSzD5nuUVkKMvm34+DfjvP1jOS5ZOx+J5Wf3lB5OkXvRgMUXqateA
GHzAc81CzCEejI8nvZifpn8D6NjGNDyDLY/mN8YXD8pdAqn+4ChqRTc0/IzkJm93JaF1ii5qNGCf
ileTnXQMcf4uqIcVeN5oPn/nmDH+BuGqpxmnHoAOAf3tnLn55vBZe/nVRJ8dpz57ShrayhupKxyp
ntQYBU25/RIInDJ7NK1+xuSpzpZgzw2ccGYm6/rzDvY92crPn8xwJFefcp06QB/8i7eAEW8rWCCG
1Ga3DNwYJUjDQl9HYeEv4aVMAy5hQ4TAVYCefoBdOkyycUmnw3eokVeRXvvVQlOCIQNsJx0mVPgE
osP4igNHlU03utsYrQ3DPjodXXz/gmR8Jegemlv2XS8QXplMZowJZewGSIWxXZGOI3ulQt2aGKCJ
JRY7GmwcQoKIkTpB4UXS5iNWljuu+1gxQHg2UGgeKPPzAAMtHHX1bQoG7TQ53VhHF4Hjer9nxWiZ
AHScEOZ25V1XG5cRLJT4YMDZJThRsNEiOLGVc8Qt+Rzn9PvJyxpIm8KTE+OvTa1EAhPWNACjynOo
/2vzta0BRAWW7Uxo00pe3MM9SFxcWnsWp/8Xpo40ycZCld/3TRtN1wHZEniBzUoVrP3qudQx8OIv
/CeEJexJbGOHmN4C0myGOtjxNKRf4IVMolV3rb2FEcrEExIKOGRXnfo4KRg6aH9lnNvWeG+/jccp
Ds3aYC6RuS3OMBaYsJG0TEMvcCGn++FzL2Rj2i2l7WnUYM/ErZPP7Po+5G0abK+raVIvyckBpZIA
MjNHZbfQauhlrukYhbMvVFH+s+uyV92xf/19drJjrD6y6oJXSim9s2tthpjBVood9A/CuK4N36Iq
YdTAKFKxCv3JejswPf9oOlGKGYGA+E3WY7ebzt/B0eMwL3/ibyVP9IgW2bX47AIQ/UsD6qm4SSTL
UXrtB+E8egPLQhcWIlpvQ8lwyk+imxxOhU9a61QeQ0EclGxhL/7G68D/jXDySRqeu3QaO/ErOg2x
kEgemhkjJTesx6etDxAC4U1CsbUONXz4ehzjxliH1zKPPjRqAIWoxkznAnYWmyxiceAawBD/0WLi
wqNF5/hmjMtZZ0JPr3jJmPuo7l/PyFsztlyLmikMNkBNzZrHmG8UqbDVO8jLgFT/hN9mpgSyg5CE
fvxBonthTTc5SE6w5S5gPnAsmY8refS6aEV6WFdjwfLSSmu9D2YJY//mAUmTpgI6N2sTSljpauu6
MOz4SN36Bandsb/pnp0aaO6P38R3vUUCpEm9juGznd9gSmuPXNs6Tk9xkhA/imbvBbvoes8+wMKF
sFTn8l0gByzJW+x+Q+HTWYGJCE76PPHFoc+0UVPzVdrjPnBctNsp8h5vIMyCEl9R2VhH1Ltwtzjl
kFGLJ55w7PLZAIGDP+/qsB7aO90cEMhZQRJrHQB0+mQxQNGtF5e091kfKAeMcxND7/j/Wf6J3UN6
vPqTuZkrVOK7fXy8Qu2EZIfdvps6h4DEQ28K5pnFUrX5K0411rahFbKS2ytF9+1dCpqLCYGrHvZK
YwiOntxtwp03h1GvLq00mHP6Twv+rhBOtNx+pfJxM8qh8JfWqDiEd2kcjS9EacniWl13JKC1+Tym
fWeoldpW0+h5aHnlV1s8lLgVBpSrXf9JPC49HYptC8xyV7S1gFiTIKbat1zceu18tGoupm9evG8e
kNLCJ3PPvqPt1NHTI6kc6sAJ30wFU42V/NQYO/7nMb6IwUnEv/Z6yrW+kkfHc8Z1Khv9Z1P95RAj
rHA7NACsl9OS5mfZPrM58F2Qp7x3xy+yoY3XLIE3b9LgYStbl6Ya30n3o8wXumos6VpMesTDmXF0
DrREb7rdhN1OOOogNTixPHXoEwhwswPiEZOyto0jonIKiHSUYU8sdMqeUzJ2ypCq8vummieE0H4s
h0Ue6bRjuT9I861jBPU4GV7NpjCdssQxXGuw0cPX8mIMem8jtcKDpPAtLfqGtfcJRntW69j4X+t0
zjcX8yE9RaKBYG7MUjFTHaE/shlACjCV8y48frbU1TO4BLWcIBL3zdReNX4Lt1HQpZj737uxgcBd
XIDdUPgTH6NBsLawfVKb1KtkxAxnWyW384cWsXWFXk4cCgguriPdFyNMmp9/p0sIlUF28jM9dUDR
e8r2tMavgo+/7XWNZVn8f45DPoDj6zhWVsGlEd5hHzcKw8PA85lbr5YIDMrQeygGpv+0qBVyTX5e
V0yYtUOXac3WQDb1Frmwbn55ZobqULABV44rq2Wxr6inte9QwUmoPg8hlkxWH37lvlk+PRboGF5s
bKPXAvp+7/nR1rxKNmjQvLmOCIsck6Mn5wgMuSeJbttUfxMkM4tNzifFnD9Waadg37sxExQLpPhO
ovDt5ZvTOIJbAFS2ddzSCN1rPeP6L79NSIwQ+g+QU0WOdI+svNVk9g/Ds1qSLgWidWGkUmR0EuCe
gBJ/5fWRuaK4g+ZL7pQhI4+V5MgjnCo1Aa187hHkCy9aWPzlUB8VUM5UYSY5sYtg29eYnGOk5rR5
Q5zyhVRB0VZo6EJRCTuJxohuFtG3dHHXTVsi8I/CNh2UZyR7AsfsvtwTO0GaAOVaE0mIPXPuOv92
BizHSDI09TS2Yzrpv7+hkm4RYF/AAZkC5ML56UEcgKi7E0rlU0Q5o0LVfAFJjqSrht5z2x0R/ux8
9rEGqaoATW0q2xzvVqNUTy2TI+Ak0RuGcmDLlX8DxgDEB0hxjmSRLKGRiU/RO3YEeRUqXJXd1tu+
dHU5lWBONaRZsvWu7y/hj38Qi0xdYk5RKjwIQn9/FsLTpWHd8+Q8zxxb8QXGGA7jTqoZjbzs472X
z64jzkVqeDEqn/AvWkwNMNQsNSG0d9aedDNZgRugjJ+5KFw7Sj39E7SHm9TgnGvZAYBf6ug7cfwL
HzPH5W4wywPVP8T2IrFTZ34E0E/fr3hvLu1/vmRkBwjiUgMdkFCwaJsLljMT3kErNV9ULgs+Jw/d
Ut9KYkDytL4+eKw4WMNkuDkhT+BbUYWmw5YidvwudvHB3q6T+0P9IkuKuuET4Oakb0QHTimjEpMh
zZgfPADNalxezUD03DqbBoVVLA2nUc+d4QylO/mRaNZe+RWIEsunXyP6S/v6t/9EyYkTDVHaolBP
WG8GLvwevwMVoCm6WBxxqgrqlaLqHD6J2kO+XJkBrr7SE4gNyZ1+Asdpw3QLlTiQ91msYsqQF9t0
c/o61sdcJeiX9+mcIx6GgiZqaowmxH7q3r6LqbeFB/32Ezze0N8gT86aHB3m/91nUskph3TX/I9B
FV3ei1ThkyBw2bDBDvO15NkoEeSZKvg9C+/wxJUllf0cAc58kOXbR2ccbvT2GCw6sYmXD+uaKy5q
zdK2y4soiW7l1KPREe7Zyn+N/L1afGKTMvrMx65+Q7MQc4i4+9W6rIbSogzokAWpL6yRzrJ8fEw8
KaG7hWP3sP72MVtDTU6APKXtu0BMlht4zrXSeUkmbiGumg053gtQnp6+KZhsu0LDtpg07MuHP3MC
y5mmhUN9riQNVpTqUdOM8Z1b3POT+dgBv/2YInM3sLT16gvtaIEp9pITaxwDuKyC939u+HBO9KfV
fbGeG1gFDjlfDoTm2IzGIn7EkPUaH0ofDnhBEvjavwzDIJWF1ddJ1RZBg43GuK/DS7lCunuEOhOT
wBqPN1/KO7dBcKApMqz7ypT5ynfYVOeacde0OIp+fRE1NFZ1lMM1LkGli4QxLxtRkWDx/XhhNeQE
nGCCjZoqm7Z9X52oC+vgdizOlX/kflDkt3csxLBKvb8N0EwQtyNI+jw0NH0gdjrDvfLUP7Fz9Pyk
nKE8TVuQIR1vEhwIi4+mt798Hkuxosk4ej/SB4z+2tKFin85i9Md2BESA0k9OJGI0OeQvCNPzPGL
KKDpQrSjPHhgt8BKjo79nGY7Nv1COCCpKtJNz88IZVZ4EhBa86bJRS0mw59Kfqfb+JfJF8wr8pML
8RPK3B79WwS2YQwKSBm+yVK0vb2cGeJP9PiaP6uEM6pJNBs7P9Pa9KXwGqnkWdMpE1P3jGiX9zny
qkJRgUTrT72F7ni1d0LNaiJ31qcRd4z97ZxAN8vf1IMETfLHvwvgMVj0Ozcp3ug4imzKpy6YQoOt
Nsket0/SLyTDuTnht7/YksCiAF6xF+0pY0cO1bABWlCYyibHPxl7qXeSjqqd3UcycJ+boKqPo5jr
iudupvH9MqNNCXq2PDDnxEWpvChdHssY+zTDUVaADUSLeJJhjUBzZkbI7YRUoRKZuHneFF+bBl2W
Kf5W8jlFMxpMj4hYwWl3wEr3D+mW5vgFIjlDJkgJp+aJkcRUFnN7YegHrW/AkE/Ppv4s2CszVIL1
CqLeSAcNMJKaff2+WVu/QRuK6DQlrTlvgPj13ewKX3A9FxdTyf3qjqhGGC7IB1M4KY24Yb3lm0fb
V+Q7208b7Mt+esgq2COPRFKYOe5nV5Rcs26AYYqN+fnOnwwSZICrb8KiO+CzPux/MIBjp0jJf3F+
mof4QbSj2aQmB/de0VuOOCgit7NFDQN/Dq5BVpGAKuJoXHMj0k10TKRIeRIu7VpXs2iogGSj9BKp
JVE25FC5m8FsQi0IoQLSONh05yVKGcMs8SaOwwq58Z4L3XNXGLtPHjKyKI7OHlgqAMCJL4Ayackw
w2jMfXHmc7O7KiSpS3sGBbp9+GuYSqXV2vcuhaoEt0keq0PpUpILhFPMDenFBlCKhf/m0l+fDdun
oOaccU+T1p2KlOZWIdNRmD/xAFQPRPSQvo4CSzh6KgSuVjYeMZmMSBVMezmRQNn2lo6eWODOSm7M
mtAyn5KkKGpzMRJ1jmx3GJaT9F+ncKivwoE+o3MjZwzYozodAtHnP5RGaL3doXFE3t/2QFwI1PFo
rRwkuQZ29G64l0ZX5PtWgYddJcaPSZ2eg2aEFdMUUY6JNGqb0IwyiB6BT7dGA7OD0k6haD5iL9OU
hZ2fa+bZyHneD52g7NTWukgOC4rkkOT3mr4R00bfyX3CF5yPbmQ4NEhr1cvJepKzt6YA2oKGzjD2
hSc7uYPZsv6GYuqyMmr+iI+oGHQwcBoEKlE3LNZ+B/KkjATS6rdkaymZK0f5UuKUw4spdpmxsVgN
HJjppivHk7V//LF6fOusoeo5B2Qi4dOc82LpSHySI4Y4/+NYPSH8SB2mhlb9nxfhIbodPYpNz0Zn
c7HSD1YVVMSAwIJrhUch4K/gHhe98VTXCeeyqFN0OSV3BslDSbPzpQzX1EvhL1/WLewlz1FXBg34
r9/kvTEOaTJHUOV/1MbmRPnEOK6kAGd7hgHpjuQ0HLSmKjqswGhkeUMXK6XxEgSEWTGsStzj4O+I
BjvsJBeTdNDoj6jN8QN4FaMYHzfq5fciqIz3K94G+ZvOiR1qVd857gfmohSjH+mXtP5cZ1gwrH9i
Yrx9NV68rZvMCKpUVrLLZIsz68oGoMGEZY+X1RHcOyXAsfMbf2d9ny0+tWlo17CwDKBP1dyCJmlR
419Is3do5RJk8A2BgzReCsML/obpe38XKC4Bf0zNzsT5em5uZgi+5TH13fpOIOfcwNKOx9lkydNO
g7wlyMvDI8kr1D61pKY9QyYa+QqYQvLCjZK/160D5Zs5oaWSC27xAzIAcft8RylJc9w0NTUrsvQY
VQxKWDHJWmF865T4An3EHtSg/KayIMsAPineQyLS2CDR6z8uapKE8cdk6exaHXRCizqY+r1Fixtb
zMCvhgBDvGGIKVkHU1KcTTVrqErVOgtJgv2Ry8sKOnNhDApzQ3XYxznB+WoQCXnYYqdLyx5eCWVF
hSdnpUxbt8cJw+gFjY4o/+EaezrgoOrJgNYqll8y9BofP6taQBvXWwrMO3rruAz0/j5YZoxom9Mc
2/dnCNX7AwSYD6k0kbOxrHgNI9lccSciHOA3Fj0BHnlAii4x19TL+OByfPXcNvvcxt4kfQjQzabN
w1fWyZ4SNV3SjXm+4eq9Hayp+zH0B9fMfdnL4H5I1GS8NMrDwppdRtixn4+UaF4CmlrK61iW4WKN
FBZjABwlIx2oSQalhepTmKriteqkxIP8p4fK+obY6RnQCgm0NlOSw2wtb5L4FCgma2l51Wvo/uwg
0GyaEiukjYR9zJJ/5IBaAJl0h5Nlf32F8fwpWOxA4Kx3/7vgVamn1/N2ubLn6ZeB+vtRXiGocqSK
z9PHK4P60fh9UIGsV2b8eZ7Wu1aU3h8mfuOYN3BnZy2ZwKnialhcVqMKOJq2hvCZ6r6ctd2BHRh3
ynrX9LG1P2B8ErSMXaB11TevP8JFVJ8tsSEgnbl8tCsBAn0RcIj4cCHkU2joL5k+DvU1+GdnD9fV
tJkGFmSyS9YhHdvMVY5xc/UKYOD8VvoELET5Irbad8B83pbRajMXmPMtSpJsTicdOQnu15iwaqt4
MLZ3/mfCd/+oeGrJqCDHxQ3rDInuF2KKGiCUsn7SOSWoErQx6Mfhk+Pz2d/de/qx76oWfy3SJpz9
mR6oV+F9cUh3c57hbL5JymqK8cvdOL5o4N3J9JJJRTuPr2R88zrRcGqcAmXHLFgWEsPSYDjPb9K2
FYzjA5KT5LVx3Y5Rvn8luFGUww9/wxiRaW2wCYDsryY7Aoc8us6fWvb7HTOEF3jnPLRgAjWsNnIn
DsUYdPxjF7QS6G7SU2nUI9zmTYUE3J14Mb3fVmpSYlRXhUV6/iC/AAp7T7PHFLfm9NCB5VimQsZq
ZLp9WZUHooseMkUnWn1IrBneYshy3wywwib2CT6KlpktcMgXseJLwkWDDP0EwMDUudkN59yLV8d+
LGozaIGYYNRDZMVrZ0iL6/H0zPO/dCLTfa0HsZBSUcFOwImJ20TRvGuYr19uiH5rJ+aCVBFQA1L6
jzM3U6CXzLUg9v5dudOjABQW08GSHayh9vMQge3/Qi0KgroXUkJMSxSSW60AQ1Ml3VH3PClmkYCp
Zy5Nto9/JkexZ6DZuRKOroVpxZ/zgvIYQL2awxekt3tPel93kiU/MxMtD+cYm0f8yzXQGomjvxBi
F2Ddv7aKR8Yc27ZQYHrq8r2fcAZUox32ybxcqi2gmvLFf/venRXFqE93wok1xI25AyRETQssANrA
sYCjLg4N5ZwZ0JjqEsmxjMmIdRMnwwZhp7Mzz0vsNwXDBgeZlx6CB8spDhiCYLtkiDKkQlk8KgXq
uFZL2CJWbQwnRgbTftTVHpDpFaAW2MQgrrz0u1l/SY5szkJI53enm1JF0FkkLTbKekGEHXwCuOe6
wCWy21Px9jQ/ZGzHTw4pBVU8SYpqqGEFCeeHJQfTXQyoR6s5nIbjXJFX41Coe1N1/vHi2jjNh4RU
qa41WVlYY53zbjaQRpIBwF4C7MBwcizK3qXo4a6iQ+yrCXA2lAdVEq72Uf7JVRGjWzm/Aim6Wt7M
CozTQsMoq8N+4xpQuGNuQWt4CgotzF0Ckm7dIuxu+6wP6nmOtQD+jsXlGmoMj5+dVTAkemHeh8Qf
K8s4TgEJzgLf942/GiTr0hfh+pLkgXnx/C3zLtfWNiKptEiE38UOQDahAp2h/g6N5wBqf7E8bV85
CdpPutGQBObfC07H/38n1mTj3m7ZWnN1ixBYpZgMDf8Lu+lKoZydus2skPEwuMMuk3KL0lWfoflt
/YUqDZhrQSwMHM+JOg1ROYlXl/2aetsw3PLbNYjt5FVqxLm6vw2bmT3O/vlZOPO7+xIXYa8eyS9L
/0FBPM8+qZwfh/oLWC9AAA5yHS6DgXcIXGl+jRnwFTsNIM9QwWQXumZmwSiFjDS4ioK8qF89yAQ9
eHwlJMgtL5JCk2zExrKmf7uxhxCGghXGSyq3iD8ecYhF5rkxmjMrvRWxMXgdjS9IpKwX/9AATiUH
GgDXfExW1+rfwFCNfWOLW1H6+hbdW96oy1Y0KSdWO0KBe3p2DdQttJ16YulcLrnJcQWqrjj7f26B
mt349vpD79Ffqbq7I1yDHLjn5S1Ol70N+iARwuhMBjl3zHSdVw0S5QC/nljVa0DvsB48pCR2SdRY
nfspw6W1x6oNPRBEoHWRAkBs4YSbeOWwV5u/FySptWotSxsGBn5tL/oVjfbvA+coiyCHGXF46kmy
ZN39u1WWPuuy3fqwuRvIX0Wd1YuHUCMOSYO6iWNhbQ3VFDJmRqRkwamXEqv3AZgLBTdWDLFNJN+l
VdsBAreVKv6N8lg1rYfqpWbbRn0xPubTXBKafIXMfp82Wqxpf6SaczDRIhr4JzQ2BAUSAbUnFbbf
Va27/hRvwXCUz+mAYOCdn/yJmGcnUyAKGW9gNhlGJ9v5clXhNNfTpjkUw10g1BBdMY7oHgtrXpzH
YWQ1HfA/UK5cpoQd92K3wJtHBsVS2lWHq2BPe80tym/hAmsphDcp+e2AaecoNu1lnHb/IVA1+rb6
TDCbWbH8nmaOhosSycvKelrnc+HCqKJl1uXQtuSCxq0BS7xN2rrLyUEwXdJeTvqd+05iPdd2fCWU
AP1EFxF8XAMmbpTjQUYJnZDjmQtvFk5FQ51MdiPWzQ8bZk0RB+yBwjXAifC07fzEIUf7ekF3aFSp
8p4aGngVzh3rq61AK00RdkqvgDdi7QX8oFPmSGAleHwZlm9mJKuM8lOWv+F8y8A3CTZW+8c2yI8W
Yy11T8g4PM2E8vbbHdWlb/EBkIi3+PyDUId9/wecNkCGyidaLHYFKQrMxTlXFpW384a5IHeEF214
nNPU2Ix7y7fsoD9kxKFRGlAYp1n36Jri1Vb+LTCiy9faQnfJZ94DW/BIq7pIGa1UUwb/9O5W1kv3
8rWcQnp5wFpzi8VkrkMepJLevyyU1Y4tc6UUSm+kKRKolL8J7WorC2ga49KpEO6BG5ynkf3kMOC1
4eNu3RMTXpH/VBEl6knxlEHuEhd3toBUcG/c8NUQHzL2InpHCXF5TCQLhm6ZFfj1TJDQ1gsWoVmC
r/w+BM72iiHMYZxrc4ZAS7hUdIUNqcOqI1daRsZf2sT56trvloemW9E3fR0aJkSyeeQDvUbMWsnA
YPKILxkKkhpbwnNOHbKYwcpvhjCd71fMa3bTIhGNOCX6ivefwhiD4TC+N0c7ZPFox5YvGZjxxMV2
O89r4VyEsaFD0A5qA2Ax1y/qic0PiRpmYgfIqoggoJZ9CqyZCHIPYSEvOW0Jas6C5xZOlFaHiFFi
Wd1uORtyCQv64nZTFZen6Sgn+wkU5UDlOBf2D/uT4VldgHufyEEE61L12fi2ArSFgheXiADf8I6R
cSqStmFuT3VzpJH7VL7Q6kGScB/esUAi363GP1offHdCihkBcSHFr3bgd/WjXbPrmOEY84Hd7dVk
CUQGV3xIcVSUcroSnbuJ6QR1yVpDV/1813JfdIRrKgnop4kUz1HTwWaj+zbGY+8+RhLwVMDJByMe
6Fizci4EKW2FzLjRewNFDoL6vzGJJqpN2j7dQAf6++jUAa45SbYZ6SzCV+X/bKHKpw7cTnqiQr5+
qFZHNB837l7hG7WVKbHItZd+ZnSwo5BWVBi9BfeZXapF8pyJLlXewtijvl6t0YgDsJMTWxHRdAVb
ktMrTDmPUTLyTBWSp4b4EQz8cBvTHNGGWkjrwfQWmwFnJUufr26TfMKDvI6TnX8paJ1Rif4WzIeR
4zTLxD+vxF3khFdMVxOM7/ZZeVTBRGa0OTFxPcfi6W/qxuy+6zYhhPg3+wuqK1voC80dLU0+51fp
0s1CCfxfHE7feozq3I3BQlmIQyrV8bPwrUAtOIFjTq6ErAtLWZKRC1tgt9QZdF/+j7Ce3YmzqEbz
Lqoo+WTceKJRqe0EHwtwpYpTEMbwj6LPdyMSFBY2zOIRAhYVXLiCXjQW2pmhYGV0Vfuh8UqmtEJw
HfsspqPTnfErXMF0dHoDC3X6TEfe3v34VuLWJcXsYsA8r5htN0F1Us767XGsMOniZo/yiPqY2wtZ
ge1KrjIEJDVaCIUM7djnduulKhv4spjKM00Dy1fbjUcoZkHyFRP8cV+xr3LGgYe7SQoF3iemR3AY
KsdiieUsVHIqRqPP78CG1CFYdLJnwLeMtzvtqunVcG2l9dHwbvEPIWtuPsY7AU1INfdEfSV0Gzeq
MPlkYAEUpd+OQNgZsaDEEnKyxwxy5kLZFAnaQASFus13Aud5H27rrz3qSGjDVvYc82P4M8JYxe3+
G5efJQVszYsG+MedoVTCKaaMNcuJsqTXMRz8wasjYnXW1fZQFePLyxsHKMBBX17cJudHUk+eHMtg
yLOICEMyHNSu7SwJxeg2ZeJMyvuWiJwO5adGcVPAnapxMZr+eLUMAUb2VkuFTjrBxH4b168ADgFo
SRQJRfZEF9SHdYujYXvdN2quavjITNvTSMNL13Lpjv+LNxili7NrEaEjABBKKvIMPTlwbiYqjKGr
dYj+i5mneSrLbAf5ExZOgOHQ6CDBD8wfQ8oUzFSEVg3y7lKCjsDH+aJlhaEiRtOFNdJh2bJGqchk
6qZxdYhVHKbX4DfwxYyuyjjhIG30e/YC6FbQuKPhY22geSSKYCn+yajyyrXEPhCMnKDIjHD1lum2
NW4khZi8JsdJEpkWkNpUJz68CRkxdl1b/zjsLxQzRKdUD6JdqDTPKr1meHyno+9+6vTb+recLE/w
U+gR3EhsuEDY6A/AektLwW5d2HO5kA5i3V+sjHMk87jOO5eoOLG16oSYv1BMnaZij6LOyt2kjR6C
s8XA+IAGIfoxpfgWHSQBZ9b6NsY36NpNL/zkMB9S+WiK1vOIGQpRXHswzX49SML5Tc8f7lEn5L1w
Kfm2AWGzxKt39lUG2Sysxme4vfLUnmfFFOJgKjywonUZXJmNByUyc6N5Q0LngR9kRiYuhYjBJ23u
a+nxJct02HfQOmLsyA9zHiZJCjGrHGP5r4ZV6tJzRlxHvZn0ZSb2NpsZ5ECPfULZOnbXI9kkEiBL
CA23pYVvSPVYgtmGmjpfmktQTg/V8P89+2fs6cusw6pw/f/MUSEPdg9YYBbehfSsbFAvKCHGdlHk
zOvCuXh5G/5clv67ClW+2CxES+V9/zCY9/Y1n4VdeJhaDrbH8fVZug77xWeFHvsLNTX787lEXpsF
cxOB6tX/FYPmNGH/25tG2vkuZiWHW3Cu2VhKUs8NSc9oe9bHLuApFGCvMjjY4vF/Z48X6u4cHxnn
1b+/9zNvOXL/5F+p2MeGB4LGMVPBvL3j0lX+SuZk1fVeUzyjTpVnEVGI8RX8bsO9apLWvi9RmgHo
aojJ0PAv8rLMDBEUyaw4JLfvg7AnOBiXwQoFEl5cgAz1FyZQLVM4gFiA0FEbEY80CPMWmGVt19wi
rYrLTvwLj019VWmm4PxcVL48EJl2/Jb+8mga2aHl6rdwUK+tMWVaSgdCCh2Dlcc4cTxjULAojEkn
JIWOJFSOgQx3B+O0ouVujRPAuQEj37RstQZuVWjwKNSKH38ZYUQkw4ulqHFYtiZr6ALlTzLusxKy
SUCD2WYtGqKvHkGLnxdQJ8x75S7Bww6lFEbkwNu30Rz2s7480CIls66gLQtsmfIxzlnbmeCKuHpu
LqR8Z2RhfM4YKr/PodtfHX99b5dEdbOENCtE+T1eTJn7RZ7snXC6h0pO56jbGEHaZG6bZFSvy+I9
+eHlGB4aCl0VPVKy7BS6PgjJ08Oa/AgKeAljUkgebnQNPTkkAboerJlAC1Q2bwBpyVe9ZS02wbH4
Dd4DoiIXTzXAnHreZ+4gUlm2p3p4RrLxFdg6j+p8SXI0canPCg9UBLmINyLPs5n3NNmOJdKA80PT
greqKjL4zeasWxw6jJ2UwYneNUZvdtN+Ms7H8+mS+8qe2IYKImrsVEmYDtkctkNICfXJUrJomc5x
tFcCm/r5IDr4q9yHLB+kZm/jLGn7wKe3ltFoTgxkUlyrG+eAUsCiReDQthGNGcbh+Q7ycfGfqJq7
zn2MZr4A45riivfluZU6Nb5JwBicJxrIcUsMJbThLUUXEfQkc25QhGwh4MDyZXUojgK470bYIdI2
KFvuwFqT1Qe7mgb1j0WZyYREad/FbL+8p9FDfN87Ga044tfXuE6Cmc8/VtaMZp7TD6QDk62UITf4
S7jxxZTYc/McWd+FDUj5BFqJtabyqqhWIJwMaGwkZ6/KWi0k8E445L0k7+cvIjoiRcNThWcs3KYj
q+R/Fdfq1xNxNxK+mwKvUwsavPxHWsjb+cp8Xw7WMjETwhkYQ6vgvGjUubxP8QlqDu6rdEfCjWJw
LFHjheCslCPwUklJSf5iwuiDcNrvb+32fG4hfSlJQjK53dtjZ2fp1bYpjf3Yfcrjc6H20MOdAhY7
lazrohqwE7NoEL45COPW4J9eJHLytuVBht8yMEEuss/e0BsOnfNYoygLmkS/HRLyy+OhJEv4xsrx
hVHC4nbMg4GAGV2uayUlPQr2YvCc50/n2DCO+1OHo+T3tWx8N/y8w5vwTpqcR6aSM8Cm0QGobpMu
CYENXutIrEkMrJ+dFE2FGBRokZpVcoT1qAYKQWQEKzQatdg1Jv+BdDvaQqzQ0M0R9bwbXOahAHxE
t3FFlX8hZA64bpru8OjgKj8xlk5gpHh2HlM9m4JeF/KV3iepWuMf7xyzsO1CyvO3yerIcd/RB8Sq
MHIO2Y6UVH425VnIYvPvqg5h2N8dLk1rLz0ekZkZWGT85VpIqFzifdnPPzLnkW3e4JEKVxE77g8Z
TNKMKYkDtjn2n+WYqbRAdiI3mdanSEKLcS+piTKtXA8ztDpshT39I7KgxUFRoywDi8+BUM9lgH+y
/nGI1jrnqM/o4VTV/DNCqi3HIRhkvWy4hSaNLaqcXGTJxFldHEkYSDCnnWKU5mhyU9gaouB49u7/
xh8T9J2WyueXfFR1hvyS36BL7popOERPdkq7zommKSc1qyLNllgYIqbn/d3TeluLeMYO+Q0QTn9Y
q9w9Tsukr5dzevwPlXJwsNkh+JFMjF/fA7OpJdsxh4KScBdrXCmIBUIjUMWGyT9KDjejhzD/e/OE
tbyAyVGYdYYjEmkEPu9TQsAGftLFwlkva5SerdShHD7rPNODK0oqoM4KyTmndr6X4zQE9bR+NRQ4
aqOm6XwhoByGnqsmrSmM5V9OefzmPbzYns1LXObs672gR+IGqI/hb6o6ak95tVJeYmCsKgzz26Wn
W4YEZ9VBpZDTJ5xFLQJBnqFgRFfLZdX6hAnnvGfMmcohFH3SzhYY/CJVA2+m0yW/FDCZIXwc1hfq
4kfLNC3euW3Z48eaTKkoMjrFbsakSc+sgXkHo6Eimyy7mH1/15+ZpQiHR7PMSfaMiGZoyTcPYulI
e0XXroz265z8MVv7hAvGL5M1m32VZ12nXheJMq4KhkJsNHm5ZxD87exYqK9v6fe+ZOQTyhynGBar
6Ka4RQsLH33qMguskzc8YK70w+lBIigd6wez3lzTiLOucUBAaLUh2N2/E28gC01a5JARmLtiUf2V
obdWyeHWjAbftrF/m9hLlifHl3xU1sKHXu9WGcaZGIJQWkpR21SJJdKdGT6CzRe5q1galJ9gvUc3
owEmnNxyQcrO8yi2xHW66kXS/s/CUiDc/oJDTX/Eb2z5LNntkLfcjoWLArC/dO63BpnCDKQxlIaq
Kgr4wAQ4QCURoZm5TIDHNeH0Jku0jc7hHJAjv1T58uLyB6jsi6byc1MNaWoWekWHMngr1lrKIQti
tJvFNg4pK4roAdreWiRt6ENSiuJ5ISJ0XU9/Iga/Dn9O+/tk0p6v3lUlckwpll5nS8qZI8hGgKnb
of4sLTK7n6etYBO5lw1S4lo50TdLpGBziavD0pW03msJxS6iP0+NKEt0P+Xbd7NfvIk/4Q0EKDsC
IPGWE+QdX3tSDg5bGYxIH4OWlzFlD+5cdftOYZOPC437LlEyn9gHjaXOq7jXnJEFAY/7QWf+cPZL
s3XUdR1vZZGMFTh+tJWrUJFqR7s7UZMKXIFuSZ0AennDqAAcZE+sNbb9wMZAqJoPjqDa+UXPsjzA
amDAJ00tqdnchbGJCf0cK/a87VLgF/ZrHThho9E+01T6zekxvdwVjZ8TkricXP2owYe/BsM9A7+B
waBSmH2E/EfnmGUwXzKNan+sZNacQL+mO2GYC12PNcYJLkusiK/vTsUmWjIRIuiQoQc1/oitgi3o
a1xe0oj+4nu4DluB3tJHtDK2vrI7wlDLoGq+t/l6y9PImQ0p+6/R7UovkHH0t4sDhmvZ6tvTQdeZ
HN6bDXTshpMg8xldUV2qg0ib2AJn4l1eKlhFtCcqGeRfLv37cTg4ihIMHGMvE/zDBU44zvFQzMxK
bD68HZozAXWaYMzOZFA2RV48j7/cTaQ44L3zJPgWYAJDzLnfJbaVN+jWutFpNfVljrB+20LnXnOF
sVzuDm7A5Tp6DW5ESUac0n7VquBNOYaUJGuJN4D50ajhJauazS6TO4d7R1q37Vfk5SNemQ7WK/lp
LJK0WThO5bnwmUZInX57V+SCrnN0cp0ul0MJ2m2vTfR5RV953Khuh/AOQa+HHAOy7KqlcZS8FLIl
rrPWF/ipm0efADIW3bLbOkLwOf502BafgL/+WOvDhlEhqhjSFdeLGT2rY6N5eLFwwnBB1P35RWgu
Dylk/YbWE2S7uZM8sTPEDSI0vuXbr5tiZOkVip5E+8HK9lZav5V543pkjpnoOnNEdzHvDd21WfDs
CAUR51yEX81jfjo2iR7C0lQIb4ZUN2P+xOwD0IZ/3Mpog8jAc1bPBHYti/KHLbIYWJ3WFWu8fNBP
jhNeHE6CWgIzh9We2znhKJEz5U8kD+veBARuNMArIrT5kGq8xXt6meFTURklaiYdOVB1R3bEDHCh
qofA7RZJyItmSgdEkp2PZn5dDvI8lhLIGj3R+lZeNQZi16MFVWEf7Ps9fDPEcXekIJv39JO6UdfT
9FQTLQdinFaJ6pbq5GCUPQYlVMrZZTx782EkSpN0egTVya+c3D9l7o838+d6Il2ErA3PODYl+Hmy
qlsbhVtlXGZCKDZJT5mxQSxJipfZ28o8qHJMQXIBWdt3OvYGj2mUa+IPBf/SP6y52nZMC31XSpZQ
T0ZZuzrUUtI6WB7YlEjuSFC/8W/aEsh/SKfgMrQKyjPYzypvAmHwEldgf6lJhuQqBG21aVNoU1BZ
KWdQqufLZm5RpUb82z36LaDQ2tXkjOZA3xAgufvy5m8mvB2Wu84HdPP91YGLULyIZdf9dn4TtROI
ZXnpoBLCKKjmj+9X9AdYXQi4XSB1tl5A79jt9xTTxY3MvRjikPsSkBycjHhPyuHMbPNumcXqpzPZ
rLXSex7EtD/YRPEKhxAD7/OgK+T1/1why/BI1oaxvLCuVR1CwRSmlSCD7VCUb5rN75TFXk/bosc4
ddX/OevMtYR3hGZ363W8/uWfD9QlaNXRimKkOMQT+zLUEOXm11IbdKtTYAiKiUIHTKC0d4IM7+uj
090x0U9mIU3+8UZ9NEtXctveZHrvT+8yGNJmJMIs6IufDjQ5Q4WKFb8Tkdt3TSecJK4LtZxuOR6x
jIggjcmTL9Z71a197sa7gzOh+Ilo9I7491C7KuUmvcpnFboYrFMX9zFiGWQ0VUmmEZTGeF09kqQD
vUp6QtB/RvIIZ0o3K4w+8R8TPjPS7gzJeaj2hIc6TBgEYQqgZHF59jVfvWv/rvRxPYLrhxAZgn7P
++pWL1ifQcRChWRETOTyCeYHudlZMWJ98e0f7i+gs2lZ8iNLOCkM6aScvp+tnKEZhV4qYFKhENRA
zuBwsscvYMd6bJCs36LLeW1jjwEjCSk9w1f7GgWoCameyDVIs7D07uOzRqsGZFcMMYLC1jS/49gw
M5xs1XpK6cFNpSuanMjxPuttNZSfL4bVM5ytZBsOZEdQ1qo+5D2J5g3L6wD/KS5cEwWedoxAjg4R
GMD2LYDdcIN41UPzBf3vr2/SACOIgP88zKRrE9hPXLoLqXkuK6Qvp1lDTrPetjUK1UVYbPipZTA/
2AUmMUhvJ2/iorwCxparBFpKmBl5iL6ENxqJ8qZuHwl5CsA19xAZTy64vUcYklgiCOBsKCqCKJ7S
h2b3GT+bx1UkJVN7p9TAYw2xv11ln65eP/iAN2SsauGIYAzBmdvZp5I5ReRNH/DPW84TRgSqRuDh
GjDUN/uetZ0ekiWDSjxtciuzjYSKGKkrsPHhnMM/TwL3Kmx0X+Qum37G2C6wCbqDEptZCxc581sp
jXyHWsJCMbfjAD6eNKpgdp6UqNdj4gd9Ewmhx4vIaUiES4qCVnwkbCwI9ylq+VtlQEF1opg4ctU9
10eZk3496hFyEfItS+BrXnawWs+2SoU9mDx5KjVuCsggobulec8mSzWlgGHug9zSSL0+MGtJxlJD
XoVtmImOqvJKjBCVYZ9mPeJ2Va6DgddsA3Qgc8DqGd145GteYQMiZKc3FdmAwmyI0jprfLbRv/2+
NUlzsy9G/ryuXs3MqwMbO+0QKCSGo58o/nAJqlmK119TjxVhEqoRqqjQeefuFMvIQ+YzVUQWi31Y
i2lynyMqvT24tAoEzqdfaCUOWQaS7TMlP5Ef4sLq/4L9lAWBrG6VSA4+CimQfjC590abwqn1llwk
Ws5geU+i+8tC3e51DNxEr8zSuWCaWNOfNwU26siXQ0rTc6AppBuZwiOf0eYvXfpw5cRGAzAPk3OS
OKGFTpZTOcK+2v6BmapeKtjFs38aipe5Zvn2dkn8Y2T6AZxO+LbUWGgnP2HuIK2ApXlLEJAEAKBo
M3iTmGsGue/Qi+QOs+1nkQo8NeUgvPaCcyYjQTvX6rywJX0ddDqbSuG+7RVNv7PHcdXMXmRsI820
g8sYdUwPRjtq1hpwx0AjerndAX3swb48mH2kgNc8FzJL8Tu/aRsc0cWro9upXGM/yuS6waCteYsx
/6G4XX9K26/X6x2N+mE4FYDaa8QlPM5w4vJuHIBcYt/2gecN0aHrd5sPtKs7+hlul1Ww88thr5c5
Io7WvYdLuKtGKa4hkFHD1jeXArasWaMD6cSORzIjofxhWRgggrZIWFQfnT86G/64/C0Ijc6KukHp
g4xyctoN2NZ45KRyrM2Yu27K7YHo7x8gYoiqAabTlNeAQLKLegQ46cS+30VaEV721zyM3FtiJ+0a
77p8A95OE4QkSf5E7zdj0RF/IsM6JZCFOS4Jp2JRqGDX1t/xgF4RD764CPHbvGYNHlhYhB91OzPc
4lKE/bdRhb0DdUbzwEQp6s3FwJervTNNtLgm0+EM0D3XnaMcO61/URkBHDQ6zbQJijz9rWS1XE+M
1hIiWE3kZYjt54htvRnhlIFI/ai5ubPp8jN8cXvQBKxp49wXf8RANt2yH0j4b14BnpXSKDVnuQMw
+CVl/Rdn4c3CeyTrDgNZApWPi0j/JwHpmucWUzH9mIex2TWEhWYw6IXAQN3SOHaFWe90LuYdbHSA
nBhMpTfucN8mrc5MgWTm4bEGI04RnStAELl5QQv1fqAyNiQwShb0fVzOoqYZVjJWBSNmcalklaet
vccgzkwm10MN3e8gAatZneIx4KPWGRjOLQ2S7cSFSXlidJ5Fr/jfYQocMIV1xjbLIEeyfqykUlXL
QzfBygF4QWo+WhM1iO/ckvbnqvCM8bSaRG1wW9/JKSnggJhFh2WqfkUhA/dzuKHV5Q66+3m2ecn4
kIJJgSdNIpDIsysUqunWcfkmxE1keREftAPM8ijHj3Rq2wfwo6+19Qki5B8pAMvIUIfIA+ivMGSK
3BF20JWt56AM/rsQzQuz52d57CG4Ye5VupHH3erd+CnXt1F0+AMoiByrtj/08u3PQue0J18HyiQj
5YAXYu3S9dyW60bDbCDrU/6oBghzGDLp7OSCATRuC7kko2idcLcIhzcGX2i58TWpCUWktNuwsdZV
b9vosIN528FNDPGuqGCqvInaDJBeYCUwD4f5PCYzDEFA+TLU5FW758Vf1vZMDKIUK5srsWfR0A1K
+ecozEa+EOx+wPqwyfroE2gxwNvPKQGgRVUDPcda/QAulxNykrqkvTd7UXEhg9ulZGOGgrmiV1ZO
OJLpVdHZo8RvHXKpkciUXXbD2um5YhKZuZaMF3kP51SOth1VLskgUhuUthlEa6wgUmgWQRSM4m2h
6J1z0GIvDyeFmimhspc/G/1ttVAHULgA5K1N/vTvF2aDHpoj0kNP4EQmToQo4SBL4dlXP3jXxtjv
VeqeRWPDbuO1cUqHkvqJuCxCamvoaT9Sg10HL70ggHjhZ0lu4h3Eb9wOPtNhkqNC88ys6/7J6QCf
kbwSFWsCK9PYqvy1BB6wg5KCaN1/isEkDeaQctVwF3ZyC7Td4ND/Bw7+UhKr2m6UELXl0oIIxv0e
YS1ymZnliF5WMXuoYZ6ArSYNVPWMaHEaAwM/osJi0a0pKNV9iAT16OXIN3YEsFGLK6PF5EA8WT6m
ng92rMmVe5WDHgtgObzLX7toC9VmH7i/dL4gpBE5kSTf6rEc4iBcrNP+0t8fe32lEp3uGzcBvaBf
v+QernHpQ4pckxOSNcZ87uZCJFmBG1OCZ/1b3KGf+1rmtsU6Q46+ZBfhkCVQlL9wvdHqqTC6pz8M
J3TGSIP52+Vq1igFweAIpDFzSYOpBJwm7umF3AjOgBSHj2xnGwwBxbM5FWeP+UViiEr8MKhmnNVV
CX4N5CPqDsthWDk69qZnG/BAQX0poZtGGsnJWNXNOYIGydrmK4v0KprhufkLarE94uzt305bvq4b
zQCgONzpEQjUKelJl4b/bs4iF4tfIoWWECe+Lm6h1llcs7I+p6yPGGm3+s8lWRyjYo4MW+YW2LVX
OxmfQf5SLAYp5gHbdwsuFifCiNR+qn10GNF/uFL52LGzCKZlKAfh0kTFCMivRdoBDuwwr6x0bRzt
wjeEwCcZjoCSbUbbdW6ICJ8alquCR2gUauosgDoNg1QymOTfFVyE63PVzKvCNnXcnus0Hn680s0o
WjlVI9UvU5M/XG7tf4ibBsW1ycaglXDAK1+BMZ2HsZl7JNePBLLv61SE/Mkzt2y+vlTAZFSgovwj
1nEnetQdCJmFTjTzqkK8u14pD/BQJe+7Ko2o1UR9LshOy37kXnX0L/dLNK1nCQe4HCU1XfNnQBvE
VEUL7dFtU08oi7hgVmDIEIoSv4YpET3/mOI0SfdeeEuOmjuiOP8wkQKrbjlP/V0MhlaA9pbHHIsy
7l9GdwNe3aWvUzeq7eLbEBQEwp50puzO7u1fg99okBoi44+VctNG6Eji+UADmO7NHbPnZvlGb6gv
em1R5RF6DOrHt1bAP0SMYysrQ8DVbMAaQ9mX9eAV2vmtkqQtWiyCmAD8E+bpVPkS/5vEEWqGDheo
069nU7CX+dtBmmpnLSbNuQYhnRjJ7yNY4v1GTjdL+gHdZv9XLUAsrhpGNrrNjaMOtX/3bLvKfAAX
XjKABYhyhzG//iR1a9gV8llhb+eNz6MdXwcwLsEAsY8R9BJa0h6GwY5CRNwRaaSGeH/Hd8Vq4DdN
MvSvzXrPxq4E98UlRXGl/WwazgXzfMrxVvLJy0LDKGlqLupZSnU1rcKC8Bci+tZZ/eFHVD6HXaHa
eZznZBb/NWc78AR4qUylh/jTPygL3RMQL3rNyipzyamBaI6BmGhFI96nnomRCUntyuI88IA3+ReC
Gm1/eWchlnthUZAHxfLz0crdb+N/h29XeXVsk4A3d6IBY9xbkXDk7V3G7YP4dTeas9uGdZxzFPNY
Vid7PFo/BNv+2Ojbtd6sE/W50M90mD4Q7dNxSJqCMw22fGKQJY2yUHGmwfZq0WbXhOV6N5FOsjnQ
qVCMIrr4+ndBhVJju4z5gPx434CHzhclLOjgMer0cIifgxKv9b3jeiy1iXoHnE3VQtelCeDSe7CA
Vi3tKzCxkCzZOi2XO5TqKAOpc4wfooSTCBZAhmfNcz0eqaQYK++H63x6voJ8HC57gJ8D1LdWUiT4
ey8ku4MeEQJrVk78djCjRFEMm9rJ18bP5TlK//IDNX4rKzoTMHch1ZN7Ddxy+Kva2XCToDAjsR5w
8mguCwKSPKINd8/cH9uU+RUSHjuSteEGz9cUfoUjQ0ipqQQe3Zcxm19ourun1voBQlHie6qw/Vu8
0lsLR5dnj7BPXE7JDYexSYCFQ5yODfTo8d4ldPGDyDmu3HCQehSByp2c/3paS35RnAu8YaoeZ1hz
E6vuWNebiL2Qr28SLoUXmbdiBX9/6WLATBy9+Q2nCMTzCoVrKv712eCf7zCeWRma7V3rQzEcPTKv
BJUyEIapZxjcDyphcoaTF1GTyKKwXCTApW/iyEW+B22AG6eglq/jc2cHxyQbKrdqxAvbVo1kRdHi
nWQf6ZG/fjKoBCvXlSq49JYIYbNP1XFYA+F3XR/cYf4Gn2ZvqhNpBIG+t1Xl5vuaciQTm9wy2dhl
yzTVdF2bKLzqjohilf44po9EUHsEMWRxmpCtBmrTMbpaCmQgW4r0kj2e+j9SfPdjd8dWSwX3Ny6B
g/1bn/gnO9i2WKC+WbjeyMeDcIk7GoZP6PEpUovdfAx/ZPuSPwMRXbjzhpS74Z95gW86MEjZ6Yin
IXmQ7zUf1nSVxNqhJfxZMiP0beytPH0ZBxApH8SS90Z8aKdR055X+VTn4q7NXqv34wNX6Ggf49DU
CgVWpiWtQHMSx48H5/D8hG0iwuRjogQ6z9C91UiYnbERcH1c09xBTnFa0t3uGmEfgqDQzEPSJmno
MjCjW0hwaX/p87yy3w0Ch3ft7tqALmaF8m6Tdd6Y07tKMGPDLAOj3wAeGIkuLh9w6ktw02cUgs2f
q6+QcYFiVN7ex91BOrjuLYNiPRQ+2kA6vO3SIkz8PC+7/XKXmP8NPSfirpaNxQszVqbpg9vcSYMg
C+J9GANy+EkYeItQpob6XzomPlpvhOh+SUamMzY0cUNG5xPe5hw+lZz1OCQR65DHwTAPcCDGnn1A
Idcg5cQgk78Zhzxv395Y4sULh4Ta1u969+0FZ+DQ73iJ9Uv0VlLkIiff6GunqkctrHKJ8UO83dst
dl3BWRIc9gExqfNiQGQ+0fRg5WSISU2FM4PypZSzBO+tPIRKgGEEmQhJ6qh4OTKj+QjejGIaJ5Ol
g/8WmG0OODHfVkMzAk3OkygS4XKkt5voapGyZexOIfY//MG2ahM/G7606ojFDRPx8Vu2YIJNH4IB
qZUm84WbSx43I7hVFUNqUxCkBaXQJrrtXtLMPk9mpE7mJo4auGRQKS6Z3q4E1i8EHyeFFdFPj4sh
ZVke8Hl4A4XSJF7ZwqbPFVFJ3XFghb75bs5/VROtg/EBT7ZLRKwji1DakgMDEfS5soqzKaGqrbzh
Su01W0eUnZ/aiCAxMWSweJN45KlPauE3MrTN25P9jpER0wAK8fs8nZ4kcEdqjywF/88+tOYZSwO2
UiWOAd1Ib7SaEVkSZxtF12vWzqXvy2rzm4ae5XUw0/x9RyqAj8JyWoehXxecMfMV8BlflNAbnyQK
l/nfYEDsdYAMIeN+gWumylmMzjx1BSAyuObIbfb4j8pcHkq2pdY/wkNU3KrR7W4UFlPHF812uR0G
9c+kUmQz+euNa0sbeTDxRmPSK40xrqjNAs97Sw6c9OPik3OYNu05MimJupZkWR2jTgsWi5onX7x6
It+fylH4D4UxsfWbjxLZdGd8oMsHWhxD12zbBNLpThr33PWHwVVBJVoFt10VR1kcPgZCzpiR+eYg
TPe6YpZJJ92HE0DUBSUG1zkQ4SikNUF4Qngns/CP6OpQmpBceUzJ7f4gS2sDhOEQoGeybq78ar7C
ebiNXv/Ob/BYGLptd/oJHhCSNV3zQkETeYayQLWkRrZuZ15egwB60/9NXA8amFgz4oifMMxLggaZ
t5PglQz5hDplaQ4TmONm7CPH6AYiztdk0WNhHJm0nV8VPtjsjnMcfmj+2Yfze/ptCUO0czDmPTWi
1p5KGw4PZqhbhG8xznE0Kod5U0Ld2GqjWHciflu6uM+1HoMdflKNl7rvS+oa6jeB+w44lj5t+aMB
/BEc0eCERZdpdQZhQ9jM2un59FN5Uh3whB0WidlAn+gT4fM0SwrPrOFxLjkIzMSp8KFzEjLxfbNU
11PlEEHUfA2mQFdVgWlTNkNcNZMj1CAQ6Xfsdzxm8US6wTva5k7wsj6AtBGKQVEKNT2wo7VAxTla
F/8/Iv535Bsbk4OyCse/8HbgUne+cHzhBwOGSoJiKiNNa0NarZgjBTy1G+T+0N5VsOk0DvWP1Iri
/EoxpRVk1mqMGfEUN8pOzY+M9ZiTLKvlZ6ZALWwud35hq2f6sxNTjxPIbTTC45Vhg5u0HJSIGOGe
3sdhtqqbHtQoEv/+6A8C/XI81hOpzEa5GEhgdJyIy8/3hF1DQgwEAF71zHOniArNB4Q4PYtQar72
4UydR/uY9jBmlhWTXG8ghAcea1sVXHJn1PMU/JulGx5+WM9/YfpVamWazybOOymbQ0TuGeLe0Hdc
hVsZGJAbPnPV1URwh1cgO0YopDioMG+uZ+J6yKE8ZwnHIlWVMa08lRfDQTXym04wKUKlJsFUIwe8
8/De6VoX1n7BEaNWlJusJU8c1SvkEeQ7tBwrpEX+Fbn70Q0AA9dDqktejMUIC/r5dtjJzbDUrIbh
1D7SqVtqVxGcL580xCrjHaVRG6IinPUNSZCWDS5XP/T+g9HkaoalzclkFUx5n7rEoUYxTvDWxR35
j9D9fkDqQjIOGdF6MHdpGJFOvj7sC2yc4Zw9y2e7NWHRcY/VsHOIft2tyH6A9JfMW63OgTOO0f9k
GNaSIC/Vhftha6d2KjoCLjLnAaSfgj4t0oWqVkhZPZIE3/HGG0G2EQLF+z9WjhMWdeigSFaEFjbh
4925D+UxjiuhkgX3zvXEKrUnTX8Y1fBh7Lobw6mtCr8MpqpgJDWrz1nlzdNfzjHAHBZfEbiylqkj
VIyBgIzsFtb7CCyYNLx5mItY19+Ug5TbyCwxFSEz8v5uNgVJB2hT2B17d1T9CJkaPeC0LSr/u03y
dXASKhqThtk4s8O9SDBWW3rGGYSz7shwmOIlBXQyLUHDU2XZTcnzB3R7EsWYmToLoQla6og2k0dZ
MuoG//16ZaN4HQNQ1iHpGKbOsROPLOXfMJ9HoTRsUC/kaLH1Y3uPu4Hqmpa3fabfuSK2or1U7Mos
RWZK3Xvj7+6LzCddpjt8bMNLGwrq8Rt24JTmdtVsbKW4E8XyBBc/NlxW9IO56HRi7V3TWvH0jYID
gVvKvpvWeR3wRI9qmHsN3+F5MkDJC7N5di68GALp0zdXwDvcoBq05ybrr+nZA0uNVyYNnQIs2CqH
jRRgbLkemNhx1KnvBb8sbCSB5Ly8wK6+qzTmIc6L4unlGuO4Aiyvu0C28CtJeV0ADuwu2XeH5+X7
AxbzKcM4RJjuPUCSVp7t8NLaikBVovz4P1tESjWlZkn1A0OJ/qPF9ON5gQOmSTD/KS38DTFvi+Lo
aLlIy9d0V+JLraIQaPHsFk/kSl5vkssfNfk+TYEikqPqFDkKfDtuLvPUF9ZTa/0d5akgYOu5GssS
SwJ0XI8+7lTft/lVwhE+p77SyXleQxwJ6tROfBPaObmvEOfpX7VgZ2ZjNnTy1r9XDQGK/BxkDWLQ
h3XLz5DSQNZpimHc8yryAruJLnDrntBKtG62usfHLu2m/PpN4yKArk0rL8Dhb4BApZGAyiLiT5lq
5CjGvVCZ23Uc+95MofzwnILsXRX4Tt7/I/Xzu0svrxAuRVpHBJyHXlVt1ysvl6XCcXp4BWb2Wnxe
sZwJmg6dtRWodXPFL+2IKBR0ezjXwdUiRlBDB1GLPLFrhkhAFTaZpmRwexzWIQcWwL4VNi1glFIF
+9VpRj/Ffv70ysgBs6CsdJhIZZZOOG5jp5nHlJR4DTqjGxgxLEN1qnk/ulMmvajs56wqWqsWm+SB
naE/uLzCeDMSem7Dg/ilwb1WNoAWRD+CHllj11RS8x7VgbXkF20CX2NE0z1Cf0IFiAF9PwBA/a3Q
EhqvbI29a+LN7xrApTWKgKgveokacaiGCJ6lqPD3q1PgzDytCSUEViSfP2vqP1+lnZJQMErbewXb
SXooa1YQ+liMP6N85mE3u9E+3+JezjbUf69AI56WCsiwnhSbK5GJKzLTUuNUumLlHIz5cBE+qQMA
e6iE4GYFJm78aaT9gQOxmiRFEAzAcb/tncqBGnz5lxnLqQDVUwDgx1X6ing8/qNpJqg6CPFdIr3l
WPgk5P3YRIJK0DQFOSi2NdzZwGk83QB+jJOLrA5Kw2LgFQV4nkYgEKYmyzr55cEUvw9ux6o80zbd
wOGkH5jlOQC9F8vVb9s9MwPXs7j8Ustt/BHojNjjW216FOCNUp84uTi0uM0ckj7TwSYJoc6l35Ms
n1v4jOfHTJkXP37sp4d5Ueb4h+CTlj6UagMQEE6ZpN/xDP1dJKGIoisqdz9VLkS2jGU30NXMJcre
J6+flvzPkaAhuQUcE2euxnAe08qrOBl9p3Gy4WEm+I0qO7ZZa32jfZZgOSEdsOQQyifTjvOYujZd
Xen6/CJ/tlfRk3VEle0jPAGrccxwpYlZQEkt5cRLKCVYM7SwDacTZ3I8W4gzk1cIsD9RRxMuf2Sy
HBjCz3jQEb2+HYWyYs0lbqQzLO3w8Jj0H1xwXfuzzN4ih5/devnou0+ha38LbVE7d549B3R4ni/e
8XfZFmFs5M0Fcp/LHzeY+kFGYov6kRmzkldvw7iQvI3C0xOSBkQDai5EwVAteB4r5OEG68YvdMiu
ZvYHRRR0fP7QBsYOdGAh6RxzDFUrNBdKqiv8ExS9I6+VMw1yRJnWy50c96mFmyo/UdF9oBuNY3Ax
kAalOkzr+LGvdC14+KU9PY2ZcGzOKcwJKmUHaQk87oySLz2ud9rAkWWb8WeeNkxZBrtEzwB8YuNO
K9sxyf5ABP452JjfJqosugdMpr03QQQweu/Y4NMnQjs8BHhvOzCNYM+iGVig7oLTzCY70QgS1fCd
YgyPVHXbieU5EKboqLmlB4SnkOQCEZbHm95TJarqF6G+tKV5LGThAZxReIIZ90/PyaKuijr8XfIZ
SVrylxv3pgY8h30DgdLOcAAQEb3uSYH+s/PjafbCwGMbPiVh1Ppx5sM98IHig/BTMCUwnSvcQs43
eVq++XleyypjW9ikxvswEnuhMuGwSb2XgyBQ2TkdwuXPcS6V86xLSPdX0y+MLJQJPuk1srCApzpc
U0r6QWao3hpL+FygFWLgSjrZftimKe9xAf5yTFy+32tYwyxLxuvSSysZ8C9qMkfra4b26w8Xxg1m
/QxMfOySNvCwi28u88BarLShVEmk6F9E89sN7yJ9Wnwv95y/L2dUdXYtA8QQMNLkWS/HJAyfvmyS
5E2RgSgDBSri6+ALAgTMnoxdujQJekjncTsBpgdTbNI6HHZQpqSpfOYNRJPEZKZQu7xnolFwaB6i
kyUOlHWjCUdoD8yHr9RA9V0SbK5mFsit3GjpZHtuoeljrRj3k7iLDV6pDkLTu49oHjhK3k/qQ06P
xzveKhF5nteHfNX758virx0jXLHSkR27o34hE9C1gPW/RjIP8IkdoVWg4RLCpzoPwrsrbOYfMz6B
xFPWy/149Y3/s3LvW+ojdD87jtIN8gqoTL/sUhhqqI8WDxNWxoViLPAuIw+gE00b3QZWNLeaPoTR
IY5s6mwhO3XhZoJ9dkm0gD/XOT7cMiER9BcZnjVJTeESVlvQ/NVAUugqq6gaPuZna8VWN8Lriqyx
nWbtmU+dGqCuoJo1hGM9ZePLw05iNXkAeR6JDQaBylVO1KKM7+0ocABS/qdzw7vFbrLRuUC3SL9t
vTJh3JgKF1aARQ0zIQ4vMN9r14x+qLJSplGqNuwFhwy1TQtAR5G10uHsOxyXkPcUfM9b8m8cgOX0
Dk204+udjRSY/RkohK3s4xYg+F8doCNlW5qH7c0hHe7gdiGZr6r6GrKtQlq+JCaM2ZHT0qbg0Z5T
qjFteu3TrFlt3NeB8knkKQmi/yPlpqYw7kaZZejg8qms8dx1DbwLYCGbvO89dqV2DuIisoI45rce
STByTeqKUFFSRUeJ4f7ISbDOrhTyzaKXLePjxVT6CwlKnpc++iiqzgF0L1/RZKgAsGCxMiQDY4z1
RBLRrmARDHjEsXBDnGFvOgaZ8ykvNrZEWNWinx3lumd+8qnpi32HECFSHg9ned90rBAsGTA6lwo7
cPJWz2VxcLBwhpglRwNUIZ5K9Y04dryPbOWRg0wNleen0kiTIm2hJ27wrkxXxzzn5wkdoJluqIyM
74rsSBlKDGUhDOcg/H5jjYxX5j6rAOTvL+F6WgW0SeZ9sq7W/iC5JoEsSwXwrNcf3QVI3qQ6lCMw
0juAusRAq7WUzcPvugZOzmAJxior4PhX+/7YDkUPpr1Q5uTSmS1f/4/ny5GYDTo/N923dQZQmmZ1
StZNBY5ekw9ibMIhs1/+jRyFATeBAkqFD6qV2Nj3MCQC8ud3EdfFRMbp1AQe1ZyflU849M3joIof
Jz8iPH83FqhQcIAnxe0zaSAYekjWYp6b0kS4B/+7AB2OugMagcE6LBb2EeKEiN1ZBtku6OjPG1ME
UR1YBFyhJqHQatRdc4iZTOqZ4zw7EM2q1LZq5dFW1XTOiOtR/M6iH3/pK/ByegvQsak6aWZbDgCT
vr//lnyQq+fEhCdZs1w7mckKKbUvsQOS9IsgAKZbLdXV1CbuAG0kpq+dYsEfUJVhu8VH1wNGBoCE
iD8CG7Y8oFVDSe3l/1PsX2ewy0buqLGUpS6gr8hLUeVRHWabgcDyl+sHmuNPzEdjtic5V2t0Lf9d
RcIhpglS66HPZF/0Bxi3ccK57XZzURjJjsMz64CLMVdR3UtDWmit0Mm3zzUVx1kpajadvqfa8YgG
D6PBChI7ufqEgqBpAUISQcAAR9dBSmZpqTJkdcJ7mxlzwfsm2mxsI5gSBsS7A/1Q5hiEZ/1DlEpa
ZkKXOFRAsdffBD+wmlSdUXn4O9qdG0BztL3vTfqbWCV7SgAVDUOdcavSWIbZVawKVw3aNl2F4e72
UDIMCqEYlvMRDmEzRCd1aAdK2xO41J5EDZ9E80rXgZIEU1ABp9tqDODcn0ecEBzeQHPjmR02sBMD
Nm5TakNoponozDg7oOy4nhcAZmm6Hl55TWTqQl8h8m4b5HLYLtNtWKR5uqgZWOOw0e0Gg73f+cjw
WXV1jpwx+sOJH6eQ1BLKlI/Gsu05iGlm8ngHilb/r+XrbOzFZiacRyunj1LYcBE6KPoxQ1kVtsqo
4uR6bf3PDj4MJ9mlBJTQzaQ+9AAa80Aj2scvfNuYBAEA5Zn2Jnh8nigZ1RYpewWbXpFPrn2+cU/8
1FDfZARqK3H7zdG7DcWOyPh1no5A5nA26DNwmaL2oFtIVbcaaFyhlaY5cl8xaXN/isUzcWmJyy1e
b5r5NZIIb2zO0SrJZ3MCCKAM+V3aDm0FQdy4Qz5l7aHRxxgIah/MTuobF7+SvLbbUl2brz3AMEr0
MJUIOubOMyHXcdLjQrNiu2kGWUHtwgxet28E01tK29YXv52tpqMBme1Dv1NEVAwh3IKKCEpSm/KM
Ds5cjMDKcfsjwoTuQLrAZmQzdl26OXkLBgEiwnSMS8rGNg8ggywbS+Z7tRvSdKlsWVS6AObxjkeF
QjHf3BM1IoH2DAJ0e71S+7wCCWGSjjXZEdWjdonNfCZaDry5Usi4NkERHtytEHLqoxEkoUalN7hQ
jxIiQ+cr+Nbj0ASnX3tP7oIOJEpTEHpnPKDI7wI9f3BbOT+YcweWtEGpYMKNq4UzwfW9NWhxepyQ
E9Tdn6GQ9b9pYAw66ZIw2KRvVILrRwl8wj+BNn8/85erHN668T7wWcUPZOCWOXk/GxNvQASJ7bk6
kxzq+Hg/Md2uU3MrITljEDO3Chd4o6tDmScGJ1XVzS0gJxtBWqtSdtffVFkB+oDfKQZKRb+WnkVW
8i7/srwL+2G37TbTJFCWo7qLyn2ySJswMCgVIMAhKWAzb5v3vDO7zr8cDs1akZ7ErXWkaEs6p3i6
Clwy3hSAiCOkwSJPAKt3zbLsghC+NQ1KtoSJGmX0JxEgLJ0sXGM4nGksDWkMTq8pqGMp9L1ZJZUM
Fi+ft84petyVGEcnn8HEyyhAfcg7S8xi5U3dhuOcuvzKcnrS+lQIGLmPojpShWN1rjRP0wSN4qYs
VVEwWcJkwW/8NXj56hI1vt3keY+6igfcQivwzK/c7dSKX1IvxNNRDRCaAcKO05uW5iqxcmhissrr
wpuNjtCefFfpslW5WsYCgEIva4qR3hURcOghpJzqRERKWRmSM96+fsO/ZMVKzNy/Tw2x7yjPqLEn
+V7UlhhiafK86pg9t5EbqQ9mwrTU1etuLjk423mW1wCWAcFo7IMvLgRZgrZ4NaTUHOYxKVCHokni
Oo2arupsJv5QafWNinmiAnDikYbrZJHRfM0GvRDiy/v/hN3Vd2XbfLVqcLJkXRTg2dT+dhghgCKA
yQxEair06555CFN8NqJxZLw4h/hZmEWE/G2qdg7/1wP44ZAuxLDxUUzV9Fl60SyxI3iy3bp+7mPM
vN5k3Ud81CmQGoZuz2fpYywoXzFg3Sp7ilHrT6BurgrGjhus+33AG9aBBeTO9kTIZRPgSoYbxt8N
agKzqXXGKGhJQUeNv8MB4PCybVZUAwEFnCpTGfV/Bafy5EoydkMx7XB+ZrDHDAfOrdpUwdN+OKfu
MdWXm6xqe+0hmuIspKo4FrtgCc9S/GuF0nI0mouLJoLmEUMSaH9rF7iIu7IzytGuNabvI/t99MCv
1Qy/88eT3dHOQrW5vWGoqZeMRrJk+2bD+W4+FzBqtvnpMYxrkQs7iiZRvE4bCHwKhR+uGeCs1NzO
oSBHioXA9Yeu5l4QePMGay2RBEVHBFvxKUTvVBXj8eHrmwk5pII6JQ0MJQkH2QfQ923RBcrU1I7k
IxBiYUPqPRC4imhkbuNhkrmZbqs8YM4V4OSHP6Yn7YKs5wGAEn/D9blVOF1mwZm+iXO+El0/8j3s
2sn+OeVoR6HiG6QB3P6vF02qH9KNh8wKJjRUYuMCuZ/KVJZ94EbfN7smRn5s6L1Gm7/VeYUK/pjF
zy9D7mVV5di7sgQbEwAFW2myBzz87tmwXTco6aEXpqu+WUrHxN2hY2XgSKPzD83fYZpk68dPC428
kVwy1jl3KR+TzBdsP55jRI9j9D0T1LSqwru5ZxKpDkVNOurkfnkrZEFzFvE8C9i3ZZI2MdUmDNKC
/gT5IpvK7Ir0lSkTtX/75cP2oId2JM8LdjDXeM9HUJUeDQHLkA6e8cP5ixlwCC80dPhw9Fx2tgBC
KpiQd6Yf8XRt5oi6wO8GC2lVUbqGnS/hxGp5Z/BPTnV6KpRtB6cn5nBeg7elSDGEK3ZnUUZheUCi
YsVsxxp5d+dJWf8vpt4iZN7UcOF5P8lPeZdu4lgvKzJpjJ9y4KmJjPp0Ad+/YrVD+eExdxCHvhBB
oaAc7IOrfF8r+TTcq3xksxS7PAG81os/TvuGiBvTLeH5ZGOtKBVN8riM2aFmUmuV3OIUsf3qdrgV
iQwrEPnKUZLu/f2RyQxgRUy7jqXLd5qBBmaG0gYfgpEE4vx+imDHTAChGBLooP8Wr56nopenhS8a
WiOP38CI1WIAeaUj6YERVKiKBgTk3k6Xye8hbay3ulzYZxbVbYTHlqHHRevwS/WWRD8Xtxe3ZLG5
sg0q7gC3sZrE+YI0a15oTn0Yvd0B9pFdKD77vETfsttTpuXVSRbej2GLvlVDg4gAHwBmP+YUj/Oa
KURCRjFTVbADf2EYt+Gled85oUNOIOhk68BXAUbza5guTH578163CRTDF+mELSDsYPGzvZshYZ4/
jVTx2YGawsFV+pTP2ZocU2wn1kdGHuCA1aXGrMb5e/StRtelIdCwKhCms/frynr5lz5RNr34mh6u
PPtyYwPet1yNRrKGOp5k1TaDRIoqaunkFEM98LxugE+tk1oNCtg7iPbU4dvgJIOb8+iGgmUDdTG4
DWfOKC2aXgDEM22Wb7H9Y7bqaR0X27whl68mhdiMrqHT4tJfYz0LFxN7kqwqToYvIN+aoap0B0fC
opx1D0zLWv9xLma/I2OiiyJdN+ZkQtHNeyO8HURqDxnILRF7cu4vWlfA4mgI/u3cTUDVtWKWQmW0
9jJk2ej1OOBX5rUJzvNq8GFJYiNrcvnUTEKBGs2Vj3T9z3QIEebZDd0zHC8o7KBw8CuhM8eD+sqb
WnnG0XFYA7K9SlkZjX5VagbwtgtVJBFFx4/lCLB6OTwun6JWeE9qzjfx8ZWpQqQu5TWTfcDYfP3Q
+exAaVZKRMtXAMoavlCy+EU0iubiroEJCYGJknWCgi9e2xLQknZMUPNRiqyxuljR35esK9t9KFFE
FGaRaWkhQjDAyMtcqwktz30dMA2TKtdeXG2VnTnDoJJTpLjM3vqmpwtLP8swTlHarb29P8Rk6yex
nWgwjp9Q2LLL9Oe8xSeR383VKvou7S0mNNO6drZPXdPtVAyGjA1sqEaR+3Re17OzLqWpmJhYXFm9
gsJjrHPI6ygAQFxrAxcmjhnuMKz0hmwp18FL+4DponTTwK61U1IP66GrhxVR+XgnqJfIVwE7YYCd
rDcYbQfXswUmSyZpq3c0HIMiB2V7KZxdXXtSeoi/lRBPi1uRlKgvLZLrQCxmTfe8MVa/lP24VW1L
kRATxU8s1ig6Fm4L5PQVd3fJh0FqUGJvpq8nK1Vg0NHiNtILVXZLM6ddkqm+t8MEN8vQrnxa46r5
Qw9nFamAyX7ndYQtAfSJ+QDaJ+OFv4/sox2RaBMGpfEQMa/EOeYJUgo0nKFIv1HHuDNx2ZizJ8MW
SBOI/40OdjWCUDrPudCF+XyeCcGKyjDuyhRuTFNlIwFmalD46eIofrsdx6BrWHtWfCSORORrJ1C9
3eA+fa5WtB8KH7SnbVS7hI+3yjLHv+Kg6N69+kNoyw8KQhWjFDdpGpeq5u+4gwWPvb9dqyI43Ecr
IT2XaotKCKygjkO4CRUA5s+kTFuMlzlM1ie5a/9EH84CByJKLklDZpMsiO29Zt2vOWnZD1S4qwcN
dMVdLTRsFbmNk8JNPA4cUI85tiWvgZE3wZx0Nb3NkvQqnHhgaHiL0Vm0fj55V7bUKT/b+NZJSH06
9wts2QTQPyfXa1dsZ/1s5cKXFUDnno45IgNQPmbAbHflVBdx8LwkitN0jclGnuhPS55F0J9NhO2m
aMCO5QpLkZS+/qkRrERrGawNozx6M2ZQxOMSAxqOHU525YrEBURS7ptLNUTXgqSDjw0uF0Vcxv1e
ps1+5fMRUK/nnRzeGxgR1+JqfeZkA/VhHek480eOsq2FoVjuDd/AbvTM4/7wa2acOffDpdvSt8aE
px9l8U25vMHCIxrJjO8dgTKW5O16IHLzm8gOGgP7w3ZySTiOx9ubRkM2CoIrDcd5WNdMD2dpy+dk
EtIkY7nd+iREMZrIkIg6SA3ELHLG5pHorxZRt31qhwTW1vcm+x1bQj/f+kBHKXkcxIiCTE5DSaU4
Vn7xJyOuNfbwocz9fJm+/r2wCwfBus70UYWwd85H88/uAG7rc2FSIEWESHWFldjcULsjNAxOBggR
TXCmHp0G6gvax/Vt8E+HVT0UeuuoViP0+pXxf1LP/6IDyYApKXoXphUWydhUiqtHnx0QiSC/zh8k
SjmH1519Fbq9gcu0mcL8sovggFBVOMyBpbK0E9cYjX/CtQdlroWwKTNhLTdNQ+sY7l08L/xFHn0Q
nRqCsTepSpZCpiDv/QrOzYCPnIVpdKg/MskHZYA+TbS4BsUqba6svR81DA5U4VeCdg41weF5Itl3
AQhcT5Ep8ZSPNmF8FKdD0mZ9YIOZH/oVDl9Vw7hZkRbT74da0fl+zUSJj7rkyxYd83KrCZNdnK6j
pXlZe+WpH1AEjqFrq+ijx+sflPXrsAQDgujtiCAswTLalnClA3QPNtyknt0SI1o5kCOPufbqTQWa
CFY/dp+XM85W106x0GiHMflWipqaocPlcxj5kOcJt8GEAjpOaSz53nBZAdRv3su9++2O766H0Rho
FfmK/fDOJNLUPerZqrNdAAbdOOUbeIbazc8HccP+Vcb9Q76FzAyLJTCfURsd7t/iLBJM+tJflrvw
m5kodMQqUQov49skCgk9vnWZvky4FNNrG+RcSvEPbKf46+kdJTluYexge7JCEa10xpblLdAV0P1P
Mw/dJco+YoR9LnEyKCimTzUQ4Laxlp+2yn1FTe8cZSJ+4E0u91HshdHvlgFslQcIk+Z3fT0vbl/Q
4LRsjKIfKza80V28ynQjIau1QyHYgbAF2U88MpSnrw5xukEfw/MdsSkVpnHfkC8hUtRTVf/X4s04
xhlrlS621ONMg/FkcaNkOVJjg1EtuVR2Ehv5VuGil/9wCoEokUfGqn7ACtes79uJb0XN+41H78XZ
hIM9TFyII4seXyab2/GWypsmynmYEBakj7x8EL1MsO2AJ8aCFXY/7yzDge2b52a3Wl8TrOwmOg6n
BAfc2TCzxZ1Lw1cu/lxqkIS/bQsynnA9ZQohHp8oQKe/6zo+fUAd7KwJAekm721D45IFdDqVcsDH
FOZvSQKfIntO+E/SIhNJed8LbUnlKWJ0hvuoGT9AY9CM+zCEwBzzS1EG659EUmi7WxI03vhOvrJn
Z17sF4mA3BGPrehYC/W4TwlcgvZM9e2EWSOHxFPdv2P+tWCnRhT1DYDRgvE0fsyrMzMQhfjR/0nE
myB7fEwTlqD891oRH2XLpNNFBgjiKE0V1apMnhqi307FA9R5IjqgQa4HkOzy9zy3eMX9MiK0X+qQ
Mu9WmRtZa2h+o9p6uvl/W3SHFCbJqzk3uv/VyQbmcSXHyqm8oAmKHzHcOmnQVxVIpDOP/+2Q7sBg
tz+rUe6hnnWGBp9qPnlM97aBXrJZOFMS2BWxMS3ijADlekAVZhxjaZYb7yUSOJ5iel/nnPhBma/v
iFhRwIDDLSQYk/7xOdjKs0UvgA3JsA5b0m70xck6baA1JxZzuIOMk6WBQVvCZq92WaeX9wWCFrny
Uy7TkpdbNh/7FRpZ8UHyK2Y5RQUtwhedbDUaMnBiYCLb6z5oxnvh8YqmSEDejId3cygba0nWval4
MyL4c0EefcABCqxjTJgMQlrWPqBRlKpL8uaMZvcwe8D2naZLmBz7scAlI/pF7gEFC9tqut4EHGRC
UWB5oK1lde2kNLObzZqcHAA/FgBZ7pxsxKVLXDO9lSNyJrRA71/q/qREVL2FY/fXwB/KwGneAoPn
7gh52aYARkil4nlYrSSF4/jNrJRt03QENSoMOuJUhS904PveJJQOOmmMn3aMsosA5wbXtHN49MqJ
W2UttKCx9uTPijiZoFUXWlTs0AJrab2PCfYWJeKymcBmvYTctYg1pHRYqBzGj133vONYvPJo88im
KSFBVGsVlTE06OY0sqAq48mPabaI+Gy7D+ELpIfr+SAPbRZmsmxU7/jfgdk3PGcqALiQuPWvaaUT
4SjT3BrxPJFtVe/wPzX1B4v9z2dNNDYRybHK6w1MNRAzxdNmJr0vPMxGUNw2DjHkpDNLol4PSzFx
lgPIslHHUM2OQzYQCDOoR2zj2GbckC6vhSrERYVpbjAuS2L08qIOgbCPmtmrHn5FXlcRUWW6erC0
aJPFQwXp3Z5igL/BUoaqLaFS6MXwxtYLj4RoS4DnypPGmrAr9fWCaxZhEtlOmhpkFuarYGW5FjZb
CRC9EvAhY5Quwx7xw6XOp4TLCViIknqQ/eEjL4sI204oJfbEQAJx2o/0cCxEuXwRkwPv0kpq2+wz
V5Md1hR63AxKtjE1TavmTvbt4td8gIhw1cR5xtvi61ydNBZAZytcuBgkDeMAtbaJUJ06kEnUE5UA
7oBL+TgNlIHtIvGultSGgFrX+4vRxtRUshkn4Zrsp3PsZpvJi/fyZ/tlJjvaTm4EWcAlW5a+g0Qn
jngzARY1vmHtxTIi/6yJB3C/IhrhH7+oy6K8X5NIc1Yd0ap26VL+4ZTjoWKCWGWPy4L3V3vAbyvw
dehj/vsqpUDhcu1G85Kz2a3FqnHWQvkLPWE3z9e6qskxySLzScLdg4AtD2uyo1JjXUJhsLbYnqiq
WbCRzxx1eBmQHDh9tsqY3E+CqquyRCEC6rncOrnIULhNjqRBS6nMQ562P38svBB7n+wHIqXQK73n
2Z8tsWWRqUgi8pqD6I4dTlW0yfve1Eq5v0ZjCJZcoH+a3CUxZNPGvrUk0OYL1qgOjIwvHINnUUN2
yVHDojxk2FBPvRw7j8F1dII6gMxjO3lszYOeS/bEOryf23UjUATgjfu6TSYRMlYvaD9nns4gapiF
1Vk6hOQuvObHXVaR1M4w4ekThDt0JAdlV1JbSG7Yg6zUOJyTjCAo9GtvXS5ZmOxZR56P7P95vy4H
Rcj18so623XQjqvwDiDWo3yzVqXY6QI1SSu8elndAdVQxYm6aR5Xt+7xoyXGFU2UZITqrP9pucML
KYydNuT8h3kAlVcuq/sOvE04waSQqgKFgwG8g83nne7646bi1Fc53MNQ0Zum4cBpFrFkz7OXB76K
9zVa5hN4Qp+FdnZ2KXK0Mei9WHeP1SYyZ5C92ZsCJoMNNpLqjcKO2pi64Isd89TWl3bRy8Fmgf1t
CMwsM5yiDsVi3lbS0sT32vdJNGZ5cF4BGUCJkm24Zb4b+1rOVI7ETg7RfHvRpM7W/NE2e0Y07+/g
cDVrUJY00tJFJp/qizXmj1SB1mX4/7xn13HjU1KdH4yMJQ8qtEfKTijp3so4IOPP4SY/qRVxrV+T
PYoUH+MEdJPQVktW8n5pOVbmyLPBeKscPPds7cMmYHlW9tV/+SUyHfJrDZeFpBfxqv9KW/eE+XMm
q6jrx8NJldmmu2yX0X85xThfp591lVb4eDzCYCsd439e3WJbYIVxEoa9BDl1Kp+J3IuNSX47ScNO
VP41z7uFPhzDq7U4+rSTGFb5w+cW1EOo90b3xZErc2Sc2BL5jOIz93U7Z4x4wiBc8yBtBVHBJpTl
vWtqs4+gOm1I2pIND1L/FzuP4gzXJ+KmQcKmkrQtDVmlibiBrZ+/c7CUXM1Xh64pf8VQM9Yq5irA
hYroWcQYAqyPoAhHF8tqg6m2FDCxoYJgou/K08xdov6h51+Xkn8dRy7ZfSnZaWTJmON+1ndn7+77
+uK5cXIAfkmtFFO8J39Ot+IZaa1l7Z52ZD5uyjH+uWSXDk5QjmNNswgpGRf7GB7I0W4z4l1dXF4/
PZERPmQhEtxv8StrtJPf0WMh4YrBmldpeiOA3CftagztiMD18ayhhL+qWIoGbWG3+a24BcwMP1Ck
1JRDgWCzp2FQuiHspD1cjnmuEwATTGM7FyZD18nxXZyfNSLUoZHXmmRjnsZ4qRZtzgk4IzGv5DTb
qZH5ZPodwr20MlYccnqnJeaaOGJb6asorAaU/2prG+/LlEYopHaop9j0gTzwf+lgl9oAW+mqP0NC
V8kaZxg3yp566eCqvNvA3Hkrr6M85DHXErwIZ1lfjnVKg7BY8avK9m/dYt3wfH8Z9Wl9GlKZDpvh
aD4WP4ShPGko+SZX/pOW4PsFjApUxnV10CMB0OhnxYYY93UNvDZUky6zxPFwRyxO/KGNiQQF47Up
i2ADsx7FTSeJyrQEVu75ZRjGsu4Xt6He8w2wJNhlJUtDsnmlaS8dlWwJqiKUhEPNdSqOxOqUrKnd
DA2UsrkdRgjQUSCAjOLpOfHH2XqHBkyycd+Dam+eR143rOrgtMfz517y9cRk91uu9F/CeWKEFVkH
q7fTUGkfO7N9o/a3i3bLSWSu1El4v2/4FbWx8MWWiQqiSwkdjU9U42HfDCX1UocQO+RnC3BPWMZi
8eQiAXpc5VJ2g6tUy0QNKUUPJVf9onKNf0a+JO8/LfI1BhnTnoVtp5ZoItaLiU1Jm6OdheZRmMpQ
nFZZikH0GGnpb28G2cuMFzjQSqz/K9xq8RPGtEUs2QPf0yT8n+lkvsTs2TKY9SWmbgs3GJtCsdUg
KFD/xIoZsKqNYVr940u84C2k4feukLbNQPmfJnJ5y1EtT8l44pM+qKRW8vyhYxkKY4c9aNjbwTu/
bNWsX+mw2f9VA4SuVWC5kbHttIJYhySF2WlpesZC3/O315XO6nOZq7LstfH1mCSryGzSC2FzQ2i4
j2UcsM50GQcbVnUBau16ezV76KygEOO7Fw8WKMHRRnkzYJM+udOh5AG1HpVlkjryMGdj4OAeOZBK
KXfBFR5sv+bzyzQ61sn2w6msFRbJwaIzqyFjPqiq5yNilh0+C0K3qcdhswoyvGcWKYpDKr19s7OZ
wrBv+C0sLaMi82p8Un+AwjSsFJVRBBcLhNU46HEGmCcBXNh8afnxG5dB1+ZoYdx3cXm8UE1muZQC
4UwGOiYCtfEy2bIY9SYB7si383nyl7COb3ro4BbYeOAOZehBCL6f9k0HYMbobof7xMstRroqEwXv
WuirTGQ/DHRvTkUc1q6J+IdRVGM2uFOwr1zItTxnvXGTFBNgEq4xifpLH5NUbUjM9pKNykFaQ+6N
izSZX+YeIfEYfu7EkZACDiKAb9+jpKla2t58mUAAiJeO7wC7AsMS9zoIsQ60Q02IHW6fiZRcP/ef
h+rxzOViXj+0QJ+HhIzUac2TPTnbCw99UCKyF7BnkGoyL5pnNdWVUF2lu/oJFf8lDxWfLAajZwPM
3oDnqozli9pW11Gg0KyVg2dJoRqU3hZvzg4lthk1+JhqznGsbzTJWHiUHluYhW5dQKI25SvTIEw8
WppWuxH4yECc3RUjtknL/qPtp8ufxdMJCVi9nlXuFd/WqXpoMoozubJvqATrAXCfEJI6j1sMjEWT
lZkXj4nrGRZt8OMaG2exS/8TItVAKXZM6iBw3ffWqVdAiaSJgFfShXXmpADcLGuq3Nsj8Y6Iuu/E
d4u2zd0DKB15unjRTKiZof4N5ojZhgh0k/bD/CA2Gbrt+ulqf8UxNtzwxL7ti+4fbdn5IxDNWnGk
v8YQssFFWO5sd3PVab/UEWCQIm4fH6sYRF8j8oWUwZPI1stN+tfiJTV5iEGAtFKMGOputltdineB
JVuFYTc4i5jKglH7hMkuM0BUcqSc5Mzv3p8UUB8WDuww/kutBUmeWb5b1WXUscs2pU28JDkHHCzy
Ar7Th/qbACr9G/lFMi3iXIdJKk/MFaw5Bmi/P9h1YcVrSPz6FsCmhdujLVFR4tcK3WONIN2Q0MK/
iPy1KsgfIgX2epHdv4TORrgk9zPSdubKqcxY/nQicpZAKPQjaNtJpHRXHkRg8GdMLD+OkM6qyoVo
HEYLZneYVotyLic39s4FwqkKDs/nM07DzLJNJ35xl3O+RxcYwexd3zBqooytg4tl6rR12xqPxw4J
y07kEt0fo8ijjfge/YSJJHhwKMzj7fjilYY1BGl+5escPL147awaoXwdqXs7Pbna6DVwgxKSAPi4
MQPoPiid5LQmPoWImTjM5lvn8IQmRMGj67Pdjo19/lemfQgJWo6KTHKgclo2J25z2PXVehYn7WLo
X91hmNwsLFW2G8yhr/GDAIgXrhifogcAi+9GBw5sj/Ol0L1shjAiJKQb6Vbj13ZJ1XVRnUqDLL+u
ZudOe601EkRAa9hlSgCJNCllnWKTntzfgu4nJr0ujmufXii7CyTmfwoqUK8FGOTg3u8gi23vVJFb
c7Ofb4LwRGW8CrY+ha0di/EDiECnvYNUEyK4e+xdbvixVyX/XPCBSA1txaRyzmh05ezQoYPk+QyI
ScRAU+RlXMLcAuFoLslI2oPbFwXbIc5i95YEu4C9h+6oNefxDfslFXsoAneF50/SGM+1u3Bl3fbp
LdQnjDh7IihoJUQD/G3jnhL7WTG/cO53lND6MiWSxYoGe8mtVIyxGV39wR6Ub9D+2yYBCv7Ps8Lx
Ndssy0/uAE9HNsB5o4MfimefnciDPqY3WCB5/z1oHKXPNPHs/QoD0RfAHRgsHbw5sZcLAyBGO3ES
MN5n37bPJcwlZOZQDtxLcBpuG8H7b5jU9G0xqTVYnnM3D7vVjB1PgNsJ0Ym3lX+vvcHelWP8N69i
zIafoNlDh+RvEXrfi9/ljKU69dVdOQDALYLqHsw0cfaFfwKtSQyJK4ex4rtPcBK3AH3o3SupSCfC
7q87LeXoCmSPv5Vp8u6QPhAkZDVylRAhzU6SMQw5SS7zH8/QPgMkxmmPIC4Hnver4oH2blEEv6yP
sOYLsnDaheWJdwgVxaaO8w9g3DupflKu5rjZAzu3B2R29BX4BfbOOAPjFcumnxSy1U7QWxUp76A1
udE+BFmcYfckpTWOEOc8U37bDLG5SWKp2+sRSTfSeB5gF9hFuOyygccpgRhZb7nbqm4Rbpuy2rWr
Whx3sJURmmPb0IVpXC1m3oXxSvcYNp4rN6AxYs+yCdVvcLy4QSBrDO0mhBbL5a5g+VsP+iMicw7v
OxeCOtKPOYzWDiGgktzzltRLcRP1n05vSFpY77Y4PiYiNtrkssjHtB1x8whDaO//3gOGDFGcR28K
9eGVvUn0kLQWD7EWDjU9xMyfgBvBeLI5U9uwjGJ2bH3Nq89NisrUK5IKGEO1PCenMGJx7Euq6Arp
An33kKavWiGOImGgD+9uvMj4hCxvc6t8RLUpecuiIislhzIZ9bKMe5GtT1J2xeL/B9gIXPP1PoZL
ine/qx1VRmXdX0lk7GYcUA6KM5n+IYNjHyV/HHhbD1zDj1mR9FKzHUFfvrKLIdeuivJ2brcDuY2y
hRunndtzycqofZkAVKoUZbF6nAvRXl5qeJB52beobeW0q1ky/V+53IgXuiYwwNY99wjBCuqBNwh4
KlflVtjiyRoCzVxuBcTrKrhhB3WB8eJQkBUXggPnYfgpJLkAoesP6xMsSleffyqme5n38QXQk+TC
qbO9FQEDqYVQv+kx+mDOeEU+fgxqwcJJ76W64ggJK+cHddhwSBAftTVvo9StxfypmCy51msat8XX
7eBhrlEh5EvUuq0KuShml7CotdeRFnNb8iDehnrXgNxtoYKLqLBgp+7qPrhvY47UcsekD1FN3xbA
l/nvELQI161rWzxn/klI9Eh2PVuNPdEuUnqc67Jasipbv9FVXqzgz6EpDsWsKvh+abR/grZRRLuF
/VsJ76GTrpSVzD61hR5tIa6EzPF0BniWTuKKmHPmlNbe1DGUuqGTfiGFluhVp+s8RVXWHIy1Erm7
fuq+zUY79T2KAMjHQhhOLFe94IzQ7ePGwLEAtTAbiVTHrU/EpDOVwNyXzXI0XtIzYoa40by9iC0U
bCWwx81LtAJzgiO8rZLHqFj3ifipmIzDj2c7cepo8Yv18hsHhgTd8Z1a3B+bDKTHPi+0pHPz0qMZ
T3NeoxAHZav8yxTN8+9tBZYcZPZp4JdLwepy+T0QGEdzHXtLIGTWhDVEHIRj23KSbyo62LfeYSsX
/Wvxa5hM1aqnwx1ce0PL4Fa0I/SIx/kGopoW84TAKnarcn1MYiaaA47aY7wI8y7Aqi6amQTawMMn
ztu81F3Vgvo85vmo7cWlNFxZMfHqgCdCpnTKFZ97RwI2OHoHURTUbiq4tR9Mp4GTbNuQxA3d+lKm
Lk1+TZ3ziBpq9LlUdoSL6nBuhFnGpiGZ2yjmDjU65VVnrFpt4VGP7oY0YD5tnz7/yJUQ3ZEzeRfe
S3IT1LWblOnyybfvvLhnNa4Id28Xh4Qe7eIGhK7dnSRrcAqWsaK3AXn7uoVnQP/BESOZMG9TmddT
+LcuNiEBtk+gGLQ4D2gNZ86lvgzCmDV+pOpnPQ2N4AzBTvkirkKSvsAIYOsLRlm0ADEj8C34WuLK
Cq36EwYFEAv1I2RzaaW+Qvfln52Pfbf9CemU926fRdIkYvMfKPiRG0UCCKJNeHhjtbhpEnAG2v/X
3OXmIPp4/kt83SpfTGvhuoIX/uQyjCCB/TIZ6Dalqpda6ymJh3/ZX1CAjXbvWV9A7dskAfaCd/Yv
+FXp2Rcsk3njHPCEcA9whJ2QUpSxInA2mPTKaNmjRUhmGZMMySNAwUj1elwKvbDWG0N72MuT6nus
LKKyQXOHp9j/iNlEpkexniQl620q8swlueO22QJVIs4FsBhiDwcORE8idtilLbpW6kD/Tn9FJhYN
4CXgy68rqLhHNB/o4TsgUvOzzcVYcTuaUmiXD0AODxeAaXzRM6EEFMNgYw0TJSSp7PeX+XEFCaok
3JuQc/I1VZhCuOTr3R6HZSpRx9beo3rwtfb+Xy8mJQN+kCZr1w94uHGq5NPLEAtj5S0lFgvFudrg
cUx9wZwdyVub8DPCDDPtbK1hp7ILElHpp+68sNYoXDdeDYvAeiU81LpChJbUA6e1mfMM+mkiaQlF
0xnf83oKgkrS+7h+EBGCoNQJ2xkLal6yHDwKg3AAJOVQ/pDWpmalwjmFO4SODlWnhncrQYpIkY4j
nXoLEHAgkTvZJHur67uiqMAz01QqTkN5Kj1xuQ9yiAxPULKo1Q36tcQMAiUEWT9H83V7lzXjs1mz
HIzLJRvAJJYCYHN6Wer23QTmqE7wIplJizKF5ceniHnD+f1fJ8my/C+QJ6Jfo7d/e67eg/pdnfle
7eI7S2iat1XaqgidzaquiLB38Fg/ZAViNe+lX2ywnbWelc1hDaMR+/0G9nTLGlGeu7zGUUApn1+9
jkK5T383D39v6fBY4k5fMrJEEvIPCvIz18VWy4MkMiipklB7R04MRZeiMephAf7m9M7ir7Cm6JGu
bBFt7T0dRN9VYPqGDlWpPyE/++hpKrVy+Ii527jpp6TebmRuZklDSISDT61Yer2miM0+jq17utSv
TGrkcwiNGwDnWRfTIlJRNwmisBJzsKlOa3FfeGa7YGBnpwjYxaXLySpvOdi9Cz32uoUPmcZ4RiU7
5gTIOSkq3uqJfdJC+RrRLwvpE7ffIC2qIjPV9wEJGKQzA+xJgCAc0J4qhorRLg2JaXKnefxJ+R07
PgtX/fhI7XAK/fdcaQYAJEJk0emTrHG+qAgo2OkNfNFHuiPKnKdcGYsKsI6+BIBMLH/D6vv6/s/p
B+VhxhThtYJiB4vthFpWnFcws7mpYEzw2XlhkKq1S7LzhuQW3MQYepCxvaFvgjb6F/Lpbyo8YRhj
N1VE8usZAmIJiaQTkKBNvJi01/AtrCaGX1cXWs509fJF50uvPBbk47SpQSNYWc7/2jM7x6dvZ+uL
WYkKjI4fIjuLzaZV0M89n8zzFjXJPQkusB7u7zIkFZnb6aE/DPmkM8eLdQMkmE3x383KsSuS9qaz
wc0C1RTbvBGnhrw942EVz34vvmC28NdupF647kil/pj36wTb0RU6QMBlFsVlLRCDj9DAT3oud60/
vCnQkqhU1XKL8y8g6isHuZHSxhfUeyTED8B52QXvRsEyB87mBOtFAiKSPqGUfBv8r2bSo7xUm+0Z
vAVDpQR+SeIqtsaaOviuD3pOuCU13NISRGS81YSLyqb6bqfBbIlhXEJqQrXCvCSU+RXL4kDO4dnw
9x/qSfDpfBaR1cPfrykrYZGV4nntLmBhY1N2MCeIFx4Tb0D4Wy57uhdPucfJD+1TvQ6HRKkCCvL4
uvtjh3su+CoI5hDCafT2ch/fWqGIz3RgSDLe4+u5v87M2DiFDPYi0Sq6UT+3zgvlvdZe8wDvszj6
VO3idPnnBvtlFqV5wN+FeEU/d/5KxtqHnJ6zsPpUu4YKShM5FoiQN/zI/35FpXcmS0nOaQT6NnxP
e0BhtqXixDKMTw3Y99uroAWTIjnV8g98Ug62QwKD4vw8QF5MxiUOv7pUsRkORkFo6qen9weobwTg
I5Bx/OuwnVq27KP96dfOxC5BWnE/u/rY6Dl7IbojRwoHfuqzltGlS9W2PRnReCjW5o5gxMOLEwxo
Bxxg6X18ckRq5+H9h3tUcgCDd87LTZWteNxHthglK3ob4T/+IZyKSwiRPwflfsb8g1cBlMaW3End
vQ3I7nRynCZy2XZx5iFGob6bqMF2qPC1Lrc1tF4rL7OM2VawoKrnYDN8hl3PPMjUkFAP7CyvkgOh
UEadXYQOaadFnGsGTIO/tpoxOqG+EhtKVA9pPtBMMNfN3PcwpOh8L2Du5L/hU1yUwUy0SAQxsyRL
eIzSb7kEaslvYmcNJTcrrdyJkjN+7tta8E4yKW+DSWzLIElXM3kjD/etqj5Wg6YaLKEFhpQgwRJW
l9q1D4QUygbDoI+UWwbXNKHLBPo8mG477uFqQ26T8cCxTGoqTpWLXihG9fvAuNlHnsv6vwuPLQS9
YZNt9+GCNLpm6SxJrfzA52nLJdP4Tyiz43FL+cLSyLmuxZiFyO2bElwrQvaaBKAIDcSDJcCDeIDY
V2MyN3QrHPiKHK80Om5lAeskE94lvnn97SekHhk5T/xNUxHOSrpu/9lz+ukg45stTcfM6r0nDjZS
wkBFVI9y9TiVHooY3960J9eyquQ6WU6jF638QyQw9/4yzKKSdmu9abdyYdMQPMiXoWEcpetuirkc
2Aixh+r9YSKl2jSCCuoV3cfJnPh1P3BlhMzVzX8WGBBigYSNJ/E77sYoTcknatTphNJVQWPNmw0u
kGTCVFtWChXeMkTtLUEMX40kvyuk/1ffuq9RPDSwrONigi9ko2dHRTZcyP6AaPQjLHNqqiWVNckJ
MVDLDim3/pPBJ2QEBqLuHidMwNg7jZlWo7A7M8w9Tvb57nI72TMtJ/ZBmH/Q1mWO+WXboLVgsUK4
z5ICheYY7pO/i/ICD7tDpFq22Uqra/Z5u3qCnt3TNOYKRQW8gXyctBO4p1g1Or6waBQFigE0WeYS
MEpHOBz32V/rvNb8ZBKosz4n3Jm+sEriD7j4E4lsAKp8WIvoSDBTcgVLwqk0SdkNPI/TKYrTIo72
YxJ5TnbnUOnjoflHlpN2sD2OumC9rC2jHoZG21eHfoz8QkxIbbFzlKTREDukitlD9yR56qffWJGB
MmnpUSrqR+WZJWHG66AMJStcEhJYlg9GnxTBB7aIb+N84+USmKcdMbigXFMbQgNj1u2nZYXqAkQl
FqCyT9C1K4QiDeBpLpw8yLaOHiXa+XalGXzsFSeHBGZOl0sPnQ5cjr9DwyYP+MRgQYIba2aHQpHb
yZ9lPzu/t1XtXCwzkI9PcJCokfmlzy0sAt72Deoy8ce557M5Jf3Gmf+ZXHhUA5NxkzdILf1eMcMQ
Qus86zRwm3mWF0htDGeoZPqujf7nO5pG2MFkIfeAHMJXBw2q8WrKNYvHiITxBZ+2nbiis/8DOReT
rB6UlQZh1C3wYdZ294/OLYpUgCxbjWnD33zfepYaU2//cG1tLN8MnZ3Ry/+2joZRMp+B2pbheB4L
Ber5zRUgOZBSaFERDLs0m7pyRHo5Y6beKBSC5gPH3rLdDNcchwCDrqqrBrU/sYNRd7PvEFBmAOR6
zf3Rd1lts1j8mG/9EmlAnWTe7L38hHUz9vF6swdFLtFj6bInaIRVCxB1SQVNhNX6cRfdmaaJoiG7
2CeX7Xas0IjXqOfO8T+2mR1ftlCVIsGwDJc2gO7XUVLea0VmKsN+PiEvm+pW+dNj3PO4NlC9lcmT
/nkcmRYf+6EIF96U4BexwNoRRdAUQbH2VuXawosY1i02yM0vlnqkvm41k6vUc0+oA0VGZ2xpzHu4
7Nqd4bymvLJx+2v6JSKA5LBpZbkMdtvGi1hKYfbtpZFmX9clqA+eW3VTwqx6TdvKsVDCxIo6D23d
S7KOJab5cy4Tu5i7ABPYwFZeUSIwWKpcs0mFlHM84+sj0Ms/dywZBTCqb1h8+AJRguBcp+Da+gg+
xXAJxB7OeOH9mRU7xNxXhhdYUePZ+/g8yGCETMUOQ0RDxf1jtLCI0nueJk4miWhKcpFk8H9N5Rpl
ZQdKKo7LTvCMLqAll99Ry0FF/GeDNBfPu6gSVtk3OP9ADMoE4+6h5SWcJEp9Cyl5g2vDyRn6WTZy
pD8Ruo/ddUg5wm/6aG58NPvhUUYDIKcGRFqaT3ms63ayckZNRKzxwXQQwRs8Pcsjpb+gxn68wiXS
xpyBN9d5d53tkL28pmMXfNTAiAqPrP59oJJsjbmblJtOR2cZ6nD1vIZvjpCqnyFyo6/vk+edgI0b
qkUsYkADzpGdm+0qWgEStZcILWGUnTpWN7gagGApB1LEyF38iG1iXTczvJipxCgFWRlQVg4lPMf6
b5PQPZBmMosIxnKKoqi/6f6+YtrFrKP4YDknL2qVQ8s75/bjfe7N/uqr+xDTMybhpKR6bWaF8KIe
yYZtEmKEkmgxoZfYOX3ReujdXvK8jfSN++O7BQXV6KmIBI5GxqTNqSS26jmRtlU+5V/ZQnvfl9sl
RFHmfzXTX76m7K0fMVwV4spFnUwzJpMp5J/r0AjnfA3ZS+JbSoH4bVwjm4Gr49FagdE0RDpNahi+
FQzlDLz1DgLPlIcbfXgLWbC3Qm2D9bcNUyiR2vNbGG1SJhz8mPFY7ooAutxx4k9PXoZTpOR9wpZL
iBKqBvwijuw8LFaxM+bPAT16cFlrDL0VNcJYx6zZ3DGhGZldYnpdUIYvDdq1EVNkJ9OlmBzXsFAq
wFPYLpnxbmE+zzKT2vx6EFNPPVfyO5CzNVRzpWT1np6iwvms/ZPK1R2L61rxJJnjkehYR9gQV9Nn
RIHpt3eiw8skx1YKbe7CRgiTVP2eDbevzCM1Y7qdcl/8ysoKG69pTNEJHbYnjiZARc6Yc7d7E95E
4lreBxUGIFa1DeYtKQxMZYpLVdakqaAlcBgDBdWhRvQdQRja4F6xdNHNTiiZtFfmYesp7+WlXK4N
XfTe11phuV5i9KKforZL/N1cqwkI73lEpJWINrczCKrKvF9BbUfixCyeR024dzLj0W3V3QBxSaeG
cZlHyfeHSv2Edyc/fmAZz7Bfe3bzW8aua5WvePGqXi78h4ULbSOZF96uqw+A9zAY+BlAJhzJVN6+
zuVZ3/XJLWxyiE33SncUfqxa4IsE8690TyhPKTl8/83p/w4RmuVkUIsN/wO5KCtDQ9NpnXiE0dCk
NdLO8dxVP84MMRwx2SrQm9UtDFVQPZCHOOK3AK3je96qIFIxFwJUyDd5qG9vyTk7MW3ccog+gz5j
wQiX2Ym2AxlDuZAkdHMoswUku/2HtkzIffKqofXL5TjUczxY43hNnyIQ/KTaD1NYR4Rl10aKNEgk
1z2BAxZcOz6xerpzXLIuFbywlbSNVcUDnDI6QZHyn8ksmnWHMjc/cOMaqpobDeo38WTipEIzZ3eh
K3JBNBxxN1YIcDToleFju4s5hurQ6m0uy7Q5n9As8io2j2q6L4utlgbasgp3fvXhiNY0rLJLyINr
N+qO76MDz29cf8edSAQYtMT9dJVjp6iufFH/P8TelIW6xFm51Szc1598yvtL8f1LqJMGmDEJZf1s
L5UQ7vBFfoDtqc3dZh06Y/+vv2dttuYwzFeB3BZXGXE2Cn+EZo5HyFEAFyDLchDbjim0602qGHPA
hw3h9xCIiC7Ts1BEsWYecPaPaD6u2XJrsj7fwxAGKLA/XynUoaz1DSy+pMxWiBLxdFEOflRF/p7B
4SYBs3yg8A8QYqqxPNf/bloPDe38Qn6yVVQ+YRU3ksexEVJ5+100flCAM1KXk28ZeEv9D4txZ40F
alKOxBvRN99rIFmWLD1DYh7SuSpu0CpOHea0YM3vu1gBOybxH0V6yQyLUN9JNIoXNDqCxwpFM847
RWdlZini8B+S1O6m1tq+F3VCafc/GHO+wOP1to7d1ilwo0quTVgOiLNlW67cUxmlZKOKl6eBxyNV
iN3o5yepx4jmCjv1ysQRBb2ztxcYI8mCMJF6U6oNvldfv+ZRo9Xw5PXuOFWbsfZXGOF3AGDZrlyQ
rvRqQiHd0FnOXfeh6v7d8pRGhxIXpypoRVd0RV91Bj2+5aBFaXMjRfQ/19JTGRDkFQRG9ALsSVux
hbAyBaLxjkHPYIxiSTaS2qfdQiT46fznduzxCtaXKZSG4+rO8uXV4IywXf8AIdJY6p1vUiTugr49
dTBIhu0TAfcmcfi5HK6TjJAEkT7x3lYkSFqwPLsQP0IAaE0PhzGIsE73HUG9Npqhvx1INrvnaThF
bVhhq84GEsqcuVNsm9IAZhtg7qADaUA4ZR5gmvtEkP50D3swZ6KDLUfC7gHiNEIQ593VGrhqgA8i
mmCUyB14zl63N1eUObPk/uPbRWcGaW/khGb9hLjNT3HzPfJjoUFB1jR+NLHyP2nVhqxu78oZFop6
qun0I+lFNJeEQjROeX28NkgiYQU4VEqtEh8zd5QYZNr6ICQ4z+2NSI5ttzRej2SM0UfjPRG+oiMY
TwkZbk5zbpgcqaD3C0uMk5GNweW8RAjxPytjMjMcSZhsH3EEqqAATrKVPFaD+8+N5Ba/OY5Ug2Ud
rlmzSumd02b2+EBAG79wnfFTXg49m7l8KGTS9m1oUx5JBJEioHHKlpm+QCnaho7semfjXvp/ejIg
W4iUlf3vBLJqfSpz52JerL/U3Sa2OrITCIHoURSWYFWBdr907yC0yVPCHEANaE3V53fuCh7Kq1ze
rb6n4Ah0a2orwWXKWZyB2rn0zGeq6W7n9WMrmwRISe5O27qmkSsgo195vsRVbwMc5sa2I31hOHA6
4tuzNrUPOKkvHG1kcWmKvgxoIHSpmFEo5chALdw94QwU0xUXZplaMTqvdLNEXS0ISAecy34ziGPE
oGuSwvwuR5StonM92g8UIwm5gbwIehqsxcfO/IWs+crdNZnIebCtLvspJv0clLEoESmlYWlSkgOo
H4tSrk8KCrsipvVYucoZ/3VkWUfKQkBN8Q0QTV4o8JSOW4OC38kpzvKu20xnSnDwIZ9uO4p1AkWk
x8M5DYq6yZnH2z8Dnr8WsoFei16QjQOMCfl0ZIK+u1WZWq3/R42SQvN3swv02YeJcGB+g/b2eslC
69Ht9x0hnsT1O+zs8hV/8nptuw1LCOYEBhihoWvcIuPf1ZL+YmYu00wu5Eg/nFRYlnU8bB6G0EK8
JW41CFrwudk4r/hUcJzqLrn0VHKCyHFeecTSSfhR+I6Tl+041JBc5JFiJeRGyInPllgmKG1xDH+9
Nhhh1KjcUd6xxBi4/3rw/2Ir+SUNRE6Pj3y63gh06uJ1I7jFS5TrNgaGU0hYcKNkudlhtkRkb8+i
tMI23scv0LxuVM3Q7pvnAuCcpjPuFfoOPh3aRB9ab1x4jSvx6l5xxUyST2xJJmuXGQpBgw/DtFg9
b4wAIlU1GFBE3nwLnXRK6hOY+u4DlZcyP74CMj7oornZ4tA3ddnaZZXFZPBMDGPKgWiHrk/43l5H
JTioHt1pRNC2ayQsoFkMm7k59N6773zQqZQfmi/0Yg1IRjnF5e7fsZmMYroPp3n5m+j+B8EdtXCv
kiYOzwtdhi2oTX1wAqxtUfgbzZaf3T1GWRlG8WabPFXs5ZUHCkeUVcA1hglK7zRVkQTB4ZdWAUTW
hPhsH9tKVWOmIDnP6PvWM2GYnhDKKl3xCD6t2wWpYsLiv7eP79PratljpeJuCT5FMPTBWxtB9EQA
TulVdrQbDUKLmlRcIpoYE9YVr38+GyDTzLxXewAFa/U+NQw7jCZAw0TBQJgo4F2Qz1tRA17pEKOr
S9CdpLqYHqXz7nfxH+hPz/TcMvsAc7dcEK+k7hCg/c9jX58vcwJumQLBvF9SaezvKM1y5lM9WyXx
6W0j61FQKZRptgp+zlJFVbBaNWEoNlKETXfzLxF79qAz9MQSgZG0e+U27gB5O/mvmTeFJ1nNEQss
3DY0NjKbpl6C5oNqtQBv7wvUMD51vtPHsAwLwpUBfDk9+w9bU4YknUgttyKZkp/3XBWUJI8MBhpW
+LJ7bx1009/ksY7i7wcvglBFjuX3sjXd/2woVCxiLQ5CplHHvcaIlxXdhV8orkcA2dX32QVqZatD
49pfje1ER/T+bt//GQ+yPz8PG+CyPineZEYf954vjCsueXkTA9P2caz3fJgBXnK9SCNAMshe/aIV
Patyl0wWaC4Itxg0mJFPeNuoRCE/rSFrsDG3cvw1N0tykiT1Iv19sWTGebSmMSCUgle9jQDMH8mx
8npVhY3suN3ZyLlqu3BrFEFq85vG9z5U2Kok9lew277p8cFOs71p+Rr9icKz63NWHYDw97RJOp4c
K/17LyXx9/TI7X2LRcB6JUVcU4ruH2Q4KgkJWdDnDZZf/Ws1IVXNDvLaQNumVly721914M9nii1B
/CtgXb3DW+HnlU0j37y1Vb7WaJQoXjY4ngtBapdY8uDzoEi/SZA4XdCOKHjNZm3LjE+2N2y4worD
eA6oKrd1HfR4uNXiBZ0qTo5OZrgevdNY/Pb1DlRqYkSPnQ3n+SBTvB4tC4kV0n2QiASV9xCUeL+K
Q+B3gLqTed+nOB4QkgFfrqV/QNjzBrVPNUx8oIBaFFzao4wyJQw5IuOdlh/FW9dMSOXKsw8JF28p
FTjnCSHmXsu7MYQ0KqsDcvyQg1zBPDBBbmD8cyEaRjHvYF1fytReh2tOxQmKjB8KwXHv6Cv8vrH9
HGfU7QTBC6QKncL7SDv5CdQx+yhvEGJQEk5EGkKqkmfL66m2HbwrqdmKIG52zL5PzDLLPRbA2+YV
LWAvdP4GpW1g7QJRGF6opEEAphTLyiqoQj4IEqa6yBzteKfuFlOyphOlzSPRZ2UxQbjFCT+j3I79
k1USuQ0YkuFUDPQvFpLemi6Vf4tNtWODo1CrVPhweqR1nP3XW+2952hin/h8rLyukVXHiO/V7g7Z
L1VtuTDWamHBJi+4rpKNA/d/9yLIUi246vOOTIeQTy682lCGnYVeC+Ac75t26Wq/MiU2kEUxSNOb
VgXFXiZxC0qKQ6nMPk1JGpMb1Cf4ekfVqlY6uPl3YG6lg80phgjGquL91gN/vHsGwk/sqKHRU6FF
E+53GufjobSOG63JQVkb+BL4U2Cb50c764hGYQddzyh+fz6oa+AssaPcfhRs/9uZfSCj00EWGT5j
HwldLKbA8LM/yCkBcQ3+bIc6qhB0mDjIvh8JN2FoeS6szavx1L8TVa57/u0Mn9ZbPsO6jg0FhO9S
6gCGRcAi9zs7/DwTcljoR0lyJW//JYApe0ZLGNPPGnLoVH6z7bg31+7Is3eXGx9j7D3ea/kemmJ1
YEVk2MChw4x1TSF7GCWki+n7eagnTRXmE2MXibFm6PF8EPDxhSRGHyMjiMR21w8bchkKvIo6CH1h
7+UW8LB8jf8DN59NPGUDdRsT3zx5KtoqLXMnybKBzV+CZjTnZrHKTDzY3GiRiQeiAp6E0icF/oWW
eAIlRMAiR4n3btr+s4Bw98bEbVh+PMzMBj7JgtedzsQx7MDmTiWcdFbl+TkgMGMDDsplZTSv6Yls
jN95oqWJjmlS5F6wEXCKSzG9Unt6HMo7+hFR4xApcGjhNKKmd0G11xDl2cmtA9AUlyJdM5BzgLvN
9AmlUipa7qCdkjiJ5nT6i2HdNn1aJxhuQJdqQggofULC9IyWkXK2H3QJQXFECF24DNtUT2jFc+tT
0gIF6lXgx2TO1tetPPkkvREdu5DbZncVkG5jXI2yrQlvf1H5MH/2IK1TLPTva90GQoBJXkxjDHZi
BYgMMIfpUNwAqUC3/CPRlHXzR+1ITFDzJIW9zMSrHpak/pRpaegSOU6CjAO/6gsEkf8XtGUXgE7n
BoroXQntfhTchVGh8Aod+l1JtYDXIMqNYZ2Y0vhIt7otIsPT86gVRdBEgngbHpK+oKiQZxi/ZjfD
Pb6KYT29KJMJHQ2uaJSz4MbaPyzIs192OibVcOMhI9R2stInJS9BZ+KfP0nMuJoWxI/jMAYFeGj7
X7ljl9R1zPGk8n/6RrhKS67Ri+pZ5+G/qUe3ki0T9FL218F2+KBTaUmJa8Hbq/MA3SNSaypkw/p5
00mdXfVInAv8y8TfRiJYTfJQJOmnRB4CY3B5H+JkKMhLrrUX4kK3gIleyotV7qhZl54Tz/w7dWTB
53XXl4owy75RgNiuvQh6Dy/FuzS0404Z47S+mV5k55OCYLxY4XFyvjgIpAIwyJ/YWuZ5D3grWMht
eND7XeDUx18c+BFhtBCFDCZ8rc/EbkxpvLeFxH7JbSiQ2erRnoDvzq5hYaPtkEmAXWj3i/Pmugh4
vjj5OJviuHyw8c09dgzd1PrafVOXtmSEM8Q+iNXebBR7ZR/rEbZFiCs6HMdYY8AK4iOdc8CbzgPG
IsEiRUl2Vb/XxI44FPScSjJ0yE2WPK8ue4dZ4AWY09It84KAuMvxz0rha98qsB/MHjW5cHIdjsGI
duS72fGVRfkn+cPWOthDo68h0kbNUl6ofhSlL+SJxr2wsQ2Cg6hu8GSrmE1cSz0Sjg8QDRDSNkeb
aXeEZXY8CoWEUBv43HzhN8QQZyHyW1J6l3Z0t4Q8rxdsMHwe+eXU5v+qDUT0zm8Sxj1ngi/5MccF
OWa1YRs+cqei5htxR2JlLFBO0x/JfKVkTC5bgYszGv8amJXXATmwQdSst8ItoQSFuX1aij6cF0ww
tKP2JNRzBntospymLWtzCv4HR/d1n9/HxSiamStCwQzM0yWsWxtBgnUxpRjknfc2pLJNKbg13zeq
FO3SE2d9Q1td/QrXvhyghCdfzWfBHti2FWSt3pkM5eLDlM9qAMW3aiWE7w970qmQfjf2vo8YPd6t
6DWld/9ja3zobeZz2RSI1Z9joDl9iQoFBsYiqq3rDIrBZIRQFYfuyLg8dW8PiKoydm0BRFeJAnIJ
ire7HVoIthGzpg8q5ByDfbc0LfbGVVHyPJmF02D7JaG+wa9USx/B+vJOLUqXDqioXvO4pYYicURW
hRQMmwgb4ChD7WVm8PEG3Dcj6Xh5wgsyZ+XfGQH+2e69FfDpXl+TFuYInNP7fv6O3yPp0nEBBOC1
/vrdReGysS0brdZ9xLikdZxWuS3jPjnUWD9W17rBExcXMG5sQnzEjBzBeE5P9vaJauLHRZq/xWq3
BF2Rzt+9gtYQkcyWLyT8fkZnIbqQx5NhwLcc8ZDb79U87lmklc7Pr0s8psa+UCBkvQaAvDeR3e09
K313cmQWS+qJZVbrFcBmXcK8cF6wKZ5HEMGklSPVkQUe1LVCePyHykQI47J87bKOdAL93aEUUGKr
TAXjtpt1sUmxWl9X9v46lMw9CDPnEV+XpiH1A0xylr2Su3FWL7dhJWG7/FgGpwAt4Ycmrvwcz31b
katUTxg5DR0YtjyBqeOf63C2R1hz61qOeW1qXEHUmrO4CeZUlzDmUGiC6ItwdHbrj8TEdh80WMy/
zPYnppt0+jMoVSswXR2dnSMZwvXcj5ZDZHsCpHENebOEKUc50J0jsfpbtzcNHktzZEM7kl/9V5Eg
+fxt9Z6kQMn8EMYCWTlCaNwXYAxxrFcs74F6YfR2o0cE9Sz2urLLNflER7TKGZ4wRnYY1zs0qwC4
KZpv7WPAor0g4XIeVb53L79suB8v28KYHIVz/hRke7cV6k/zF3wr+FV+3wK7nS7r/jPFSW+nTHyQ
Wxn2EZiBlctWXdDliJnwhi0ijYMrnncTeKJny9cxDCE7BztBcNX2UfaX3dJGgQjIwkwKyWQyQNjA
wY9qprIaFY+kOeNHWBqB7G0xnZD0CS1ekWyiL2fdC7Mwm/BU3hTTGs32IEwUvBmwNipx7xkhhEkD
hVXIgJdi3XiUFEb86hkhCTQK6Frxhyw1Qbxp5X88DmuAYXgQMpXAwG96DadJL496kYVvkDHCbrFD
1i6Dj+4u8DC1+GsNExyk51VACf0vumNrN4fSYusk7Pj9o0rc7wBt5fUxlNI2v6z3mCs9aIOE+w5Y
eXWpmnYtacb2XICvE69F9nmxUuXU+QdOZrUtdNssGoDioLLY11ulXj47GRkQVFlNhuJYAiSHUGUv
GO5Joh+pp2dRyBiHY0ZG14Ok/J3XKj8Ir5dtPeSg6crtra2a6BHrslhHwHkSY3eCqm0h2F0XPEs8
/O1Aqf+crBc/59plsJIgybD6GYb7bnIC0yQsTDZIXYGkfOyzNPV+MV1PYNsEMRgYHhbHbjkS1bYD
QnNJbMFm1qgMP1fklBrdraRCgy0EErfyAICyCXLfcOO3vaziKNKIaKoOtz/ThP1NjNIFIcBJ583i
bgWYVgnl+4jimIylQ9PrGsYk7dVL9jIjsuJ5jsQiZTaZCBKS/nh2+WslHNqOfVlhrURLzU9dangj
sGSPYvX/5MlZyvx5YNey5ydtuDuvWoPxedLBxJTtIgjC9zdthEWgXLDRGPQ5LMANtHSAFha/k8Uc
lorLvus/pHiC+ndOW2ZVf4qt4Z0UXtboqVvZICC9pdQ112ELiw7Iueu7UDB8j8QUY2aUWkjM/AVS
Snf1UZM2Q+MlFK4yTID7WsqXjA1WramHUIOUUZAhUYla5zYY/Jbto9YAtd/d7peDlV/gBpPqhEp7
LRkVKqcyUK/i+BCNsILOGyYOi1YpBUdCFWUiXGYhCpzBaqp9kBJBu9E223L/BauOJzWKTDQYj9Nm
Gmjd4IdSZ0nk0aby/yfESsaNK3Si+S1WDDNbO+DCdD6lgwuTStgM5tl6UZNiykaOwdimbQqm2e36
Og+90XGk8aTGi/hggXQzOXZrnunbzBG6oZq/aoZnOP00GooiCfzIEfTKgmeeN4s0quowQiIKDvwm
/J2qNfZN3TIQG5isW19zvnZA0Zge2YyvIC9Fxmh7Xyb4X/DxZa0aCUsygIoXcuTZhYVni8XTncEo
TzIAHMlcPJehF3ScxvTD/km3b6qDQRHUEBT7fb55Xy3zvO63TalTvF9McVy+EskMRCBvH7VCksKw
0kVjB99YcWbWr/Dm+8U+wfJN5Go+PHCd/YTwL+mo0VxM59OxpwHuFHO/PR2W4O8AQCkwvIjc0Uf6
UBfN0a4hTiGwQBbgcT42aLjkkWe3cbbDvWb8R8+CUSMbmDA0/pUaVQMffitisEnGb5B9Gg3KtnaU
Bv+IE81AGzikH/3fIql6j8nIwuEneL69ya41xLtVN4BfppI1//fejILsS0st1nhZWA0oxeNezPGW
+kT7nJlBEHn4+XCnGPwdsXrxO0RiSokGeA4VIeic12Y7nWe2+9f1rPDEHotZJeZ6t/vQwH9UcLzz
kS/7Yn3uaalvYwiO5EFCHSeGKPZ7ucEFfBnFvKXkKPF++Nz1Qzt5yPn7GuI+IoUlw2UQAqFxtTm0
6GVnt6MXRI8t1Da+YZzCIrjR5cASrpQfMO5PRnr9Tk2CTmSrfIWmKnLy/mH/ebfzTic+ZIeLxt4v
ZYlghk/a9dXWZudOFVuguU4nR4gt+IXq4bH+PhOPJkiw/OkkDyjjdc3sP9z6O1XqBhow0+wwz61v
3a6jtt0Er2NQiBVGCUXQtL2OaLfjjdKRorPaoiBZneGZJvOORm2ADlrKBd0uS9OdGl2U/FCvWaRN
BLPbB7eb6GFKZB69Ar8EkTmwti3fKy6vTjf5eXsOxsQh76AzuH4p3+B/kYqBjZ7NLHaD2Y4GP/cj
5lzX84eriy8KQ9GPCd7PJAqVoE3VhdpVnfEPi72KMhn4074doiB5qVQM0cF0UG8SiRsFs3Q0+Wus
oApSLftMnD7w2s4mb41d6gk/XpKTtzVXLuo5nzNDFuS4bcZSeKIfZca42vFsEGCaEm2sZnmMEAbR
OSW0vOlDyEoJXNut4hZ7FP8WAyVXAMyjsiRqRIsWGoUbuNjDJdKOqVu4HpX5msVXazvzm9/AEGiY
ELE3X8I3bJkb/trKynkjwBwYNG5i+Y5y6mOE61aqu77JkXvS2sRDddMQrMSpw+2bKaho/ewC/xFq
CCG7GpxpaBkYFtv4hj41yM4SY3MjW32axrTepBjn/c+R7EcdyuxieZ4rFzI4MAM/AymFs6iFTbrS
uZeFAleKOzh/R5wVZohtX+ta56zZoIWEyUTep+SNQUmu50rbOFBiKm+2Td/6V75NdfMtnPIMPt0T
N+8icinuuJfpZmSt6kq6JsNMxS1Squvlp58GdBQzgIVJDqmAQlL5OXNFIY96fuoYF0TBmCZjSsdu
bL3HHQwlUB9psv66pdqHvt6oNeqPpPVvDVJb+rau+JfQc8ZQt4XzGo59qYVVNy+iJVrSRU/rUiSA
kQMgh03gRtyxGm+yFtdSKDeE/Oks5gYLkXrgxXzFGYbP6M+6Ugea8Q8iUQ6UAfcLQ8rryRJ87SS2
ly8De5kgyAVvIMSSJy4k/q8VFwyl1cDMFEJ0ovqbKdciHeXpmy1lgHVHW0er8UQpdiopPc0BDsAq
BFTLba3Zd0jYWQpM6H0YJADXDBgJyImHi/6gKPpDJeSd25HVeT7m2EdGs6utudIsgwaUmEXfY2Tk
GvGyx38B7Q4sdpbWFJT+CxptZlKfd7jypKQrXcQgEcHqIyFJI/I3pB7noe3NLqGiKEnRCMje88Ab
zM6vuduhmYyI5i16BI146An6egsPl0uDIMClGLCzaI6qsC5me2MQV/VWklxRPKe2WrNoUuNE5nM2
SA8LKfy64NKzPywdWCRoemeAvGyQpwlD6W3hGE/jpaowsKD3UsP/eslVnT3p/FB3PHnxDUoZSRxb
hKp3/2C6xcau96lQf6XChdWQ0HCSM3/x74PnAAjTZvwCNKWmqBgTX6WJg5drWEQWSd/wSUbE68N4
r055XLgbTUjLMAJsTlCWB03iUWx7WhLtpdifR0TNsNi/1BxueIyljDCzBUAK8Fkf6hEKwBY91dmx
W6jNH7uKsdsQniZqkQenIZY3vY7khQnY+Ftu6UVqIC0Vh3HyCuWDY3DzyTFG4KY4ut9wqSZNgn2b
CPdiBzEVnSvo2W7nyeLBYMgDpCh7C7JI6jKposNo08OCNS4B16CHZIMO24TGudXA3D8T/vpAIZ3Q
JSrUYt9qd/DAV+diW6sBqLOJB6XDTT/reiHV8NUt5xBV8TnTxzIbVwJKwgic7IAXbQeTKutnKxpH
u3C0sllm4bJCe/u50Pc8QDAcSl2sHd1uLSVlQfwNyHOYBrhHTKxyT/O4ILn2rJUYBknZUU+lnOTs
PmVqiD3KrKSuRf982t7dLoNu7faiTT95LIYRdSGaTqTDqI/JEMOPSCRQQ4zTyjq0TsQkuqO+w/9+
7l7SA7lUIU3c9VpA8UtD0TtQaTpuIQijwbtT6oE4oL/xZ0K3l/yMK+mLVqvFNaIHzc1hHV7VNsQv
lBKk/VfErEGdvw+sBfrnVkWo5ShrohVREc4NDdzI7UKDG416rONUh4L3p695vKDJ7ZRQYznOL4zd
A5aCOzW/QFfuzrU5jRXEnUVB8JSCQ8agFBrSb9c+EFbVEAB2OLBERyKut99bglKAEqUi9yRetOnl
RaM/g/Kt/zLFrADFlL6k+yjebFI4/NSxF2o3l91qlUsW8za3s3sKa2gF7gC+qRLMy0HgwAP5qg8c
BUe69i2jZ8k2uhdmS2f8/actmgIJVNcrVlNBzUFRk/gj3gZSDZIeUdUYGDzGVTVxJqPPLZuJLEeI
1qPBTVqWnNBVjgl4vFz5zX5VTixkGKm85Hhpznz8D9+ehLC8v/chIbdEOxhpZKs1xM5xU47k6/2L
1nX2r003leGRCec4Ke2kkG5atOyVztb9X/Zqgkl/BgmN+pPXFzILMX9QyqxyEwfQe3zlrWphrpyS
f3xjzDodTixMl8H01KjSdzAebDkdXSGS9bypqU05qR0QZAf91ctpKN08tgNJ/vE0XrMiGyBjvVqz
qoeGZ0u9miB5aRCc7Qw0cO2ZerFdEX/CMHul2H1QO9FZyWZKlnZy9SMOtL9hVhCNmzoK6lGMnOUD
pduoqhHd1ZjkLCkT3h3cy5aAYI2iLTo+2TbqQKz+dQAIicX29wRWCmDf9rFS5GPt+ZfTSsD6J07f
27fU7Zm55sV/wogtSBTNBOCr9g2UJKgy9brWZcxEOpNXHblvuJo9fttT40frKTHh5jaKmVyQo7zY
d91tNK/+MyW1rfNVlNxa5y3EPscLk4itfGJ+A+64D7Xg87CNZVpJY6xC32Gx46oIVKEVE6HyhUcU
0TL6X+8cMNwm/nTQxmaPzg+Qp8IaMGCs/3NAouGayUqZf5EPUT4iQQOiS0G7OWJ5LDpVHjjO01ES
J2Yx7HDRs2IX5J/MJv/lFJ6/EeYJ1iHKkJiDGiWSLj5IoQHpug/uHQVDO3+1hp1jwAViUFC7TTRA
GdpZHr6BJfrq+w9bVstDpmR3A4Klt7ceIg9r6MnIWbM9cACioxujdYd8Tyxm7rVb5i9JhbjQBAYd
bNP+ykce8sRyWBCiilxR7r0FjIBVAtqTwEXSuy2DnSBKUAWIV9hz7LN/pkvbqer0vQ/ffcMJe/wi
aJn9Z2uikbdtaNSeZJbRMhh4/Ko5jMbA4XxKIGf0diW0/NkDd/xiqgZhhnMKOouQ/jw7RlDcTXvf
f+xW+E6O7F+2hjZ38OKNg3hu76WbfGow7mrzTQVG2PNBtKAe7dCrWEwso8tqprMeRfvZRm5W7QgF
u3om3j8qJqdUytDIgTFkmFV7qjh90B8czez6eeI4OBi3QdUWtY9hiKopY/spw0rMsKR0QvYk3UZo
ceWBTMqHJ2Op0u49/B/2xbB8aNNonC9Ds5NobqPhR0V4y9NupPDfXAOmG253sP5SI6C82V5yEn/r
ZUb7aG/r2O5Z0uDD+NptcZX+alKXB/D6HNySRXXFyF9MHxTuHgV8Gi+JOzxZiYVZJ4qI31Zc0ayF
DLcL2UqtZDr62BZBvOCs67pS4c6UnBpc07C0luL5Jd927hs+5pBFhWmdcQRim8QRMO+E1iALk2BP
wqgwaafz8rLn1U8aJMG0Ww+ODWJgTRS5cREfKbS3w6i/FOzEsGQhTjYmyVSVuFrGqGTJ4em60AHn
srqYqB27Q4ZatJZtUk4Vm36TNBzxVhRR/uFxxShsi6zqDIAHnN8Lg92FCyIIWb23gNhMrpKNB6oe
roplaEZDMBXhdEEjZX62yFGpOK+rsqweo7KL0d5Og1MzP7AS6o1xIa41ERopx4VldWHPpBKg1+xg
xAiv+Y6b8Ek1P6OSSmsQWl5UKtuXCHta7fh1x1DW6ykN4hnb4bJHs2LbIkalLKr8xqRXftgSUSYe
5Pujm8aMhn9aHe7THLdzAUU3Z7ypiVLgqvO5BSFRPsFyMmof5AiZCPZcE5vICuc8v0wfoNdwzQln
BUwlElfTvvL51uhQZjZcEjP/UwexpS1mEnWrtvvlkMs8XogCK2zWmlntbVv5942+vnpVCL1Z3A0j
8NLsHhq7mQWHe1epVTnj/I93buC/ofgeNxoDKM6vT3GXme9z8N7+SOxY0XlNWC7RJ1PD5jfGMu9G
wJGnL71rlgbMi/UDb3OlZThE3Ka5AHs3mlktxuMw+4p+gW1A0lxOjapvBfXAFSgXeA31hOy0PFgG
Algt4OtJD+YTdXdZnT/tuZS6Tc5kFJF0URRJ8TacLKByUP4k62yewPlus7JI6qlUdVyUvZyhSm1I
d6jsoFmstHeiLQU72Pp3IwAAYCUKdNte8CE9erzOceTIzuAT/SzXiz/YSs0zaxMl581rirVU5M6+
/RSJQpyap2+wsC9Xshqe2kKmtO6pYMJu0yBNEVVH6BJYhBkcxDRp7BPkiN1eEY/NOKf9MFI9xQat
UwS8rc3thBM73FnphbhPBfQqMENEnevYChWNNMyBppSYpZYg70VCOoNjZg+UP0rpXlwA1gvLCIum
TGxKUTRKEvnBxayiFWBgYc9uYfqfrjOgxU5c49DcYx50Q5ECD88bvMBdydJTE/YwHRwBa8CQcKCB
9Zxzg5rYnw12aUV+g0uZO7056GIWXEtxi5+Zo/VxveyhERDyBSPAdHPqoyOFm8iSJLnHU3mVNOpc
DAyfvbpnZ071MlYz7vh2uc55saYw2tEI0GnNYCQPfkcoL/O1mIJs6jUlAkGl+Xlh+g1rjOagdfrP
4JnhH+Elx5KmC4d/TsbReFDS2fMvtTTD9Rdn9llxduoR5vRVK5ST6v5YTfmbhTIgk8sFA5FwUPGD
Ded4qMYNfmyBHxEH6uu5jEN9Oj6HuQGgyQ/H24fki8TxOM3gOTWqv2aFtXaF5/bb0x+eVbB7ZDxp
TSuOh2VgtSHPhriqyEQkM2ttfybhU+MfS6PK3Gq8fE2DVV7dq+ZetZ85YMVEfY9zlVBBENi8s7l2
BTP09Jsgu7q2Ax+g8a7d3Wz+9BgNSYEGvDcwv5O01oJmP2z1MmtehJfXjSx3+VFOE9JOECdHZZr1
fF2cROl8oKYucM8WPLzdtKB6jtf17UJmRko0st7QfoliFdlCEnhP06Lu9VSeUKY/gZcFbydlNYtL
wDUF/K8vbOf/2VY0gNk3gajv4BDJl7R9tfR5OkOI4YlVuX1vzneOIOX/MsIf66xjDd5jcN/vXtIH
hHKNxwzoT1vTPdvXKVjrDM1Mo78WqZHxqxF3xwXBCYNtez2C6D4yU+j0Gew/aG1tjRMcLtDBtZVv
QEJc3wkvgPDR+LCJY74nEXgnSlY8qqnB1duk3v8x5g2gqRXioCHaHD2yCut/8buc1g5H7Tp0sjac
+GreX1LLfwcUjq7ctg7QqZN2j2mZ/leB43q6gKFzeRHUrQV+umHC2ECcB+tVgfv8tCWEPoVHBu37
md4lgEskFGB9JcNHEAjuc4spMjm9DWblPx/6x4SyI/KyuGwFSisMO2QuhPXzqQZ8hcAywunWrDUM
wgfMog+AvbsgpJhF+6tx2JJiUcBRrdus5fGMcSnsuvvKr05l9kYUzCr/vAdakuDIegEYz5Dxnp1+
yAyOj9zfv1YxrmL6offnkPaYEoH4H6A8SasOKABY37Jqru0FDrURQInlMVIQLJFcblyPFLPByr23
eY3x2ZaZ0JVk//KyCMNWzNYZB7ZYk0n9WAbfdPBRXRQvYLTca0kfvKY5wYex6alD3NUkfnnk2fnV
0WA7JRKPhSrm7yFwqQhWi2/hqGg2lAi7M48r04k8wnD35JAdGbTjnhycNZDBEOQp76N9d8vXd909
8yVI1k4yCP0cdM7oYTp6s0xEYeWxq0sgZTaP1nSHwJC8adecK1GM1ERxsMCH7o1iSWU93IJdJJhc
Q5h1LKmPNv5M0ruovyGHxg7I7PFigTbxVOGN1fwhkWw2p4yFa9JDYFSFQv5h05FEdYjd6zL5jSca
9EIEYu0Pj2tjSftIIgjmfhcDGjuBXI0I7lqa723/AB8669R/nQuMYAyzxYd44J3yC6yflZ/kKhNx
g5OywNCPqs1U8/xT3AFYKXLXRF6jLYrpOcXAJFvPrYgIZy7ISQ3tKp8E33roKsVaYhqww0hCOTTK
e8XQfDKx7WkNk55H4jO82PW1xxBLQP0ZeQY5Ymt2A1792lJH2EAbEGOQTzASdNRZdqvStdPAaguD
D958FfsIUmghncH8T1gFy4ORaCTk7/Cn4tnbJb/r4okCxDI/xJu/Nr0zClosfH3carFyFqUtBQ9m
PdwG1jWuzoM8WlwgKHtpnkGnYlQE2rZMbQQtQs3zOhZiqWuHFFasUaioEY9LfkFKcjILnRv7huTX
vvQhaDEzQvujDJwg56JhQOse1IPx4QXkpDVtRz3NKye/c+//jQaHm+tgBxFes4jtS3k2RbMOc93q
cEM17Wm2NDVAHiG+zr74XFuX/gbQaM2LRZEP8EJO9+Xf59LILKkHf6xuzNqnfyfaVTtLEVSnj7Ep
1JbQSegdcPD18sumZnVHfq1HhsxqutDpC5tahHRh3sqiZ2rIREfpLL3cp3NfYHAjulzE4MXog3lZ
/tnaA+GTkztnXn/fsuoRBAWi/ACKts9+np3BOIOYM7DVa5xTsE1fesIzxoTCIkjsBZeACa/IaUMq
hdM7cJvhVQzjDQorjdSHM37HCH2E19KsA+6185LSl/b7TP85PoW+ByMdIcjNiK0kD8CYhkCd6QSI
cskFrVTVAOtL6w8TBvSEI05T5fjUhpMGThUiq2Oj0UOfD2IUiOkdktCc/9rZnlZ+URZhP7qEas5m
qDjtgO2ygVR5KIW1QXrvkjbr2VFxrnntN6f1mOqR/fR05b53aSfJ33/fY3lNPWu2ifhyKqXiVvVG
g1o7Ete2a5LiywLTPYGEm/QnqE4VHfA5jjCJsecw0udjcCJd9ENQf/0OU8HpqcqR6CWBMm1TX4eb
gt8NlIYvs0/QAIcGbAXb3PdzX5F4G2NKZWxrrGY/dHCAw1CGBJywBRLJUnHr7Ukv2NIPYRhkjonk
4BomqKr/Xl14pvHI0nOhLWcPqqKNDrD47x1Nfpenem/p+Wfp9wq2A0wyZyEofqR09kEjerbBcv24
+e/Y6oG8VKEi8Rog+uQN/A5SVA4m1HlFLYZAyzXv3f2werIy0IgsmwhuylNlkKoBg+cvaGLPtPne
2A4lGkrcn7h6uRN4ZA4PkGxou+28S90rUQmOsl/V+yaSUGoqMqtdxZn0DuxbG+aRLgnTGN67JAdD
HslmGN6eVgqgLYNO0WTSKDBmu94HU/BZo9GhWiM95sY6xA6VTnpCoHH4xx7qRY4bMC1ZlpvItvXS
46jNPB9EFTSttLh9GIOfgmKfi5neGKkDGTjzFSP3Mir7sjpA1p96z+5yt8Dm3vurViV5o38+sAK2
yolJ9e0Q8vLQuwHwqDJzTatw8vH+xP8fWr8B84Jz+zp4M8VRy8yiCEoqrP6GNHOkdAY2z/KlvuOB
D00cEddf7ZyfQYIjEZ26REjuN923kdcWbgcVXTDJ5LDlROLFX7o+0U3vsJVxcPcwoKm33+5rv35P
EMXb8RO7IaEZSjPe04t2z6xQSqk7MGTQQexmlz/U8toySjX8nwuLLKGj5CiEyRoseK+iDHaGQOaO
TQ6+KwualK58SU1dFLqgOJvrY0d2LVXVJIcXMMqBDUloUDe3AhovW8q1gzLDXXveeb63BhB33lAv
lIu7IhS7TlPYjsDmN++3a0iakw4oWtaaOb3YYaMM5GeEzLeiSfuSNqVqOk4sWbwcLwZt1W33C1RD
GuNtJUCs+dyJDWOPO+J7pOmIerAEvYcGlC2sBA7d2JgY5rVpG0Z0tAKR/EdAp6JG0FoUy4DjEw7T
1x5KVRlWU2+YjUwA5wfJ9bOSqrnsBlRMsNTC3Aoa2QUKVbrX3hJVsW/mVt2i2DA6d7+QGBh1dvm8
JuUab3gAIIpvGdjHpdSrt5TYAGRMNud++Flrr2rHHd6oBxUcs94kf0LR37L9CX+9zG2MpQpu1boF
jAHPME317XfRHaIOBcVyb5/F2yf5inasFZ5WB4L0MctIiMNNpqaOt0HJ1xeTJWDSDILPrpGUi5uM
k7Fc+oJ/qU6m9W2IMiTmol7pYi/Ru6bK9O612rvVqNyO5kC3fdodoKX09n1d+8slV28qjpYrIF75
2CxUK/NjMrFLaGXLswTI+Oer3Jdyqyj4qCXuv7szUjNOtyV3nRMxrosMsnmYj6Lk5kG95RiUD/CJ
F5KQHAKEyMDlFSbcMwEoYqQecEQblD5UXUmqvQtt8BWz3Vsh65lLCzsTpxHOcL1BfvHsXLlVtna4
kiP/vgNobjw4jCnjrrd8PJve56u1U8a82Hxk8peH3fXJK3DXPHmsY3N8dOXf17iLbvS7gIqr2XN7
ST2HGkOPCE35yFYsYhKoTEWXbjG5YmgqYwWxxn+CXU3WBlDqxLciTzLah5S9OyiWaP6qBEqnOLhE
iiyQ3wyJSplcMq6Nhp8XPPBZIr4e7nbwAwjySLyNPSb0jERYfyEyOD4ZjWlcVizRC4Appg8rN/AW
fKnNj4DY91ZMpY2aS9iXZ0VtMSikKKmUp2YiSSEl20Bz20qdVFC4kivBe54Oc+sOpU/OvRH7w+j4
Ab7DV5SdNdxTjw2gYBvxGqi5SMEO1TL5wv5OBJ9rcoJFOSfhnt98b9NClA3l0isoCXMkespGnZj6
ZqGPFY0SEGhMdoHSLfiZMBhHMKoNKglTVatfwLDfqfs6iJwVAVwiFfZYVkzwd2S6Qq+cNY3H7fbp
1fJg+Utpcs1UImsA2wVUzfoePMPH5L5ekFGzzU3x/vDLQn29RkkABSgGoqiscl8k18g0vurk+zzl
rmmlq+/hNXTvWDOI36ZTZXxChjdHgTHoFs4tZtK3otfn8PikoLl8hVygIJXNC+PRaZBLBOsPL/gl
TrC8kpicuuxysURQ669E4AoP4Zo4aNzjLVE+braBHkPLjHoxccOoQHKMhrxo/kKgmDiYLiRFVXNL
ktOe4rcwlsCS+bw56h9yDTtn5POsYzbtWNLmAQSWTGu19d+VGLf7kCr5fY5ORZ2+0KeMWh2/ry+j
eisL1uFnefxpL6OQ1DXXlYrc+AARaSBOjO0bOI2StKFz8XpIyLtS9Q5AyLkftQIXnGm/L5SQA9rY
Kn+5VAAaGnJteLaEK0ogbxCY4CCVB1XVyWqP6nLBev0HssVM3iqm8qqXnSQGbZDH1aRnYVLlJZL4
xMLSaWQ6vaJAqB7St7Z06QoHnaxlTh1WfyurLdshQtThJOpgyrr1gMS9K49SI+IptjInjvVtjgTA
A6Njx+xCo+1noeODDAPRxBL3Yto0RjPI951UblHY5U77P/ewVvGoHkePiZttcrl0/R3okq2kCTkN
tHxPXB/aKZYxMxjTKxRqP+Z3LHDhjiAKE9jwXDSHfcYKjBGxFsLv/HhWiKBT6y2QPyHUEIXTV/yI
Hygy0tAxz8iEPuI9PPrnW7eGPA+sYrxFBOXfLPYWiteqMCq9R4Mww3tDqv719hYLQWUggbLssCcw
uZl00myWLLCk+2hUMXUUyrDOhc2n9TkcSswPh1hMjPS/YKYlwgtEukxgJBLmZatd9hUHONqtBUku
3lFdOEQGTXArYWPazoMAvV6yx9hwrXxrRXf+6EBFNravcWQTqzFoN/5NbO6Gdm5qCFXgA/iOzxwQ
aVRsGtlhsjOMMueJ6ds+nX09VPqZM7ZGEylR/A8BJYYBpWx1E6CrVh6lrok6G1vgC+dpRX9ZzRFr
Fmf1S9A1PtrUhS0+QM/9Uv+13jxbVzAm7EDHfTze9JwzF/KS/1MAR4giGkq00yzoeyvq3oi0bZi5
Ob3DxEJ5crKwIWqEF7Q/gi7V+YEwxAF9byaJeJ0avYt+hNkUiiCS3v0XXkSFh0YOOaZSf51Woq0+
Hnpn3BwdWierlUbDegFW2sC+5DO0lk0ShSIO5TnfHsWMmdQ7TUAmh+pGoiEjh9D8EKODH4j65Gx+
R3FsX9la565HG4dvh8iazvLLvbE/dDviNQU0VFyoQk12YQNcq4w6vfP7GsNRyU2y7BCKk63OcDhA
6T6Ou53wVZp5INfTDLKxnZNWmg4FTRGLPpdbHELkTYpTdAyx6/YtfQ5fCSy83cvGsKAFvjMsQ8Xf
SkCgR81df28M67oE7rxhT8D9k/1mbvm4DdnKkDelS60bgwxyn0WT4spLOI9ifE9CRWd5TqMdvBem
8z1Rm7UpCwEzbGZ3TWS/EB/a+WgkkX8XrmysOKGqWuqmxGHsRUdH/wXuGLFt2aJD8BCYpy8dM9HG
WOsf0x/kzoiQ2kPo3kmsvChla7YfkH5MuTKHPaZUdV2WRL7uQCRKc8XtAVBxvdxRlYI/B/mW+d3t
7UvZDBT60U1kVN5Cm7UpluuS+EPH+lRXXJMryT6fLXmb5aneMkmSz0Z7MLIAWdetm4GKJ/FIZ4/N
nV8kTeTcknacmBJkCf5tYD21YXGghzf7CiI4KmZCVQf7EGAm6K5n749xsuw6inIf9liU6hb1qaKN
FT44RGgZGB7gW81ja/7gMItwIO6GwE0ICkAb5rGVIQr0ezpyTY2prptmyj1wh6efxkk4VqZ4djIK
zN3fPD2VtuaHtH+52/tSqqrEuFy6MGMfKXbpF6ZfVGsiJONggO/djgb4ZdBCpB4Qd0cDeHY1tQqR
Rdnfl6qAistC7w3sNJ3yvl88nlJND0SGLns/ni3nPtHkN7Xm4tf87rIxC3h1hFAGTWv9fgMP236B
mpxj+glNsn8HzCaP9jd5cfTaMQFq5GF7vD087p4QwAFpJKlyB7HxxElV383gz43TeIvq4MkpzmOQ
sMDT8fDpCUbwwEOKHI/6S86euaopO/L8Kd/Y1NpgdrgRyDILU1yVcxjZn75ip6AO8gIhru+fW3Ci
ShcKVRu7JUILc0eKVuFY2bEun+vsfo7c5WxF4NFA/Dso4SLkwpcQr/AFRDK2oMMXt/vff4AAicWe
w01TQasuOkSbqeFjx57t3EoTt7uOu5KVwvb1snWsrcL13GJ6L+4F3nWTOtzHRxH2lY1rV4SvJFpy
6Pl50TEPXlru0gAkT7k6ydoNgg9h++Jf6eaRkj62QJHYuCF3tW8phHktrA82LJCWpyxWDxKKypNd
Ye82ycmqurFtyZpAqRS3PVWW5hUqufw0SG7ODYN+qB76dx9QI9qs6R0KLQuP7d/zuQ4q3KWa475Q
fV0S/QBloqGQCZyFvbwJCWBeyMWg1C+7FjURscgQRr86R/2QFJYdlH9EtS0FOAGDMeWrY69t6Rky
5r5YHrqCEuiAbOZT9tGjAy888y14/xVIO5pnWBQLHDTXWNL1YsJ+gwIJeupG/Wu4FVP+zqebpmvx
xdCw5JSJQ6HY8gRsAFoMCtMqUabxKtLfEgSCkjsJMnIuuzY94exhl9cWFjIrfSIuNNx0PYZuLEYV
GPxavclYYxnQpVCzjWNDo07if0vkwHGyZtVrOJi4KXUxWINfrZnw/x0ZDz225xhjiH4giTBCtpVG
VHPBreY7aUlcFc5vvql92lp9Zjh9rH4XAs9N9ikrrREEr/Hm38U+wXQXU/Go+m36CHc/+NiMpktV
zp4RK9+TQNYH6/bp8gcTIO16Qz+jcRt4LIDr9337P9yASvgpwDnK5v6Ba4u8JYc0OAvfLkowgr9Q
x1aaRo3MvE1OP7FyqMMulnlVuq8RWugt6SbB4Y3LSmqpw2z9mbSTert7vowvcPzsGC0spo1jhvJ1
9VYTOxAPSukyWivP6sgS9xBteofdVTT66b64V91RBvmOeuXaGUtImbDr/4FGImbQUrwWSB8CSu8S
ubNWJIQkwTpP3/xWRqbYtihuRrX8gHU4/3Bj6LgGovVTaKwl5ZdSKLmDuRjLb+dkMuAjgr6ccHXy
l6COf7exx4QJ4dPAQFcQEmkq3fytDWYVjHXVCKDmXEW1Mm9Y4MuOS95fvArQ/4MIFs6qID/yOtNh
VCE2lX5qjSHgbeNI8wccNyRm+UppqlahYfwrcvNV5Bmjy6R9y8Y6TmOdMbQdu01Ud9eSkqSweW0/
AnBDQXJc+V742AxT/aGq4wfCWi0e/vdl+8SQua32ruulWcSPjfxEfa5Mk15YShe2R4sJI955SPKY
Lu1TeRDpK3WhLZgPs9b6kmtLRmLbYIkExEjq1t2+B4PlF7fGI1GHJi9g8bAnWNGEZlFwSZwMUHqR
YekVVh5QpAw/gEeFzoLwggdAhUEYZW4lWQZ7EldhJ8teqAX1TMweRs83kXGygcz4os/sXXkDHT/k
U4FrCAJtVMrNyqPCG6exZs6vGjsrXs6yT56k+yfcyHXGLX9YmzXf+lG7TXUKLrbdgqPTVsqzghm/
f+WfFhMbDHurQmcvVofLmJqSt6NKXqNk2VcvpEOEjyXOW6Ps5/hEimQMYHjbhK1OWJXugR5zfVfv
PAF3ZRnkw6NK4kYjSUNP21y3vF5kfiVRs53kl6FwtkilO4VSxOKlBJ2VVpLFRxI2096tifWV8Av3
dysprKv4wRXXSpU8o0NF3apyeR2CKq9dr4ugxWH4Kosi9BYnz3Q4EztngMNm6mVyzhjMBtIuBTB1
3a+cls84tLcUH3/ZikqjqIkxijMFscWvW6QwPXVh97fdm9hhl8Gr7nsQRGKiQOSlHRe/rwW8O20Q
5HZPq3p9iotPcjjFq8/IBmW/y76+hc2RMERxGYgXk+zQHSVVaRjpYDuR1iPF35EzUKdBOyXCJltL
/F+2lzFF9JY+wz2EA6bMAnFG08pYOb3fbM6DU/zMybkdGacqBR+LWeR7mDdNlCjuQv+WHnWQEQHQ
1ayPtYEEGV7CAc/tUCVhthqx4twjBj/pljC8MiMPjmTU9Q+5rCCBzpmILUkiG/tSFr5IMLvERUd0
opJ6aMCZbsKHPiXg1k8EhRfK41ap0XGP0+L3WkeaO0o1TDPmB1wXhxUIwviOvf9Gsd7bNdM2OCWZ
S4b1iJs9xq9IDBJ2+aFqQ8Ix0XTcn5wXr+w1URG5S3Cs7lrOHQxPdXIj9wJ+YBixs1WqcC31LImb
HxzxdZjEvALQyZQar9+cN6MKFAXOeyiBvwzQm6cTrZjVPIHz55h8ztDT34FGtysl/SK2e6Xs3gFF
9jxC947hXsY33N1eQV0eqYtYPzlTPLkLV3wiCndIgOYs1FjvmUrOp7vASDnWiuj1CA4YDmCZ0ooa
RgLl6KvzpYkw38fRpcZXJCyodl/HY5J5TAeoidOX0iJ+XiZJTpAg+QVOiiAKAbdyaquftsFzZY6i
lMlQhB8fh5Uhoai2fHd7h6b136D+ORKdkSYIM8daNwUtR2O3EMCyiPOcFPxtEc2nPMr5HVX3i2EY
Bix1dh5DZe4+XOf7gXD+i21rIgWtYZjcGh2fgMcbu6OUxqCVGkjHI8KaIB1LvSNhzxscPPU+2L8n
XkkN0TPA2gh4JxVNBZ1xs/2xdqpSbB4VPrJRI9FqNdhMxwwvP4JUJ1GSCGSg2giRb6FpnmWCRqGe
jn051LOUY//FMTCt9otCPPGjMx7xnQBboYSIE8NkjtD53xHzwiHBfFyyPYaZdrLppPGZblDvOqlC
PmHVZyJsxnoSbjOIPodh1/ofNmICZ3Dzcvrwnk7RH5yyWrPvq3YyY6WGCg32VzS4SNuERvebySnx
JXsQeWHc56xREXXeeijNC83Mm4fO5cfd/rOMD/E24qDitDEjXsZ5ggCY7/c35cUbomRt5rN/aPZu
D+OTNnaoRFSn+A6+r6ygvebPxJvDFaMUNPQf+lRAJ3uhPzcmAj1mEWL9Yq4+dzenlG7MXHmYmTBB
Mi2XTPXLc25HbgK8I09O1AoIk3sJTFkcWbMn9qDvgDZe6+WYKBFtLFDT2YNZbTmqO9jh7nH+l6cn
ssMGTG8lGaP0ykkVlAFz+CBRod8YSDaVAvvTHTFdAlYHFoSKXW20KINlfKJP9g310vwO31qPRLi2
ZP2u5XG8r5WECY9w1qt+xu9vqzK7PYp3jq9TOZOUW2DaHFqu6qYyl3K6MWS8LrciDWMlhzQ42AIa
qw7gKet7SOErfG/WfF897M7GMACCL/+Vz6FsFUn5pCrkdpE3Dz+b/9Xg1r0vdlICdnw1BNzFeZTH
D9Ywd8opZLiTyyuDWWW0aRYPBHv4Q6klvW/3vQKsqA3K2NQzmIsyTa1Pq0SKXMDllrbqC+loiNSY
HtTWM+30vOC1NcrbP6dzz4Wx5d+3FuNSJ9eYxZTZpRl0taMGUUmi1GyX6XXC5RdmLSG4VhvibxZ4
jJTxf8pYTouqmIcx17v/lppwJspxRgtgF5/u+2wrX0CQtLA+iZ++I/JVQV1r/6oGT/9PdEJtALHB
xshoryaxmOzQITBwHiOTDSQsASlWF2u9k8RS3mouD53QzKYXD6uCT/U+6JRr4PzInLFMMiFfO53M
yUy8OOLEo329EBAg9ARzrP8cUpkXtbDLYyguw8jxEGckv05QGE09WJn9Z0MhXNNzxBMwTydAaJcX
OzUMPRxB9sFubC1+0/TRlFePhHSokL1IIksl7ZvSJwOflLuY1a+O38gS7/zMHd0kBepD5GoWSvW4
uW+67zstzuPGKRHGQqrIm71LhyQFTaPbjv+Ei91GM/I6d4SaYrXgh+jdre5gJpHJCAdJqEKs1KMy
CmebY0YX+jbGTNaZCwAfG9pBBLCj3kAIEF1fH9+OUE3Xak5hK0RQddPRYE/FW5hSFagSLy9gMrzD
YjePHmIEAupVg7lFBeitH3WtzDgmbaDzzK9QpvKXJYu3PuXlACGpCq8toC9QI/6gFL1GjE3Zq3hR
Awc4y5PeH9hOjekvo+Hu2rOIKv4nJUm+Z90y+05EjFRgWYUk1yOkCo2FIA+JVSC7zklJebLNzzZ6
smJkbcaqKHl9z4j+SZhs56SHpN2hlQQgmxykUie3t9BNz0kCSZ85wjg35VVfS3QQhpehaP1VHvHh
TThQwrJwnjqjPa17AK8mHPtasDVyYcqhEvuFL9j+qTUAtGVXI8vK1JWmgX3VQ59NvCsr3DQeq1eK
pnsIIRxxlmoMADXfaonz1SCENVZoQxct14nxqBobqfSWEwvwFRM26Q6Huu6RTTnazqaA/6JiWk6Q
tDqmqSKNUXyOOIS7Ys1Y5+7nrz1Ki7vwlyfZQErnvQtdiqF2bMPXyLYSDgYzi6piopa67WBUzLmI
KYv5tXgvFHN/WkVPnLVG9Ad2KeumoujhHDv17xRhjKPpD5Bo0SGsamT+h9AoSF4Sm97v494DGAyh
GYGnbU+VF6DS62maY/62LadQDkKvwoT0wIbEXiaMDlIXdeseuX8Rik/IsXlcoNW+kik+RzJZF+td
h/mbuW4r8UN8TS4WYPiEeXYJ0LVoCRIkbOP9TWuQySL1KJTVdE5e1iBTGk9lNki3+N8BT1JOuxNQ
6U7KNeXCoDYSC6xuzXAeP3JJkFsJ7oxlUbt31DA2cK42SMhvqlxORFvZS3DoTdqCdN8/T82vbHtc
/3VLaWgwEA2+wK4OdtzEzEelvRf5P5Xvu74HD2ClhAQ+CQj+gbW/TTkXw4qvSXGpRIyP0jBo0JPz
I0KD1Ca58Ew2zqaVHlQjjWuFY6mVWDAXqga0tHuhXkmLkHDV4+nsrL1PpkLB0Cl7FeiG0VtFuBqr
2GeWTpOwK39+V8W8k28PiSQYCtTICPZoszJ5uQsBPvOOuAhU28dygG2fp676E8yDJOVSBsX5O85F
nzd6cM9UVPIjeCyvdYGrezPX2K+2I/zO4CwMnEwMM8mqrFiNXLXqp8sKnuW6Cxh25Vjp2OH8gFEJ
IoWamOoTxZzm+AlzbLaH+iyiQWs+Hh6mAiqPBG8F0TuIMvZHorpzoHYaIXeR5JkWxGaU13o7Bx3O
qTA3xBePyxgnrcNnGKk/YrxjJVnkShU4BztZtUUmNiGCsr1mG9IjllRJYkAySHTVgGovsgQfXINn
UwsK+PHcygLwoSk37scDeU3eRQ0+VhA8riKIVQuiavoyxF3AW/izUpkhxtTjDiHrp3WMHubeNB87
5WhHX0QhDRLZuj4a9mlpl09kdLp3eox28a4zLa+LvGYY/nL1O1ZocUvNHfdgZp8CwFTvve5SeYWt
MHfISHfMv9WDMR7w3CqKin2FbRamnuqBR8pnj9dUrKOTBopZHNMeMAaFfzOhqSfWnDYdWJI6ThvW
valcQ4/GG51Nkkh+j+YySlvRk7dFDr1WNPUMtc+mKKVzEc1refYAUteENlhee+tTTOPIG02Hg6pX
TXxVAt/b/1JtE8hTSrf5+hCNuG+h8eTA+603Ybm2fg1d/B1dvTDAGghbK26fsfmLp3ntDyHe9rOA
RFe38b8YroOuG2aGf4QzbkwU1CjJreFBFrgjT4xffNnY6lj7PJhM6DYr3qqMyWTxYyPpJ7wqgDhR
3P6FiQ/ZPP+0aLQSP3+5Y03cRCcKCsMmjy+LuG179HcUHem8BLlP9y89jzZHu+BX02GGa1hzFlHh
d5U8aeUN2C106CJ1cPtvCWUJBj/QoAuLwS5tZgjaSE1p4KAOnNsllfuEUjkMiHive6zzf9gViNrg
j3eNgQU9Qv/L8SAM4nEAtUUM4o9AbzyAUtkT2kewRCpzLvrfYrfl6u5n5fwAgFfxNWSraqmrh2Mt
yjOhLTK4vp++3FZ7rgi9ad0HAsChv6iYf8Op7sEw698TxsZtI/Lg7xpYnjgHCzzkgnKj4RxP9xWN
OlJq+cDY5AW6Fu39xml6iVDR/jY7d3NezrigDRNEO5GkDejtKGJ2u4LWb/UZ+J3FHLNvCgUPNif5
GK4bsv71wTUJDO9DYOmWj+c/M+P2NWExa6A6xoBYZq+xo617ZEooJOvlpW1+FBgIrrHX7goenNFS
4bBHuOiaE/fAnzU+MfD2CJj3bMnVksYd8PYP9ufWXhSk2GJ5+WogRHZ6FuCwu49DdxYzrmObmkFP
KLm4wMgQ/wEXDrAVEWkNfSjI9VE7J1d2NOEmF+FfuWNUqdHVU2m7/wt1djFRsVQDUdZbv6JAIQek
HMPy0Q9rWl3mrK123AOmjhzA2TZszNJgTcAsqXKHQGkvLsMD7slliy5lQ2qVytJFd15bKH01lKII
1ZRVQtfKHZxj/2ZzVBtOlB9uTxKfLrK+kg9xPyjUyJWnaOZGlPzLbWiPBOPVqJJZxC1KtSqEhBY0
TEfnXOCWpNP5E5aG9GwHYWFzinGZCzZtr7BVPSLk1WGVB50TfvVc8w3vzv7mh325uDbMuRvsoReT
YqOsdM42ySNAvVS8aQS7IwytEIOVFrEbc959vd5aTImEVQB0exrQa7IGAhGk6ZRlpdXqjHGIt/bL
t4eRsKZujn9FpvCi0r4dqawx+t9iRFysURq6t4cx8ejxGOQIW3vAxlX6+VP9jynwadkHv3njelgI
T9ty9PqJqbl5/lcy2vW1GOa/zOmC3YDNKakt0luCKWr71K/8qYSJ0CFazMIt2IzxirAr5JjtL/iC
RbE0bvU5N+DW2aBtjyQ87t7o+iEhEx8HWUhCA4ih7rLMwKnJ5E5ksEfDmU4SYIcyqNP784x1qH7b
Qcqz5s3tcXW3gpdLTC7/C55M1TM3tPJ28RB8xO61JwN57M6+elibKjuUfS86hj73QIGBQsAUb8gv
nTpIar6sWD0KV/h8xrgLkc/7tjCrDjFnLH+81xoZG+0Wpdg4PIIL/gwNWe+9cJOYLqMwwohbYA8W
7S21ADqC/hTZP4uIHe72WGR9zN4218esIHC19HS691CD1Nia4h5MHVDL+UF2htSWVUtVsPZS96Hd
04wLZGijs2irel+klM2yKYk21oMfb71EAXL+qLT84GXCjpQR5/zci6VeD7z1H6/xqwGJYkwBAi8o
HmdP5T/RYsZ/aUtSbSpTUKbOSbB8aNTfMubtp4Zdu2sp+71wZkoSHoJX7GPovlPicl5JfP/yeb3y
dHwGvt+72QSG0Rfdh+dsEUYGBwhutI/ZSgcU54tJG7FiIjiD9k2rqFw0DZlumGase1N4WlWmGjP5
b3Nnpd0yx9Zp7eacT514+Zl7kyUEQvWOcC56mOxcQ9G8Ju8zL/pC4TmeoE2bqXVHeYTDC6+MfhRl
AdX247rjJcm44Ph6M7BDvuC0O0Mc4Oa6Rg0000Ly9/QaxzSq32Z9hFnw30vTIQNMKzFnl1KUFuWt
MnvNaSPUDw7ELT7bkyyhzAhTtDJfCNSDhFi3S8Xdz7LCM5pOEBtwtbSzelhUhU3t57hVNF163RJ9
wu15Lz2VFY9Cr1f7jtxtgPL65/6MWJqBVDudnuYKriXtWJxQ7kpUBxzxprvmqRLDiy0ZMySwiAxl
dlzUesiDZeNsqgY7PWFz5dM2jBQYAqracuTGBQh6uTPt9k2pcaYCh4pVSrSVc5TMJyVB7VveQSot
oocPsS+iUp5Rjqjww7eV7vY+QgRQky9CoA54HE3QCstEuxzYLzOSaWRjHThk5lFDGZdSHi30qnRU
5C1yvdqMWksLPhNFm6wZWU/xaQljy8L01xKvNNkrhNVV/K99uVBOdBWQHh5BnViYU5GofxyEMRVO
KqttcLQxRm3TmweuylWUHwola7lMdbkfJ4pQw7kqfJax1uV3yltKrFaJT1MwK3VysDC+hqzso5uZ
SFM6FCrnXSS3EVgR2zXtSoCzKQhzmTVdyOtcSPShgqzUuz9SIjqdC00j64ocO6DnmoMhVfaivE9V
dzGLLJfPzEAbGPU1AnKnkkDP2A//AMCbkuiPQsjfKA5tGKTRwthWuWw4bflu+e/rrUvwaGQ5oEZ5
JtGMQU1xz/sxmLt1ghw8vBW5GCoB5ctt413ftxVZwl+ayPFwScrFi4xVNmo4peAJAKuhcC9Y28fM
iX8wlP/Bl4uLFGbQ35kbuCWxOp+due0bDm+uNoI57AMaTfzR6oWlftlC8QVuNK+khnyEbZ/0S9tO
tOkdMV6Xq8sHYVNpDoKa2GHcF4X5KZsXLwk0ybfHMyFv3kaDlzeERkApZFkzr9zzOt71P/MewAyy
eNpBp2PQR6BF0pXpQggLR7b2bZ8qecdFe9e4XY174lkwk1mRIMz/SZ73fGilTYXOKwv0iKQPE5DL
OvGt1zkbizaBVQxUMdiNKURSDtXdBi5vcgv5XIpJpI99IJVcMOgOorfY+hYXBW2aF6WgTNYXcfKi
swkyS6gdBRXCo3ZVrb+oH8gPaaDA6R/Z9oD5SiYxzpMBq7LOOq7q38N/Gk2pY6/1Hlwyd2fl24Dg
FYHTYWlVD+cghug7Ihm/IvsY422J6WMX81gIoSXworwpTy8SgORhAJmGlRKJ+/Q7DlHsGGe6vKYo
K2x8TDOOjRBj6CcSIfUwUXP3S1a6C2IFPy35TrF33yzuJ7Ph7ejXXGC/WADqEkzwgzF+5el5tRYv
cM+iwt9eOYNkkGdhzP/SzxJdd2T87wYG60fh2xiytijVv++rdZ36+8AhpASFcEXYGwNA9K/AxvjH
s2kMF/cQMHQUtlKhpUM3P64P7guyQ8YFZ8knxhOPYGwT1mO2SVTgHVvlsxhqx0DbDF+JDsiyxNYD
Abu4PaoaXoFPvM5UTnV6D7eVuuTonS8dmN/Lzmjk9l5e3b8ttjJ00FKyEDMHGtpo3IAwabrHonEO
7rsGdUZ9EPz6gHWYdyov6qbHtrMYV+T61arxoZWDeA+B72ZTeV2BEkkobFnvq25AZFpRvb2KMShF
kIa3GMYyTuBRJjaSK20F6MLA6ZA/ARPVzC8IS0yjPvXyn7+lbMsK8aKTCAUTIHloQd1obWG5PPcq
NceZlwmyRbElI3POuQhMVfl+fhsDoRX2f0RO9XmZNt/HGTtaAOz7IHs4xOzUbb/e7QbisCSM1JnR
QSM2le8gfMBNPRh0ms8K12dHegVCXsNlSO7/eMPXrrMqyyF7mONK1o69C79oqRJ9QqNCrqO7iuHV
/toWmqjfPC01KrZ4xv4FIuLhFiVreyw5HR4KfT1R1JM6elEh6wtyOkSz2Ptb1lz9KjpGhhp9pKJ4
P0CdgSk0aq94U+RCwwi8/Qa1rwtJEapiEHuiHSH/PNNC7Gn57R7sZgkqkEtBZ2yqwlzwF9amEtai
AA3RL4Aa7mADPq7tDWH+xgHnHC8BFpZ7KaLdsx2xHjVIwruybS4Erhsi7r3N2Q8n9pRfRxVn8Sn/
Gxonu1UXVAA83Knq5veTxgIs8H2VFZu7q9MPHvT28jVlUf/jJ4ZNAIelW/9w0yet9qFULv2pMa5L
j7k5vPzS7M9bNPO0gIXzUxG1vPRkIjykxxYrEzpaIoTPXmHnzlC5K6dWFCPzZFsLkCxP1mC94+6f
vli0AHD6cUvBXUSHC6uRJcYg0lartgnTHwAl9CgQaaNf3ePRzuxp/JjkUdrvwdnCd1JHIdFVDipx
aSMQxw7RmWNcoLEXTROGztSARGH1dyWmg0BbzLGH+/VAoqYQ3Tztg3nlmj/zi3xVVr0SByfxWkIn
kOq9AW9vIUkNthEet8P38GM9YM+ol03e0cJ0Kpzb1hJHuw1Fr77XROGf07bycQVQLZzWvKyHWOzu
kgBYYGWAYdMScaKrxoeJ5h56ZfAIidkaxXvRQfE4VcSyN7SDwNRb1A0jW4ikDZppDJFfhK8H2rFG
gyZdJwnxFb7eB4pVY03ta47M4n7FI3uDk1kVtmfdk2ObBjWgObtBa+EutdB2fP/hIvhe7BioU4dM
rteQdlskvWtUHSCijQxMuJGnvQemjZI8sV4gvP+BA10c/jv2diThMsLeo418l/zQ+s1q4eGHFbns
TAFg4YZ54QVkPJzidnLiNBUgs23ZQZl79hf8cQsvbr9sdacnwvOD2lVQt/SPnFZZIOq2wU9dx4nu
wIhagQw1RD8fxIhZNeZiiSO0aa1/N2nCj3tq5vilzsqUA6WPYD273w26mbQTJ92HdB7rCE1fqMef
NlOIzm8b+j+F2ccR+GHfDivvf17q6wl6gLbgomSzFg8DRw3H3/+Iml71oOWOnuepGqe+rGHxxU4F
cTch2fC78jJeWmGz2uRxXZ2aztOqHzoFaVshVYG12ZrcFF7dOYhjnM5joL5EVxD5ybdtFo7TKRkF
W+BC4t/UJEmwiJ2049AFrlcOgIh0qBh+eIpBLwNyX8aNzPWwwL0A+zpl5V7HVlEr+LLG6uOsJVS6
lTzFz1sW5qHJEBgNPJ1k+ogkdjAYgS8RCzLb6kdR9897K/+OYNOEg1q38VTSEdnMFMGAE+5xctL2
dSsGee8OEa2ZJrzAA21jH+b3qb1MC8OLVj89avvfgtsfDVbCZMYamB5b8sGlsIusuzV7hmcRWvBC
uHQB5lr97OpiN/GKbjJ+VyPOPceVglEh96z1yTB0kpF9gd/mP+dBp8upTjJU08eM6IgmW4RCjQ/0
bjQUD4L40WE9Rch8jgDXI1NrbrTt4qpG+DKVbS/v+4wQcdEtFgMMkfo+hSqOaaq25TfyzUP3UJgw
bvn42TuH9IvluIEq83LsiHFHKL1MPWnso+wPlC2p0iedun5BtMydmBD6UtexUiHHupkKtE5z+CXC
ibyd0PBow+EBgMdUhvWFw7AdmOKqg6NeVZNnnMPR/oVkepyz+a8gE7NNmbjzeN6nfREeXdijdd6N
uEFEBHrFUC3fv/81Xm0NyD9wkUqSzhMZyNmAvbsQkg6wtq9+vXAWKi3z66JqrRGP+8TbOJMq5mcE
g7kqwcgvvBZ0HyvQFn/mUqOFznaMqvZtdcVedYbqGl7NsVRbJtulj27Sv4Ao4wH+vEdIcE1DJ6Hc
Ftrg3BIKsqjzQz/E5Oz7GgNRLVYjvHPOTGzYy0enh/vQS1/IcRfnzgRtKP/vSTViVdY6La+DoXKS
INMZQT2PZZrCEUbmOF4oRSMRQ1NWipSYLQXwcdfvaergeWKYrHppdwpl75BpmRm9NrxWiJSIrMxp
9S7D2epDUdceBj3kQrOjwapf+LGlHBLEqzEbFPkTRcx6/7QnG7jeISU057vbUQicVafk2deeg5OE
fCsHMd+TI0iE1Q2wfYpbnx3FZHe45bGcHM5tAfwpkFO7CC0dZ3w/69ffzP6Aa0nRzea5ePofiZUJ
s0KnPUuZHlvcKgvmxqfpwiFUv3S9/TR0F8OYjoyFQXzOWPF6BJfs+wj1UAhuDNC6C9BY5caQEMIy
HlvAF9f0ZnYv/jC7mwv3cc3BWKYkIG0tQqfGqJdUQKYwX3l1X7nq5lwDjXjVGqgjE2jLQzIPk3pN
/9abOoaXagbQmnxoOdreFE74BotbJRS+dg0r+AtWRCRD9RVK5y5iHZtI7DeM0CX2XP7oGwFmBmXe
i1deFuX89MvQd78i2rf5rcmlHYit8CL2t/6f1y5DGVPR8C8HUxFuw32pmZM9Jqk5UWy0pruhQgb/
MuBe9rxLHLqSkyUnutk7F0+rnTCAvtZI4oeX0ZFb1xRKikTDa0zWnBrkNWURfsOBs6wZutb6ETp1
hBZi1GUpUp5BVRlowtUVrWugUHpzo307ZFEYf4HER8U7R8dfUDuK712159HkfdT+S004+GR19vXm
uyEtGyMio3Xupj5J839lt4EDzhkt3DyKhZPLmUbPUDRuwWkWvUvpyZRwT4L9cgbbWEDkzk0ML988
0S8fK36OH+v/tP4vqIYgXSV7WjBIXtq5dQ4Ui5r8djhh/OlDzwUbBa7lVYIlLV77Rf/6LnD6n0Qd
NRSbHJXJVRB5j2LAXi6hoP9/pGs5Z1GKLsf8Tb0C2Zq2KqRhFyCqRkGniTY980J9EySuBgMqyS+C
o7P0EZw9IW1mX63EeIer1m/G5GK0AANZ5v9hwTgzBRNSNj29QTjFFEUfh5cgQWIBiMUjDSNm3yNA
TuoxYLfoqLKTDDw4odpIO7wugJsDl0cAUNFE8p+pjiJcg6G70lbWnovsEJ65Nvy1u4o14eiQVvRs
FsPJS9FQxKwTe475IBvIvGxFaFMRFhiYgS2vmNDZGJx9FVyYORxzA89oZkZU+8Sad85STCPFVYhD
AMHgzoK0I03tn6jdE325YjA1nWS/Y7Qk5ugTqZ0zfnXzlvWdELJZp+/jXML06gIYBCmQsTAf3+8b
F0RAsFmifsmuhUr+aIv4iM+xV1lH//clpdD9+L8wO2T5h+Zjp7TXT9VmyR4fhXJENDGcOGx70aeW
spi+Hfuiy5xu1bLCPSBW2k8O23zcptfJIbwIcUTIwZXmOgVzG0ikXlNE38MhWe0QqSrlK0a9lJRx
IoEB76yJErTw4yUiWX52LtH3ra19RQyN8rD1sAHLI1HlZZ5kDvKRYDER91iAKJ+lo0IoTa6puQM0
U7Yd/ySB6BTBifJb+O19ppchEqmGj9E/2GNqxUgOsmT/8CrErEN8a/6sck8LQXLZ1tdgfCY0uRbs
X1vr3wWW7hqmdkujINLs+U8QtyQfQx8Sv7XMeWgUcODDk44y8djrAZHU92iXX9Bl8rpE0esaGNlM
GUuNMIupgA3g4qdpaaNh/1DszXT/kCeZglH2Ls/Wmfjy/2NU3JWAJpvvvfl9U7lY1HOq8aRhYL12
01Nwuf6IYuSq4d8hM3zth5yWplbkX+r5frm3B/ugOasHWVWvbkXPRQ/v2qn0WZ2kdCyAoVc8DBnt
WQ56DMOSawUrwOCZysyC+XVDH4q3Ey+x3/iU37WmxNtq2P+zLrqiai0EUdw3m6oW49M27RnvKsB7
DxwbAIArhwYdPV31wCEYBw9dwqq0j/TXDDVPQgKoSZwN2R90/hi0Bqlb9BiBh5PSBeJaSOnGx2un
Im/1eFFlEWlAfd1MjZAbO+QhTjw6QEl8l9Urs8AaTsJKOHa/iIPtkGlcoGmMaag80W0m8BEAuXqS
SD8GQ+5TZTLo4gjtMRFmScfMMHrtim7BsFhDaraMJdJkl1SzK/1Iblqc6H7UsHAnyNT+A++3fyUS
xXsJvTQ5/RdNRzq7ihT8QO5vC4uD8KlJiBD/K9kLWvDkZ54skvcMh4UBaw72KwbdSWtTv53zV8Tz
DXAm+0ndtIQfk7OhRjBnEFQP5bqLXd9IcJyT+EqEBGSkj0jNwVIGfGX091jEzo11dQtJd1Bd5Pmq
NsFxeJvyXCmOFVhi5ourNBhMgvfOe7CbsrVbtpEnUKl1EGTde87uNmwdbLp5XIUCEIaq//JjEQRa
jV1P72F2z5hOmuNuOmq/RKRz0HDWTGwu7Sbk8AqeB7+HKaQLduos9anMDjsYhE/6nO6kA45Gmxvu
wumgxFiLzSmgVR9A10JG98s8baAKQY2Bpv0z1nZc+6okywVaIA7hN7KzdCbaibUCX7KwfvyQ9tBG
anAVrFbA7NpvLPdjCWFCk/Pgo4ONnkyYTMaPkjBHjqAenmv+GfjGMgEGedw1nVp8fUwvsaT6KNzV
Ur0w70++HS8e3mO99TvOY3V4O/36igqW7eGQEdocvdddmAs2f/bDjfRJ0hzdqPbSiaCflxeLbdja
hYmbIw/5jGBQ4xLZfDvqUDfHVhShvtVnsCmkvlK7wRurZP29BcWaJ1uEKtfXPjbmjCzrt7HPtf61
RJQ6KdYTVf5ic9nX46CeLhOLI+tdLwn8E7IoiFiXUpk8E2r/2Pv1KkaWeNzoxApdPTDZplty8Y8q
g3DjRjmAzyts5ToBiJ9YktCgfWdnwPimwEfplu6mXuBxGl63tloqPrVdl1/s2UDJcQqIAL8FvdU/
J+W9ACAbx2qP3yg1HEcbPgBJbBotLJtPcig4bTm2piCrHV0e1Qu/l+e0c557GEyetvOcUKuNDgQb
p3hoV1NhhQJwqHHKMLCi7inY+eIDZLW8qPFtJwshxTjSwggw1h2K10/4o9uDoOOVk7DdKXI6SHNm
QvYpL/XJ6Afm+vRuui5VcoAMsbllhWX6lTu0hDpO6kNBACddlxPD3uiK/pD43Pq+a3BvK5LtVTdt
k1/R3bAgo2P21ViTKcMJsTYLRciQtxHSQZPh7rst5VHiiFRjY8Z8W/EGAaPdA8oSKbroYBAGInCx
RMj1oZOy/B4L3gvn8vWtozjy9jbFuHYNd1VGQ0QH2tRzIx6tPPKY/BbF+N4b4uyde/Ezz2cXPXgZ
63rZ+ZWSMroyOJnIb5p4knmgCmaRJzKtzUopDa41fg++1b+zf04DvQgRvRHMpq/+/UzQ7u4SA/pV
vtY6virwC+Tkqg5Oh2vtcV1/dPf3KLdp4b+RECDgsfoF29IrR96D+r+LzYlz56nUwiOUt/FwLMRx
ZLwxot5vKpocMt91vpqx5KSq5AR2tlUHfHpCip8ZIQWFrZTcHF79A/OVqsRIrtjtOeHaJ8YVqLPY
r6PPP3JbCB2wndGSyNf8sLWHl3azjdvtjjSNRxTIHvl1gmzh/dkSziOueWsIMvu61bwy1fc2AowK
7muxrfl944/+vY0BWJQUA308p2HneOj2MQiN1ffraTkrsH6Q9kMw58z5Z9ISaWZUNqLof+kIfENo
JLE/jP1+KYQoa8L23hQ0rpX4f88NDdRF2GnkDCw7GVW29I5/0tJNhGr33hvC/nFDGWZBph14AaDN
WUU/jJyBe4wm7n2UQ34N5MmSDA3oJ7ZGnGJh/TqzVONFv2EK5Ld+CwNRgWi95p7x2/kxSVtzsWlp
KRco1k66XYd90Vzm+3uGuvnTlauGnPR5eBTxYcHjNJXuZSHjE4M2EXEh6iK2kiWxgDhv/Iiz+joI
/9TSdvusMpQwYcwN2RNY2WmDZ1kLPpmbzspm9w1q1m+qaTuzlSJeQlymxRtCoinNUr9kbsS9yl2m
Gjrmvihw03CK16KXdDo5TuiNJ7ojpcTVbYdKJmtrIsY6w5ZQKlrXO6rH+3CsCnMQRVm2c2w7pJEV
K6vUcY2vjfltjAXQITofPOAsdSdbAm3bOXpHhiDJEh6j8iJiLoBP2/yd1WUElQ2LWwDePhybeCXS
CEscG9rnlYLgNGQQ1nFaXMY6qzqLpkOhJWDUL+kSThp5Cp1Fj+P929OA6HqQGGCinCzAoEMmdFyL
i9vVQ9dFmKd3lY8d0lefpk/7V/c/04voXMEeHZRx7lGO7cPQJ1CrQe6qL7Z22cBKbvv2CMC0nmVu
JAuqR122p0ukNt2zJLe9qlmZQD0cdQlTHIuM6NzFwozD33RG2mBZqPP/IZLl4DHBdTzvxBop5wh3
8urA6kyYaVcTGMivIqjFgJbOuzPcQbNQLaz41fh5YhUemDohOYZMaV/+uJXguvDsuxWXke0+jy3T
zR8w8LSNd+9meNeFbVxaCkobumOuFkyWYiEtn0vG+YK3gxx59YsaWNd0oWbOp6Y0yNf561G3Rme4
eEebVCgf98jR5Rv+RleXRTeNGI+mAecWteNnwSrgPNPHQ7JIAYdWBWQWjdLZD6pp1UsqmX/HvzXu
UDpprZweLKk+o52KaP4VgRsStZiH3aEDhP60wDZlsAQduBrZp2CWnciibW0LUddmCFVhK9eGflNv
gaI5hyWrrB1c25RugaC5nIzzacoXfJjjwVVXdgxtyl1mbj+hQiKgxrKMgvKCg+Lee5Cmuw2zYcPS
SQaaet9FaRK7J2Xl7+ooMEWxHfjWJE6j81iXfRkJt7QxJR/RWO/18IPr6A8nGmDH+5CkrAdUTsBn
5YZj5t62bs1KhUHNZJc4WWqmSLuNejChBuQJ+m2yi2VuUF9W6TXKtwHfGHUI8Q2/RQxUA6txG96q
oD9yzlUPKrKNb1JJCPeDwZTZAbPlmEprBkEMj4Q6J9NAqzaQcCBPfPIsZUZ3+WiyC9GNpCF6XeQz
VvO+J/HBSRSRjGFzgbE1R3fvOa05hLhdTYCc1jbtB7Yeqi+ii8Ha6O4ia08oBqpPpU0ZcLCT5qY7
Zj8+s7/bvKGvxefUu+CuS+BtJ/MbzOsHfOXYOcmC1x7+N8VDyyX6pUR2YDTq07dELeClcCzD6ZxG
0sfBqKqNqBs6M5FY7SE9G44JJT5DOOUx3WutEAXhUCrRm8MGV4hQjnysJdkpWKINXAR8uG94/mQJ
QIb3U9PATB9FiIItU4Z8qWDrFRN4Y3W8fJsyoD67HnhPbDYqIq8cOPu7G4zpvpqWcB7YHxyAsO4y
T9gChddhLoAWwR4RYDztrw6JZyohwulVRVbZajPf5qsKaMtHTrPSQHd4UVG3JJd4PlqlN+SVRWUP
wHhmJu8293CTTZaBQjky6Vv6mFK0iBg3xjiKiQJzmSD/XfH4Wli79hFOA5knypG5gSOzpAwZrMTY
yyri0835o5nPLahAerUnseI1mwS54gwXAwPH7j39lHzcsgYVeU54VnuChUaS3fy+fZxug50lxtN8
tIseRiCSCbpYzmdUitnnm/CrZMxnxTxmrfuDjHjdqFwgGCjl3G//J35diL/iq7I2W1cLHuEM3l+7
0oCy2VfT/jHRpenaNz+r0SSkQaUWvBnNWKm1HLz0i6ivuIkFMqxGBAArKBpww+2Am5dvfbNyhcN+
DrshEg72bdj7wCbCVmhfrd/LTHqO+WDVJE+N68gQzd1UCbs5Jt/psX84azsgf8LS7U1/dsFlzIg8
cvMBMxEPa8IgPZfQasYbytlbwTee7tKeTgrjwsI/oQRd8ipNoNza/cUoGrlV/AJENL+llisJMe5g
i6Q+wAEh9dCQFsPDQBVcrpreZ8IyzVidNxcJkqDLLq8wvt53gkLUb4WJUgL1RjoQrPGfuKt/nhBD
NZAG55A0V8MA+FrsQNqODsil6oLgTyjIFiYnNqgl0dG8p6C5O8hKFo82HMArEm/FsrYG7HWVfrWE
RW353ZezC5CpR97zROw8amcr2Lg5XgT8qRkLvzc1nFw0tnZ/dBXTI2qPBypP+HS83ukaAgpbY0M1
vykZQDfgR2dRx4a5W7Q43JN+d2yrfwWZ+yhbIxshQVZPKprDRg+o9ww/O6iGKyM8vIC4VmrJXyUq
7VqMRCEcw5nXnjUKI0C1M+AmAG2kmuiDzZ7gyKHK92bsDlYMtDQAoMaYMSqF4aiY4cGbnS21gb0P
uLy98drVCPEDLOgoz3QHEt1k0+5Wi3VQ1QvEsnO/H76RZkRvcQnx/DsZAUZovBveIffec0Vm/oav
H1fXt52uDX3WtlxjNWrlAv0/kn76fgIACIpTHdDiSo1OwzkeqM8lzJ3DhCr3/6yBPQLkAAWzPM6H
DUSRuHaOpg7RCtQMLF1FnzQNtiec3Viax4YgqBfVB1Y+cRexpUbOgVviDxcd7TCXegiqw2hJK0Bx
dlu1ucgF8lYzvfpPDNY5K3QMUGUj1OVxLyKhF0eFNsQAR5t5P+KECH36N0WWpfnyCBZxSJCMv1pY
Xu4XNLtxUTMDiHD9/PXdxov0Ov1jQzz3Lv7EZxHmeB3wC6lT5jm0PaZuF+GshgjxCj9EWOjYqasz
HDKb2wfc/5ZV5WC+5XZ5K+W0jMcMrjN50Jm/vJPKJocqmnFXZFOCTIaJLhRYm8JrvKwUJ3P35d3j
EOVWbv6nn+UfG7jTwJl/me9GSHwzLy8I5um9bGBJ3iL7pCw7cNZsYz0xXS6tlZ+xriPJf14d7jC+
wH5y6YyPJ+ctNCLPXOAkLg4aglwCqh1/z1J5riBOIKbXN400c9kwQ4hBq83ODIpfJfiwD1QGTF2a
egJcmsdSNpdunCKRjB1MdjH+7FHRcZ1mbPDLXr0HK2c3qBIn9o5CjsMvJTLLRXDy3ugXZ1eif5Bb
i0Ug0CUQK2FAbtPpGA+JEmGnayZSKCaI5Iz8tC9VATjM+JYszXz3wxZmW5L6TftHk9Sj915SldmC
NoJy1/UpQsX/r0BUL90zmWqUHjm3JZOhoSXlH4UvwDL1g+qVIowCxvPg5c4qViDlWfa3dDqCoNeV
cAMJ51xj7YMmd9ch7g9txDI1yo9sRpkE7jC7wbnlPCwxHf/xGCKEfqZeaPM16ZsNR71cw1XHDcbm
Bqzz7Teu0VoeZv+Ei4gFp8396uBZISjuntT4gMTqcL0FQZBlwm/Dn/LWmoIS+X7ymHCRukeveaau
Ndn+d0mc2Bxht9fFMZVQUghsXnIEs63Zb3k6Xl3n+bEYHYSlAh0gtHfnroWqOugs4UW16QFtceFt
Pr4aIZeCdaPBNw1lCwNAi7VFdGqN9xSi/WwwQiL07o2gUEXlBUeC3AmL/Llf6h9d8W3vgKhtFiP3
BYsNzPytrqVugWPUD1SZFJ4lByO4G2USCnihWs4DeEY1A8/ur6nBMTNqsprse13iNUENAeeaCYTf
Z3sZ5MM87pjV+q2EzWSyNF1M0Fr1tzYEcNPYjN3q7TD7AU/fTA05AbguLOLSmwWUFnUT+matYnFV
QaUYRZJbNidvgDfV+CphjD4BSbTn2XI2tmhasWSn+BRYyi223WE9WSNIwcZvgjFcG1xLfVZhFxV1
1B2QXjRhU2k6PfEQJHevGXcis9+62mp/TdFz3os7AIwjYjbDjCiQviEFLd+bhoS9tHrXnmjDBVtR
WvVqOdUhJeyQ3nO/ZtOItqOYWXudTLA5RPvQMdP8Os8AdUoozoSCOvFILPbTvOd+i8FZAvasa9YD
KSm1O8lhOPSIzqGELvpRLU/rVjnkISKOVoxLR0jNgmAl0TGI3ryroY8Dgd+vWgOk2cCy5qgUACjB
dYRMPUA/+F3iIQm1yuqMKmhkJe7NjPjfzT+Da6M8DthzxVq4iDDLwsiZU+bsTI1kBTi+kQjlrF+1
13Fm8reEPyB/PwsS2lQA2DJzMIoIJCljoCBjVXKifXElhEDQvhw3IB3ZEkOsmJbHEHVk4M2XUZYr
noOcb97hHVKXCMUlW6+S8/LkfFzCtFznW9lq9Lx6LjVXA8fOKsKM3eqqj+8UCb6bdaWgyuKxYFI/
qbs2I/VJ3l40Yu08huENKluWXz0kZAt91HMxyWhH5LRJjWAwzdK+ubgMinrEVxICRwylhZIWLPns
V9FNoNX8XIrnUT4Q1NMEHCL1gr0kX4LtzC80fwp32IFjCRrISngapCtRCaxvRZjP+g3vSONw0nf8
VYUrDa42bjgVZNjKZ6ETPw54o1VyKvtKcd1oozS4ZOMCXPwd8cD7xDLQI7Y11BO/EBadE5kkIraJ
p+pn4HgMvkPm3yV8G9JAGdly0RjDNUQ9iaZ2EHQG/HuwIe9PiNwWqq+UHICwey8IkrgZNIe1B8mD
EMCnMSt005BWbRnYgl0kH6xwimeQYOVSstEoMZ+j9JrMGt7FjwpyzNITjIOWWgktijhaGA7aeNYE
iydYjUDJMVlWhRlulAS2rMTZY0JzA5Q71M4NKGZVIVc/oPC1wQ72A3lIJsiZXn/y8OfI0ITyoWlW
hT/7TruMPcjvcBFGD6Q9kPeuHqHCx3wWXL0C4YAHfDva+ufF635OBmTFrJGbwI1OlfFaksBAyElU
LpsIReEEkgd26qYjb+8u29o319Hc4/f2VdBHq4yaXwKclb6Ac+6PQ0UFQsabK5S2P1wpHqOUB9Cg
CtXEZDdlz/5PfZg20jYPLJJ630Z4pymSedjigmuIHzSNPeNl6faMTj3mxcE/9SJstRaLlkp3nXZ5
BzcdhWAONS1RA2HLgKzkjqLQqYPlhPr46Tgt613L6aekmKVY2/ZamFibmaciqLfOylSU7Ld4skiy
LMgXPg+q4vybmUxA72E3hKXVhfiWWigDfVtdHRm/cL3Goc96QBPDJEoehukZQ6lTN1zlwF1vfaeS
NxZF8TW7cTPVK1bI9mwPQew61gAKdVfDT1FjUgTkZrWAz58kGUTBWRG2kRLWHK+64xKfzmrsXaK5
OabVuKytncJ7g3lpAvdON598U1GIcCPFb73PpQ0qVSR8E1f+kqlHf9fkFNU7y5nK86H+/Rbe1SzF
Gj/srGo8NFvqGJvnyoKdYLvqyai954YzKJ5rVUiYGAqrUXubmJNF3fbAfPHnbiRiTXMctQ7a5av9
lJljALL9QUT6oy5Dj1meDbXW2+f7nArqgdfzK0pP+Jo1ktTr8vfs2ojTYMSmffNj0IMuOMcVfY0d
jZfKbHpn+PhlnMjk0fnaUsKsRvY1JbbWnjlseAmJtpG4c6Km0yEucUdx/F2WSxVSWCeGZa/LlOBC
aOFCRK4ZV2MjAWQo1745nLKIWGoPZGX02q0W97uJIzv952fiGW19qmAhoP2/LsSxj2KRyK959w+U
C757NBtz3cJzboMmmgIuDc6C4ZHkfxOJSX745PKqKlaQ52f6/i7cxk++m5SB2fekcrHXed3M+vFt
/tb00u3CQZ/aZJzaBj9ACBVS0wUyy7j2IEGS7YZD7//Z7LNs1YkIO2xKAc1AKfYlELBCqHuweRol
apmS3efvKiVzdSTrj5/2odZHsMQm9d1IA0N4uUwoyj4MKr99WuiT4ywBr5hw6H6ok6QJvSE2omPN
HZ2x40ecO+8Iqt0XoLKsgSwygXGjAKhFwdbrc1DXDBuaDc7ipPynOjtEz9AjW5PSCcgBILkTLf7N
RSIfLD7DoIJIvsg78HUa7x8eXHNCr9bHu9Pk4MoTwd4yV+35fuPXKuBeJry4YtInOh7l+Q6vlF9b
M3XxqDiVnjt76G3dKwJLxjLYzKQ/Mq9Da//RrAdoFXxvdz0Evfec0DWBqLbySEbSSdFpd7zD8rR+
zO+Aeh4iTkM4OVAhsMue//vS1wLaUG4sSmDSgdIbSaOpai+TnV3+ZJas/6BcGnSi1tZvIqPv2JDv
phQYZ7XA63d+GZtXVhT+EimBy/A4+nZ7VHKo5UfIGD2N1r2OpPzBwZelEp3XdF17zlrK1s9mdTFI
ZKSDiDY2z7OuhbyAhOQiGLIJlMXXm2JahlW4K/dPDOvyWkww8Ojiuh5Cz4Hy5JZDVDKturgmd/Mu
HmYUwTqCwz8TQgDalZYIlJ5/AgkLC6lVNvw67IcCaHKxQzJvCbLGvY5w8y3Wq56sV0XDeK46FBui
WGPiCXMgpAErw0QFzXy4JlRJZaPRPMDn2x0uGuUbuRLqMRVcHduN6WaEOLS3dTbN8AMIEZDQFifC
NDNxwwSSapSEoiTOy8Lh8EffZ5SO3EMeudxEZaz/rx9mSiCQHcEkabecCrFhwvo16aM3T/H+KO0/
eUqeBigXyCNzu4SA2CK1swqSeby+BUE7H1tANKeWYDoIrwCohQXXlhcYhF6Wc8lTnwf0aozSLiZY
hCuvzB6bBpAn+hCajYCLNtbJlF/sQPVovHbOGIO/3bm/h+dBx15glQ4RGImjaxatUDlL/LDb6SgY
qRZD+xFYzJFmANMJB4wXV6UVceuZLIVUBifQziwGU7lDYkiaYFgFqXT1Dgz+kOGdrgqJSAd90J4H
t1c8fNdP5AXzJ5aUG0cEnpGEMhu+ySUVirfWvJ8BJ3jJK9Xi7LP7+GxawK/et4WHGX0ZssgUuUIv
yBvPWEclnj6QiG5XqdRm6EMU4wKAaWL0DUJLrcxFAJETqCQ5SnP0PWchryuYLQS7t8JytBv0CDGl
ISAriqg44UauUgK1OgdJEF6aNzlQ7BRJ63Jr+xQLCnHZpiAUyaBHPU5xOIIpkSg6BS/FPXKvSMaZ
647xUDPobSJiY47vI8Xum2TRSMzr0WuWfN1wg4kMr3KlKpp2yTDlht1sLtpUoPGHJuseiqn2ckq+
/nvv9Nuf1EikfsbDGwN/qtPWl5CTinhVXgEfD4x52keqQBtWxLwUQwArUq3piwhmsNgxSqkz1NBa
OLw5r3LMuykD18Mj0kteqEqZ/evFbLHK8towy7dM+pvy55ScyJd/jj6nxqLSYqyetmHcBdRxVdTu
JhB6UVsHpRIiNaGDR9TRpil3Adp5RODhfmgtv0OyT66NQhu4c7POe6+z048Z5LmO1BoUqFx5I9gY
HX6UYzP/T7ah/+S4xw/MSxKdtvwgwg1O9oferzr5p2rbFpJ+tf8z8Id5LPyo74SlPqoNo+hg6PoO
B8EeVxkfNCfUr7F8Vxs7YSZetspHNvUv8maAc2X7uC4C8eqhEiQGW3dz35cV/5gChaZCocfBJupj
IB7BeVm0wUqZ9IZhsVqvbEqWMTpy9yMVZUJa7TlPCTOOdW1fF4vDEdWATuTiLXgKh6IwYDlnqHNy
tjwPq+rKPdO4T3+310qu/3mg1CCzDMgmJomlQmB+7/EqJkMmSNY8qs1WGVl8EkxChdAJUNdHp+0U
jFyhLZHQMWIHCQZ7GeQZkfOVLDGCiQFzZMjDY2xUSvykgXLM9qB4RlkDlVlkQ3e5qP5mGvBaFX74
0X5xX22Yw0vD3DrH4aBqVpUcM+Du8XpvRH7QypUVWsLUYTZ/bm/jnxBAaI851YXqcDc6fe+rrQQK
+6ohp2F6v5uc4O40l+8pb3hJOHm78KF9IsNmVa5Mf3gMI+pQwrekBFkTksaZKzAutDbTohl+6R5a
uiX984zTCLmZmaor6OuB6pdNggjWlt8laAkL4ksGQ1xyKMlt2lJw2IIOoAXxLYpOfbPBelIIWudl
zysKUhbmHGjb4Xbmi1prbayMmMjbiBqVaQRCNAJzujVVlQchi8LfIREuXB8Cdtp4wFHxFU/m3wFN
gOG5IloXCOrGg7mxb51Ehqres0olLJlhdQHhVp7nGLTWOHhx//DjthvyxFeE1/sEMHnstY+xcBWq
mOLociaYNYFWEyHu0B4Rzi1vVroZIslZDeMFavA5jJVO8iWiPoG4K9YCy2FEOrb10+TxtTkBqVnH
dWXnIsyy7pKc76y2L4ENoYYVT7Q9jGO4VJQDv0uWlHfTgJLEtUPnt9uDBO0kbMmZOHRbA6TRzy2n
IoJZhR7hxHLIHh5I/uAFGYGpJ3/07ZXb496bnO9QxzJdZhYqeqEbnqwiszm+f6PaR9YlCxQextok
rHZumCWmLGewoF/jIs6hB9i+gAcOJtJ9TN/ar2bgPBHtqHxYRaW2hcKgeX4lYwRTL7To1s4W80GK
LoIfc87oQYVH5yrs9JINWA72yYhhhCh+mEdo9LPHug84TfW02sYgN6ZsSs/lEv1MwDqoGL40KXWq
6aOKf1Te2MomoQcenuBEBIaguB65eKzlJlHZ3u6BlkJUvdNcSKRkkviAw3urodsC+8itXcIjHmKa
OfqEcmT+B1+yBa/qSXpoDYsMcfPOYk7y2CJI78BcMannDk7fwEPWM9IzK/RGMDignPw7iEJp4p69
I5qDnsmVoQAugPdyKFfeIDltmvTsoqsCyVWG3g94bHJwFyre7+qp9Z43z96SI95KQMgSXxSjfbfC
q2btqx2mCg9/n8F2rbPvmF32HNMctycLhUALSlGCkaGBja7i5lq9nY9rap0Wz+rhXksw4VX2Eox7
0FJA4JccmRmUlXqNPCIQZbq8XGUbE3WLecDfz6GpJts4jJL257CJNy0ra6QEJNXA/8FlL1nlxPP1
ciiUdrGv30CZUXcZxeV2lg87g62beceLw/fezXHQXsMBxgFqGVmk1eSvvcBWUe+pikhpfJbWOmTd
XjKXXT/ytfLvB+eIo+xMsjEoG7sHh5wQmilxXfT9Er8586MQFCtt2BOC8guFbSixSyUnDNd1EBmO
/pIaUiw0T+K7TbP1mQ8nur3tEMbLl5xfN47ZAlBR5WDjWVaUqURuEVDOmA4g85+uXGZsBDUslcmP
X/foPEomDEkJoY1CLzbF0DjOsDwuJh7SKcyjCBgPLdRr4CXrodyX9y7PV0VovM+GJ+h7MyaRVzSk
kNjbaPpIfjf/E1Ge9UsJLBCfpmhPvnNNCsqKAJX9JinfqtO5Pw8SSnmYZjlu0AWdqtju7t3Z4Tuo
CLgw7pUP/gv6kyoRRjQvKDc8Y08ggD0JPjVxCFOsNU81MgvA5oiYCjK3Itk03+joBjJ6i5ZetPKP
MkCjqC6SJrey3XeHAHpb9FluqcSZG0cXpq21RF5V5x4w885G2F9pYg79HNeOhImlJjxBVuqTQfEG
jKCaPu+NmG0SIux+M/1rpCVx+UO8X3ETHA+dW+AL52NCeAAh4G7ltLuSJ4TU8W9CuEMXHJljgz6/
BCjseOVpU4M3ZJzkRFKkXKqfb3X/Ki8X95f1GP6Jjua7bkxdOyJa5M100DcF5lvuV2Mu21nwHfDB
h9NGYLJMGs+Gg3qibZbsiS8CfYgPQZBW7hJVuFh4jqwox4bvtUpAvNQow8ywNkCllJ1/utJ8bNQu
vQdmCooMNO2hSubfSJf8FBMRgLl/GDTmrZd+gARdGCFrJ+nINf623Jo7a80dozctLiPNv/sLB5Et
9Z61f2BTjGsrDOV5ZGRv1KRdM+rG9SDMT+dQpWKJLVw34AtwY2CONcf5n3wi96KD0npEWqWgHbns
yu83BjyBCIpEPCxYzerO3xoPuqEd/fg1nWj101Isfzi0ESEsyhzrYkzKuO0Ipr+zPt9f78ys212P
4M8gT5p29nKSjjQhFnykcXsrE5pYGaQu4SO5Df4zAT+32mgLrQkqdyO2KFAMCQJeC5iSDVGi5RWY
S20da+PqRd4s0R+QTafaygAZoZQVHgTjiyGbAh+SeoCa4FexluZgM9XuxQbwtU6rFe6t5R5PTz+L
1FGatWr2hj2DihgdRBhDVnYqA22qI4Kpiu3U6tq5d4uz40PnpDOZOKIBvLt/9wOlSkTeSjHi5tf4
a4rG3sz/VhI6slkLzONyTfWnpbvA7f/r/5k5YfWOHHeMqV3Ab4cqWbue8xpKd+Z2nC9amtcD3ujZ
dFbYAbxauRRjHADsYG36fq5bp+u+mghZDiX7PKdZxOIbu95ItczkGZyYLfMTi/gbFDeZc0rilSz4
XLucc6jztPGnamrCi6mF8D/Q2ymcaSA0O0V2yXKWwrxP8WMWirRrvCwUgmZezUmzIiZafiqSgJYV
yG8uftnwkRT28U9W31GnjcG+b+CS2jsnuq8fRP2srFA8LzIdMz/pc8kSVPFFltgbuOljWq+gbrSI
RvYIc+nYZPFgc45j+mRvfbcG9GtFkZrCEepdVMAImiHXNkK7+r0GAnGJncVfub3ZsfXjYUv0DH2d
5EyQub/pXP9GLix/bEYZBkSIcSnoCKrCSX8UM2UyXk3rUzY2wnFyZflLGrwwnF7RNFVj4NDBnzRy
JNVD5e6kGRyKWNmpS9AMKqRKPY5FdOZaSPn/tNW1IY37peiKjLRP7FQs1nbewwqfJbAtEUcVuJPa
1yxA8aINQwkZrOyJWnFc7pLOHeB+aEV/uzogcrxMweGq7MEvx45NmbaUvUIIDIBwYanGUSOYMgxB
GXOeAo+ZRVRh6cq5EEgWZbwmCVdc0g6+149pIcRAw1oR41jq6895e9TovMQowD5vGggd2ZtaOPfJ
0TJ/W2ScppjvBPm3RtNy/RrKc+yOb9KjixYe1/U8+GCo3MAy3Xheay4kYB+3EpKZq5qFhoZx+/Qz
y3lm4YehpZ1VliTEXFfwMTLrZMZq9sL8bgUc0J0kjF4UBzMCrQ7obX9xqBOg02pZvCZBrOp4NvLx
Tig5huDVyP3lX1DtRUzi6VGcvrM1C/RCH+yKHcCW6jIA3FjXap4aRC+2dEzpFQroMAzUwI4hv3bW
XTH45/srGeORTAjY01Unt+lwC1P8WI20p9prkW/OheJSm7Gy5N00sC2X2IlRX7BACUslEoJXTpNI
u3rvtjC5sBKvzq0ES07698+wGLXLkEvK3mqyHizGqEQuMuJTjYQlAYJXb36Qlv/+gySnrtXVbDY/
Shwvf/bxV+zUWWYcwX7TA/ws20yGaW9wSytV2mqQg8lT/jIxJ2L340o3L5A6NnXBttjSFyIq1n5S
OgijH7FCnZgsSXIFYQ0p3c4P7sMo0fIf2WMYAj4bXcTBYqJO2hIDSB4THwaT2nxk2buSqHzu1YTn
Ecup60kmdkJcKqNZ8vqiUcDJBr19xP/xwfSMYQbmhzDUcDaTCE11w1Pj2Jmg1Ucr5eITOd+sykQv
Euz1j/vfrZ24kxr4cjKN9rGrm6jyV0VUmhftBlhtx1IGEkUKBDfGDd9vDJPoZNjylOBFXjnXfIk3
drPbb6TMKs4TzMW+k7hsncMQ61KdmGmUOwWEzpYBwdNeBIcWj1VOyeSm2YArlXVvSkexFMvqOaH4
RbyDc7YNSBK3lOQQnK/T+qJjKRtiqhksNKK2043Sd8sNkLdkpvy3Z2BzLGU+lVRLLXLZHO3FV3u+
c8WwIp2nE1LFFZ7LkDmdESyOIImvxJc6EN80zckUbu5YjdbvTyl6koEg60niFQ/qs5FH829yNgP+
3zRUAy1KC+28VnCRlHl/X0fGkn2dD4naq+ep0N7aIb/Iq2C0aWgV8ilZMDgcvrU1uZBA3GFlLdUJ
UHgpEYWxK2B9Vkmh3a3Uc1nJnT+/wqnO33loKAo1LAYXgBolnPdDAouv79W2Ahj87lEJnPc0GfP9
spBZQpUcZBFMVzOoTzPjS093sttp1vkkhntGuM9rxE78N9RepF9jX2gZbfkxdrd2uIpoCpNIJZ2t
FiuzY4GGw+ZGKR4B7SFrA1Ns8szxzMmFo1Idhd1Bp63mIYlMv2vqQ51LKlFlYuq+c4sKzquXrNGl
+pmQuAiQgLeID6hwetvT5ApoFguajygtevG+m9TJkNrXluTkjMlN7M4saSbaksSyJBmxvAUzz3t9
yGRdP4eYFBI3AYN4McstdltNcgvtUyBr7Gm9BdtftdOgTGsi+efpH/khW/4qn3rL4nIF85LI4RgK
p8zZqNbjg+l6RFPEcseeCRwC+hpQNUZfARq7Hlu8fh3SLytoEQ589NMbYN+Pfhuqdmk7ss8f9MYt
0Cs5bb6WzMAf7KMA+p4ei3TnEPuqO68YPeP+vOQzskV/PzX9g+i1e8AYPhB1juR7Pg0pfDziDy4G
U39r+FApCmePMv3TFYR7jJyK16S+9/EKAaOstruXCG9M30yioJkScF7wJZZ4CYas+M/Wr4ZuzOfp
PKE9SQsi5zwCsSyB+NGjdgqNcmStRNUbF2PcWQeFsOW+1yT1qubnkekNq209ELsj7p8JvFcfcrDN
93xO3txPAl5tyzVQghE0kXZ6Phz07+In6tJrP8yWbSDM4Wc+xhq/WaTqypQx41691/E4br0msHwW
4VvYZdm5zXOvo9K/t/4MOVtWbKOwKpSKBGcHzCiZ2if403XrKOeo2F3IaEBxY5qpN3GfPwcq7OTi
H7qk8qITMCF7IcDnNL/bACmQdcSGtujnQukjinVkwhXq96vm/G5kxzGy8L0zjWxn7I5He+kCv9mR
v4DNxBCgbB0lpPXICCTGCl5BXAFC8GQG/m1AJchoZdNM3QDA6VB4PqiK67wt6qaUdBzR6M98lDPr
cfCBo6tQa0kLqIdjZtzyuP3D2NPaXqcKnjOHUL8ZPVVOlp3N6m4lmxgiT2Jpa7A9zL2zjqbU5Ux2
iv/shqxcJ+NwW0FLxG6jOxQ9siLbbAJUGqcxTHC0wXWSPM/eMsPL7Lq6s2CPfSlHN3Atgf0eny+8
MlUxMJgpnFtq21cynUCdJV7FlMrRfJ8Cjvkno5n6ddGHW6RCyvA72Bxuc/b23oghLAe3SizSYxMV
WhKF0AArVVEVG57w2NYb6o2/RIZx+gEL+0xI2ETmG9prrOCz3ylsCGt6DjOiUcF3NIm9oF5eh9Fu
9J7VfOdKCKbtx7bj2kFdb70mUUH/TjeRvRiCy3nRTyO/67cqK7QTJUHAK+W9Db2t3KSQsgBN11T+
+TPvYFVkjxrJd6CxvFNZZ18yCp7DxfoOIeHOJml8yUAHHzoWysFfbgfj8Tr6sAxg8nxfw8Boeiwc
vhmI9PBWyjsZGqTnhGmkJR4DZeTsHtUKuQRCdA5SoZufyK1iaEMSxxxyuiPjh89u30Fs8+w/k+qV
bNxYfv8Hpn2elJW/VpG4DKxNPsUjFawjR6CM/hRV9Yy7qcnWAUcsmEVRcnwGP4fqdvcGeaJcIvEI
LlG/O37ZoZ7feupdmnugOuluQZm0HUQjTYXEcu4ywPkRLfcDlyQDQm1TznL8vsma55Dlr70ukSKH
Kz/yBg69j4+LZcImj0wlO5eVxo91Y+2Qp3MHvv5gnjmualXzEStm+kA6gOnAQ/NWFQWnV3crRP4Y
mkZzQHscSGwPjpp2UjEGSl9iI8sXBV6MtHdUM4t4fimPlGUgCk7GVWEcGu1xspPPXFagOEeeM777
f2gLvVJOCERDlTqiO2bamIy2CjoxE8o0mWxC+Rlai+pclOAVarZBWvnqOwn9IRKhPwGUhjnbAJiG
yh97meTFzOeGQkcIUZk4vz4RC0lyweBUM1fkw5jdRQLda1gitF2pZcI4X/a8co6ARsMk432GaI41
WvuNSoPR0HFjl0ZH2/T3KKjKH+2EpcSnPmf+BtRnPTxRkVQk/HC2YZ8+2EEdQa/d7VXpdbr49K7T
VNpnsfW7G7SVdetXvgmVF/fUCUiemujo2rDIllkZO44u0JQOT8wttQ3MzvWrwP7HGP6w1Wp4W93F
OpDiV2rvHkTdq3shCnhw5BuOJ6WFPFeROOoKTTpKUPXLN39sHoClBY+Zwtfm4IqrJVapYPS9WaYI
4G/n53ovUjKEAMBZNj3LfyYgJqmuQpfqMt0PYrrJxZjYFl8ga0sjl/x9S9igqlgMTozEL2BMVjS3
0zEywHfIwaesnjGg+CCS25IZ9+MV8nAVyG7ULsY7PLvpQlsgv68329W8moqIaaY9GT/vIlBaSvFx
0gy/Ukmu2uKWNaRkx6S95Hp+7xqjjTvMSFr+GWGADOopIuj6H2VBfEBsmYi/S1M53rt8RxhgcAvk
YaX39v7GuVUFn5m+7GxM3VBwT6dsxzMjQk3u1xLZGBtfUyKhJjz/z3oFU4MjPkclXp9Qny7D///j
v/jgTVFexq2iF3YnUllBiInw+ocZ05yy0t8LH+cvSiJn9qVCtLmNMjKPV0uKsUQuT6lioFsRN3H4
S4tb3Bh0+EoytU93JwGL4PlPXL07MqBQhtaM1MRVbJ8l5D81zgY+9dE/JZv374MeCjfeF7t5GUdF
wg/tmvQOK5hRu5bponDe592z2X+0hc142gcnejIiddM+IpoTRIKFJ2Uwx80Wsf4Jab1xoLWwUvga
C5cNxvGbua7JvllDeBQLhgMJvVlYHjuhffemUcqLouOhx+1hhj1r+WFXIUEvK8LVrc4OtUvGthVl
0yUGC13CIgckUyJia5i4leFioapolco4tYWnVRCV1sw59MP5KwfOletWWgzxCoXhYsgIwC+78Jqm
lKSgguXLizrKqZJ7pSxDaBlVLmbZ4hXk7OpXji7iy2RKzKvIHRzZrBYO+Puo02gO7R8VkS7EpNgk
Pfumq9TPSrdLGhsFyWX6NpQt0kdzKGGXlwd60ah5LLP9SMZwlDoO2SoVjPT04pmgJDNboen9sv8d
0lXk3cm7Gm1htztHyst5/q7MQewyU77oX0PJ1lxB8VirxYUc5wTti19SY8bhQU9fF4wSwHW8WHHv
0zvwXwxkY+C/B18npOHfd3CivrBB4OTgbTrEqLzKGMADgWKWkGdmTqtMDoPhIt1LeW7As73ogp38
9+xTZozrL83IUVL9zndYYJWZTlP88AwE+e3OdrIKAguvRCy+LEXbEd4gluEO+u28h+QF5Jr/m1P8
xapltLY/sJLiij1MH2rssYfRfxIaPd5eNdFdIdnwYcbqplWHIcOLSD539RxERPWjEaOgWgds7FNV
gcsMxa+98Vmu8VdD3v9vDzUhcPrs8FRETWeIsyUf62PNsFGYefiTJMap0hJJ3sNFbPxlTcfR0UgD
cYQJqjsnnmgsScjNFOg5dBfMAtYMPnCKE2mN9R5RU7X2aU0C3NIKe9ln4QyCLBQqgRWGYPo8t5K6
LzKJ1aaf3WmRIcy14mWM0OS4tsZKFVUIdf3QLKnznQ5WFSoSNjMaF2pBf19psdqEVqE/zdAdYPGr
J9dm1koc/0lPzaFuRplZR/aSHp1p0VCBdW0oj41w+EAW+ZPhdP0IyfcIGq5yLlsyjKw5hPNu5hu6
4VOhnogmhgf56Mh+4F/NfcKh4CoWsrzDmGFpjGiU10FJz8IIII6jV4frs+3hG8OCrYPh6XD6548c
3BOGTvVmjw4T3k80aOzVD5BtR+b+nVm+YeLC5ruYLwZGhtVH1/rr27nWhpRtNbYrbs5WDh4C4abo
B8JUsPXm96sHi0ZpDttDaqTChAYUDSrbq1/OjruzBdkWCsLPj3aeihgpfSXeZsFKxSZHKSiGNeHE
Snalf+Q5GL1at0l4QKfd4MNlbU26FSP93F9J78uXHZXEuHjWaECja97Jm4rkcWZPf24/VV0Y7u3W
y4hFyC9wELeEEW5WLVFlLq+vSuwJMVbfcr8WjxT/v47yWHfkTWvBTwqXpJqokYiUKs0WZnf15Tk4
J07MBhZXI6/YAUB7D9TxYCrKsefKtYPCCndxPT4AbVfSrQ9uHPtEgWbaraYjhvu5bVl3h9/WcDVf
3wkXNLcrqcD4Vwl/+7Kf+laKOGackI/kAlEMiJK/nClH6fggpqhZr3OUrn7EIBQQHDammz8a4eNB
VN2/cpBOzhvbx5Ph+YW4t2ef4q/qzdInBnXlJXALyHA5WqaK/Z10TKqRG3bq+gH2HjDlbeSnHEiU
skGwCT/SOhRJcZjGXEORpI88MMSa31w/htOaR+ZPmBzAMv5PxmM61tY8aodtO9W8YNsSSHmr1Ipe
VZ+VS18Mf2mdEu8OvVO5KP+95M+lWMmEintBrXeAgDjNuRhxXq5mhDL3biacKfqH/V5E0dGEVr6+
NKPFGTnkblueM7ePC0PHmXpaB8mVSx41TodpDQIlC1FpP3BJzICvVDLZxZ6kPvc1INt9RO1ySIxP
g8l3XLBBgQ9FPOpkDK0WfxAyW7HHW05VjxjooUPGhmavtTj6s81OaDM/12bOdW82kzPxXWdfbqgM
zDr6ebXZLSwuHpfr/dI6RV9Am+HJunm56qVOSRb3qI9EMu5RRPZzuILjvlaIrL5fXMo4Cw/7lsk9
CtUNcy6alL1eJpAHEmjvnMn6fLPa3ro8yclsiaPf0ESGXaccQ7Ycp4ohFI4YdAjLIU4bMOd19DfV
0X+D7sa6VIb9j/eFY8HBFbyjK86t22maSCElOe5z6DoU7rTt6xNxm13Y5rduELjnDVku5f1+4TNU
xnI7F7h+dO9wl2udNZQ213TPCCWYcVk5NdBqxdNeSQUQHR4ua2MaIhfMz/TASJuj9ljma3iMlQlG
+8TNnQ2lGTqrPE0tfw0Jkdc7ai4bVjkLwq0U10KCLVD6tRHMb/jPMRMG92zGbS85dT7ozkFpLDOb
9zboTLEUlsUcs29IGUIe7moJMGf2r1wPlvS6qnhZHgqepKLgzvl54FdwT+jEEst+KMZiYJPhuJuR
vqv7OEOIp51igVGs0JetxGNWbKWOACqqycx+kis8EikXi6fzDyEJvwcLIGJg+RtPa4bJrKz1GGO+
2j1v5tvTdWTWXEVVtd71dfCdIL/FLllFJQ50l+vL7yixet0vxcmUhsw3rEQP1Cm+xvHpxlP5VXVs
56UZgQsU2zi/Rqt1XrinDnc6A33GXr2g0gP9UFX2hHT9aZz66kcQ+TMrwJxt/tt2wgjOy19+h8Td
FncMRSxVYPqRGMIRnVpAukkPwR2ZhmF+cMg+2JOaUIdneLV6UO3vlCWVzsjthwqzYD1wOmYEzcU5
xyzc956hDPL5kiB7zaStH9dDv8h3wzXj3mZ3+NvdAuv+RIvqZ5KIc/zk2RnwF8ffYNwXTzLBHJb5
lf0X0qzlBPostP3xSyFq3xUXD6vVHfT8Ey6otnM8HSFneYBmJuaNOyLDyAyrE2amthEI+If22GNS
b08P/aATuTMb7WjK0foXAyUKC1WWMZJna4qSfcGMO31rvp0mpkfsGAHKmrIzNUQSVqaemoRIpC6C
dNsCJYcOUap68VAxSk9IMMcfIkeUyW3L7UsuQ39MeMwALB9GiVIzLSdzMGE7fNVQo4qkg5Z3fILP
ORAfXx91jk8PtDP3kQLjblpunbw3lGGIGNl2ActRDw4fUDcMzQeTzn5RQHP/xSqSeXXHLXfVRgZr
IIGCJ7HpIhEd2LjBOyCyEQOJRnEXZDdTSQQ5u7Fmbah0lpp3M3WFk5NBhpp/YqHcvrUfgzkItr0W
uk9neHxtrDd96OIpqoJSNZQRFzYMtL0L2AGIHAIMAHkr4wIpvk2h3qAkRB8xeqZsSbO01Mz2KHQj
3phUSY0jKNgtXo6cbs/rpSWZZ1BGQjzhJO97WB3ioaRFJNWOrTbhcoxdbtrhqFr5/T2p4uvZ1wpf
UMWLEOAsrej52V5kE4FGhz0YkdyvxTkyrNkVzW3Oh7SNY632xObsbXQsgFm+xOh6GeI7wvOlSqp+
UKGIBeEybvcMRvUaD9YTEUl0ckvzLQmIL4pWppjVB9BV4s1/49i0wz4aCPq7+MEeJme+XGf/hGAB
QzNyKmegB2teKCuBGT1Z7g1YA7CVHQ+bmmkwgvFs/dk8xVGg9SFuQOp6emN4RHYPNukDUPMTFL0y
sMEOGxV2tmASvO8FFwl6przyQtk4n2RyLM9EOKRZo51XdaOHmft1HYuGxzsEZqKuWGI02BnFck2j
OErA81C3r9v8L/fgzewhel/FRdQng1MGHUBRaqnquM28dv4YTU1733eCHnkPICHV1oQWN76Pyeh8
OGzC6vov2jLIA++vmNwi/UPTgI/jlfgmygkmc0T1lcTZyuw2APEuFtRVzPac5vcW3HNE0QqKPJ5V
qFHCn3+InY6VMq3vgeK5l5G4mokAHuo0IRz2Lmw5+zVa6YkRf6QYVnCDjwIN9GA2oqft07pyghL9
NkShnIl3opFO40oJhz4gYUAoYA6aAzLQ31zNT4MTsrsnr7ik5MtGMD8raCQ3n2qLav84TKb3PFoN
W0EhLIxngQZrEouvpmFZ0j7ec2c7CNpwGF29o0g2b/P+W+b//RbJZkxv+Yu1++vy95UcFmlX8Qkr
Wyq5pqE0ocJ8mMmO/b/MCnv/1CexxHMAbPR+5OYD2MjUYpWcenUt7L8+6XZaUpgociYZeIFRjNDm
fQWG5vxpTIANOP0eTDHVzUJTt9UWab6BZuzc2a/wut4bkJJvY0IEFsqoNGKsCXupJQ2o846pYH2U
ueGhHkc5YKzbXIJp70BEM5oJ/QgW7mvUoUSmDHliEHe7hKtoYs2mhufZEaNh68XYBCUQIZu73gRh
OseZGsPcQFcfRLYugGI1ek16BNr1DhNZVE8A3grIF2m0iBO394z4CGPTc34f8NRtUtHJUkypbnT9
i9aGL/R7DpPdR9SsNUhw6lA1HXKHMXxEjw7SkG07mjLvkmd3/jrWqSknPuWF2xsnFKSw0Htt29+x
zC++cMovwRcPWcDbyCA2rBE/v/ivJDtGQiDhunQK8eoYgZSYh4NPqThB0YWYKN+k1KRbBfpZIXzc
yBsfOSkuv/h9eONDkp3s8VRdiqhNSHtNK93wSwZ1DlcsevxbKrTv8rnhQRnMgB2i2LtBHM2i7JCj
HDeXuaScODOkuwVwIW+4P4b2nqgWchkSWLYTBOdn9ts/0RQPkl+9FGwTrFXXs0qeB1FPwLhQ3wTj
qGbwm/Rjp+6ADHUfI8EI15JdCiCHdFbLAUZh6da8soxZN5VN1ApcvM0l+MDGrNSrDDmv84JWAIxf
htu/Ex0kLyEXXfN7s3c6dOa7PwL4Nzsat6kVWxMf/WKN8M3jmYSutHgH5Lif+nqYEXiyWNP5Gn9q
VDa27awm8FxA3883quNvuqiQ5zSp5S10OmNk4VaRvL0rx2o8Brl13SErwOlHEXYTsvch6L5Tmskv
U2jwuOzyllV13iFRwkAO4jwF/d06MZo2yGgt0u8k0QQ/nbdrfugIrOt18b/iOX6V8ykVgUPBfvn4
2531GebM/CKPn2w6Jpzo4qT7bKshSzc/HijIb8QCEStH9q/CGJ+BluZUIdEQPbaOVJzsT5HJ23pP
4ZbWaCeMYmd/+Gvc4AFSM3y/3Xqfy3YzoxwlBVTrqjcOtSlBetyusyyiPgOE1ronUc27eq6EZBwt
9dFFNBmo0eUrVRuqWGH4OFnVqDpFzCXzS37CEKsdbnKSiQKGSDTsHhpvbZzUerB+Vv+P+ChfGHSj
jKaOUDLHCkhGpGni7egKhrZxJJ+K6L7+NK7BdoIL4o1tBmFZSGiz95J2fS9y1KiZMmEbfHwfp4E3
eylihaZD8TvhfLvkeIQjAE0HbMvB5U3n6lGr0dUQl4IwVjjT0pdiGAGvqi4pboVRqyyr5P2NhkPk
QiIURyTHiUWmbOP/YuOP90dzERVKNH6u6DQLgJn6OR6WGaeiequ1Od27dIwlX37R0ZpDTYgNGwLg
JQpr8wkAaedoj9m2SXnbMT+M3Z0mLPVRl5UvGsrXxG3cUx3CZzpXp0wI9gqUB7TAZmbzeaXhQFHn
719uRs6orA2NMOEvlFKRcI3pedkwbPpoQ795Otoq8vH0y8x9aDnnYLRPZjxnjvmIlEg+AmhBESke
i3D/P0eh2ya7RuqjO08HsbubjYwJV+85WED8ZZTnMoF8tewRoY9GUY655w3INvc3smtk/2JJJzJn
ErYwJhAnJ8eUgEw5j7tZPrqT7L7N40Ia7UYZtTHOCqupaDoreEb6RGXiLzM2YANgjKA0lehSC48d
GYyvyXBRJyVcv1MDBBm5kqoAQXESYU1SwyesfwY9ag3p1lHJrWZsZQi5BsZBRf14MkyxYpOmt6WW
BQgBD+zhAvNWy1jxA/e3Btcvx49dqol8tKvdqJ9d9vvIzZwX//v+Cxs54Zy1/w0rZKYSociN2NLU
5e17hRNVKBidiVn4kPBAuxa98U/TOJOPfezjIm+eq6NZgEiZ3x60zWvP09L/SN4LKVeKKppTpQtd
Lb6hp6Py0TpUrriJFFsef4g9l9VziLMQe+3hUCRWtFRkirnX47L2MPfwmfFEYgkWpJKISZ4QAxOY
s+O9CsicfDKusv7IprKeZVFuwqV/5J677JIDGltHoKi2fpX7HNLpOsJ4cNjlq6UWwCD3ImdtA92y
OO28TauPnnkUzF5uPuu13y0NwYFnrLokiL1H0IgFqIdmaW7jufRCvawW0gVi6wjISkP1SOnFqTG/
3rTvKvmSl5eE5jtjzGEkSBMWoBrtYPHjZUOvigywIOhapp97h/GWTptAarNbrJceZmnl2kjVEA7/
tAWRqPsDzLq2pYhJW+/7bR1JrRBybxxsh1Pl99cNgJEDSoAwp1LAgn3Fmg4kFTKTgOSwuVnBggY2
0ZrnLFqrCJCa/IQXUVsXaLpHhJaDZQf05vVnHdcXZSvIMve4B5OZ6eGABRNfMYPwkC2OmABML/Gg
Plsn/O5KVrX11wPkq4gE4z8T7X+wO5BK/0ydJBuR7sN+dsqn6lhrRL69qy30sPXFuCdl5q2pkVFg
bVQL+VvGXkEszCV3Kbgsp34LP7pz5EOIXPLCKK/L+41toz1MVgSNrdrajbbCPXT/5CGcoz0w0LcA
F+lJlLiEXGaS6dzD9PrXpojGhYsGSMJcr+a/2i6ZAZ2jcI64i3ZPp0qNAS+Olt9IDPJVHoWLf3JL
EgU0sa88wiK2MvIbXOGLQQJJ8zx/mZRZOoSgbAQOa14iNFTQw0P/fM5wxJ8VP4iunlUFxqTbrOW2
UnV9KnwUt6k6P/hF8+yTXybf4w+2hpUAoSk4mmL2PKOITO0+2niNnEo0mysNbEr/b2d2EtQ2Fq0Z
UNlV5pKT0VVc+ChbVbKqaBmEvTdMNkrX26e8vD8fyOuoU+w3B8pRO2Fgp8hGU7yRFazNGkFUQYFq
kL4NPl43eA0FEiqKIdz2pR6HbcJmddzPXzWZkzzqQnGpbmRoLzYFj+rZ8BHmDmj/48rBfjyshdFy
xAGxKWJNt9SO27ump9blpihU1ASD3/zZzY8re+C8dpdmd8tAtcnxRlJcy8rdXcZyAsXnrvtM+d9b
mBiGYtOfENOJOqAHOeG5wVBQu01gIh9/jKRcjgYAYkS8+MAUBieFGuiPdlSzuZqfBFbmpV/SBhzu
XwKmhrbb/ha1XWN0+MCVAGjE46CzPw+eqoCY9u0MIFBqJYfxhRMQOFowZ2T8GSBnNke+YfDmYA4A
m2f2knWUfdSiaE3KkomOf6/kNt2I1gFU0myiZ+utGGmPfaqbVGYi2f1zbEoxUstDZ7apCAvYdTHd
T6Sw8/Qhd6GWkR1AfxM60yyMe3tR52PjkqcZwIRk3Ix9KCS+OOX8EFe9byFtkB+rEyOPU3xOMZHt
51gDJ1XPokmR9DeUEQetRulAFy+U2SD7q3c04mZaL2pZVg9z8tjTRj2WzuimUxNReLHYEBeoZ2hH
KDBFBmYEd6ovwFlameYvZ7RDIRC2h/AmOrG3IfvauHqthUCQYxItp7hmE1vsQ6a+LWt6Ln0KPE/e
lolpYNXegieflSYj+Yby4nwgWs3OJTGNzBBeesTo8X4kr7XoV5q/Ghsn+QgsFZ/1UEhHKj3N2rR5
hMIBaiXGlvlnrg9CE4BP0mcZL4G80rhfP479ySe5SaaVgRGrt4hxkKoXTj95ijBTEjz9PEXHE+5y
BTOUY1Xhzy8XX/+KOeadhKtXWL5gdmNYYFYKQvOIDjlQhGtrt4Xb8i5l3frBXPpWpWQzbH5Atoc+
506KF/ya+e/SpHqqnvvMLmE9so2LBdtzlX+MvYbexYlxAICtupgsydZ3ZAj5GNJTKIhSc/Jeblk/
UtOtKa7QfR43Ua3u04GbRsofgk3r8QLVDR9xrs+w4Jq0UL+IQ71IPeYKbhkFRyK5BZK01shwfdWo
3FWwsgRE+gTPEzOjJaJQD7K8yRrwC4HuoKNfwx3XrLCZ/4Jeq8GtgiFXPRvzsYtht5X60oYJKcJ/
Gk5m9JEx4VKA/kkXYxbZvwqQeKid304llsGXrpzVp3j23TkzV5ij0g/6CViCEaUrzGNqB/tfZ7o2
+NTeNnM98XtzLHQRPwVA9pNQL25v/Sh4EY/VQv/dOQfMzEx+W2MpiRj8aGjJotcqYba/3escR7Uh
Uc5cLLIMcPISgHNtHF5ELOpFVr/c3rIJonoM8iMY7QV54tUckklr40NeShb77JiJgXk7haFYiJW0
EbfZsA4x5GxTZt4c4jzFbjuyrvN8pdlNztoehSXN3Oyt9gKEFlaOc1BRuOR6H9kV/j1lPCGrpZsS
vuH/x46qWRrg4tfzzpnJXLDkMLiMpaXy1muivgFCaMYfKkBoS5rdnLIErALPQkn0JNCfh+R0JrOm
2FzpfSlMdDmDyPeiOqh2DtRUhtYjz+XDvQhPCiKv+ymClEMAJ+AyMUqrtPEm9wNhphKYf/LGvpeR
lGzjFGxwTKX/hjfn/5R2d+Q1Y7LkvpbbqFKiibYyp/hJ4zUBIg9CNo41Q9m3gygl/txPkLZBC3YM
d4ftVMUnQwAzr0lEqnQc67G0SMxYniyhCdIrRw5gtgwCm0gbXtg0kbPHwCVCiB8PLkMdsmU3yBtG
NpuxQniy4cpardCLnqRnHB2BsmQd0a6aCnIZeamJarjUI7968cQST5etJaSX+YnqUSDmUzrPty5T
U+U3tpuI6HTW4mPZJTp+WK/tZgrZb8x4ENvSiyXNahAOxFT/FKc0iNwNrdVW8y8q7YiBix6aM8fS
vKJuzfyN7Mq45r0cLXsSbMuqavibLf3myNDafBNhe7BYEUpdmNXZXem0q9KcV3exuhxn4yc1Yz91
oXJ1cZ9ZZ16TVHYMKj8pEbhWj0ONKz7qq51H73PxiZRTvIHIOWCZ8k5iacVgfC+1XsymGDa7SWd0
6Fzcf0VVn8QT2I+rnDqodCL9rnr6dgl9z6QJcSqjUCcwUGQcnaCDfkEcLenp8103r8VSFVIMPoO4
0M5pNSYstgtROmvsdFi7BNuhLYYxxPUQZ0YsVPDJXxmg8lAFuGvNVycpcA3lZj7/21cRKezWKTQH
2C//ngjkjJxh2bBwX9tybPMAexe75bsH+WbpmvHupFGVcLRqAGVqfVG2mAkl05EchztMbt0wBTCs
nVBuLS8vux3ZkHtDkEusUgIf5JVaY4+uPqd6LzAKjj2Dki2XwWmYX1HbaCOX2kCATWrBm2G3DZfn
VbwYogbzoB06zRyvd+AQ46lUoNEL15nKqHXk+KElAKPI2ebB80uL1+ut1NxejbDq4DrBmIKMfZtL
emw0u8iKFmtasLuGuFEbNKaL5LDkhS2d/eLTdaWtqarAdhr06KqdCMcqjU0l6Z2UnV9ghIIhv9im
/rSltOuYNrYP5wB68h75XSNM0paugSO/okuVr5rcIfo/gT4SzmiKiyITvU4brk4kfEcO5LpjvFDB
YBDjSVh0EFpAiiW8tx3stKGjBdqCoVeYIqvFLFTPokHt4u2oU5SsMB3qLY4XWG7Ni/L+sbCoY1yA
RPrP9YR5FUPaJ2SypxpZ0/OzQcSDl6Tv4ymWN8ZaK0vvbBqQx4Gu0KUfV1EIJzPtD/9TodBzZMex
Mnmhx1/lPWCvygcoiFwb6n55dU964EZZ/NhrfGrRDkviEcY9ZP8pAyiJnpW/ak9AJLljwtA4ik7X
nNcwWgNALkNd9yiBVAZIAjUqCwbaYX/ylUQyWujMEpsLnHCXXPLJg4nxyPMNo/AJSnIjx+A3P+FE
lWckp3oIJSVZfOgTiOT4CB9W/8dMQRvq7XGApOY3Ygnwm1m4+2+JlT7hQQdPqDYOmgHMngqcthbA
uzOFJkTiEr0DFrdar26wdWW3BnQaInnHi2ttuXLwn9fAFf87fVMm5mxvQ+PVNHOX84Zx425mB1Sl
RTjG+snA5UesORQODxwwbljoB4jgw7zmjg3HqU3/gXV2O1pMkSWWeRuLk9jQ1db+yO/r7I9gawxL
8hkHhywDHotZQ9zlIIOW2Mhq7kEthL8NulkGUWmB3A8cwgCbr1j3bnx7YrVbd7jXPkhKX4X7Z8g0
0LvqnHIXgPQVuN2UZC22NmVh8P0+ZIFd6EwrQJnLdg4GQbtvBNmXdfJrYQ+FpAYLJvcEj3I+wAEy
gbotrn7TF2OD0kNbe2+un6hQwlWUJbB51/MMdQo2u3twARipbT9Q4Ea/YGt50fThfjelBc20aILr
yBIj6xXkPH3D8BVQgpjraA2ewyX1m+VTIG25BKqb2AtsUJsg+3H39ntByyDQSzPCtaaGowhgBkBT
8V2J3b4Z+ABQbMjwsa/28kvgIQjCuvXAEaYK+8OFY0JNXPOhcHGUMBFQIpCIOWGi8AYC+9KjEAJt
tUZ0ci0ixDS9JaypVAO4iKs1zZJB0HCaGUXRK+htfXuA90O09vov5q+ctBO5ctWcIRwblTMRi2Fr
2epVs8wo2Qj5zPjj8zcVgYXOKs2Q2swCvJFOaFg/TmVCeE904dRkY2KdrvOjb2SyAISpYcBnNPa9
62l+TZbcaqO6ftBrFo1VuzI7VT/hgL+nijIpKLuEHr9M7UFqLWNXdZJ/egQ9LA5uUO6pTRrcnG7/
OXxaUqAGLf84WbD+wv1a1ArZRmeJa44w5ko6cAUkGGktj6jj2ICTcxeVrUvp0CV7F09QrNHKGVLj
vZmcYqX5ZG7NQG/WA9uZkmL/oych85AY9reMketM957dlGlXfmYcqJe2B56LA2dR6uUqe+XlypIq
N6aUUuzk7Mw3sJFQ2VAKZApAWUXnt9PMPvuzQKh1ePtkoX8X2hjTHo/jFfrvj/Sg8YRVeE0pl06m
TYpOeYpXmzdZJa+Lnr7QhTIDcxJqW5+LuL0KrEqJPrCKoBJkJNHxdTR7xuIHy/SkS9YR0nCGLAVB
XYU6NJKvNpXvERTpm89W4n3yjY1ZdWM/TKEd+/5+8c/oyWxdXwOYQOTB1/ywELb9Tn814mqDpOUJ
yiObZyo3I9JgGqQLHBbVyr3YNjS0RfWb11mX0wr/GO6N0ORt7arYBV7pTM6PC80h4D3cBAynHW2W
VtDDLDYJWFPY13KAcmbOB6NLheBEvE634hg6IZ8G5+Dfs/zVYRcns9uvfdCohk0KGDvNGArzJNBG
Cb3IcRt0yDsBsJUU1PAEiNy2BH55ZA6qSpMvAzfME1Z0SUD0tq2LgqmaWVLnsoZ73JL7UoPKVwL/
lUKboJDsJ2UpQPMJAh0tsZVY00eKF3uePjb/Wtr5DP2XRlZyfjmZLufzTmUJV9Fu2Qf48BS31/R3
oftN1gVKevUMZ74SzyfgfcyPdYdsYY9ka6e8xAy4zBNt7Gg42+o+ycsPec3YZSRAoM2TOZ//onlB
XOkcSJ1gLFrtMcdP+akCFaJrcDAMn9KwH9qyu7T3R+MUuyFlZo9z3kMuVrjIXKG4yNE4Gq3gTg20
cpYaHK6ByrDdUtGEBKzLsZDKLv3wztdGKKoWILNADvp7dfhbEBIWllPquusFx+gTNqmQZDuI1BNJ
GXxzbriZWJqG+anjT/WIgulAZBpoHlK9MgKqpTW9SPIhZe6Z/DBf6dmdPX/pccKebUwWB/gFBsj+
G6TT0NpGVfKM+DzboSm83JTTjLKZAQvUBuUGhsdioRjILhDqK9z3d4Y64ZrC4WBz6HWSz4gpOg6n
ouBDKZ2tvpmmv8QX0vN2ccuby1khuINAGOzFBlm65HygYG8YKzQt03PDDQnlOgewXK6SOcJeErik
0ILlMAhd0bWAD2Io6bW3rBX4aeoCittZ+Em9pWvtIFadu4wfMR0NwTnsHsNB4/5ev/JZYaCuRlTl
lldH2cTL8lFDdgRI91D9qqY2y/nP5Wyx947v7t3VRlnfmnq4E+Moql6MRF1osoPlzQdIhh5MNmE2
UuRbzJ3cUCNiIZCggrbIw4AHt2Jotlci++jsIihuIclu71bbXa58KKewMwzmZF/cOFKiXckl978l
Oy9dZsoE7nfUgdm+OjICaw1JtIO8jSt97OnHmGHbg6TaHeoj/cN2IFkaoM1C+O4/iM0Cvn5Kwsdu
ALW8FpG3B0DU/PvbkFMbEmrCfnCHkHPF1mF/kaZkMwX3XKWcVmaZKf0BtVwW+4b6vCGPOXRaXnDp
UeI0U3TUbBzoC78Nu8FX9IIl8VxJSMDWWB8CYt1YwjH2lPwhhco8TPnBA5/r0Zg+9XJ+V3Pxb+ly
3e9R5xYbqJw7t981UNgLGFARZ0yK3DM02Ghm8GHjuomAdbEUCFtmkSYNY9aYFS7xJh6mb6M7NSKw
4TE1tp4z1o7F85IchKeQgQ0HwCrPFXn2EH+Pj1lIx/Y/mIe3+i08KQlavxbBI6/fBuAhDp5Eke5F
wO4nXCQ8F8BLMoHq6Qz1JcWOh2pzPz+dnu/o+Ilaxp2A1ShJUn/SKyVPCcf0vREU5d3n0n91xuX0
WcdnM5JzPOmytRa/h3ANZep+1CQKjwRwQW41UIKhqN7SF5O++ZxlimUfYczYuft4SgkYIjHsb4gK
P2Bag8K7w4U+C86zOwBrlk/mlgMxUgBTs+SnmXmtJ/5G8X0gdKEh8kObMmRShXFXbVtD5cl7Q5tv
1szOdDyIFdRnBJcY9KkjK7exc8UmnYgz3jR2VkV6pa146ZxsTdmWyzZGE55GScFIqF9eby51bgL8
mtyvDHFTdEYAI7TrWUn9p3g8ZEaI3GLsBdqP+MI2QdRyGU0ejmxHTSPSgsD4Ahv/aiSVQK6uwF0Z
lFBhmVEB1nSTSeiHKk7OfcdVwhGVaqam3fp4v+Tb98EtG0wzKIFKla0O0j24U0Wtz98i42262/mY
WXMCKwuIiRDIaRb1GugbNT6o4FYokNGB6o4od9tNuy1wC7QN+8MuTvflQ1H87O03xIG8YnI5pj1Y
t4NsDx39fPj1R/RMU3K4/fXvntaakF3G9H46fhbIKCOgh9L0o2EgbMYi1fuHSc4uiJC0JVvEjymX
JpqDMnLSyBT4Ppj2xczEBaSVw3ydFGZ/16ZCIt2kdM2dE4lQxW1/HbTkYkiKfF8s8JMQx+v4D01r
6LxewvZOfksJ1P3w9ctCH6A1S38h6Dlb7ATsu5cEvtsIhdL/MYdKf5BYdZZv7Q2fpC98AUbiMzXw
LKDGVBdIC9EFVjmhyCinMT4fxFHLOA9l7NBM7xRsPXjXm7uXjFjX1wK+92HOtlfGpnf15ncOw3am
hZM90T2u2W09NRL0eQD999kciR83xPipPxUgo8OwAikbSkA+wOBuy7qvV3xhIoAqSrNE+NGBQEdY
8MwNaa9h0UIEK6PIJPn2J/M6bJ0o8+up+5PSFEV5OzW9Jf38QPM2yEOMAEtIH2Eng7QmBVF+v5Kv
SSO+qnrwgC7VbmecFESYi/h9g1fsEJGIUAYQhan85pvFFf9iTX8IlFVSQQ084+gO3dFoWA9VDk6N
1+6BbjighuVBQuZWiLOzX+YDzpCu2tDqwroZD8514t3q2OcJ4N5Jjb5AIkt+TR1mr1CaZoKW8hfi
/pcf5vJew8We7Jl7S/rpT6Sayo24xBzSn+X8Ybbc7+sob+LOD9Qz+M0YXiTUccAWBlUQdeNbuJc3
7lzkrX4eSLqblgPfLKjPM50VbfqGttcKH/3Bdqee1RiSnieICByKCjxn1dW4brkqSOGPzJV0Ol0h
jfcUtglQ9aPuG1ZCzh/8WIuCSPkQFfBsCmn7+yPepZJDjsYCe5DlqUezrXIlI45h8XdGTVISpkbB
JhlemdSh/s+cEiMKJDwarACVGWfT7ZtSBqeKtdEvqIcgnPaoIph4YS15pApA0ZUybIv2/Au1+2pf
ndLuGKWpDtO84QW5dYp39hk6tilVjomSdqhB8/5tOu9a8tNLMu9WfxdZuTEccdajr2wtjNiC/hue
sF30IPy5qZs8EeIzWPRhkBMk9opI+XF7GVZFH/66xYtzKYOgLlz/W7dG0RyvyygbNKXvqcXkUcIP
ajf2dZMm2nSZC7vtseAXSvqq5dNCwO9vLHkkbFX17F5C3qajDsQf/De4PevVc+CYpolJaI4K5Hx7
XDmZVf0rfp0frHktDy2wSsg2Ot7qWl7wyPfuMPlhlKHw8trxpGq6Y6busnXtxF0SdVfJe4HTe8aK
FH6tJiXYYE4dWcH/OcalJpkfKH7SxelJF8QxMMggRzp47NyHIt7/z0YzwtrBG2yzXoe3NRVPxHrr
dInUfg30wQxYQ7L4rHm5pFInyTXwogt4eGgQNEPnJYfDLwqARIkzC1ZhSAr6ByYXh+pq9sRDiZIR
mSfYfMRsqHjPOIaG33o0H8aZ8MdTYtitY4IyfvBCOYO+QwlCOhoxfnj/eTCTCXdr1QUvegKAp3bT
fFpW9/7aXpcf+88W2u0Zoyc2luenBs5MDLoDOn5S4ylH8zG67/0TldujjgZ3DF3n5M4LJ1wN3N/k
Sf5zXxctSnt9JFqyQSmludSLMvxIBkMQOmmZz/0pm7bTtV+66PFxZTsQ1CHbOmrCsgzJp47jWqVn
AZPV3MKNf+BSl4suHep+3dpedU75BB5mV+Ed+jJLto2OG3R5+q2jAvwN+zSjYk9DdMI3JnE98adJ
6zWeEMahTq2yb9UJN26KfSszxFVLdv2EgD3MK/jNjsPM4y4Y/BarZII25ArKEPhLyoVTSwKN9sXz
XT5TCTU2jopSuDgYKGIQ5HBYKtKTJbPyUrm/gr5Ym2z9Fy6vn3aBmD3maDQAGv+oYJqip395NuRk
pO5AukH+lmSgYAqZ9NKi1n5pQ3LZZ8QXrakTWR5othHszHrk8D+TVAXY76sKuCRzZixNr6jMW36V
uFw+CvBX3nftYN2SvCekLRzOr12LPvew/HAgHHK82FAAhGfV1Kply1XMGgNwLlXckWUwf36YM+dA
2mUYNr4192CvlqGZHK4nv5K0y4M2vaKH+z6SYcQk8gu8cvA9WVF88FDXEJmbbhyHMrjE9TgTRpJ1
xTcgz65jzfyC9Vvo93MEbZ1y39ObYA0RERO48RJK5Gq6xOmDau+AsYEXm4JLpKP14qkp531fDVyg
3KvPosmSeLWg2wtaCtxq30q/hB0dfTLouM4WLBObyczhK1ujLwHckx4MMEkw8/JbQWjM4fueCZBC
eoVDxiH5bueyMZ/5moRWZUeViIwiiB1uPb4snxHRDq/BP+uZdUQAmXdkgNlGtsTSSZy9hhg7351+
B7EWh8GMcOCSH8Okq+9MCDLAUiL+x4vwU0BQtDpSGqc0OXK75f+rRLOsDp+sJ7tdKhU+g/E5Bl40
gzOsMEDWVoqP/tZSLEK49w/P7fkFKbnlU9Y3LO7htHJAWB46ga1GKIFzk3EXOieOFBqYR/E3ESsW
FWTr6iH38OhZEHq1bJd37OGv2ZK54RR3AZ7anOtpZ/x3OiDvV8nzWzSJc+rQyIOa5VKNnMAzhDLe
xFD9uSYh4oLWWNaSupoKHJOXgtZPc/m0mgDmcSdbjKidygoPc0sDCMBXODUedMZjgultqV55+28m
2c9ZG6pIWoQSiJTgFKoDj3IZ0SuF8wYKCCiPf8B9RA80UsDEuWFtre98MiZadaBgySI289Fxtx/f
p6+4m9ZYrw32phmxBfQC7v8vepFnQSKnXtYU+Ic3IT9alQVC8M8JU9+kTveDiQyu89lVyK/mgEk8
mOIS/2bI+gke10qdvUbnTs+WtEUWTLW8kibmEj5ZxEAgli3R3PS5GpgZfENu6R4HgxIX+Anv9PLT
2XTf2TCq/pI6bhjL49LaWQBBjgXZjJ9AiYgiP06unzCn7AnixoaE+6jrCnC4DLeRilyqnNfX3QMY
CzVPyp6rUJQUvSIjutWNatrE31qM3RcYg32g7dmqsSp/1quxNnhu4VQvrEFCKaMApn215T22JEt5
PHCb1W9PZR0YJQKVjMBHxHLk5XIlzuZ6W4K4icgXtFWxXtp5HxgfYTUDdaqG2frcX+0KwLLwluFN
DpnDntQG6vcg2g3bI+F9/rjPXBAgod2sKjCaGzjXSewH6UvgfXtMUiCGBJX3s85i9/AAotRZcUVx
Ut718L9b7TFgYxxcTUYIdoc7zKQGkH4aqxkWvcSPheKez8aJsVDgj5ILIJ/kO+adY3VA148pFiJE
lQJRC3MS2SVZRbZfvipbLeUQus/h1quWHY26Q/Hp8ASi+iOeyFnmJf1dFQH9DTtOHNQ1n9PiobVJ
P46EEr5iQAAj0c/TzRcpKF89hoezAJT0fmT3DiJ8tnmjAuaKUNXm2rWXkDfBOucfo+De0ZEH4LTu
JP0bt6NvRgkmnTvOuL2QGoWf/dF0ZkkcvP3NBzPlv1DMbH/COohQ8Ib1rQZL0w+WeIpQ3xqiCoEm
hZ5uDkWyGYXp+4E1hownRj4L9DIsK4rGI4D5y3rT4OFicl7ByAfCVhGmkVzXl6J7QdtES2fWgzG8
jPSWypoONm/DGeIn4eKugOkACCQ4Jv4+Ozwc3lWEto73F2bqtUA8NOCfdOfFpbihZWdf2V3JP80f
EumbAZ9P0IiCxISziXVF1SoTCn7YVCLrDzwb6vU1EmXnsPmf52WD+pfEEH3fZ+1Z2DYtkpMv4v2D
IzTcDysC5rvRp39pMVC7bcE03p6wLpe6qaELgnYbCMejA1+uUum1jr3/vdqr649RpmzHcDQKasvM
/yzWnRZZzKoyXMBc44VetKbPfpgxfTpdZdO7CTH7TXT+K4SefLQpGhsJ6uckn5ttD2cflmDTJ0vr
IeGL26wPOtRw/SSEBrHfj+F/hxf4Jfzuje0xlAgoidq+RTFJo/VJwsluHeVLVt/sj6vtymw=
`protect end_protected
